//------------------------------------------------------------------------------

// This is GT common file for ultrascale devices

`timescale 1 ps / 1 ps
(* DowngradeIPIdentifiedWarnings="yes" *)


module aurora_64b66b_25p78G_gt_common_wrapper
    (
     input  qpll0_refclk,        // connect to refclk1_in from example design
     input  qpll0_reset,         // connect to reset out of TX clocking module
     input  qpll0_lock_detclk,

     output qpll0_lock,          // connect to &txpmareset done from multi GT
     output qpll0_outclk,        // connect to single quad input clock of GT channel
     output qpll0_outrefclk,     // connect to single quad input reference clock of GT channel
     output qpll0_refclklost

    );

  // List of signals to connect to GT Common block
  wire		GTYE4_COMMON_GTREFCLK00;
  wire		GTYE4_COMMON_QPLL0RESET;
  wire		GTYE4_COMMON_QPLL0LOCK;
  wire		GTYE4_COMMON_QPLL0OUTCLK;
  wire		GTYE4_COMMON_QPLL0OUTREFCLK;
  wire [2:0]	GTYE4_COMMON_QPLL0REFCLKSEL; // select 3'b001, GTREFCLK1 is the choice as input
  wire		GTYE4_COMMON_QPLL0REFCLKLOST;
  wire		GTYE4_COMMON_QPLL0LOCKDETCLK;

  // Connect only required internal signals to GT Common block
  assign GTYE4_COMMON_QPLL0RESET      = qpll0_reset;
  assign GTYE4_COMMON_GTREFCLK00                          = qpll0_refclk;
  assign GTYE4_COMMON_QPLL0REFCLKSEL  = 3'b001;
  assign GTYE4_COMMON_QPLL0LOCKDETCLK = qpll0_lock_detclk;

  assign qpll0_lock                   = GTYE4_COMMON_QPLL0LOCK;
  assign qpll0_outclk                 = GTYE4_COMMON_QPLL0OUTCLK;
  assign qpll0_outrefclk              = GTYE4_COMMON_QPLL0OUTREFCLK;
  assign qpll0_refclklost             = GTYE4_COMMON_QPLL0REFCLKLOST;

// dynamic call of GT common instance is here
  aurora_64b66b_25p78G_gt_gtye4_common_wrapper aurora_64b66b_25p78G_gt_gtye4_common_wrapper_i
  (
   .GTYE4_COMMON_BGBYPASSB(1'b1),
   .GTYE4_COMMON_BGMONITORENB(1'b1),
   .GTYE4_COMMON_BGPDB(1'b1),
   .GTYE4_COMMON_BGRCALOVRD(5'b10000),
   .GTYE4_COMMON_BGRCALOVRDENB(1'b1),
   .GTYE4_COMMON_DRPADDR(16'b0000000000000000),
   .GTYE4_COMMON_DRPCLK(1'b0),
   .GTYE4_COMMON_DRPDI(16'b0000000000000000),
   .GTYE4_COMMON_DRPDO(),
   .GTYE4_COMMON_DRPEN(1'b0),
   .GTYE4_COMMON_DRPRDY(),
   .GTYE4_COMMON_DRPWE(1'b0),
   .GTYE4_COMMON_GTGREFCLK0(1'b0),
   .GTYE4_COMMON_GTGREFCLK1(1'b0),
   .GTYE4_COMMON_GTNORTHREFCLK00(1'b0),
   .GTYE4_COMMON_GTNORTHREFCLK01(1'b0),
   .GTYE4_COMMON_GTNORTHREFCLK10(1'b0),
   .GTYE4_COMMON_GTNORTHREFCLK11(1'b0),
   .GTYE4_COMMON_GTREFCLK00(GTYE4_COMMON_GTREFCLK00),
   .GTYE4_COMMON_GTREFCLK01(1'b0),
   .GTYE4_COMMON_GTREFCLK10(1'b0),
   .GTYE4_COMMON_GTREFCLK11(1'b0),
   .GTYE4_COMMON_GTSOUTHREFCLK00(1'b0),
   .GTYE4_COMMON_GTSOUTHREFCLK01(1'b0),
   .GTYE4_COMMON_GTSOUTHREFCLK10(1'b0),
   .GTYE4_COMMON_GTSOUTHREFCLK11(1'b0),
   .GTYE4_COMMON_PCIERATEQPLL0(3'b000),
   .GTYE4_COMMON_PCIERATEQPLL1(3'b000),
   .GTYE4_COMMON_PMARSVD0(8'b00000000),
   .GTYE4_COMMON_PMARSVD1(8'b00000000),
   .GTYE4_COMMON_PMARSVDOUT0(),
   .GTYE4_COMMON_PMARSVDOUT1(),
   .GTYE4_COMMON_QPLL0CLKRSVD0(1'b0),
   .GTYE4_COMMON_QPLL0CLKRSVD1(1'b0),
   .GTYE4_COMMON_QPLL0FBCLKLOST(),
   .GTYE4_COMMON_QPLL0FBDIV(8'b00000000),
   .GTYE4_COMMON_QPLL0LOCK(GTYE4_COMMON_QPLL0LOCK),
   .GTYE4_COMMON_QPLL0LOCKDETCLK(GTYE4_COMMON_QPLL0LOCKDETCLK),
   .GTYE4_COMMON_QPLL0LOCKEN(1'b1),
   .GTYE4_COMMON_QPLL0OUTCLK(GTYE4_COMMON_QPLL0OUTCLK),
   .GTYE4_COMMON_QPLL0OUTREFCLK(GTYE4_COMMON_QPLL0OUTREFCLK),
   .GTYE4_COMMON_QPLL0PD(1'b0),
   .GTYE4_COMMON_QPLL0REFCLKLOST(GTYE4_COMMON_QPLL0REFCLKLOST),
   .GTYE4_COMMON_QPLL0REFCLKSEL(GTYE4_COMMON_QPLL0REFCLKSEL),
   .GTYE4_COMMON_QPLL0RESET(GTYE4_COMMON_QPLL0RESET),
   .GTYE4_COMMON_QPLL1CLKRSVD0(1'b0),
   .GTYE4_COMMON_QPLL1CLKRSVD1(1'b0),
   .GTYE4_COMMON_QPLL1FBCLKLOST(),
   .GTYE4_COMMON_QPLL1FBDIV(8'b00000000),
   .GTYE4_COMMON_QPLL1LOCK(),
   .GTYE4_COMMON_QPLL1LOCKDETCLK(1'b0),
   .GTYE4_COMMON_QPLL1LOCKEN(1'b0),
   .GTYE4_COMMON_QPLL1OUTCLK(),
   .GTYE4_COMMON_QPLL1OUTREFCLK(),
   .GTYE4_COMMON_QPLL1PD(1'b1),
   .GTYE4_COMMON_QPLL1REFCLKLOST(),
   .GTYE4_COMMON_QPLL1REFCLKSEL(3'b001),
   .GTYE4_COMMON_QPLL1RESET(1'b1),
   .GTYE4_COMMON_QPLLDMONITOR0(),
   .GTYE4_COMMON_QPLLDMONITOR1(),
   .GTYE4_COMMON_QPLLRSVD1(8'b00000000),
   .GTYE4_COMMON_QPLLRSVD2(5'b00000),
   .GTYE4_COMMON_QPLLRSVD3(5'b00000),
   .GTYE4_COMMON_QPLLRSVD4(8'b00000000),
   .GTYE4_COMMON_RCALENB(1'b1),
   .GTYE4_COMMON_REFCLKOUTMONITOR0(),
   .GTYE4_COMMON_REFCLKOUTMONITOR1(),
   .GTYE4_COMMON_RXRECCLK0SEL(),
   .GTYE4_COMMON_RXRECCLK1SEL(),
   .GTYE4_COMMON_SDM0DATA(25'b0000000000000000000000000),
   .GTYE4_COMMON_SDM0FINALOUT(),
   .GTYE4_COMMON_SDM0RESET(1'b0),
   .GTYE4_COMMON_SDM0TESTDATA(),
   .GTYE4_COMMON_SDM0TOGGLE(1'b0),
   .GTYE4_COMMON_SDM0WIDTH(2'b00),
   .GTYE4_COMMON_SDM1DATA(25'b0000000000000000000000000),
   .GTYE4_COMMON_SDM1FINALOUT(),
   .GTYE4_COMMON_SDM1RESET(1'b0),
   .GTYE4_COMMON_SDM1TESTDATA(),
   .GTYE4_COMMON_SDM1TOGGLE(1'b0),
   .GTYE4_COMMON_SDM1WIDTH(2'b00),
   .GTYE4_COMMON_UBCFGSTREAMEN(1'b0),
   .GTYE4_COMMON_UBDADDR(),
   .GTYE4_COMMON_UBDEN(),
   .GTYE4_COMMON_UBDI(),
   .GTYE4_COMMON_UBDO(16'b0000000000000000),
   .GTYE4_COMMON_UBDRDY(1'b0),
   .GTYE4_COMMON_UBDWE(),
   .GTYE4_COMMON_UBENABLE(1'b0),
   .GTYE4_COMMON_UBGPI(2'b00),
   .GTYE4_COMMON_UBINTR(2'b00),
   .GTYE4_COMMON_UBIOLMBRST(1'b0),
   .GTYE4_COMMON_UBMBRST(1'b0),
   .GTYE4_COMMON_UBMDMCAPTURE(1'b0),
   .GTYE4_COMMON_UBMDMDBGRST(1'b0),
   .GTYE4_COMMON_UBMDMDBGUPDATE(1'b0),
   .GTYE4_COMMON_UBMDMREGEN(4'b0000),
   .GTYE4_COMMON_UBMDMSHIFT(1'b0),
   .GTYE4_COMMON_UBMDMSYSRST(1'b0),
   .GTYE4_COMMON_UBMDMTCK(1'b0),
   .GTYE4_COMMON_UBMDMTDI(1'b0),
   .GTYE4_COMMON_UBMDMTDO(),
   .GTYE4_COMMON_UBRSVDOUT(),
   .GTYE4_COMMON_UBTXUART()
  );


 


endmodule
