`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JxjGnnmd6LJq3SXIeY6qlNkJsWotmIYRzAmIW6gYOA7dCRJVxAetxNh37eu6dltottLKn62zuKa1
SGH9WVveSQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FeCmbFsuyPSt9zPMXTPPWEazv4BGe+0S+0aNSx+PxIS8ud+EtxhO1LZM1clsm/BNBtKVB7aP2X6+
rSANUcURhwYfh3j5q+v4kZSZZe+EnOner9iM07L7X7WBv7zhvMEJO7NegXjiucqGnIW9msZfT3Jy
9OjeAizAsuNmZmfntJg=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DMTAPfPsDW1MQL9OHleXXNEYswdWG5kjbAwzF+iYLog1ixoqKGpSY2osgzCHQlY8SPRYVV6dtJ/c
Fpl4s6n1YQIfgvnzRGQkKSXd9HJxem2NNhTzRu8QVikoCtEXcGEe2qn01nXHftpCucAkrSOfFEdU
eKki5oM7ER6l+RnzX7t/u8pRXAZ5TyfbHJt2IYT4/PUjBYtyKHhtLCZaDgyUSSmbbfCbLPnZrqgv
pbK1PtaNAhjD5OMdGmiJrrXZT6SQevzMDYxPwb/k8yfcn8UY2PeXWGHx/zqMa2dDy8PGUjGkKWzq
mhc3yuGhkHDfjVj6AwCz47IifZ0mytnMH7syfw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g3XK6Bbke46LB1M5tPDl3Z2IL3aWinQMS9k8CWIci8FXUAnGQny6Wj/yAu0hOAnrgLfF7CDW9mpt
S+uKY1RGkqDI1201D+PVlVkzh1AYwGdjl5V3PiNYoX2DLg1SIy/D8HmAWYDguX/vkiNN2mFAZPl+
Grdv3UEWcpCbJySGz+sl8+Z1lzTRRYuohJMLig1aQTBAk1pto8j1shys9eXrIcBaAQkQ2Fwuve5o
Kov9THat1ISs9gavkbfUv4Z+0AyVol9VLMIkjE3DQvHpAiRzOHwRFoclOsS5Pu53hrofzBnLjA6b
IJ8/1hlrlnAsFSSAgDTZaWfbTCjILBFSbunaow==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cEjC7ttWioNxLTCv48rH/kCgwmooGdoWoFlNDl/WVovS3ozKJuIp9ESR8ai/y/TV/atT4zh8KGyW
CipyiEcrqOxGzA4GvOZbnYRc0vSehKTm0g9EEZG+aaoFtbcVmhxI0t4vnGSTYErISkYillyz50Oz
GZnwnkoDYDrM+PPRSXs4e10VG2N6qXZLIplEFxor4MDPaWtmnh3eJPsju77xfxX4p463j/pxXUaq
8coIPxm13ThnxEapa8DYsBTmDlD2oBwaYv0rLUKrESX3r+7I3pVROwOZMwGgB0aNaZsVhMzkV1+C
hw2lhh4D9vcmmmUx8gjYtVeAv9wKO1Ey3WYWCA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
h+zlRM+6FU4PIWYLeR47HHRzXI0SfXNcNsE8KER+nct3NTzY0+0an05sOoy7FyogYtyz9ckQ4tGQ
TWZuLTlOumOCFDs4P2S5ErEG79HvtUWX3wKEveRgkRZcuirHbbdJDtma+i08mEDkQd5Baf/36JTC
cmBTxwQo/tuUqh5taic=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jtifFEh6xFFwW6B/VeypckjWmrS4PykwwFJGptGJQdIhJ2nj7VMyG2efrHIg0Q8/RHe6zHlBuQX8
YGCFVyszzkTxsSVHNWPCC8tllj07+PWD1IIuvc3VFQEzvCOqlV9b/9lzNXAXRjx/Wy7kuqSY0tGr
Rh/LUwc1JHZsQ5oGfSi+2/wLiuRRarqnl0SfxIJXAbKEa5KsjZOwqB1f4PjKO09q0lkIBReLEmuV
5uwuA5jXowTbAI5gqhb5X6Wtl7Pg0nHZUP0GJepC0dydhQNHu8DAUh2KjR+cyx9y2LkUQAM0b6/m
njmb8uup2ybhMkfpPVzyKxpTV74f7OvrbnTtXA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1814000)
`protect data_block
Jn3BAOp3EQwhXj7sKmBXXiFybcHSyKrBpNrjPfIdH7FMjVufBZ0hnECAD0+OXLbAdxdS3Ru8xsYW
3OwnoaWV13MBuYDNglvrqmzLqRwCgBA+p8Y6UIUdDu17NuCtZiU4JycRwstbkb4CJOAUwI+JZmEQ
NgpoI3mteDwB5qTlwEKxbIOZD3N4Kso1FL3tup/6PcFWmetc1HzsMVJyhZlS3+tvOLQ+AipBcFKV
GkreyY832SieDNQeVyCxrIxAhlfRgZpn1EdU0+4k7J+hUzN3PHxbsWh3HKMlP2pBLGSyK6ojNlYS
JWIovIQV9ToMEkeXCiTgYMYI5UtksYHMinoVhAKSXjHEcYj+nGIIEC6m5XTdCZHWyG879HxWRYVg
TN+oo1SWeOt+n6UFOMaThpLnFEhZPP4malHGtNN08yHVW5Y1eNM1HW938FNZlq4pWxjCS2b+QSd5
2jlZojc+qcdoMbbOksvSg4j3n+ttVYGqr53NFlySg1eWuGVkXA8hpjWI1joHsutmZIrdttbpFKWD
wJ5D/6gJ3DagdiyAacxv5B+o5nLCx5nvWMQeEn3NNw2rASGpvfOnx3BErbZlbIYP7ZbAlCiCoaT/
xjgbt5k0T15FP0zSlKiv4W/MF0v8KaAR0AszqTW9y/4jWbf15IGs8GkOs2oZnJ5723ClC1NeyntB
rY5bIhThNMrGVAQPNZBxCnt4ChsgEbPvW5mKKFcNX9jeS3mvtQQ62FikFiFFaa6hR+A6LUiXJAAY
GQhCWFQrSXajcURDOIg5PSBNhqkxRv47VQ5OhUM25RdPR3vAyxVPwvQ0G+ItL5iHDOrARNJ4J9UQ
RZsCYNA4Js7QXQOyH9dOInMCpcNIaO/rgshtIhYB0N5LL/lX0iOCl6foJ7PzgaopKgFEWE6Ea3gA
bchfe0ryIOL/Zbu9LdHYaf+6kkYuBvow+jJnKuXfC04ZY6nlUHzccY/q0Bq2FiqFXKYZabFq83mb
cZ1F1ScLECKWDoM+mxb5Kk6mmjnI07XpVuuvY8iGe6k/NtMB0jm6mqkzP/AEqKD2fd4wZNBB8Hvh
OMkNZ9OmpjklL3leZd9M4CXiwiIQ6AnffC/UQMsf01eSWFxoNOBtRCGFA4dDcSWHAIf7quuqfy07
Aa+3Gv5XaSr5SHqRNo56q6i8vVY7l6dTj2VsuyMky4uXjmKNCv9q02N8Fh2jI1RnO6BPJDWwps9q
HHKJIt3V+Ceggwj70Ug4BgyNPh4HmFo5Ld54Ow9BUzRs6C2+q1NQR7+NH7hCPP9GixHPhdzm7AwO
E8+1+cG+ydmgKOjzpoiU8sxSUJueDcUPLlir4O00z189Lp62GBNtWFehobzGQRuRxqJ6L4c68PiC
ASfPkcK4WWUsKuwOYhOzL45BzXDdSQDUco8jP8aG0YdD4x+P4x70gei+33phuCaim1XQPpzy3X5u
8hCWgjZNM1+gMn/laBTJ4aenCuPJGTj/5pYa616t30QS03pFlHB4hsh36sTfgB5v8UJYIGz8ngWE
Dn9RmkvyK+/+ATfxy7hK7vLweaOwquFNXgL0g0bs44pykliEl1hNrVE9v7ntN295BFvm63uGcPlR
tz321XnENQ8l+YWKiKVRBXTewY9pAd71pDB1SoqVyosgik3RNvl6/V0hnEZVLVfMfoI1si7vYycQ
gjVSdrHZGTv59u0Lov5DUf3cHU9wdCV66v4P4oCYCjnXMiFURxm0rRZnqnokdFswZYBjgP5n5UBe
OY47hVYRm4MmvtBiySjR3sJYV67Z2PVNiWLBAaEZkPqJbkjhLXp0p1yH786loSW0AsA9C/wmU/uW
00hwPmET6Fu9bB0NwlKXqjNZbv8nnhb/L2PHvh7wWcxXMTSvDhWm6eILGlhn9N/jdwUZf/GnaPeA
FmuxitBLKiwn/q/zed2HQHbHhDMC1ueBzARYQsEq3vmYh6NhsUxin8GIJ6e+v4ADdyFEm9U61mYi
rbDLu8gXUj14V5qUizR3veTK9RaEw4d4Lh19NGYS2Z0W0aOjy+kc2L6lBfaiFzbCXn3yz/0mMsJU
n7e5SrCG3RMLbGh0XCgqwU2+UAP4Q3P3M2sN75AI/HItlH1X9TELBD+LjFG8CUlIEgLrhhjbr6SN
Y24wtt6rnhLWbsONfoBma//Xls5g779MKOw9zmLjSYXCO34DtrzKihIRn7gfBRMWOIIJKd/zGSO7
DLko7u+MZvSjBvrPUKk2gseCPiAehChfpQzr/V1fCwl7l15dvNB3FfG6gaxMaylcYwu3H6s87vDq
i2vpkD7BhWm+kscPm5IGXguDlQLzRKnX5IR/jkNOkfclt8t+E9gBEijgu3QZZgaG2DmwotmQ/fDC
+9vQ8wt+VQuFWAedMbzPg0fT/sno592/umMvyzwLatcZSSHNc5inPe78IdaUvvQYLf+tUmCj7thf
kfU/qQCeNLbwYUyHA2MtBCS+0YDkMP/wKPMbkTp13fQa1cgoxy32AiQJi1pTji4ats8utJiyVMDV
dup1DEKrNHElLjF10sD/aknHMrsgQNu7IpgvukwFx3ksPxhNJ3lahAQ1b6lF6gBe7+VkK9hPZFbl
523ZWkRcGXtewEo4AISrBsolwuE/QfU/VJuUJogzCPzkmVLzEcgMnJdRbvTNZnmRNAZlK95YxXgS
j29hlXEEqliQNrK4Cmt+QBB3bGww4lnPUfhzgVj9WlNg/L6OBSL4GhLQoNrgW2QS5Hhb6RzTtI0t
R+ctJRfIn2rBOCz3EgnWoIhyGePJKRubtwk06/Jt9SNJQHM+zoLA9opSznNFZuj6yi8zNP6Fc3zh
TkJ4QH/tzQCzX+LNeJkfXfjIawEJMXaUu6kJPMpZHGM/sdfFfe/IzlJSh7RmFcepkCe7Nfq0nCIk
SEvA9OoLuqGYNjA9JhlNSVT3vP/ZxOodqIeh4S/pvphKKlXQEYF2Qs8C6FGS+LQaPzR1zE+Putvv
vD/7LyLQwW6GJCssWahi5Q1r/sw10WOwSftbsgJWHX6qtIaf3gTwAsHiMeV+JQvv3XQW1YlGgAe9
/0oa3U6SG8ynsK89ZUgkpx7tNHvXN14huPCx+M7S0+Lm/nFBpmUdrdLvBY5M/J6xAk5+zzEpFkFh
VTRxpNjVz3Nnpp56+DB9Jo9cyV2S+WJ3vQn4hLmLNAWVriW4Be87vfDe7/IY1QZQShb0wq2MZOB6
hOh3hnAhi9yzxYiDiXjVCD143Wfo/FHG2nhyqBoZ8ASnoX0ehw2uqLjl8JnQJBqJWXPSuo8ytO2y
5u516MGMMaTpGGfXR4W4ZLktCKS0h4TatIzK2QFFK2JMTQlXSJO1xEZCIjYUgQ3+Tqe91Wmhf2RL
rDepaicT81vTz7CeJXHSDF6CyopeknVsm9GM3133R31diblf9fqiRT76UgdZwoeBpl6NUYxfD2Hu
qxRRbvTNHiMfHewJxrCgEobbRW7/dcagq6c4UOrh41kaBRNf22dQ57DO+JRevsG+jtuQ6rmJ+otb
2srmii6mZeSVNrWK8qS4U20ZxKn45otgsLiiTdpiWlilZ4xBHGQziQ9lk+VpZ1AebLxVCliTJOgv
IRYzWfniRemQ6ffJXk8/iuhPVbEmbelah4SRhmc6ajyrOhVgdOCp/+LW8Fsl5LVAK5GMr0avMKS0
9+IO1VlMYv/n1gTUxNZpUkSb6bMubBTbKCbJkxyE/FBaq/EVLtPlI4qhf/AlZtz59RENcS/Tc+73
W6uCr4OEEvNNqXxlH3Z7SREJXSAxp+HQJ4FRyIm50CQf5vsBkY09TD8gh6SQ1Cfev2evwzSzMolb
HkHl4VN5zsOXzikYq04R2/JEwgHgrq8ToomHLbkYfBy+Rw9N1BpuGN2CT1csasXj7FKWjqVQdcPM
XKNXc4FpvqKiFAQRfn3TE3Fd2qjnlx0+ka5iOARagAr0QLjRXPDtMRqayiAFQJyWvm8y/TS9sEfo
/ostLz9u7NZ0d0TooQ7GqP+8vFFYceHjoegPY6WRJOT4i9vVhnKAyt0NBZXYOHu2Z8yEKeip4z0/
s7Iufw2Kz23VzaEIR9zZ2u3rFDBopGmVQ4y1oW7ta+gHN7H6+t/uB9+02LWnZrdIGgBs53wmGLjo
sClDX22vmJLi7OZruFzshzJPlvhZoXr7WV/dlmddbOysRJ2ZpM2bWpQ7RQ48TLM+1gTWFtJEARdW
HjA5XgHr6mImuNasFkqYk6Jh8fTFExREjlY30e/AreuqeRha+2axdU7Y5wZ8boC49Ak4k8rvPRIO
OK0CjeLGg1E48Vj9vYMZ4JQwzLxD6DjrdesDV0mdXJTtnSaFmV52k0nI+ZP4Z+RpUlRY6sgQjtKN
nODFiBuO3vUa0xKQI4gtXFFC8krrNpBaOi4gWUBxpwkrrlTrf0kCeJ7SWZ2JUm2DSl8u7N8M/jjI
7waHG6uuWuX6+68fBMi1bOKu/jVgq7YWL4vTLWK6z9KqXIIA3E4QDcJ5uw5As79clZ8NVNqQVTVH
JTZAWfMHfdntgKHWPfDgh8ONCrjnIIqaSsjF8q7HGG88levPSE6dTgbfYgq/QTuBl+OFyiku9qN8
A2834PkPEJhnNVJ6otolGgG+Ml3pAh6nOZ4fm3TkWrkjnF1mK2rQ1iCNagYvfFiGe6aUxHHHe50I
jmQS8EQoj+Jl5lzJch2/VsusIY2ybk7wnCuMQ2X22yHUgcZAVgeKj4h4uC7KhYhJwpCdiy8l9EGh
qw01YQV2hTsKUB1dexg+SYfzMIWbDTfPDzDyYwE/NP1zgx8XbNOWiAalGt/IzVoUI/rkCvW5PmTp
axRTlclMYCbQcgk9FQtwLGH/Eip5axJyZfwcFDz6zTP4A2IMpIVUSgQHDfa9pZMIYjkcjStLlygc
VyMmB+fU+VJVWjfz+PdtauSWj4Cn7/jPmYm2aLYiTrF9xG/IoBgybo1MgMN1q0HLzG4RundFhDq6
xBOfS1iXAST03GHJepCFnR9r1/pV5EZ4Ya9xCVLZ1ZoB8v2iwyevRtlYKGxrIwtzSY9AQvQyHfDT
by7TDg0PCVtVf0yzds8HNLdOLKyaa1/Ne+yihBkESyCwJNhFJbL3d+1DTWntDUWNm/DabgqVT3aW
XqKB/cD3IPKmMcG2LjbGgL5g7C9Mc+SnBcRuwxHUNJp+KXxwcRkdjyQv24PbmsHv6d1YxwkhsBlp
SIPLKuh/iw8XL466JN6QTJrHINHpyfM+PvNze41DZL/3aon3yuOukzfJpvZ+QIcGorh4FerBdoD7
Vl0rs2BwOHAl8dMIFRs8Zb8+wamCjLstBbGSVMfD1LW8S3EQj5t+bQ1AvemlaMl8a0pS6h+10fyc
nC/enQfGsvlCLSBkA3OpHqespqX+l3tg2t4d5BowXjUtKVrAk9F7nhEM7+BXjcYxMgDS95ZcUU0n
MOh8q/PV19n5e+doW9PZ9nCMN7iaCdOSGhteLLD4NQc5caPjae6R9oawlPZTbG0OAE54MpvntH2R
W9+oUex+dGuFqkWijyZUImI0GQnnLYnXaQ5Y8cAILLBeTigP1Xo+XIiIvyQh+ADMepIItgquxWnt
HEpuK29eWGErehvpWN7HwmXYVf7kKM4UC+vjIPpCIjSmYWLT5+Dd1cH07/wgLqjXe1W9HY2EKn3g
2Bf/ALc/eKOJZicWL/yu7B4VDg2EDhGPopHly/DpN4g3PxfjypUHLtyW4rLPmdH4/w4UkzOSqVrC
Pxt1BWqBL5+lvpuAJHv3oM90UzgL4rpp1CxyB1cic2DnSKTbQqT1Bkr3VhpYVv5LfyuP5ftjU1t8
FmfRpd5Y5O3YkBAmoABVGe90fZZ3wfJ+F9nmMoHPnLaj8PJDHhP/GargJFCBRIUzr3247uZvxuRO
1llwLuUG+q6Eze53rmSISF4Yh7enzrdXQBTNkc91p8DyQxE2YjtssrUlVGiJjSpkkfrFcy7cQcUV
QTF/4zRXel9CjZbAuPWeza12qmhMYFN6q0fFmH+AM0ER9luiCHrdYxoA/FU/GhPbzzJUE43saiuG
EXDAJEV0loeizI4/qTA46/9CFoI9c+UWf/G3uF9hHGgV/OFzxOolhx/eFQndE5nKFIgL1/kNRdTm
Qb0G7YqVs1TKy6jZmBaOY5Q38a8o34suOykNeD3I0Pr/LjF54G9EVmgh11Zpl6cqy60TJ2PZv6da
JttBX6/IIixEbB/Qet4r3rUjh1VFpVHQrUxBOpn9Y3P5eMhFw5kVp7ndrHIDk7+eIO3F9rCfuqJK
8dezdsskpGrhr5q5NW4GP95OJdDfbdv2UQhQc2NaU7FeDBjCOMvSm/sgKYHE+qg6cxQAcWhXe/Cu
DOXfZbYc7aIA3GmVdorVUdStayTaWSNRpmtK7HeIdpqW+GXXHtEp6xgo7kooGUT/TbhtQKvvRZya
bY/KfGMpdrpvuWhUwDrtNdIV+qFDMV973/bpjvVC3RKsggyca0BRB9yYRDyn2wXNUOv9cQY3y7u3
SqccVuTnh+BcgTy6+Vbluqn3J0F0pRSQbNrXgtTcXso8E02GYYlpH3Fmq0MJxME8CmsviYuO2BRa
rJ6B4F30OJ44zVnGmzK1Ra2/e2iSMBBElQxL2vdPtLEK+x6zUCfEqVS6sGmXYuHMhEW5nE6sv1mv
0ou0MsuF/1mAPfy4/XSlcsUduaoEyXOMuNLbPmuIDOaXMYOz740pRwERMEi3aU7wgxY708aZ5rFo
in+Y3ALdieJ8k/wh535N3X7d/D1Ode+SHNgMOTb607IvMUp2Rx/bW5FOuOE4nC6Fp874Svw+trvE
h8ULTBK3f3DynRY/bQ8LRTbPQEOzO8sJl31XQ3IHs4IVfI1+sQ6SpmFz5F/VO0uakbpUnzqe569J
vIzwZNDXphUQWUk5iYMhyMvpiZP86EjpY1Er+ONuCXmZWFmjtzAR0uI3z3wVZx37ZHEydapsBo7e
rqmwZqde6hSrILFzga0OLuNFCfBHWYv+FHhaSWqBh7lTFdcphmbU+2z+qeXb/D/ih9eecHHBxNzL
dMtJE1FHUnme1usHN3VmFuFXJx0/2pxgbwGvARzz+Y7ukyCPytY3t8Ujl+5cAATgBBCMIxl4G2uJ
khZucaHdjezVsJdRX5oWAzsPhs/q2MFW6/+QrN/4O35giO1D30fhzp2QdGzITrk+P7CvNXrzlGQW
QnyN9/f2rTUDFAQi9rOByZnaWUKoJOidZ3JQSHac1E6v+QSFaWrD5L2YiKFTJ44f1gyuCZW0Ohm+
dMTmSzYySFhIKSVlnLltSqcu+N78JOPYQTo3Je8PARHA0aSZZXDXX9DF3C12YKKtzSCVQQVtw+DT
T/VkSkwNIXKb8MAYjNvT8pTeBMcW+JNZvd03vNiMzQ1WdEcZonX5YfYeB58BQeIE1LSXZvdADcqn
mzibShoJ3UyHgChc+Q276XRB2HlXNJYAOznMHauGOZatKPF08ND+SKFwvqZrx961z05bpnpMsYq/
ig4RX9R7Zu4cHi9FqnaoydAA7FWw7Ajs+hzjzKGWDOA9KXUi65ipGwnLRG92QD2tD6OfrCefn3+W
orIA/MFgE12sQ1yTp/WLMBPx1Ax+FeZkK951ByDmJcjPi8VEfGWrQbu2AGIHJCLG+2Dd1mGjIcGv
0Qy4QN018/oi4+uMV356bEjbSkm2+67Z7uF6DtoORhzhlv0/0jJNHBmXVnECBCrkdKdYyMBrLJFg
8FtvOSGyFo8H/++1cy8IiQw9Nh+sZzyoAVDS0ngeEjQdNquWSAsznQ2qkbqdBgVsRRZ86i7+FPl7
1MyEE5T1lDOB/h5oX+hGLtHQiWkfiVc77MZ6D3XMc+qro8XpC3yapiNDlBiYDjWF4NfENULoL3Ac
mrJZqgKZt++aFfehVHd6B978EBT5gUVZWMnZmB9EvvhWgYK8TSEagADh6iy5opcW9VXriJDSk839
e05y4ZvHF9Y9J/9y6+hMNko2zL6p/3QXNhjklkruvmwSUDGCT3DZ9MjjQJ1TnvUI0hkMIajfPuoD
RuYsDzB/sY4Ev02qkARtbPI3LmljkiuYl2NR1ur8dS0JXBO2anO6VusKr2PHp8cGeHuJOQGRlzeb
pMvWl8H6d21aY74W45CkwvlCan0B5kw9LOsET9f0eThKxh+NhBWC9pTMl6LZUAJKMwxNhJCvbrmi
PhuzmnPlUB1jY8Mj1qQ4HIUPcH4E4Y8hpN1mU4xrxhy2EmGiJ6kdI3vxf0Dx2VwKcH8cF699uXDu
we21WvyLlJRUiGGwzfAkgJhPm/4/B4axNbk4dAU7EFwJ41g1CHZVuOQROFPvOTNt3GB35Xj9+gNo
GafDD3/D328+i30Qf2ytNb3QGtjnYy7NtxiMHaA70g3RxqOp1mU5cDTz2stkeYY5eC1uHR3XZzlL
8kWs+uyJ7aq/NpH7JOibbaA2kmA3rerAQC4L8Fu7MoZe8kpCqGAYz9f5l6AbGDDN0AcYAw3mpeHb
VgE1j7GAtMfHjNMDX13UDWH+N/E3G2uOkJOfob6BXRh/BuJTcLkR+9kY+KXFaz8EWrLIoFiMycy4
kUtr/JNlDpoYMFUq3RHKdaOlqOnEaOhtkJcWinLoQ+lDKv85TLKYCwjSgZo/5hHaep5/nasO4lZ3
H+0mt8WssqzyxSI9wYcB0YtnrpECg2RJcA0HuCQ0iKe4J8m3LKtiv7tdBxQ/pkEB3C0LgS+381So
H1DCuKMyRHBnN5lDjmAdZnzIIV5fAqyDky9SH3If4DWaEPplFYiM/hRnOlzGXN/XbOvj8XREQKNp
EX2txNk5AVOLO8HRuVM2uRU5OZX4VMUbsL0dgCeW9KbWeV8yyYaYk0s0GYFhc0+OPp87W7LgjVnG
sDGA5LRyDmtK30pWu8QtFrlc+OmmsPw9vwCVE4+9ZPuBk3aSpVRUBmfp2pJA8KDuzwOLAFkt3x5v
cHVYKj1E3Cb4lCP9PI89+/+VZ1VjGhL/yX6XM1fEs9fDziNIIEXiYjEN4LbMkUTE4KTsjoCABAsx
ckr9fEgGgZ0PPB+Xav+xPjrHnHxilNghXENLylGb4bOEVX/jyvlypdQuUAUjYV2JNO8IHzsAkupT
lIRJ6QPceY5ZhrtOttMVz91tRE43YXCLCoNUaaqTggrB0HMD+lkDgSeuB+HTyoT3Wr51RYtQB2KV
nwq6JaYVKnEqD6th8aP+BQyg7w8h3E44rXWAiR7QK8khBnDAy5PsEOx4sJI6Rl3lwqt1eLH3Igkq
jWdvNT/pOAaoAWLAoHqqtWewOoVWxMWGmf3NQAQrVRFm5FDOi9BzmNudBO93ISmij7ZUXP7GwyS/
LrQ2IK/qIEENC/OCXun+alL3TjJBSxNlUjk2uEj+VTfbcAacFBcYtryeQNgDiFY5DZUgcfMTvVYU
HSuRXBcywIAuXes9kNWMrRKfd8W5e26l4BIuLfW2BKq28T2wsZcVCq2+tvKLRw9YijNxQ4mWpOuH
+P8Y28H/OALDjom7BeRz00+xeR5YggB6spjyHzI1sqqtmABAJyafRug14CPExeon/Xstj1VjyQyy
NsH8ul+QhiHezbSgnU4XwVJU1dT9kvZuOyQK4EoLNKTM9elH+60od5fL3xCh9vsr6E57kdgxpWo7
voojkqTX389hdp/ge9M6IuLzETOpgaRjZhuDOEtbGpkfRn2J1V6qbDBQMvxSUk7Xo391JJevwKms
iUh1oljeZraoSR8Gedlrf+j3LcsG4LO50JqHnqZplfA1WYSE3k1q9skMS4Gc50YVy2TSAtne8Vc9
BCV/6HChCchM4ZLdtIDb1bzo9NUCA8cEjfwyBeeey6IbMr+eujAgSbd/m6BURy+ozY5IPa91fcel
zHfuPHFzH0uxtd+fbkhduc9UVHkQWnJi2MwmVuWlbvC9ot/70zLqS7QVYEe3QTsXlj1CfKV9ra7M
kh60vmhAQ5E42NiL+T2/y5xy4i+SSRe165z0Q/vcX/V9xGC3lAgloVVgZ95B1MRtZT+DBEWs6gjF
XRomagOLYygXRQ6nMHAYLGbzrv1QizlUyRzM8FNgsYxCYjmSttjd71Ieypw7sXs/gyGz4vCHVhIQ
GvCZiia5lFgdqL4YP5Ratu+l3D7+nv+Rkirwl3SfbYEWTRY/0sK86NYuXqtnTzAcrDI8pqBEn3FH
70THM9QjdYXFro7QlhYF291p/oU/bHj2NyH8cRit7bVVp7HHTyibFPn5/Vc5/4Z6BVELYldhLOFD
I7u+ykTAJ9A/pzmO/2TgkAXzvWlwrgYsBkzb+nMPeMT3pqpJNY/mjE678XdeqUrOu6ROFsET/ZzD
Ngo5E0aJKqv1/tn434rY2Q7eskZ+j72VOmXsi1ZrpNjM6o/fTx8JSSfrsIeLyvGDKdZFFfJvh1B1
Tu0pQi1bLgRWi1uH0pZF8UkwG0dDbhvIxU0tdb4MHXEPQHXVc84WUtVbXg7reBQISe82h5Ycir2V
BwCJ34dkqcQNb+wg6m2yMWqtriNOpP0QgHwi9dqS2S0M0/B7Xbu+uFDLZcPBGoCzK4gAJddkiIHe
/WSoz+yQPM8z+TjHouS1vUBtyJoj2pBc13SUESxmhZPrHfnO1Nzu9vrctfWVoIwNtfYM94AmpKaY
6mnoiyh+QJagIqK3SVggHORCZU+SnbdK6opNRVwTA+IiDgqUJVIZTZBMYyicmjQ7nXZ0YtQasQWP
3fNgzVpUia+fweryyo4LZ6c0oBFMJTaTcScNdwybgGYuxbljV78r1H715wEXEVG+Y7Qafutuhl5P
knBufgQMa76ZcIjgwSltw0GE1KF3V+RaTgGnEPVsFmfk7cFtuf/MkmmLdkX9UtQ8itvTwWTWE/Ar
OwaHEk9HDnnVXG6ToJyt5VJpqFNXmgccgC/JmbdAx7L60dkd0nOpH85mJ7+QYB3Xo/Vn8ZSsqQYp
1wXDtuoC3DPdOUDhVOrMonsJ1E0JL58c1hKvMhh9fwYqJSh14bDPSBD3F1EBnLyDKAgZaSL17AlI
9kdp2jnBUv8ScdCcRcga3YGoyPbi3BPLx7KE7HMcQYrtGpZUQu4334ImyDZdlk+hFwG/KMfbCws0
aYeG2g4QCRh5EmY7342Nryn21nj0MjuW6X1n0IEyorFytoNwrwmsHKcRIv6/hhDygiQrWrWb+uO2
r78bRnJBqrQqAIGN6xxNRs9B0NUhd/uX29owMpGih5TNVlrNKTvnn95NZOGTGSJVPdQtNpFWV2Y6
y92rfcP+N9Ycsg9dkLgpdaj9MimA+mVf6VOwlpqmTIUG7IBlNJ/DQ8L7h1oWbslcM4+dhSbztY8B
eSVMh5HFTzUcfXrt1bUpoc2VaFrPqxhLegvfcR0MqDDY4b8Syc5DuM/X8WZVPoOg8gLBKvpEDSf+
1FDakBuM/OnKzZBRr/3WTVJeDJ9nAox6lYcSU5x3z46nYYzslXvoESlSn+waSfWML1lQ7On1hPrr
ieIIWJYMn7Kx7lTEN+rddpHrLK5EDo/st3Cy2s0wuNzjl6Xj5kb6ReSHm3e3iFjsuWjs6rG/NDg4
B8ltk2IwnDohcj6BblQeI5EGISmQHmnfdZqWmPLQba31wBJbnW6oWZY/wkwvEgCPX5jLZD6hIzG5
e1U2lWxSezBs7QvXOlbQhpL2aLywSp2GWnoB6Bo4tjyIDD94smdQitNQD8gd3O5sEng5F8/CERlD
8is+AOcfIUCaDYM39TgwwT8EDZp7pnTG2cUY2U9k5I260gUy/t8KvJHxeSEIV7dQcrS/PQ2jvUwP
VXphNOOoUIbAmETBhA4DmRpoogzch8LKUcXKCypwIsSuitiOi4Kofl/VVv1bbV4g98IfKm9DMfSi
OwgQd6LKzdCbHHiVWCk4xIfvb19KK/0eFlTXiwhJlGJvB3SnsVyH+OveRZA7GIIPAzD6cYQs1bsk
KgNWpnh4034zS3ktt0jvZBl+fnd3GabfB2ibxVaOY44K0Waw2SileWdoiTr/ZSU9CZxUklH4m09H
YKzk7gjmJAMEpUmx75ddQRbupMDXGRyrJTnyG2sqFEHb71H6UH8fus8tTaU2AhgRGRT8joDvnTBP
RvkyPjMJNYzxaX6/XqMH2YakampCMNgXcDmdhFltiQFoy3OZa5FPuR6iXgezElxURHKbWpWquPuc
IH1LvvtkDS5Lnann5WO/KwhUFTSea2+UHIwGPN/ruCthx0Upx5oe3xg9pMCYz5NzhrOTJLzV2BPY
0ihL7inh7+xe6N2HrFlxNwL1iv13wd6LNhCUQEER3HgJB8ZqDeYhtOrb8zj2R+im9ja/XFRJuXX9
kiJSv+pYNDzIw/8WsMzz/Z58X6eewpGnBngbYQZSA9kE1jPSDYupYmgP1GFZAWg1bBajtpwYATcB
fsPXjvv7pZSdleLTCryxiOFDuKWEprJbMcqCFhdlsCZImibxvZlw/fq/cdrOQ/tH/iOht3DTYMZ9
xXQpNsKZv9MvFpjaYCpb3Xq6Avbpou7tE90vU0Twi4EqSk8MOSsIQyxqDTw3rr5itUwIZmOg6e8h
QAYmEHCPog3DTbjKXF5WUsDcdxYkvBHOq96mdXHEzrkOQWx8QO9wq/V3O3CKfTkNJU6junEZ2kVt
t2EA82wcaWNh75tMVhKz9UGrIIJ3I3nsvrl/0uzI/ln22TTy1Ms0+UZPg/nMppLh38ZqkjZU7G20
Zrc/hnIF9ykDwIuDEUr/4DIZcZm19mgBZZoPmN/2NXRV5AJBRBOTuY8jqAo6t/rkGEMCGjLnLwjW
nJvXDF5d3muB1y5jBazyNNkvrUgS4jpuwj88xY2VcI95CQgafmpUjYMj187UdCncn3JBzU6ncfqP
6h5+pV/dNczhdiXxjjO667s9okz2PEBKpfIf7BYbENxJJfloLkcz7ss1dXGBL3Q5kA5uuy8XRnNN
lYAissRmmul3n4lPlnAWOlXDknHA91sRkNxcjcfEK8LiwWa70Y40sC9SyQv/GfEqH6qMYXwQsgkJ
yANR5KmyANxH2JGY5H3TIplU9zrDl414V1U2w5ADUSFMmqRS4wIvco1a9nXsvA+gUyqksgZ7g8W2
RcczI1I7TWm85gdy1JnyWWr0uzQmnJgkp66fwsW+OqC3Am/lujKNuaEv7O/aIu4aOJHW5jrA8DgP
iasdF5z1q77O95stJm14dVOEe8F6Xlq0r7UkP922+WafwQBXvex+Q06+TWjXNECbCDH9YcThESKB
W1USjjJ2kH8o2JFYg6nucthR70Ul+e4nzc3REach6t89NnEOtAlV5oehMO9+BzkJ4qUFQ1wFbJbd
Se60XyInxiBzXintuDTItYkVhpwIc6oj70hN121pwvYms8eXPhIoPtEeEzAABp9Xmos4lMyiLMq7
grMRa1q0SSPgZmhgUYpjIcKCVn3Fl80i0cB0Ujt2StvmUrnIF0XRZxzAZ1I9BMTdonp2hgmX6zDE
CuVxyFiUOi2k++ACLH0hP6LYBs67Pihc4PNxjUmAaqkSfdU/Z01BIFHaZU4jzMoYr42UnPwJbvOx
aWax9qvzff5Pf4118jOHycrOTJSQpnX1yWuXPm2WYjCWUdBLOS4izlFW87U8BiEMci8rqbAnpbZK
S2MSt8HEwRXdCvm6bJV9dlFrjgXvsEVBwmSn7MlE73AWvMtmsPxaS+f/sCdiJXf57j0yGNF2m5nZ
SB9SZ1bjAdxXLZ8ciJI4MhJoj0LGX5ct5TyKgYB0ZCItE846S9jeyoRJfY0jkcgM1CpZx+7VaUPF
/Ykp/T6Xwbi/uCNuzgoD5MtEddHGYYG+j/1om7ezzNhJ76wIDcpOW6ciJuDohOdd32JNhw7aD0Vc
h73wUozrK1Hyel8h58x8majKPxSnOEpzLTcHzVmwTk6gZK0rVXW93ZsDWgAOm8fyC+3lOu9ZW6Lf
K6laZ2BTVcVk5ZObdahBlo/aYjjULIEI87EdVjhFfVuV9QDF/tcyLUMjmyFxQu1WJ3tvIQzeg8cH
/A959fH/M0JXkwAhC2nIuCMd4wuGOd1oHMvDOT7vgIA685GC53NoXrg+n+SueOBy9GRdnoWjK8nC
gX5QlvFfoKFB5iKnLlEzfgfT8roK2+JBS29buxGbftx0rPPVvd1aNUWUekfA2A7jFoJvBUKvKg3a
OJ0yJ/ViMJ0oUuWdtZLOdtRR8j35nMHmvvE6PQAgeCAJwxriVxVEcMStpxfprxVB14xd7u3IPFhq
9jpKmKss72AVZ5htYEp+gMgVL8otuWR87KbrhaPyOCKLsWbW0r5qXrleDqWgA/WQ7Bpk/UKIWNMR
P3twHQoOofb0Mcov5q54EcLSlG3oobBxbb2grYoPqXlJMeVIZY4HtCEi1kAvWO5L1uT5qYeAok9P
6EceNmbLOknsi3mLXfPV6I9SJiVkogUhhkDJffsbHGfGzgWKNQK/QhHUKXs78Q77iTvnFYZeHGZI
/qf7iH9EMbRUd+Ju+Y31iqUUEOYjKp2BeB95IdbVxLbEvGeHqXWQpLSzTJeme1HInS2MzvBQasuD
aVm9ODYWeZB6mQ1Z7WL5JjTL7qQHPGJ5CWNDskaNs6QSEaK2TZdxdu1LUyfnTeu+LbkXjIuEZyHJ
18I96bNWJZvsZEXD17G+ybCJZZMhUHCp21K7d+Pjp9e7Kay/kNnh8hjWc4j2Q1OMHGBV/cm4i/KT
ugrrPBWElQz7YbMrZzaOWu6CRCUMSCMx4oqfnPxaht0nP1Y+rvy2p9iISBaku/w1k2j4g4RqGeij
fvsDL/PR5t62i5IMyo0Jj1WPdJ+st/dg1w0DzNigRqNu5v5pG1tKkJiDjJQnBLtfUDimjG/mvvL9
MRpA2/SpCUI1YdcVkbcikl5iI8eXabtsbPv3JjFzr6o4SrDT+Egzku7+vEHj3IqN3D1AG2zE7GpU
PiBYeInMoka2Th6OG1WuPFad2dS1iKgWbWPgbct4tLhPG2V2yEZKUnPM+SGbLbzI2VFialQqTBbp
0ged6V90AktkqIIGLCknqpTkCmdG7bhJtmC2soeREfkCOv1CP4R394KcJx0KLZ2eEbyh1qCsod1k
wr4nJAC69tqJwkJ6oRjzS5OpltPBdCPjkoMGcuUXOytQP0zVGihR/LJnuC0oJFEOAKiJf/4SWoLC
ISlwTUggPmI4t67fTsDHZDr/4FfIifxhRXzI7jIyHZGd3V+S5DUYTXobsvTARmZLBVfp4ddlnjOW
bzKni3PO3mhtHq500CvC10IHpe26MrKfUGbJ8reMQt3GBhU2HOLmp7lIEYzGL9d0Pg32BxEIqZuc
8zhoBJJEHCKdGSxM3zrRhCYhtZPROVvZJt69u4o4ZbMDRe4VnQmx+7iQtHKjhlsCXl/nf7RQQsBi
uGYJqXcGadAet/DjnjIIw/4yDD5/ozTgQsYMnhmFvn56m7RhVeaqzl0Sp5Jr9llE+CHsR6hYXNFI
Uu7prASCV9BypPvN3YkeCr9Zr2jyp3bYtPYt/bfBvZZvkBAd1Y0sDis7HNddkTUEgCChTVLbVUzj
oTr4doHWYlBzAUZ3t9jjUJDWlCB/nIb5lBuqg3u2KlTnZuRzOH5MLRR54K5wpZdALoEi0CiLOH55
vjp5DO0DljwDKW7CUErpL3P6Fep68/ete+mI2+lpw+LFZQSzQ66zW3/2Eqtdh4W/mZdzjzL0Ouun
9XOjeX0QSxVqBcOkmvcqfKyZKgumPFvAzsWor6ErnUgtWHA3/g5QJC4FpVr9kZIBMndqDSQuZRvo
YGl6v0Cj6vfFmFqPv42QJw3tC7htfpZvpbfQTQsgte/Q5KDMy0/UX5I3ZeWZJCA1P6cZIT74M1kv
1uIEj7JztFeoJ2ZPG194o9UrjMWD50C1iQZPax8IEIn2/jpujISUGdsRVHfaM03RIF0vbJj/lwjV
upGX6HfE57yfZETq2OXy9SvRJ8jBnRelrKIxbdq1yzms7lsXobbIjVhexHqpYgZl7+h3MsyqOrAE
fgo6wn2Xaf4oDCK/xI40sjX1JPwbM+4ug2UmUlGtjorHIBrqbR8CZc6/4br6SIciNnEW6CvtjMVm
gf2zOnfaWMOigRxtz3+8K9CryN0iVke0B2tWeNkr4flRgGUtVvT7u+rLs1GaKxCXiZmSGQe33qvW
w3JB1BN0YaMRzriIyuEeZ0b2ppGDSb3ji2TVJUndUQlv3H5TSuT+DwE6D5MQZsfdhdzQJ1ehWfGP
FZsnRS+/49+MBCDiEcNkUMH1GWoQrNefFTjr+jODXEuH2IRcN7Rmcv5VMkTJR577s5HxlLaAkRxb
d72IuK7Mtl8IOSObAZppG1VX17apyC7XDP6PMJi7h+6EtD/8vPExQ6X+ckDwi5EiWZ79fXyBNURM
ZK0IREmujer2kpa7dlQAaGvPdJVsLpWi/gYDj9x34inny73uI8QOIQNDrz6/tvIVpRxKrKdpFazj
VHo45uSaEYB6tFZ7uQ1we/lkvSr0A4K7lyxwB2jLlKSW51Yjy/NoDXFPYKcUzZMQzOXmuTgLW+hG
/S8dPJ3aun41VQS6b5LwHqUXlovKU4rA62R801IQf9xcMeYuKEJtH0wMEXbHTYHGSRQ6hXGgfG11
eUGWedcscF6ibcsQqz2KDOF2Vv66lBvHok8/X2LMoyDA1sHxlhmde7MrF1JBHYJSOgVxHnfjltdg
xUcUAz8kOZ3IGy4CKhu1JY8G58DuqZgS8IghMW6m/nG98itwpuGn/6Y7msjQdt36pN0cLwRd4YQT
2ta81In0VUo8AjY2WXc0iFDh30fMLPNHsCk/EGw7wBjkNIPlZDg+uCFGqgmkjf6pcBcMF5LvAR3b
NPQc30ajTJJfBny6KPYvuEu2Ro7vBwmz/iWJZ3DuBhbrFLi8xf6YLaErK0wo1LAvf2RJbyVSWn1x
qz96JwUGtkjfMCOSVdS14IZSjxJi+AueT1+DgBiVnY5/IFJhfB+pKtNXLY+PGsvX5VZepwMnJbS/
F6KZ3pcPnsiX4Da1xIL/ggtryT799jd3aWWevgQqr957/Dacu6Y63469r7bdobLDuoSpLOhBE+eq
AaK4w8Hk+NpZcddK+PJ1Wt5ak+z7FG9gJfq7RZ/WSZ13fncwP5mbvwrs64YwsZQSPjkgfk6PP/m/
xyfh22cr5ae96rNdFAcTRWC/+DKAxkaZzLvxW+VV1wtxLt35P7NtEyIy6NTxHS9ZNXX5yXnd5pLg
x4IEI+9EVNUKKs2K3bDogSFknTSSVI2jYXl4I14OLh1JHAUIxKTZO9sJHw071Myp9Zh9mSNqkbya
Rjo3w1GkIfAZAHFP6+BhTmUvcNddHhDgfg8RD8FL4KkYIIqa3yhgAIvMW7u/VE+S2IeSZj5fOERu
wu6JED9NZPPT7Mnzz94DM0eR636+u9uDyi6bUAp3MXofAAEhy5Tl0lpZN8svwIDMba4K3xfAwZrX
Azm/IxIzJMZ+7HBZ8B2HSVrJ6UdjXRF9ztz1/4uPI4iLJD2519UqapaZfLrAzOPKScOaTU+1/xep
UtEbg2j5sIIq3AO0BT1Z41Kck73qNp/lrxKifDM5u+6e3i8umzOUjayNJZPaXMnIeX/eisW9qHpe
I/A2apK1k6SySfd7m7gQG/s6odKxVnGK4J9CRij8mBtM8KUvg2MfNIkziacoNgHeTEPO/m7tIwnL
2PDxxTvlJLet6FVzJqY4lkHivcQ90I7NEKzuytjA2dkGgzm94t3DTwlnigRqQB36Lcgrlq4+LRgb
4ydiMtxeuDC+dF8UgHfxJjsSej/QF8d1fgTCI4hFiihGkeA7wZ6u1TAI6N9te3dJlRw9e6FHNXC/
MG5XlV+bqkFSNw+PjfSM2FYET3W3XXnzFzS9uIw4o6HXoxNSmlo3DifoU71NGdviuPh3fJLjeWgI
LJdkZuJKRPzX5M1BvJj/syDDHOZblo5TfiNM8/D3Xas+Ze7jAJOH2IM3rMzyYvtT5uno2qD91S2A
U10zWtBMKp9cPBpBqBKgge5t5u6VWFUXJu1z/OzvhsjWnm/PQJzg9p/w53EjBOJxz7nERAghatd6
ULRE0gRLCJUFY127OIPPmbp1CWPc+WZ4JhWe02wPUxBi+2WSu7eQL7tREvOKn6L950v2U6xSQpkF
N4TMoQkZ09F3CGiMP+sYg/j93IeFUgUH4Q/Ue3mTwuRSrl4Tj0ZMKUvWo3LZ8bIhJV5eegT6VUix
UtddkdQNtblNFEuRzjoGgkcIiyRlhAodqhxgtccNOBb3WqKtjetzBWk4C+/ZCMOoqpkO3VWPh71o
ABBKKULqI07F76SgtaVpwbFrx7FK0qXyjzYZrJnuPR1gCbxELBiEoeh1PsXL4paS4WBryexooy+l
Pe/w80w8brUi3RKfPjyVUQErRczFEOqUmcoxKowYvSChIMQoD9kmf8/9GrTen2z9KobR+cD4N0Cy
xNSo5aJRWMXC06eYLqkadDPY2/OsaX92cPPjSN55emAZK/R9zQWEclm6LvLf3nyvPKry/0u8n04r
yoFH/XAeptPM0aE8HuUYYBGB7M3Ac+J8N5aMlHwp48sz7a63fEWSPAjqIj1Ba9cp4V4vZmsjNXeH
H+RPqjoeZCCrjN9mjiHRJsPKAufQ+glqmtaILjAjADKJ+eoHwnBqczPSNI1Mm5EPOCswo1H31xnv
fVr5npIlS3GSLNnDu8p5HG0JyNMefx25yglpaPM4XHA84dl6A5fXYWIm9/pIDY2pWlzJRGPeWjIj
k+/Fgd2BxqsNLXTGPW+Mt1heQeFjx6/o7n7DbVIoB1CpoDXEzLt7aHFT1oNoaQy7Lz7rAUsaU0jw
VF733hhA+CI0lhN50EFE8xQje58z3wydvIbmvP5RFHOE4RogrD+/oiJmdGUK4/luC4bSmcF3tVbW
3X1j6on6V4gfuhUG97XjuVxjzFwAN/XWl3zjr2vqOR/UrrAA7JaITGbivMNNc0W7OhxLPxTgcN3K
ZPxWScUa7Cfn6thgIdu38WEHtndx/HNzNkhTwbsiOVQcZTrPU/+1zC6vTnS9ctbTOzRQPUvuRiUr
hM1oR+vFjpU6Gmd7vRiPKU1d8SDh+oG61dPUp9uhyzu6Q2cWPBDU7+Fgjbz4uTZPOQPDOtHPt0GB
YwkomsgBlGmT04LAQaF0mJmQ5DxVWRwcsP6UZjkkPQjsDHcVtDvVzj73wc3rdY3UuS5R+xGd3+GB
GftaJMoHElvTWq8v9ffT+fYA/e65tyqNwBD5CwYzgO4tVOQbUDqvUAvko8L9bMIcn3cmNS9YgJUp
Jmh2Hinn9dbvmr97wtGsUSJiGjXrVC+DI93cd8OE++2lDYaqlMsfMEVEi11ZSH/RdMiYCZMcf0WC
gaHCGhAXzCrZnU3ZDWdjbHPd3WpBePSxETOSG4U0Lr/c14Z/GuQSpbYDufypo9lYQokr9u2z630K
6n9O9q43oq3jFAkdntHYBITLm1N6tBJDXz5TUbNOwKGqLptXeoX8gyQtfZ3xOkEOWxfpU11WFgKX
3XGFogSzfp+lcfUd1MQBZnkqWoe6+0i8DPSedG6RF359GQq4rTtus095jW1pkwZHO3amzTW9fjuY
2/zfUE6N6rZe+5wW16Gl1y6EfMbNIaaU1uuAjlMpUB4NBKLrObwzK67SckGoxHyKBmC7XvmFxZMc
GrAOZ6upmLjVY4x3Vgu/wZ6BoSx6fAtEv48srs4RqMdCiJHpXTIzEAz0sy46FABvRI+Jn+XEIcKX
9F6GVDGPOtSU8DEvyVZL7HoAs1Ke2tDiHzMzH1CsvJP14A5QBOWbp3ajoo5QcAf8tjRg6a8zsuly
Rhvd9683S5SPjJlQsGbKCHVs//2ZFxTpNl2//f3BfUJ7zNuD49jtUVv0Ek/Ikh7KZ1wwSCY7CXRW
oORxbWgNZYOqBftPMT3m5O4ZQkNZt8xtbC22FqwjjU6yBTndV4nQRMpJHaT4gJb8WGmWJ0XRS/85
8nPD45fTmNwfNzw22Ft3ZTlAfy4nB0iy/3GnTvGkLnhuX8ImOBnuoyto56WNhynlUGA0y8Cp27PB
ncgUc1iqtEAG2cMvUJAjG87bzG8piiFr31YrNAHZEViWwaIw93QttOHrZkB33y6J35pOnz/+NhjC
i27w5OOChGtdS1SIbUIuA70XGkuvRDp+zMVKXEX94DOHgffJqCcV6jihiPhOjPULLsP/mEFhpEFp
IFB/QNksQhmmWi7YnJrkePM4J9JxFadKkpMpELPUAjYLp+R2mzsTGBku01etp2INrC/dCK1qsYoo
G8xoDjb8qJIkcTc+2NEbdaD+OqGv3q5HmGeGV6nWgG8E8fG1MDMA7MASqfLFrcrDZ0bLi9XvXHsO
+XROG91QuM5nfryL1PCTt3DVCZglX0OC1TDf+dglHewAOQRBOuKty8/fgUZLJQmGeQyrq5IWEw0n
I2TujyEHnL3IOaj4lgoKplwUJzM6oRO6uP1I+CcxleS20XoKRymUcvCtPIVngj66JzZzQQVxzaiK
eI3zX6c2TvWjf4OajK9qLBLT1j8oZECHhywx13mB4LvSeFeJt6AM4agxI5KwRT9KGzz4sOCS3UFp
5DMVV6z2zxWf4NtwCZDdu8JZQhnwIa0z1/l/U3dOx+S+2nSJWOOtbXAy72nrd7QnbdQyt3lda7XT
wueF7Xp9y26v+cZIXpLy72GFPb1K+GJSa+kui5oNqIO09sce+4lHRKuYWVfuaVE6XnRaBEEJdluR
2YBMQvTz031KUM+R8k9UFEyul2yUAfb61TbSzAnqBIej2zrUirSB+gsSkLJIHtEGKmF101pZeQr9
1UFyLJUvHxvbiI9+IrtDQzZjzH+BVPhA7y91POYyxPly5jo1kC+fUhVjaYYqzm9cq7FGPZMpNooC
DTANBZcKuxQbCkdrueVB9fIPHpjeOLem+1xphrMjMSmKvjlrLRfafKE4bMRSerrjstoaWaI6ZLrt
+9nLW7ax/5MexD2G79B3hNHjwHk8Qh3tdHK35ONLE7jUhH0djOWN7o0kmQRBcc815N8bCdgbUzfC
3+gUhVf65k8l7a/NWP3aKx60Llm4sTT4Is9KXOQS4Si6SUaIZsqeFbJgkG1ojUuN9/0JI+IFUp4E
qocto5kCjwpBS5hLaBa/GD0ovdBoJqWfXn7NJiRpZNHpD/J7W6eJBEn21P5ZuJFBrOpwflvDctu0
SOWxqkzGmwOu86Un16cgxuO9tmQ3RxqWy2nqwHskxzD05QLyEVuYZRaHFWOdi/e+ebMHiKMxn0mh
QsUCaNRbCZzBDL0j8/W2b6Sxe6on+WW6oDHjANLe4CKbMDwHRhgvaj+hZjALre3Qpc+7mNkU0+5/
WhOUL70hgIv9Gozy1pRQBTmRFmCDs1lMg9yja6zW4Be64J3XrMec3RPZh7oKE52YuidDXjuBAwO4
7lqd7luac6zmovBC1ztPuMtAey3TRVdPmNmtqXYUX6N3bt4QU4/MfEN3Xs2hjrYaX5uTxWs1ljzV
+bFULjUn6vcUJXhao+dulz3AFHxUcmF7octEHR4jE4HI1COVtNl6ouXjClVGvASlIs4avasJCTkl
Uj7ETEYr8o3/vIhAvbcF1Ds+Qh5V5YFz9gHEGhCPgNRNEpsRTb8H3kGe+97knSzQMpDEALqiWk+5
jgZtwUwjRMRrlKhZkbsnXfEIE0eIPMHHDl2SMgplxYjSjY4HO3cjWa4dVnz+MV/mg9ahqqmSkcb9
v2UQkNFrMcEtLbvfDRJeenMIsjtsnwS6jmh64j07XAWZc01cLTECQPZXZHJg8D24QyGC2ghTJ97G
OqSadCZgMfiXHRjbkQT8m7H+JCDAFIdysDFwMim40k6XRfVWtKCFWlwPshMLPyWXGM3RnHRHeg6b
Z9BUa6+qQYsjjU5MMrX+la9EU/0PRp7ZvbckhrfhGqSfKCs1OWBLwNk9WgFh/gH+wUM5VBzoLFo1
BFpZKXsWYHAwqR8tluyeJ8f8j499bzN6HOKAlAFTuuaOpU3amQ8ItpLvfOU7j7HzEWSErWy6mh/J
7/OZi0y9PPcZr4a81hiZF9WEgxlTCnQVNGpJxNZuFDb7LnMWuEcjkUwN2yCm+sELYMqPsakfi1/2
mgU7vCWojbupyy6wqEwRjEamvZ6Mziy3OMGj87S99N6eo+ZfpLs0tkecAKgvCuUmi409DLyI2hJm
keg9dMvD/cSfOknoMOlrQwcTmorVXdd/tRy51LgbO7KPcUJchGwUi2Uduja9hkNX47eIsJe7SIoL
n+drd3JsRXJblKZjWLLgr+xDA6NmB/6NaR82L2BycYD1mDDPjz5Hfn1vDoODSojvjV3JQOKOj4U4
rPZKdrU9XDqCjBhhWx6WyXeNYreyCOLsDxMoA3Ih7dlrMd8i3xtWbyJYK52PAeILoNmdJ3METsrT
do6KHCdq7AlhirzgMGBglDF45xgx4GzgTONt9IhODD3LChBvkMJHVOgRABRi/0xfSTf4NFeYXcix
zL3RXoHlMHL2xgRLxgo+TrtBHWi6Vz5okAcFkyXlIjX1bUfIzmQ9aDY/0ZljBGgRlGYbM9QqWsBk
sT+p0VgMK+G/k6JL5VoZhYAY9LgjB9GTBb+zcWBmskhE1m3Vufzny/CbjP1k7XXmkn0+2bDz2J92
489KX9pm+bo3FBtAVnH2Og3PFUpsBPY9e7iHEvrNXHBDbwDmOtlGlhy3ybTimSzbUOnTWIvwwcLO
SJPNoz0MREeL+/WF6Q2FDBMF1pkr/kh1th0tj/wdoGpdSZhziBq0Q7pGw/joAUOeegnuIr90KYDf
6IvcUbRLQYhORFTAfL8v6W9Lj76GB8GhvYSpTt4ILYoUu2ljCIPdGqYTbFUKZixIgiL6T5ZHaVHn
hokDFp38j4Z8XRtY02kxe3a6+JMmmRiOAiYLQ5fWMJALZ4Tw1q/eig5tU5Xodm4xyLRny6kGJf35
REfzWziXgubqu77KCuGzGV+/mxFzRqSe/RaEQ9oPEWVMRo00TMyIYB92hS/npvFXBLMj1SbP66S8
M1gCYo847ym7UTGD/fe8rbYnyZ1n9xYB5OC0EnpcLA8Lbv9PsHAt7vRh1sRc7qcFRpBrKKHjU3wj
zspb82BT7o3Hss9Oyg7dEplf2TEa+m08OpqBIvTGcAsaxdbLBlYkUmEziBcCVitC2evHaVEW0f8c
sBIonUsy9Tn+EE9nzaZXz/ZS43ghXFLHxSsgmmiPjacDYL/rm1AMVMGaULCjIXMfvyvGKAaGUnBK
yqMzfwtlNkMmmAD+a47GFZ77V18uKLmlXh2RMQctEA44AtWBc8HRGrLjVnnzyc/wCBQq+0lJpnpC
/2ftRplc9zHV+sGhxEmZNuA0h5nM3WkjF+6JXC+tWmNxQrSSBni0SFL2s2H7KppesKbP5MGTRpRJ
b9EbVLhXcD85y8zmQbjx+Akcj1kleraO/BeZpTP4xYkgSE0QnYeAdkPt0wpwwkdc7r3tjeaRff7r
bR18qYFpeV7BWaBIE1lVD+y3sV0vCizoarHj1zmoqbvXdaIY3zHqfJ+asCKMg20yOKrWvQyu9o1O
JgS4kK9jIyuII219VaMDVXLM1t32ldEYmRO2I7jWqIm78NfOZyLnZyNOS0AH+zcvg+HYPrvlQwRG
ui2r7QcV8ZBReJMhU5KLgBXJJDUkoHTHsgEiTbhfu7iToWefPGhgR4TlZopWZQ0RXIECDLphXX2U
yEeXz/3wWE8Zs6/MfuzOEIfke/alYGAC8SgE30VDekyDGDacqal6f8G7H8hgB/q81MIk65XmyrbK
qk/9dJUHTpeWwAZ5o88zpmBUBvUI7pdtEtI0zw1PTD8Yeisljff1tyEx6IPlnwB8FNzXr8ZlXO4b
BtiXXQ1owd/Jf7prMydIDe9tiOjpk0iH+0MpCaQ53Zpsx4UUJdUwKvv+wtBrpj2jByuLZr6kkaUx
Ac4BjLMIzGBqW2W1NiCYKyhX7515XC27YeoS1EgEk1M9W/NL/LyBDXowyWrA3LM5BFcB88xGM19r
TdByTy+nk6lY9U+rHxOU1zw7tDZXr91HZWtezihV/UQAOks7D21+bLKMzfPnn14/Vh+BjOL14y9t
dCmsvzmdLLms3ZvxN26n8gO9jn1/GakWgt9w2ZFm247SIWo4C4iMDxn2sGhQn0cpbZ86C7H2YqSh
QUOXj3NroRshkDFrIrgkirUu4tu4UKNekuEQKRNewPCp0P3q2uoajAhsfjKoSiogwmyCSOH76ZKL
mDQOyTjmW6JjR9NWowSzfhCBLkXtjZr9GsbnzvnkWxny2sZvQaqeFy3DVxxlY5v+zfwK7k5bgCBU
/TorsX7jx5ArSoAILmBCSFwBxXxRx4/YnWML3YWwEi7ZXt9d+FpJ+QbXfwR8x1pl/AWJKJEOAKDr
oQoCvOEuE+OBwR2LDo7k06GMY8hnh8sAgpXeP+TifDzKLu60qNFyk5NGnpZGYyHQGHoKPv+H+ONA
Z+nHaMTyyy2BnZmNRwZeO3z8WGH/iYzYdaqol8mb3sYxG8BG5pMScqne4n2eBFT5Msk8xd5r2izH
zzeHPqWzVHh4FHWg6/PqMkKMTDMIo8IC74EhH7B6xcKzmpwQpFLwIb2NBiggOFKWrRPy2NAV5aHr
Xd6ihPWznnLJHH2Ril8uxdsgem6vVbwDcLoNXha9it08S9oGqaLpXmBiRVzPchqBnKKYHkJItbFy
2u7F76k7AzjzSrNqRFx3ZPP3MBoT3miyuAmlg2L8/fYCO4qQrW6zT6CC5/RuuJHlbrG4Xz5gMrEY
s3qXhlFOmbU/3OOrZAAa71kOQQAF/Acy16yd5JYRbGidO1uCPbxFy7v8EQsTSb0ok9tqrGdB/gkV
1DJIEixCKuONbJXgk1omKkgQPR/R11B+2Ar85OzE3BNJhwZd7ydvj92QnE38MUn+8k9b8nQsZDI0
1txka0rVQaiqMM711BJPIAbCrconjLFn/XgMZnh4umK2qFV91CabbHjqzdSteBAea8TNYzeZl+PD
H1WwBX3Mr5ebB94sKyAGbUY9pbUx+N7Tn7WLN+Cw+ZG7CctdVYK8HwbkYqU2jkw/TVaAPb22Vw7m
MzScNAYo3/lJ3Y+N0MYpV9tl3F8ztycA3WBfurfkrJIK1yaQCuruNmU5f7PVToffA3UMjKY/XTjV
p62MhAH1/dIBHHUUNBegdia/+C3+c0L/U4Y4WgLxYPaONnzk4fDoMXka1ZYwrMkqQj8wd8lLtu3h
WVkHsTaQG0++LZmBDoZL+hdnYDc6f3llbKpOT4b7T78fFiS67ulSZ9oJ99iAzMofeoEEZp9Mto/9
cpdIUvzgprwOzS+inx6O6iHEQUCJ9PUw6N4blUQAAdBhMYpH8L/ejnMBUVu1MgKEfNwnEw+bG4yN
J4YRwHAF7ItEZ4mqDwXlTB9iymSUVshjETii5SigtmBOQCXYqm0PZmhIs9xPZYpxDpbEmXUhETbj
PURzmp3z6+uaf1DTNbPFqP7E7S6IyZfdbOSiJnpUvXhq6FTmFC22kcnOwzUzQUB0YpHsWqW4f+lp
8oW5rhg1NZsrDUZQ09whsd9Eep1y0UEl5sGkfV8Fy20vvbF+Dmr2L7IO1WEbs+UOvLL3Hjt6LMvt
3s2vmhUSUaZrT3lpmkJJJpoMZ1INHHt54Veg8pvsEkTP4mNSGtC6frCVlnAuhCo1REq0m3pNhNfa
Cy16O3vS1UIRTI2aFbYMROgNZjlo69HxFUvBNoFxEMazYaofXm9K07azHjGLMztdkew+PDvgnYy6
1cXUNbXSLoR4LEOdawC7Ck5c35oPpYY3xhV96vFTZMAc8PAv6STsr2khbqeqv4C+B7ROHmqjj2i1
PZuz5cJW3Rb1r9ieZNRq/cq2FyP/lisfT7PpTm75hY14Zqi8TCupiuipGppfhAEB8f6YKAkzh/OH
7YvF/rePA2zeuEwq2lUa1rQOTuryl/8/L4sVa9T9/6YC1gId4mDeK62lEeVcOka706dn6qxszAGO
LxhbXN4BKJ0+OnouaUasT1ghyA8UP07NIH1bvSwSsmcWsGxq8bLXEzzKKZwgLYbuf4+a9la4B23s
52OoWFEZIDWkjxojdOBYcsmNMA+CMzIpbb7shNr0o85P1xpXva4FPqxI/V01Lxe2DwPIQZHGrtUJ
miun1cY/qVFWD/+UwqkNZ8+ScfFYh6JP96S/E1bu7O+w4UZetNAyYtxjjIdGtXQcyI8477tjuyc9
+rFwoZw7EKW2zgoUrwuAZh5iM754Ja0gOEfuVIZpNMHAwdLWin5dCv2qejEPD68MPmqd6d9rx9br
ogSEpd//Ip6xd+j3RLidywfRJATn81/sG/4vUL+4Ty3urVlOSb4Gwx+Pf+vYz9Imp7pyEoNI1bwN
2YWaW4mdBymAc5/vDmN21v58sNhMyxjkhw1hAhav0sdzxk4S5p42Kz0GXAlDPlY7VTCPG6iT7CPc
d0uZ6VpiCNVcfZnCIeILB2BmmD80uA7z2W1pRRQhJBlvPmYzp0QWRLBf3KfimS2PBis+7NjUWirk
zKZouXyJ40RdIIUMZ7hrKsXGw9mG3o70oASfGPkn98vfkcMtjBh4qr3SG9WV16HvzCmdpiu0Eibf
LMC8LFd5HuJPp8dANeJ60hOrp0Z4Q1/07iiBJiVlbwn6wq48R37qW8t7xmHqBZu2wjk7nClXT2W2
qxCz9Mj9KTcC/cUFxdSN/xLTOMBOO118L5tkVi6JoAWYAA0WmNaNNuHfvPjAHAhZv8ojXCBW2CPD
bg82O69xqL9fPu8bplden++79l760QtM5Ow7Pnz2+URXPdJ+zWLd/JIB5UUOMG3F+4jE4zNFHQJo
kQYS2GXaL2V8msFjxB+9+hkQ5kllgbYnGtGpvpsAzoA7YPGD8mhMwlOF/0kp9X/qPaMti+OXSBRu
FDY8Xc/StSXTiCMlXRuyncsTdQoWXguLgU85IYJJIv1+50kTa7YRaY7ANmxmcNtMW/l9EU+IZY4E
CaVSoPZ/OlvDnX+S1T6sRDePeg8MG8pWsaU0ZxYaWpyr92ED5Dtvzcsz3Vb1PBkrXi3MNdAC8Saf
IV//qS8c5zU7XNLctf6kbngCqCxEXn58ImK+7S3rRs9cFTa4iUJYWFHxCAz9df5dBa6d6stzJeJ1
VuQe/WCgQ/qfQhZ/4SZk6PNh7h2dsub86XRhDQcKgn/u0i1y0EoJHy1Nm97y1AT22KvTfPNnw4sO
Oa9EKUH89Fg0I3Tpw4nWjVxunv9lv/fP6Sw8vI8CR1zr4FlaClTIrtkwf+GbJdWSnzy/JuyowUP9
MFTNBGwMrit6Rcrp7u3OwKzqXemsZa7edyCCTVM3TVQbgoGxc8d77ax9xeievLtiwTJW07Xru/pM
eMdj4FxMHlrv9/ho+xlHopgKQXCvalwzO4gh0z7O/l0vou2vFw5bUuMpJw4jBbesmfwh9zO1s5nw
8JMQOHM72H4rNwQjly4Zdt6+DmhvIu2FEqnLwnBP60td7dJZ+Pfsolv6WugTiXNaFdVc0b7G+0nv
EIY2tER1k/4cfn0VLRHz0L9p4//vuoYFjaU4iQgoW8vL1NB3XI44zzhY/XdCFLXPgS0axdEWTNKW
V5b5Ktf3sxkn9nZJKHWzeH7mH0Z4GP4PUR8cHGgH95CXt7KKlUCXTosfqgxQ+Jgzwsokn1YI9pGd
FvPknmLXiIeeN4jCOxASxqPDK3hcFCt3huHx3GHQt4bnaXfKnOV6inyzpp7U7HKlIZqE3mUnkPUK
H22lGceRbsLLll1Aba3mU05SSUp4qVJ40yuiTJpy1Q1cW9qdN2irL5ff/m2qyKpn8Fo/EO6d6syi
wu+wml3+3Q9pC02FgsBRwO80PrxBpBcfzk88VSj4HYw8HwL7pERcRGBAtSsNp8MSvDS2LMedwnP6
OjEd14Ggn+AWAYT/FsbWf1yTWqKMTtW0V+YSWcsRS0Ft6ktLFkGMpM9Y2m1Edk3VqYbcMuJ7Y6yq
6Bie+88sxpzs2FF2UXBCXaCQef4PDMihe4Abjd2QmZDg6ZMQXbAkbS42D5Ex4uHKR/2cXmT3zcck
+nK4Ix6hnCHS16XNJ4UH8J1Frl/BPLj0Vks1pPl3kPRLIUcONtVPKkzKlBGTi3+xOrU866iP3/XS
8qS73GjIP8iXTBLOVQV/l2HFK7relQEtMhZDXJixA/N23GUdXofvUoOyn9DE9HdIC/VJ1hA9JJVf
kuohpEtAROv/1vmV/JNyjmKUFjSE2URE36OZuEQLM9AEyLrfOvBwQwB08ma9H3QIAmWDyOgggHwT
SMuYOKvz78OHuio+TPPwEJrpoQvdmdTp2o+9ofO3dP1MiexNIjGL6FEVnkv1yxFBhiCSLzXp6lCm
SdoSsv+TjjlfcLHjLm2auyRuqcut6QZC3+fOmDdtlyjVhXkX4TEZ2gaXX6zCp4SIau+yl8gYP0g9
SaNnjI0mDOIyWRrXmULXPWSDWosZMVMe5PWh1T0EiHcXP2D3k0han+Gs8Y2ok01BOEpHJcRuE8O/
BVcoK7Acbm94mZ4mzznAKorX9cuYWpgd/S0OOpSfieiCJVyUyzHJoPku1mN/CFhMZGBMU3QvyWim
o3IgN2QnRO9jjG3U2BQXF4Q23aaU0TETqpap0pxqBpItWahFExEEm3sEkY8dOjDJrWHZbEdZcD/s
xlWwCNIIwZZMfP9juIFvpwYhjl1Lq7juIHFAa9+J5xCyxkk6IEVhamwLSNadndlmanZvQH+Tzon3
Urzjoxwk4CyAT24PWlBPHgfTKhLkn1AcFMdOSu3+B7jBf3wTnkr+71rpAFkyTAFc+ntJC5W9VBbh
3EzKIIa32aYzLfwIExSlqxrTglDIHbbj7vd0ihY6rbL49/T6TPJvl9Phu6RiPKg58tv/9mgwfGll
6ktgJOOLh5HuGu2cMu+1KAehDLK7mJk87ZzfyoJxttqrsZOLp3L0TrfHuLQO4QNypH4FHmjF5R5v
LrKZqYKWqEF6WbIuLVyR0X9CvSySMjv2NCASzu/bhtF0aCJaJSFOTesJCtpxTZsi/szeHb4ZV27Z
issJ4zOuhxQa5xlm2bhQ41tpm3T+0uHrEn9hvyMFJFrgM0swsaoqgAynjRTrK+d1eGdUbfBUb0sI
dAgIufRrdl151MMS3sy1nFciIv9eGyolU39BUdb9+5odYon4vOsxbiRCZnyc8M2zwjdyxRJw+m4y
ST0qdpnzq5FhLJ02FyxgBQS6rptJCiugGbW0rggYCrKcmHYtimTbh7on6NdM+sbeD2mbE7JIAiTR
pwymO8iHZRWrXDqkMqjaXryax2rbuPGASe+KW9I8Db+H9pvR8Jwn/dzyvC+7QBLJq0BCfo4y+Cey
Dc+yYiwlQdIahx+TrI74svnKn42YJjvNAvVCsWqEgeQSgiwqs+JcWBdEz+yrD2HRkvoXMkddMes+
WbQCI7+mQJ2Q4kFhxQEnbho3Q6z6OporiiVRC/Xo3NPaCgg/lt5cpJJeLTeBE90bv+JIkEkcfJnC
Oyyvd9PEQgsFBXEDX8qZei8VdkevV5O0yGL2zH1BfsGkM1AyIVO4TnbAh24jylaZpkDGtqZwf3zB
JHv8L79/dTXQ2UQqz0Yhcj2SGkv7+pEhepd45KBMOm+K96ry64bPJXI7Qif7KzV7OollQ/2+ZcYF
CeaZUYnQ4N2qZTOwXRzR8pu+1WLNxvaX7fSvJB51FTfGiUifDRDKzbJ/TGJnfAs4A5M9RkEKS0OK
iPfs+Uxz8J185mICZJ41u1oskq5zgM/N3hlkBBqBM7oz4c+puxX/bhU9BxDQyG9lvgCbPBIR0j8y
+HnU0Inoca/acNeBPkkgElVXzv6iwI8MhzxVqCdkx/3/0gqK66+VUk1nIJPvrFScKK1vFuilo7GR
jX3435sWLcZ7Up7fvK5njbbEO9yUPtjcfil/Nz4oBa1rTD8nuosni/ohxR52wW+vZHUtry+LrVAC
wuIUuG6cQe2yDlZojtu6qcFtkgaZh5WcVFZC+6DFI2iM/z5nCJEGsk07UJj1+7RfuewkP/9pvm64
NRMm9xCfWgkglAY2n+B2zUs0bpmuPRFwavxHx9Qy7NDqeMvYeJXmRgLVf3Z3EcNjLXLz2fyKV+9c
/phkYIikfzvbyfOz7LLjFl2XAoW507ePWTye8o6TprFi90Tesvji8kabqb5/ygd4IHiZ5470ox/p
VnKSJWPa8zl5lEQShE9OS/3h11FUceMHAcc9TcQlNk57HbZVAaqWH5kQAFKsR3kv/8HrYFxAJU4n
6kWDoO4P/C8HRIw8EuIg7BnTeeMuOQiRNLlA0JHjvbfze5FwHsxsFqXrrVZD68DDql3ackYdgPmX
Polq7txBODiQ57gBnMw9XdYqkwKRhvKzFjkF8Gk/eKQvQnfT+pgistMYMJFQLcxsswrItCQtuQXw
GHqN7dByRjVtv8xSIqwuSTN+G533iYG9fAJPBtBwngKX+RndllG5MKjRcN9idzK0QH8e4bka03BZ
s3sPP2ogd9l9Em1KG4OW8iW+jBS6itlrZcKrROR+L1+suJe2UxPRa6VKqErRxRlXMNHqkUL9ZaVQ
9PcTUhT1XChheruBOc8NX3s3hQDPcUnr4z21yGl7BLN1iLHd1WYiik8+nN3DFtoJHFfVwnpQjkH2
ZM6FxgaG7OgzYtKYCK+qLrYeUTfoVgPToSwvVZv+GP0bqH82gI5GGu3wO0X7ldmdV8NHZNmvkwRx
HlXsucyy1GkauG/Vy4iqiq3U39+T+UlraRuTR1nguw59cJR7VmsxdeQYoLALJu678XDO6arlvGu7
kGeVMaTGW9Y/pIzoJ2O5sa2JjPi5UKxZRGJNBuMCcnJvjQB2jLATDLr6ZNPSgLCIdt7uNKIGyf24
BHQQpms0l7cIFxlJjkR/udvc/fT7qILKlHYBgZjz7aN91e6+KBfqGo4IM1V8pdafPdWKbMRnmH33
ynjBQYnaVphbyyODp0++UqEkGelvPpcJwF9bmTpO2KWAPT20JgPjh81HEwsu6vKmVLGvvj8zr0YE
6w9Wj4Z5HzFzwFJpY/KnwMrybI7YY03ovq+f+h+AixJQ7hxrVNoLoDer9JwAo0IYGDLl6dijHydS
W1kutf7n/bQfQ9ups22ZkRb5FGn0umA1uIpd7x+Mgg7mJTDlZf1MMFBDfFEJZZIcbcY80JrrOHts
A8SYIeHaDHs7ZS6uvm9/EY8VKqPxEacB4FpIMdQaXr/XXJ0C9PqOEr+LhBvZEsQ9dZ9A8bEPPL0e
vmu87K1EGUOQ5g8CWzOjNln8hWBoAzZHIu4ezChv3kvu0Kdy7s1ryRFFYNcUOqd7nGvr5L1GeKoY
qnQvADSAf6/CRS6vHjuyHkniaWRP2v7pUIfAjSl7+pqS6TLz4UtJd/aigSAe8d2m5NYk/N8ff1L1
M9EB1GuhbDbtSp79WWc00sPdjMHBWN+FhVqeUpn2asnfHy/ZWIsfyv59V+W7mbxSMj7aUFiyGOoH
UB38+miNopQlTLd5k4gu52SohMjvqNhWCd0awDNJqzDKdOJMF4U2A53Jg2cWrO4KFb4w7X+YdONy
DiFoROiaH95U7mTBljSCDnm53mo+pPY+95/rBRRkIHFWatD0gQ4lXV0tZruHVfZl7k4neZJUMOpE
hPYsVHVqI8/E+cZyEEf8Gu33YUd2tU2Srpzh0AdAcwjo7Dm6LfxloKoGQ+Uf+rmP4mQJKSgfvbNN
G+vD/dj3dUQ7uvVR4lzQCJYQ1gBn91dSRvdAIPQ/tbkL8QHxKt7V/UcqLpe60O3v2l6yLfIRjWMG
6Os+qQgJ2gLl7NAwVFolkx6PWBm4A1S/c1bkmoXcC3Gm2BIYT6Cuobv/0rsb+Oo8dRfusTZ6Rdco
RabSA8YulE9+S1U9H8IQpxfTjwYkzJHIZqLn5tyz1xNMYz0g6Od9eEiR9uUNOxsLPRkq5WkHAM5T
ULLAZFzMt1QlEPMkxstaBqgpNj4BYjKmK0U3sVPSlBNqhhD1NP0aezkx6PsFcDOmhw0tLf5I5mMa
StFUXRA8Z1FcSqAmpwOLYufiPvEtSq+ggqYf22OyEQBc2vmS0JVmh2oLu+j1NjYoi6Ss5NdbWzNW
YycwUAiDzPm/xi5FWgDUkO9mZWRleNz20vixP62FzfPSE/qV1DDS4EDGAhDG2ciu7kyQzDkVrdk3
tdkpSywhftoltBXaf71zqtOLBcssOubqTqwGEjoOguqQ2QNucQUTjeqtC18v/xJzx6yjOC7cvPp+
dJzny2Bud9cz7bV1HfmWAfMBc2ncyl4+1hCzvSsBAm12Ggm3gcl/rq2QrT0ug5Vpw0h+MAvx+6BI
RCSfcO1MHe0xIxBMtN7qYewaZA+VksLs3p+RdZSK2xduJURAKrbXuD7+dpKljjFsLmSBzQcTYC1F
PoWjg0lSjs4wYchBVr+tcBb9+o8Ve2I0aFU+otf0QZXVc6PNBfO+527Q4JCED033zhX7ph/F3Ckb
1gUXloKD09WWx1vGJt8s+JVh7DZ/+7YUqqmA5bOWmTRzOFF6NUaolrNVjbnGw4b4JrBXoALp9S+O
N3Z13mGOE0RhQxtJwlPmTINaPmuP+LbLOgJJUtytv1ucZ4EfQNJzPHGVe5GN0K8wR5VvqfCtV/o3
uCRKeKSRP3ZHIShArGwalp/SyHaWn3b9byCB+p5rVMWQ26uY/l5NOWEdxvh6paTJ+DdvaW6O9SSZ
GICnkgLCV28dBajHli4M/j8bnZ1GBjIDVPcdNf2VGpRpQlEbLbQVq2+ZHwpXyPx3IevJG1GTXYI+
NrEff1UGO46gTxpGX/gUN4A+PulV2F0Jo/G8UQaAGYk5iC1s4z5K2JHtFmxyf90Z1gpDcz2RGOqN
t0wO19m6Kdj/9K+/UguVNv6kIyTG0wAzL6ufBY9cZQKsknWBsDoyGDQsBOshaps0YC/FiVmPe0W0
lY4gfsf4rcZK+0ivDtV3y++0wzAE/Oj4l1A5xy8YjDxjTvRC7D8XpicbZn73rc1BjXGLNBl47BBB
o7PM+LQ8AH6SMUbl5KyNU554SSGV6urlvysKWzctTFux1geNeGboBKMoTw27bhQH9LNq2NwrV7J9
uey8XhI8dYRvUUE50nFblVacyqWpK4EhSQKbBGwW7aFl+33FYJTepMUT05ACr2KJh4J38J65Ybe7
TWbJ4kpKHFszWmbxOalRRCCxdFiEcDOnmAPiunJkktkLJqOyJI16cFm28wWiw7CdCWZ6O0qHh1Re
pF5a38uvL7gR+5eZ6ZNpjMXmZLIaN/oPSsZFOfpzZ+FXPKOEPyDCWZZ8XTvjaS9RRWIIqs+iUpIS
8ExQlIhl2zHdYGqtIzLlKlLJ88iBk5FK4Z8dYA3EJOBEiimY1OeRsf+APxk1RO9bjkvgzPCaXxdm
tzToFMnQdca01p/ePPIbr1DZLvhYKf80LcUuYGiSUdRgH10Pe9O6M4Ys8+lyodqF5UABbRstmAGp
O1B+JfFgahVtmRrcLKh5SLmmrna1S/Sv60reGwnNvmBAwKoP4qPhcSH+W2L6umeQUtfW2CG48b4w
0mtoi1VUaGSG/KCzUV2h8KmLvLqkf/fx/TWVOuTfTU/hsDHvl8V7hq/Ee0VKJY9omVbclU61ANyu
H4kC0aqEb7NjHGmdeDR5kZUmYq2VERWG/TPRu+TTh8pgS2/cFceXnpGpwWaDsZfTx5KXyR0giyXA
QsJRkjUm6U3/Y0DN0a4fw5hfuiAdbHWt9AyAW5H/BQn1G5NlGloa37T2XphXKQkZrFluWpQgSdXW
BcoZHsSQJv5WlnsRgrdlRWuQ4VmysuT3e3XAJdzg9d5IXhjXm2hZSV1lHEY4CapqQUNUvExRirqy
5OGZmNF3RbMtIgQJJebXqc37voFlabK/plMmX5iwuvF15YnsQxsjrln/T/gvQ46cntBmo22GnEs5
HgfWBVaD3t2w0CN67+TI88hVRX+MSjIkCMN3pUD816YM07U+/VJ495VMS7JIR89dHMmtqqbhW1j3
ZbSbxzuIed13QXIscxWbQEqvVxsaCwpqcExwxCd1m0RNiUuxVVBWzjskFQPBOR2D6iWl3QLCFkRL
7S+RQMNnA9y7625VfRMx4q+uNeP8+jVYb769KU3c6oO+hQMe2Oeul0zunbL3vOsd2CC7xTEyzLA1
VxECCvJPhB3zQWPCqhMOjQ1JevxTpGfBDAr/em2GnHLPUWSldswi5mAObrUkXBKr8MmiVEyn1wpJ
ycUyKvx2gycPk7IfP1atVBju915XZc0+5s3l4LCN2fLoki6bxP1/2f8zI6u8oGp6XSMBSqE4mxTH
7ZxH+0j5azUS9slqX1txvfoF3NeE9YGQyx7wdSOba/GG5LIXYVVf6HtblwguZ9hBNfdIG2+scM3c
H1ky0Uo82qR4BmjeH1z4kmsSx78nDXgeqRUMEsZxBN8YSW8dVf3PH4i/DRD6QoK6tkutKA7YVkLx
d+/UPZpcEHr+BX5TLW6oQGh6bfxgiwi6Sgf9hqmffH7e2tSazxy5oMyzdCRgyfNhSolIcrCU9qru
wtqv4AN0hGHA78IR++86QOJ/UqKHmES6PtMf04WiyCbwBEki+OXcXjzdc+5YJh2iHglq58U8MXhf
SgMYoUUtyku4V5UpG5+/yw4/Bd5ySHcuBBelOFvtZkmOadWayR3sh2qQHMg6yV7ZpwLrtGycrtOn
6lbZnGJNEUY8nh4c+Q9OR2wAkX8P9IJrMVM/DQVNYX/XtFZGHLNVmygOQMt+0lWBvoQiEwVs7/fu
BPyfh+4MtGacnzUzLMjeS7z8GPx+627fV+o2stHOFZeFUIhsIoVTVKRj4XNVMPrJIiMF3s5SEVJ+
uH32IK162aDPHV62a6UTxQiGwKSMJJh98fxhi9xAFO2lrHZkrEXkxyGJrnAq7hAP2HZjKgmxGsT9
rCivs+1+79ditwOwOD/9DWk+J2Ms7TlSRjWkuwqdRKdTDD+Vf3t58BMqJRq2lNyrWfQKNuVJxYCO
ZxvFrrebeE9dzC0qvLjAfPcvmgapU/OTx9AYhwyS+IY3AOZlWg19ZfRunJl0TLFfrCm27kundi/d
PJ3bblDZpkhDtCAsj/7xSbtTUbEXnhlgweqwB+Ej676amwRzAA0ZecQcR5rc253eYT7EW3ndSmYE
3EM9Ysfd5LoyuLm3eqPYbyZzMdQ6ZoZaxKH9c1WnjJ0pFGP+JSocFSbqrbPDt36iniRgILwoJFgE
iL4MnYpFacVC4/kj0N8ujhqTSPxQpE+++S0jWeqCxq4ATvpWKWcqRCzWS5SEdQerDYq7HPg3n8gO
Va8v3a6p05cYtPMY+gKJgSxPr8WENGyb0Pkc8NmHouDJVDAmyTrOULGjAU1yupRfK11wV5d3YdQg
LO0JB3Ob5YGLPLrG2IHzbGf54R4F4XAHi8gdwdBDXR2clqkKx9SoheKjjEq13lWS4UifdmGTB/80
TX4VpWvTBKHFYomBRhQ43zeCWgkjbemt3oVThG6BzUTXNIGC3q9KYYo5VaN/zZgnelCB0XR3P+WA
KTvTq4KJorm1TKJBOvgqcICmh3EvY+5ahugigNHUGeM4kvE0r673WlbccLq8A2s7i4do/dNDMKIL
PcSxDWCmqoQyRpfQ/D1NEw4VVSvn2bkSk9LRu0EVJrO9cKEnZYrgo6z/3fSdxh0kDe9VP4b3DYWl
Jb3YJwe1E+OrQ5hVa9O8hvQFPQpoHWCHqEERohMQxcahLwh0YYroFZmHtHIeLtPkVYIRG/WwghrW
gOKpzqKFWMJ3UGvjWoLu0W6Ofl/ZeXC8F/CpS5xyGc/7zHV8PqCuM+jIsVCeIi04m2seTrrAykjU
GaqrG1lRSbbKjU2y+vwJmFajdF1TD5R0/ujM98VGme6TBW2P2BMPww88OHi3CXxHjsBySq2kQHrk
Iby35W2q+lxnPL2Z5CHYgjz9i7fE0I9rX67TPy44iu0l64P8UKwjeo4tdwIkBfRmKc+3A7Wauczv
c/uS6lv+KA+MBaoXYFsEfos8rfNajlhVVBWXuFQBhIJS64/fOjK2OS6XHBSgs4fO2hoMBOYo/ofJ
rA+ooWfqTe9tM5iG6tOWAV0xgzFohCpTyDN9eC7jtzWHKBusQr0M21i+m60Ngm27eN/HC4u5N2oT
Yn1FScyk+L53LlJG64bDn2pHuYzz9aEofC7mw5ly3G3qK7GPnehZHOInpvpoF+dwzLuD0zEpQXib
eNw74jeisKmSqkwhqsEE2sTxjh74Vai04rASA3Cz94TCQ/gGbAyEvlSpQis9sfqMxMa2E83zny9c
nTBpNqU8wEn7p2z56VGnVN+D+ooRzcZXihoOpr8cDkmbgoqyxAji9GaVTaR0DOzFMmjXEIx1rGiO
lW7OwQgodmUVzE1IEe4bf89HmNrsrCUNwFFcGHzjU7nmp1qlXjqiC3yvpEkxc1CFDAbpAKKhA+nF
Lu+Ttg2ISlp+UTdgUnn1CiVyZPDWXcgeU4rlwXDivJdMjJwtSEXhGDAy+ni9M+A995fms/oUIjAx
cV+RhRE9Gk2PHf+/lkmtuXyHRXcr3sB8yN//hg6oXU0tsD4lsqWLEFiCjCfbZ5rcekI6CgS0/K/Y
iJOKzn/J0dvxdzwQi2tGFWRgtWJeRAf7g6Wrg7Q8xbCs/NOXCX/pJO8MH3682m3DSGSA7JOoJhzd
zWrbvuyw2DinYIO6qcg6MQbRZJXCA7g9XTu1ZhxCDXTsNHAr5fD2mhgzMO27ycSOK55JihdcZsLg
vzxdsu7TSt/D8ewETQinXrG1FQ0w2LTMn9odhhDdzdBItv+3nPq0AFDPyf0kayYXCV9eCmGOU+W0
zwrqF2a9Yf9hh4Bl2qxqGl7fMkYF4ZtCa1L+QMp948kNek2q1SPLOCOCcD1nPtWTo6AgKdpjhAyy
7gdfthVbS6OjzGzxCNFiNTUyNJYndcOqJ3Q8nioP//Zg7RSdm+ewdFCAmQG6B8C4DCNsNM4rB8/0
SQ0Vy3t+nmbM+Fbh/8OvItk2LoXxkEGwkcg7/oVh+WNLuC5B6E9g7QsfBlO6S8vZKq4yfOUVs+la
HjxbDTlZoxJ62owhp4lCivKNkvqH/2y+/i9X07Tem/Pq4zr0wL+bs9w44yjoFYHgWF2wcQF/0frU
4mz+vyJQjx3basDPHO2XpwuIRVqvsqh5zNhCqtpZladpXLtWaPnPSNWFJ8sxNKon8lRywRmIMrlg
u2ivDZxxav3S/dr6zddHYXbaufgmarTLM//LllSpnOQ6IdRm9g559XbkzInbhXbMbXb1LV33nX07
FR5joXP/lun3W8kQEtg+HCEfIlQ7cjepSpNnsKQUlXE7cwJkAN6XJE+y09Vxyjg1dSC/JusstqWd
5RSQgB3r8s1Xbwuv5HSofLl22+OrMNETYLcd5svlaFXYwXPdHuPawMMynf5VCOhfChcXPLJHmtKp
zZaL6AAW/lMB+Y339xyYZC9Zyvczf2UfDbGjLqWi0TWMDyBhgrQJsvh7HJNAC4QD6khB1o8MYwKg
pmXfi8hmUJTw/EI5eFeIYVcNDExfpsHneMliTV1GJPeRRyCROnnjs8JalpZf0Z4qMNCOHYnlAMRT
3XUzWmGXwgVicnumJB5vZ0b4I9U3rbnqZszP7thmQkLQpX6bADtjopyGP7maaLeJ+pOCPKe2dkxp
819/G7oJczvsaDsAb0FIu5nMl8fa/tHup4aSm/W0UO1IbGVaR5eyNHcmiwNGP07bkf3nzmnebI/S
gYWhVBREHZFd8hMhyFre4WbIJbMYjgTbZYzJZKG5jlSxSpz+sPugaTJ2T2HaAADQmZAaHOTyLu3O
iEkOWAqqZYsyjshV8qtN9wt121bxtDNbQZyKTyA8rHM4kwWvsJG8Abtr9fjwIXJ5Z+FtTfE+xZZL
aPZlP0zntuPP797gvxGQQsgZd8WULVlM4GSTsBU+0aaDRbVFiGxG3SH49Y/UPeDg61eVZyhw0hrw
IahdluBECRxL8t88R7HqWIClJuHM7mR/cUpK6vUd/kH4ZyIs9o5o3M0CxsEWne1YplpA8rQoTDcN
QlU5TIwccsyvOxrwbOdCPDB4bIZDuepmu1L9VeDmdUWqglXOHzONNNhQIYuXS1IM5or6RvXbOtUM
pG77SR1cM9IHE3xpX3/4uyt/YA1Nd3bWeyvQaRhxVEKeru7ePd+p/nZaTY/IPMhHASdkx0MdHbJG
NMBg/JW1KZG57dWSjim3rW3L/kdwpROsC1Xn9xot8fZSM6VZPNfbEtLnoiSp/lpTgivv/eOJ4Mql
WCtZek0S4cWwzwdSC+jKeojm1L1vJpOAwdU1r9dPU5SBrK777h+Yt9BBIPXiGvhnl9WY16c5N1xh
UWZLcUqAJkaZXBy4ZX3TRwh36POxGFd8lCYClNqoJtk3ti1AzqRJnVwyvGcHShH/1KclLHr9PJ4S
fKb/MHj9KPjmbq6gCchIqr7Sz4uRmQPIdHOXoDv29itlwmYKwysIZEae1sTHYbbNALoSosTNIekL
iu56JEOpzkeWka4voVDKYjg1vd8OJvuh2okTgERg3WGQF7jcFJ1s/meWvf5Pd3stlsAnOXLlNtyR
lKld10+0FVDEALY2ZOc0vw1bybl32n1HarKvUjY4XFJ+0hKZWqtEsaO10WVARussjuCTk9z5LoMV
IAzp2mHMVWVK4hBKn0M6c0u4DyEqdWiRX47LRuz26YBNGGSg55/hijx6/GTSM7Se8SWLHvG1BI7d
B9FhIFP6lEshiiddbuA0cxOAs+ytsnJqVeSKQU9i/8Haz+COQXnD3Iyc2i/dvRo1E7rV/uTDLE0m
AC9Ah+HTXR/OF6u7WWOvNguo1KLjfnnfFKhZZeaMjpKGLJ/sS04L+0BnHQmgD0ZsKYHftow7/2oi
dgD6ujFFKh2v+8hIniV3RQAfWgrlAWO1t7NMwHi0GfLAkHVb3St37WZmXzFVGlRQFfwhNxslQsUc
czC3VCPA3DwdJ0H/ckfvihHvI9P6HTzErI3zvG9jdk9Y3jtLqdYq9WCYlj+1upmGxrSK3O5glyO6
vk3LQaOJHN4q4Y7qharsaJlk1blPQtVgDg19bMUGSKaRr9ZHAKu/LJ/lY1Qd9517mG9BPR5zGDVD
yhsprE3j+CN/JghD3wsNy24H3ZXSb6V6VetC4wznc5k2qo29SUUkSXvt4YAqXMjmbS3DkBa/xfWh
xS5uTkO2CRa0WcHlLVbv+4SMW5e0FSl3LM6WC4iIDCevTl9xQa+mVi3iDPcYtuhxJrSb2MCCLhdT
lClkah4ECFQY0OBaPoLuzHUowumiH4J7DIe9wAkID7csOWUl603LDpPM98LGK42XISs+Gaq7O6AT
rOrMidSjP0At17f5guFT05+TnbrmF3cQ5TlJmO1Ql4xVakI/ZTjuGzuHxAI6Bmt1qzINHmJBzbdJ
lOcY+iuGgygoko0TwIon1ubNm+bxDYLbObM0NwWlmSrnlVmxJkrRssKHS3b3+pzGFt2AxSq96eEq
JRs1g4NXlsG7BbGv9D/U5uuOpRb0+Cv/9B6xxwzz/CFOt84OuQtNCYv53aekMv9B5tG03F+gJkgq
oWYEgvedZRds3ENRrfC1VCNdQsrl9EhnnmNuq2UqJ18I4/5sMqJ3W+ZEG0UyEXT/WLL8fnMa7AgL
oQRxTAR7N8qMC2gU9LbeQ5f7uZlNYPAmUX+2o1b5CosDds6EeLyvzwTLYCR7sXIgChE6XyLVdkQe
1strKibjy7dk9rewuj1jpGK8agoU/fF8eOogFFXFh/39umg/TjMusbyONkNT1QMJvFmuVl4grpOs
bYoHP/CWh5y7KrjhV4cZaxjpv2XPsc0Hs6U1zphYGFOWAo777nMkCjVfc556WmlBsL6NdHEvd4wM
KbujQ0bf02PhVetRdmGjO8xKPf1h1a41z3/bCi84QRFWqq5Ky10f/fNn8BTZ9imqHbf0gjf7LfTK
2l127Eod4tCJOQ51YepUrg6wjiwGC7AnN+IvC8O0Ipb9yyzXQyDM3vj0NQLQOSZCb4oMg4bRqioH
gAbESDeU+M11SkQScLTih9i0no/xRzmxg9aonehIviwKSwS+VD1l+dJGk1q3QE9nNM9zhY3Ya0CI
jVVRO1HXgoB04qkbPW96o6S1BHb4XPmzEU+6a/QfUBcZ4Qo4wNJz7Tb6bU53Pddr11gBRt/+s6dq
5X4iZI9pF7cWjdrwqLCGsClUWgykGj/CKWUVFWBF1R2Ywz7UJncC0+3C6KjISF+sECwc4O0w1n8y
l6yydD5C4AfZZfhKzSV7bCjC2NUORi4S/hEFgQlJ4WTmv0G+gCgBXllC4EfybW9FLPnQmXVJWMqU
8b/tTf3zRkA6ukT/jKG5OKyOqwy6MGOYNiG2ysfN50OfZMsFY/9jjbS5sqXhnhufca+YaRoejr5o
JkOSEpAQ9ShWXyteHtWmMKKLrhTqRQXpPqtzlCGdzTgbEh46+Z7/VorL/UfD8HaGxSC6ayftAdTm
R0f+MaNgt8sOcUpaYOpy5kAspWychI307xfFSZ64hmaAJhSZkrja+XYNp5apjqjWBtij6tK8fN8N
vDCrzL5oPpA06DZYJYeWt+dmxB2zvMeDvFRgDu1KOG3beCzuFeyi8QDpz88Ud4Ac4jVlDIYgfdf8
zZTtGLn14NPmtT1OyXzlOoeEoZivn3OweTGlhApLKi7z99EVSMMNuqtZnAjxuM3TNdFHQuRR7S08
ptu6nbWN1Uqv+9eT9ZS8gS1C0kjLk+4bCtyjBzsmZlLB9IC4PftmlaRhoCRcSYjwmMnDcLaWLln+
TR23q33T+qRszAVdsGTONn2WA/YgPs9thtjax4CJobO/NLGCfOJaJdTXNJ18v2Nl3f7uuWewTcbK
+xQ5HbICS0OixnjLVutNQIqnlZYHYHivOZIlu56HuHMk6DEBP4O0gvQc4lbi5BPSTXspVE99ngd3
ojkYcFyl9HcQ4Z+BGyMbft+Tpyo79QsH3dyZNyPG5Ey2QRrv52pYj2fD7WeVzIz9KLC1CbC97iw8
1GNymzW3RAmTV7Kgdvg7XUKPcBbuDGAf6RwOxrbmns/SwDC90A/ZNdkIANHWkSlsriKi3e7BlPzr
s7VDGpy3FoSBLleiMrJBv+vPpg6y0AfO/yZJ+9058lhyrzdBnwPC7yxgb088R6VJH7q5xptvrQsx
7Dc3gcBmPp8xp9l1BIxgKRgaXZhd5g8MuARjH/Q6SOf8ys1IP2FBue/+KsU1LIrGkscE46tCcnkb
zDQuc4WG6Mr+GadIVpnIqMsHQsDRTImhzzyfSw+1r1PLmJE7fNbx6m8GijRZ1C3FIXXg3awMNY7W
xChpIbwlovZgprrCCSR2phdX7UX487ckZHOr9kD10SG6AiQQTuqsbCa1aM00DZsqTQ5j+VfSIruN
WWvUvmDU4ouFuDfSJEqYi/LkVCEavBo3VlKNhzgdi3kWN+KJlAKhAk7BadH8IszXW5OT4ovXL/4L
ZFrCPDH1oV7NVmcJ5Gt5rCFb9iqJzx3v1SdFsZ7sO90TsmODwHS8vjZbH+YkWiK+z4NlATrDq+FG
27N1Z48rJ3Omu0EHQcRz4r5HHGm8ZdetTsFaHqmkl3XfEMmkDpU9fUMDcPG72uyoYceY8xGNH9NH
SLfLZYowVr0jUdkwJ8neUKTsojlDxV+GIOfFXogOKsOxuar+PGtvhU0M7Bg+ZBhLmr0xZlEqUjC/
F/5F1/Jn+tSPgBasvzsCl0QwhxXFNduNzc+H5kg/vzpY+jf6Uj6TM8TOIJKuathj/7/KpcYdKyk3
puftjVT5VF8NJfMhyvHvqyGjUvwjrwGbQz2szkJ/DIjAsOcxhqSTP+vlNmcnYBSLUXZlt+StIML7
TAe5S7E1sdKjOpQk4w4zGJhmVfq9EcHSMfxxRJru8iq5KaaOtrhFis4j6ER2pr1wnSWMx0h/sFzT
IXzhEEbJ+u4TyVF4xLyFCkK9AxcPmjx8z/PtN2ZKyoDID2qdexv4orFVfXuWd9dSmJxouU8nAqVg
d7uTLjaES4IlcWJZR6XK75AbZhJXIPYDSFBU1EWi7jhij7sZdwKv3S5JDO1MBLFPUADWY+bQ3Ky/
x9xAllOiHzQ0vkJ0UY7ilSOQiu+aTOdf4DkA0ZLf7/9TPhbROEBp1peC4LuyHI3ZwOgTMB0XX0ut
/OiBPBZJYXwUV2IowIvB2mz5dScw5hlzQBj3OXWm2hx9YvvVCV6wHCNFzRDjEYFmyxEPbpouAmNm
YwqDjCALH9mdUeA/KgPPh9FT4MGgHd+O5Hu0wdg31aN52G3bbRxE0GYZgiwZB5iEf6H334hanUDm
vtFF3KyUMXjyZmq1to7r7G2b4NJN2BfN2ufgSEYMuANukd6jQh56l7nBTUd6YDE2n73269GWS72/
gfqTrF8V/BItrmlP4GiEiHVUbuo1bvrQlSnrqts3cfyjH7mjSmU9TMimLZIT0C+z+b4aGPWGkeW5
4bRopOQBbc4EC0Gf3ZzfI4pYfnkGFmNwu/pW2vxLJsPq6vOH+QlEiEZ4pych1MpsIm1J6opbDgET
ZIDjkXa7sVAiUdxNIzvTvSsyWr9IzWNUHKQuFRInefl6ApgjQiHKdcdlnWscwJGZ6uBzo2UwJXUk
PRc/Qyam2967r6ntkfR5jlQ3JYJ/U3GCV0eCgAHCjKqeSiTo77FeVp+LTzn+h0F3UFad+fsel71+
NjPLRbONMGPtjeVNrTMymx46fMuNOrBd5mwuiqN+aICmZC6QZDz4NSeI2nSrVVaPsHY3a4hJyCta
kTe5blvrSsACFx6f/25dkhYUWVc5vMV4ZcJU/GpixyI/DnV3kz89iwhGRdH2VIae4UUT0d75/VfD
ov1iTrLg67kNb93HC78WEomDXpDg/4rvdH6/NRuF9MiBiH7vW/hsSGJwyecoY+rPJPkBKrkSYRmz
PyUYlMt5Tv9/ZMWBkUIl19Kw7c/Bs8oYcJ1Fj+lAM6dSnAXspDj2Vynl9ziXWs5+nkwR3wP5FvX2
b0QF5T3LydfxFuNROKgj/VRuE5CbE2wqBcmM6eFtlo/l50Ldxzr5YkePmTtK6I1WtCyzYI4o61uS
U0oqSZ59knBFo2NK+P4giZQF9Y+zjlwR4XUqvc9k7ex54j3Yr1bwD0krxCIZQJ2FyF9e4TkcKbjx
yAo260RmKdmIMFPt4OShZNmFh4RgpfVQPOgC19W+Pti7nfBtGKsZ4L9Bf/SvZfVRezsPV7RzH5gw
byQbJo0k72nR7HnkgQ0bFBLDnuaqYdbMbpmEALKJWIm//jzpAFkccMH7cJsqmYsmMe0mjqMibyaF
rkcNYo43NEnA925tZCWuK/oNVeWlR1kix+K8/onKIxdBczuOXqJfJ4XX6gIcLd3W5czQ3S94EAbs
ZOSkRxuN2xWQOuy44l1JMlvU+E/j86OBJYq9XFr1k7XkgnLXmIg9n4qRTIZx79r7TqwTHh9uUGuQ
ClgwN0NEkro3nRDJK5q6WFq35SsiiE1/KEbYSxVMFOiqRy6wJ1tiLOr+n6vzzsn6WfGiY3APUI7H
Rs91S1gTHi4dWYsrb8U6xU6n8TTDFNcQypkVcHBpj76XWyXotwc+hoGZaog6HeA8TRKIYENl15WX
eGy2awiMnNw68ciIYdnJDywjw4rRobdzJh+a8Dvg2wtLwA8zBWDgdbMtFa3N+QeXpWx1WktJgUS6
lQIjBgUyOjS0LyxbAS0+Ga8ej8RqZpJgZBfwfhKGLjwg6CV8e1JzamutGKKd/cWaEhOeOAZzVxbS
8LaQuvObiz5XMaZMZAo6hItk8nm0UPF3QQ3QRo9RiIrikw7hWwuoJ20k4HYyin89KScm3sjumM//
WkF5WwPE8XCkJ3q+elFtGFnhLJV9oQ7HIxL6ESxa9ahQhDhyG1d60X43HWxhrlvd3IMsn1od+tUv
RMtAknf8wgtNbw1CgflfpAska1O9zCXf5hl3YiyYzOJ/19mNyyH/CnLxdfhq/mjN0S5VXAKR0xSS
t5rWjWgzLC0Enpmv4n2aqdJ+FgpVuin/1nqA5OUG1DtMlQuCJmr9IBhoFDrxl8itSNpYV33HClJP
2d1WjnmhQ4XBF6gZUbCicH8QUtA0g1Fk8cN4CARY78ToexSFxvOu7urskU2uKJYy2PuLaUca9cCF
F2RbtO5MMfKlv2BzAB2yosZBPJJRUHA7dbxvK6BvujmXcu616nGKYsXGY4ckO8jE1Xidlc95AO4r
MWzIp8m45pxHUstdGbsy+dNfJIhMuwsJY0v3WWkYh1upA8BrgZhhQ2D6yZBcqzoslJKdjAKcj8q6
Ndvzvqe9IuUtC/mO4tFbTpAxNb0RwrXuzAP+8wYonnUrD8V2hKxL1Y1gmjTRrLqaNkoPs+a7f0Ug
Cmf5ANsWt7FKsSBf4lL5Z8ykj3g1ZghZcYfr2BOdLzfWWAesyMPGvHW10gieeolw9pKeg1g9EcxZ
rENNO+Cu7AaOz0NRDhL/fumw3friePYHp5mrTLU64DtXUFOERc5aT5pnVqUIykwpsOeFfcXSixlW
l+hf2Yt+3JlzPMBlIl/pI5wlgJFV8y24oWSg8LHxhayYJMCmATJ9K+TQa2i+21Kxi9mTjyqWB0dz
Icqqg2GCvGyY7yvBiZJjGK+8qHjgLH7lAnHD9As20eS8lWIN5ZzPNZLYcefpJPMDJKAS+I8T5k+f
oQM67x3iYg4SLAFTvpHcpSaI2N2UvWBgL7xfe8FJ6XjwTFXOE4t/CmLdkqWqIj/6dfVMfbjm5R5h
NCumzdo35Ei46s8mnDlegojMmCrRrtWOxx3fEgQGe0RyezdooXWQrxNhKiDIOIldHPLit8XRFVk0
J4mmU9uHqAlSqJV9Hp4Bgem3Lo57vOFWoa4FB2lGpXR9YQA4f3q/s1xhgX+wdHj2rXAE9S6/RQ7G
v5CR+ID/lx3caZ/92OkEKtRf0N1U96xtsEECElXi11myvG4DR2TRqws3cudHtZjLu3A+d7x/uPip
0Zbp+slwW3cHG0Y6BwnEvZ49TzroXStOQ+Cns0bxdF+rFG4ONVmpz+t8DYvpWmIqT2cflnt8OClT
pe4EFBTmyDqEkjEz6NuvZJwDPWYVo0Zf/w8yoU5ly0Y9sQQaA9qNqwFRWf7u/ecmmGY7NFoPmqHl
bmZmjusytCypRapOywYicq63EWHN3K7xMxQuZYNmTu3Ia1eVPOCq0Uyor6HlajXZGXp2O/MBDrVx
Nv/GdGEaRapVhJL5evQc1cowRHeD6jL7idCe1ryNAbXObRU8wQXpxHtP8iBrfK9/N85SZTr2UD6w
303jPbhQWw6UszGexbIxp1B6O5wCbS1wulFgVm+PZXd2sE7XYn/8pFWqws0HKQLfhp1NoaCVvO4p
57xJ5E6xZFLEdqHJU8OHk2z2vg1yPDjHPoQmGPlD/jHKu5w3kA/BsSs1ZJW56ei5PLnPxTO7Hg29
XiOFw/Pww8zKhtSGWD8T71dJKU+vU6Fb2B+DKHFR7TMYQrKk/fnR1/MJR89c+rggLzXLP/xsXBE0
zr+CTX3nQw6bFHdwdiFpZHl+pSkAVNMdnHV56RspNDWkzRvSSzq76jOCVAF9P426s2kWav8PFwac
lbw2+TSe3hIY+Y1LEM+FBisyVCxIKrNOmjbKm3+3e1sR+s+pfhD7Cn1UOaK6IxFhBMtGkbZsLWCX
1FMkd+ZsPTTiAP/0NDDQX0fMf3jYs5D7Rtdza+2Waloj8tPFxVNK+Jlfu9673iAKukcwPif4k5UH
nLFNz2rdBILqKJuPjQ0o6//Pc5BW89GhvttrNW/bvySWcRShHR4Nv+rkbq7BGSVVN4XBNg7NFhzC
z1SGekN/CIvVgPFtu+zXr8fAbm0ZsCmxP1Vm48x2iuv2OZi4aX9dzHWgxnSIZH5atRFlQa0yA7Is
GpwChxl/OWJezpZztt0DK7Z1NGM2Yu+zUVxNNGr+EV3bnzSiUjVvXNbtf6ai06/f3595QTFWWm5o
T7c84AkCdHEucVmtKIkYLxm7SvqHdplN/5jWc60VqEACHORIwngQBqOPyVl2qlGLlcfTCEfGmRti
/pJtVGDWrjdsDkNrwKiVVFpl1MygMkiLBwQW0qt1gR7wMUjR/ehdidI8+RrejFfWigsVH8Wt62u7
Lbgizs6BNClkyNYQ06qhS4TGXFoU+cgt8lPyVqmesdYVI0jltgaScFKwnnLAaXxkbnmh7tcyJ0QG
/B0V+UuVOS8eyjSi7ianHRy7tPLnhyY3dE4O7U9KeCueR4Ro9ZVMVenKbUp5oaP8tFQbOUNzPptg
JMLylTFmgn4OGkNXZhi7QBHpu9erGafUZ8kK59cY7f71xcf7vb6TboSyz1ODviUlv1VTlRoc1uol
a06afCPaWOGdYPLfPk57ZtWAMW0NYd/0Om2ew+lEOvMTCN2DhVSxO866Qpo9Q9WOkxFgcR575Bou
FQ+cCxccLFmIHauwMTm88Oa4gi9jqVWEzCUkOZwfmBh2ETrIDBcqjqoOha3pvktLkpPPqr+rMLXh
V7NIiDwb6EqfghqsG6jCR1gzrM7uW61IWCP6BqkfKya1YWTsIMRmCSbcpIQgC7GiPClc1IZAWxmo
636tzdWRmGprH2XhCKYme7IJDZt8JwW0d6zYKqw7jKCdxm5IOR0NQ1AYhnFQZldpj7H77F7rJU7y
EU0N14NHaLOzDOZr8CNcdSASNZNCP1mmPwMSZtqD0uyUf8BLZtxKQmmkRJEultdbBhlLKQO+qD56
9SMwxg/KxHt57drh9IgAVrzkvZMMowIZA3u+BlFxoHkf78Lks6QZ7C8y03yquzuDIPOr/GNNotKM
fbNc8yu1yFt3IKdclY5WAnLFWa4GtB30E8TCEmcSDAm9qFTwlBlmJNv2wwCLArSmAu5V7eTcHz6Q
Fd9H/ITXl1+wpoqC5ca5y7SRle9mdNlE7QQWdOS9ZJRGbyfBXuCB0kGZNLukQR8VYxVw85wm3/5k
CwNl1eO7/CVTIY9VAJM3t7XoU/QfYOR6lHGpI49Q677Pv9qgj5tD6S81+y0E6+kdVdZP1EhkmF7T
3Yofw7xSB6adKvUVIMc6pV0vrOrsajQsBiWtsRAlGy06xTvgmdWHtkxpW5NtJtthMVvFzfP6BlFj
SNjbtGzl+LHbz+KA1/zwQ5M4egeD4/Wz4ICIQXDYeZ7kfJ5tCH+AQrbBEN5gd+jdX4m6zp4g915+
0Uo3e3ba/OUJOxe9pmfoa7xZm0+AZoDAMuwmCtm4cT/OYsZcmGsos4tSAjLrosmoaurrmamji+AT
pXxHdGY6yr28hDYLncgywalfC2nzouenqyETiZw50kzW3txvrzOTKsZYWYRrBDrMkdD8VE/rE3CV
i1zGAdxt/t8oEGshhXsHPyk2L5MYswYabeZC0yjku0aqdOiR7tzrlys7kJ5jRAl4yDDax0lAWDZq
LPnxaIeHmiyhJB8BdRXadCidWvKR8KnyFmFrpcS+qbopqLDqbWnKj2v5NNr0t8fNsMLHBuozrdhr
ZsW6fkLsxlw21v+jZe1CCqitmvvNXkSZ4R1zh+7JmHe2QAlQYdxwt206FDmBL2rkA34ITzX0cWjq
b/UQJXr3NTGpjByGy9V+aYOfD8uAX94W0kE03uZPx5cU39QD+SvhIijtQd0XmvdkZYhTMhK7KeJk
E2J9NyGPjveF1qL/qUNoPtfdtAdxgkU8F1XNeK81+gxbuSLkypp3tdDQ0A1MUaSrSqGWElvptZBX
3FAiGELE3of/fUVgjRH3Ti273zKIL8jcncZxf/w/LZ395nQw0sEArpotSrJPYQ0f8wY9wThemlVf
YofOOJaCuPTc9o7YfBT7ASMisbTwcjcb0hp3ckFrbqsBOd6k3jS2/y3BmFnpz/fGQKG7OhDTCqQ5
H2ZnEseaGmK366uBLARlIoAg/j4MIm/QWMaJ7zVx+oI5qZSJ+eH1r4AXmlt2qxuZ7NV1MELL2N40
FJye53DJ3ji8QW4XIilqRevjx/5a7IFILdglhFUFWEbj5jQ7xN0/HJ0RMPZ7wAAhwsGv5Sy91uA8
O3EnX3Yp+o99OEOx1jgLPuq5E0jlELJB1dLunKpxzswmGNP/N1OrBxu9v+4FK7gXlFmu571u3maz
lOWJdq+U/TwmzGXaM7QlqgUV2MeS/Wbt/aWPdfG5R2fCIqpRn/XYdYuUPf0k4B+9wvPrBTIA8Suj
k+FteodSbJnov+f6EwUwyWAb7cmuHFYSUBiNBx+3mjdaS/1h3orQPAMEXm6TTfJCfAmoTWfXunYr
sR2A4e+9vyE/pX0TJ0ZsGW8Ddfs8ZX1ApxuzFXwe2MTFgr8NU7mvPB/Pw3J8hXZVfArxP2GbP5Hx
hdEDyalLgu6z8zm1BARXZppEmnHFCGJSbm+qbQvRKILuKA+sqcuFu7HIKLuPfMZtPrOAryJOqAmb
QzQRgPel3qkV8p9+OWg5yZ5VFXONH0rO0Z9Ei+G+ydKp3LE+n1Ii98h4hkCKfHMipJgENUSOwR1W
sMfxdAWHFJLgQFggqCGm4K9T2X72kKLzHOE2bsOyWzQfFhzo1yvqkLyBa9PHYqtmIKBLZj7FMhLl
CbcimR2N1IskGsK+U6EwC0WmGTnReKDOOQjac3iLfYqOKhAQ5xVZEmpgzuGPNHtcdaL/WVvc8Heu
Ca5Yl/obRDPDkI41IDbqAysPnLvvBtwbFSezd61HCIpM+xATrleA/g6RIA+w7oG35EMr+0JGHt1t
s0Skiy7v9MEiRGgP3SH4PvCRFrtiil/LQuVsa59YdoXWWky2nkoGuiAloMHkntt5Oc8zCAjF5g9q
wwGOWUwZf+jDGe+jF0hV/iQEDc0T78RmxeAJvCavr2kXmkF7yC+H5vUfYHtb0uWhxtHFt3Z+zaXU
l1AtzkRD1x3ZDRtiKGPnTVH2D89alvuuXpw/C06JC5wXU82DftzBCf8CsEfLhDJYEddb9a7udNY9
seVXLSHILDiQojS+2C7+WwUa7UbGEyucJI5hli0FdD6QAAt5QTacAQRA7VAxO0E/kUAn/6Mymlq/
flTOZ9twCNWRN6yxbS4qFoytfbRvG3rHn/0Jy9nJ4LAPAkeKpk+x2j/NpWZoEfkIJNJxB6IbFGTd
6WFpqm5gICXJ39eext3Uc/7i0guPjoUGnQyikDJLrKVDZ6I22ovyOyVMtJ7B2eXY1bXXUMSlm+aA
2/g+nxzKlra2wk3SNWQlFh/CWEdZvflJrOW9EGwJPYbAAa/0G/8jYQg4OWexdnDBfW3aOnT2N2eK
uAGA0gfX6e57y+jpvuVv169oACP9ubDTaYNigL6PApWkDQL78wY0sYJIQDeYLjmvxt5WvBtOtu+b
YSFXmHuQTTDbxZuEStPx4j3jnSdZLmPLSw26RszAobjUlgyoch0kVriNJurKGf3x3TZP7Blh1mXL
UbyKISDlDycs4lCOZpedD7vl6mWrnUOhMuRYAi6ztBwWh7+sVAdvH9spntMvkdsUPtSwNY9UZ1+f
hUUN0KCxQMKZl8Gt3zWky8r+fuZKuHq9dtT7RXiVcTAxf6+asRXDsyq1VXO1hr2aXa98sCxkIEqo
CJWWd7l/EQiVP40mT7hHOclc91GSsHgXM0JoAHAeYetcb5o7WO86FU+TSWiQWftSlcdRrNI7es0i
K7ntMEbX8klh6NcubA55/euBWGntX7C2uLL3qWNu0IVrtqtP/M6K7EJw3wfkMl1oqVLPstCai0rX
XF33vxo+9+sWuYQFheERIxuPCajPsbh1Cx0wU1MuVxs81aZU7heN48vhraUIuxlaylbGoTd+GMYl
65GDJXMOcmtG8/bZjNfa07E6hUuW/tMsP2sx+hc3ARoGodGRRzKqPPcsNw/FqMDs60+572hfPGiS
joQVAL1u2japER+W7d7z1TJCbMASQKvi44xCdwYCEs/IZmUJoGGOfpeRcGVnNk7T8tVkXuv0luUT
cH97/Pg/cpNNtRNTIvUCDD/hGH35wqgu+aXQ7ZNMatgNeU5B7TtKpMxm+XP/a827oJRDjbuCUiHg
ltI9RRFyQXq8c89Rf+jq9jq1tQfXjx4yOuBm5lvlzH0ukQJ0nTnLhfAte987/ZrvYvDUxe8q7xQI
5AhnC0u/XI/GmK5kf2e9x9B+49oHREHs7zOeDKRq/wlET4XkwwWIc1j1kIkYzNL6m9g4xo8ZNuNN
gTiPlMY7DTwtJwqt/GOx0vL9EEJAGEbNBHrGoBsnMc8y4GrF3GfT50eQerkBdLsC9rX73jRI6mMZ
/KCngsAMjU7Az74xiYUpAzYQnhMPyOxa5AFLhVYAphDxtqDk9+lASq7aJ69BIMhq8jCMaVWa5uO8
/PeyTjrI8tfeIlKSpEkX49JfnCyfsmgoikOxzHgmSnaoUe7HpoHnxXkeNa+GSYIrjhygFgyHt2V5
ljM5ISgn2xT2hx6zFThWgyAGYeVHC78aAojR05FpUKzVe3lHSqeA8ZTsr2Iy5hHUm04Uxsms5DyH
WYTOXDYNY3SuDmSgs3pZPBvg9tcXbQYFOTwiaUh96b1Wb9dikerfOvWChlQ1pj+wWSiyhBdTfSSv
UNm/Ho6+gpPVfQ7A7LEXNjQybIs0oTBLYSyD+/ZqPqdySvB7CC7Lb1V9ppW3bNhOw6f0sBXA3oFm
fA2u6NwT62yXC+8Pjux3xW5uLI/gyZkEGd2/ij6uYY3GkQNXobkNJc/MkITtQMFzkuPtKARYQHm6
Xad4S22CAyr2k8deZQn5Aj8jF1QtWgtHbu7mCRL5L2mNpD6L35bTI74RyIDQWOb3IxWxC/PqXdLB
Ec+eb8J82sKT+5o3SM/O9aK1nfRqoVWYs+yu0WikJcR3QeNEiuBzIZAofdmIojt/iKmRT6FaIj48
8Hu/9CkFry2AHX7H7rHgXdbtCkFllldQZyOst3N5Nsq29B6A0Wt3zDrF9gMVN26Bonh364Z5NNG8
zqBtAWr49SR84JwqVazD9ZzcqW9yD41RGTsZowJI5VqcuDzNT72/QsMtvFGGtN2Fp30u6QPyQH/4
+nHmS1ol1tbQ4ijew6kzlIoo1jJnLL9mx2vcOZIwtZ/mqo0/sVNqNwcizmSkbpbqDXMa9+zT1exs
FuE0foca52PPWSYgeVKSaPqQS+q8QIJ3Dn7YlME561g6ggF0M5JPt+DSBgWxaPXt8MTz6RU5TEP/
Ktp4LkX2fomQY02StbvlJwwkC2Vksxqeo8CUC3mX83DlL7J2erltsly7gj+m/YYMiOkcoLv/8WoL
kXbERFOLOvw5r12f8AtXxGGJVSYoURy3da9xHGnz0WpXx/DbFQzcv5mZXqwwbOAUKg0e9H/OsN9P
N3DluVjMFKDse/j2S0QJ+F/+Jd/OUR524MaA0aWADcosonrFqtj1pqZhFfv09I7lsLG0oE0VcWLm
ikmD1x9x94/PuyiHd1bsGW6H/pwVl3T2sGOE2A4ym0lRdXbhfbzanIAM/e0jNKg1xvyY5/c5enxG
VehJFyRCoPdRKdDQ17Gf3+1clhz3H+OSuX5aja0/axHwToeH0uYtLb4egNLNN8hPtw0eb/8rC4Zo
qhe4EQPpRAOnJ7kP/4z+GnwMY4Wkou5e6o1h0BpfXHV/47lpIz3uX5/fXG2lAiGcQFXtM7ksKQKe
Y5Bv/mZVsXpzvQLK/+7cvVoSipDukXbXGSH8LyC2aoWgD9m3DHM9JkaQjdpBFzo55hXPc/phuptS
9rHCVHMbjjbowtuFncZHsF+E9UJdnEd2tkDuJ1RAEFdXbrwmEiblQHmbTO3h1lz8d5Ixr34G6eAc
dTMebMNwYQD3s+EvSVkA0M2z0P5myIzZXjTkAGw0o/g/4iL/YEr72Z6p0+jI8aB95YCEfQQjEdva
Spc05S64lQxEYcvDSX3yVteXefpU5glPYGGB0APSfuaZ7VsceV9A2FpRacpx2ArCYIUMxUA12+KK
MTSilD1vmVt82YTwjZllihYQGHNlXkrc+Y9wkOcs59f1HLn5f1cwJWUJrARvXDu/wzErN51bG0ub
RKX+7KKZPJ6wu6aFdG2bbwCkt7vHOnZFnsdiAMZL61L3vu7LDLdsWE6QWrRErd6RaqU0/v7JwBUl
birisi6rSOXKgQgAQOgvFP0RVJsWZSPQyoctA6NVVeL3uAoYrfVIJerKecEd5TWWuwUZbICE2nXT
hnAMqtGdyiXxdhwNfkFXq/v+27Jq13q0wtZY5fNxoD+Wiefoa+wj2eHZjPRbgrzifDy1Cs6JGBEA
fW2r4TXrEQMWus0KhOo7RhCgOibT4Ntt0suyC2F7Z+daokw5RKnEDKV0E5BH8MuYF8MSps0RNLS4
QmDFEmjQaKU59Tt2ZabBv2jnvUdnQqkbyTDglxuEef6p5cHbxKu1zdqe/GyVNkkOuFI7NVxOz5ty
9WYCVNBEBPJUX47OrDrjU2Jf07dRipaCYGvpri5j6TnCkmSY1rUPmW4zjxs/Conyr8U4DhmHLULR
hz81WpHCyH3CrAB6sN/IsaG+GfUYK3Sgl5iVpmnV3aLP76LkGmA89XxTkApYK2dvM/i3+4g+eI+v
2zaOWmIumtWeIcYnDOdbIMXWUBepVcCTPkbQKuRRRQQ86osLKSfJB7cVqGF03nHDB3SSLHh+1JFJ
bBR7Op6ZI3gEMS0PaaiH8R7q18Rodw2EwyTTo1tHbqzppQATe6FsdzeZclj6l4P0blmQK61g07IJ
4BI5XSwTxLm5Z6oy+zye67eafHUGd+fTQsix2+xIOhcBfYLHKCl+dBAXT0lRp9ey6FTnDKnIJBQ2
FsG4w5IPxmrazHuETGnmCvrnDodSfvmzLkMWYcPDrSwqPO1Blf/ECfVRMZI5MPwmbzEKV0pJ0b/R
9t4NStHhVva4MTQHEna5QgV2cn8aBkIgY1al+3uncWZm+h1sb2WsAz64F0L/HjC4UBcsz5RVJFZ1
NxvSMdnvju041+G7DzXW/MajyxYcVhE/kgixCqH1oHzGkGTpNicpGxDx+5GLFVnAFfGpzl/6nvf8
rC4rhvj7UpjgdUrf0HYYdF5gJ6QSflbAX5+UPQbJ19xzRU2WtKMURDZgbKenlqNTdVeGjAaHjuaI
cGYXLjakwmKwYuFbXJCDzP6+yVC0SNxp0EDS+7KNHY37cCm1tSpnndjdjWQyF9E0HCBy00TNTDp0
T3RSBBPxQ8URRJ2qH/p7byuEdaMgjrWUaUL6jbsHmVGxJ0dCBdXzJbZQ+OdiKRt3+gvdsIRq0GC8
nMA5FEEreZ4Pmce5NmSURM3/fALxbKwpLOFd3Wv3uT4KDEVJZM/G8fISSqLyl7RV8jMNuxsALFSx
KyPoogDcKrJG5BwNDO2WqdO21sEjLba3xlIoELBpMuEcIsxhjw/Qz49yhM6wZ8vsEKvYaqMWlN5y
sdh0rL446r6DV/Wb79Xq/00ujUXmaueKOelDmtlf4LOa1gHk1lxdiiYfzS+1xXuTPPESowq7r5H/
80lnU7qTVKCuigbs+cKo3CHAOpuLeUmbuKHxC7+qh2mT4YUvDQ8ckOHRg0C3BCsIyqMaROTlHcMX
vEKSDIEsLRLD26LZgQF08Xd5rcbP/hPT1N60kKvrBE5lPactbJGfm7wJDMKEyXUjbPS6NikxsX9J
412z5cKPIWpUpVG87x6ns4CZenotPgLtE5GJGcut55OqTaSVnYh/MHT9iJzaRD/pP8pJDGdu7O3j
btajCuDDG11+1Q5m7kSYggd1wGoPeo0e+Fq3AlQwafBXDUGSG+QvKc6hyIoQQHrl79jilBzyX+Gd
owPlQjFYeAgl6/j+fP+cdLBN58464Nr+gcK0zXq+XLEt6/5uc97p7b43+QHTKVmgjzA4VCpwIYyl
qSs5oUwCTAovnX4QRrGlXTXauQtLq3ctnLTeecl5TlEWemNlAR18V+zcddWn5ToAmFpAR/z5DWaG
8Jt/OX8Omm0ZcUcPkKiNZN9EbaCoWZbQGw3/qaSTCHDFp03KWUmCDSQF5Y39pOP1nDzt2a2xWflP
oOKEf8re2IGjRDAWr6Il5PT6WOPYXj1IpFdaGKulA6eWQlsvAfjk6d8I7Q5cnVxyewAiFDHLWDMj
egeTlsqwb+l34oWNf6WSwcc20I3jx1ZzVQzGiwCexwHRRvC4HgJd2AKNWPbSSvPuWlTwBBJMXJMn
B/XKq64bpRYpe4jmXh4fl1rWFAl5rwbHAOnBml2eqGswTZnKhkuakJZnfHpHWOqvJG+rGTlrEdov
AJWPCs+Jm4poW4/Dx4Tnxv/O+qSpwt9MSdb6izBvJhr5YfCLdHJMFiFhSpHvai8w0NSDs5GKPUAV
ov2qsUczDqNZLBj9GFYNToS5qaRz7ehDheYT3kR2b2xJq9A8ANX6SX5UXhXjJO9OmqNKrBZ9GUBS
0LneIIPh/2wLM98RfLHmod22y9qzTvZELie1RUjaA/R7OOGlEXbhkrkWB9RvcSxVkp7mX4YP4h3p
LLgFz8AiUd7zaBVTVlgHfL1UltNGrm4LE2Guzz3uAL6j70Kxgs5UODm9mfEFluCQmtVv+O5P8n7C
IKYSTFRh7/NTV+OE709oqxrQJ8khdIBMIFkNI5ylC5wMOvG7iVKe8D1ilkdlv4YxzscCimswnK2T
DhoNqUz9sq/nh3Ytp5NW5+HtsH88LmCuR3yabHl9RPaR2Lv801HBuCINI5qw7ojDI1L5OYBkvyYv
vV5NQoYgA8e6w8DiK85Xan7YrQ8iD8dOiajsPlkANV3Ee0JZDhvCXEu1iqHwMBdfRGl8fYLwgN7c
LqK7IFiJPTmfxPOaTrDDksWOUmXwgk3F6sF8hUnVa8ulWzvAix+wRTpiarwMoEo3cFI/WGiyfwGv
cQ/hU1Xp+QlanBMh6GfHhaMwjvaBVOCMdtbgByGDFCGZZV+cNODK3/pw36tJ/PLsiy+QFuR1elyJ
/AH3LnJnonyJhXRdlLYgyBH573eQWwMD8aPaUbZ6rrH226LVbRJ9bqwg1qaoOJofZexqMCwfDuXS
w/ZgcU8ODeCvmmdf3QzedPd7Ld+2ElamDIhpX7acHbWUpc55YroeqQhIaUtu/z0hnWvcH6N5WFiA
GAJzrLKNo/vfvsW29H8aOdwckzgjF7pd3htSugltIa4TYlnskKyQdUlRLFhr0gYkQcyl2QTv9MB3
Hk48v4QNE7sVU5UyMmTH1CQh1NQ5GLLGd5lOjnhKnldU/zb//W7r3XEpYEomHtuFx9IObU7zQjCj
T/BfLGFYuPy+sCtSJmVtIcCGPyltfvLxCCbCt+Rm1ztheMzxTmIwjvflPUJQ3yC/Ug9K5jVPGxKn
oGgH0NnFWB+gFBMT94iYdNHKKidHy9agdDN0VQCvfjVeO5k9EFGJjt6mD9xu2t2sWuRJqWXIKfdG
wfZsiT9i2jffyYyDpJhTi/avZhomP2lX81cDucVTVAC4eyOEe5Keww9ZT+UclsgK6hsvdybvIvDv
Ehg8ItSPRnWTkagQnOqXW9fXkzV6nShWMxHbI3srt6UJsqSqcnB1TfcFYqdn5hhTNkdUVWobPzKq
c/75ObPJL5lJp+70iv6dUmmUsvAlNX1UUIZA3a7sB3KfiKWE81WU8aEXbJeuqVRuFMSbBDcT0t8Z
rUvs6q4jsMjuNqBDktRU4G/IQW9FA11hipEYMw/orTFEUsDZwKJdFexipDcQV8A8lPi2mbHWefhQ
sVt8XNByzFl2B6dsHpDViz/WGcDsy2LpmWnpfBuxSkwkaFOjez8UY0ZHXA0DwDQo8vI12KTIx8Ez
+aQFLsFthy+i6fdTsqg4b89J/D32Fm+XYfBP8Wwybh4KI7mLdZFIrt+qZF3aPyNyXgwhiNu0CYv0
RFcIAE4tI+k9pmx1GxclnCEWBYwTCZLZutoJqxSXcfKB1xQBbSRVL3wJRtZJrw3wqQrZVu3TcQbi
2fN1DUiy38dy7JXjyaOK+tpSSXKSPsCswaUtW8SYgFNnKRQ0hn/YnDv9RVbyePX7cvEljheAeXid
q8AFJsXiyldbsvxVCXDtzBX/sdhntd04ONQ4d24WG6iHD86WrO1t/N6/helRPPmLfcEJqjsG3IXP
njzNKF5ZjuXRaziqjJIzazRgglDBCpINzgkd9J/MEhkdVfDKONeYSCANc82E0uEfoK1EvSQmfaOv
HK+ZfzEFe/16QLkAvc064NTOgnQvgLIJdl64Vi29jEojCwjRDuLsnwobniZoGGJJcHQ3Q1NJAUOI
Qe2Zlmo0j3H1o9M533b5TnhvUXn8MHADoi4tNU2fzOL5KNdveE0vBingP0v8JbGLmFTwh1mYO3Qq
lPe7qnUAa4Yt7XE69VlkQNk+sn4L1xAiMv0gG9BNquUtMfKRtaUb75604/rb4EVyvmwzhAds2/x9
W20gJiKGsF92bwiYsqTVKnSfx4YT9g69XoN6oVCZErTZw0fUPYEZ0e2rEf77Hv8791Bg37zpR749
Kp+SeRwn5AjQhPh1SgnaWSrrF6hz5ovWmXiLB/TciUhBAXhW3sCDvSLnS4Sml3EnIEUB5WKjI2O7
UVP+uWDnf9JcVieFcjruow3AcLtVApEYxYI6YV9WHhGCBabEVaupybAax4MBIzdnsEEytGMBhJqn
I1JfkNdxYjIAxwxPsX8f7fTZ0zSBr1/xL7KhYV+jWsIoPPIXXQoyKEcSAYqwwgjsdaNvh6KBJcHC
0BGzyrBER7up9DOGetVQ6l9g3KpWuvLFit3qMpJ73aO8hg1w2wtv5nn4AFtsMycne/dbDMj1NKX5
JRhR4Pb9QqNFbF9hzjD721ZHiTnfuUdUMe7COrjp1AmyR8TaSxUUuYxOm+6oMIIA+Zl6o6IrB0A0
//BZ7iH1loIzdECy1CiamAYFIdJ+jjBzmPH10xFVC1cAk5MQKropobv7Wzokg0+JDRDBit0PX92Y
XArUFOeZlWSEI6yRVOFAKifawIDFEJdxAq5RODRF4JLrrN6O3Cz39x2wPxQYFcPuKYGROD705fEK
SfJx4J45Ekrsz0/iNfb2XRa+nB5d2cviJKl+Sp05zjhxoyzLxPLdvUGNzMkjR3I6faLzHaFC/JiT
IxYiXK9/UT8m9YHxrtCUffINU4t3LgDyVgiaJxkjH7KvPqeOgznhBeVRimuZoCLVqSJvy5ORHFfc
9t/9IOIk8KYlzwg7I/hISr5YiNVnr4pC0ovYsjeGhoWTJbNeCo2bLUsLxD0XXw5b0zJLQs0SL9Jw
tWinre7JNR2HxCLQcu4me0pJQphZFYKfUbS5lLBbf3mrdCaaeaFqa4mntHtq2UoPYrddH/CHt53A
pX61xacXhUCjZp3DexrqbiUFulSSzJAsIqsmoIO6ZI9selNl01M7c968m3ET+t0OpxpQd89mrssd
1judslt9tCRKBEFUAZapSjXwxgdEopBzh3zxFinN3kUgm7XdmL5Pnq1kkrG7SwOfPVAEkhDz/fJs
+wnLGARjCoMWvCdGscD8qqvFZkdQsLJPBOFcrGxZY0sdyf6xBJiUiF1gmDDyryNoOE8SgqAcn23a
D2cAsXdlW15MBAmcmpbjANOOKMT+MKdf0Ci5XcLrg6MtZfPIO9ZFYMaMrhKtt9m+32XjuU6OLdNh
RIVZ6BEnAPx8JNaHUD1oMN7lut+bXpt9CmtAYf7aJGsFcaKSakaAkB72pNn30frx9bzJ9D/RYVT2
9jREQ8d7cIntlZgLejcLJyZVoPT2IEWgdnb2CN09PJwIWN3DoNqPuSmTgK+hNcHZnmhyYNcHWacN
/5uE0wEGUlKJi+Lv2RXUao6WReJE9rCZldZHxQ16gpvMPJRtfkYfebTjPwBntNYR2ZW7nFe4ZQIf
B6Q6ke306nKwnKVfwAXYPiLTGstWktFeWzt/yH4Kd2RdMaBW+Y5f5DTDoUx2yzoV4k35uSinyFLC
BqCW/NLDKzzCgk+eA+0YHZ7Zff+k1dIrj5jxf+9xcVD0JO2KS73OkDGLkGD2CQTiKND4aiqS3X4k
fB0wHPfpdrGGPe+KSR/z4vN7S0PhZyYx1EGU8pcoxZe/j7eh8SrDv13tASEPWpOWwCNak70y2Z44
GB7WeAL5biEQjDjx+FU8efeXiTGT41QeT1ZWXhK+/rnPgZ88q3j4IgCG1M5fq7TlO3RqCVnpi/I9
Kxs/pzfLmExasckuWyHD+6gPr3cprKJNuSylJPRf/NL2z5Ov2yTgD2H1koyr2+05gsrrr/j2qoMs
BgUV8W5/rMwnhqJEgX/axTgKzhRS+EIXCaoqmBVWEjsUsLW1ZJvL7uHCF07GBIMyaBAMYqiklWHf
TkdjI2NfR4Ry6GItFgdthdBFBinfEspQaUhyQ8rExqVhwA1fH1RVlttvQ69pBermKOUqG+amWpUP
JGH1xCa75Toud+GET303GNLyQbDqKShLzy9ubrZfPkvuSSp5PE9WNWEi0pIk8uKZ7ZzXNao5VvOy
nXpa9/acWxr+OjZL0UmiPcKtfbghRxBJJIiWZgf5N5ctAMJdzjg4iav0Wf0vq5KD0teUDGfHa6iO
2mbeNPimxs1/OOQp0j4tEZOQWK++p1nmdQ4mT1XHywRPjNV2zXSNKvmC2OjIdD0f2IrITLanWTdl
KMSJRQ4MPATWNY1mxN6OK8pxyUMi3m3dLAMJ+dtFxYVUhnJTJzaGyKUyUPgJgEDheiQy7gX0bhFl
+ZVeut965oWbztXBlqlihICuMlKd+DvvmCLebt9FgqJuD8Lx7QEr7FHiNm4mjMuikDoG5FdKpbWa
PpiGZxz7czuZcw5qHnxgRZ2XzHPX/Igp9Amwtj0sHVpa84LcAgFN+1tLR+AXSWKjxp3gSPmNC3tR
8ExJKqHrQ/B/fKefo9u+hJa4/yo6T5IcxW1wQEyhwN0Y44IQuEIVlSHqSO0bH2tFt1UXvoD1Icss
me+M+aDk+oMb1GiPeyfy4b/WxQU5Cl6SZJyI1zGnnm1cOkVqwDt0PfcugdhLERPNAyR8f6gMXagU
NnhyNAsEPSvFF1hOcB/JxP1vsCt3dJ6Jlb92z8byzkGV4nj+3gHsCt/WKCB2y/2pmSg4thCvirbI
lLU5xchliK1FAAKzEZcIKWipc1CBPSaEvQsL21c+AU8KZvYJZwyTNEFtXNT2hYRv93zFP4lir0Ln
5y1Y+7jEd17E+L6W4tz/cVkuoq6ZA2DJZQtY2XlvrUv6Vyo9ndnxmpXlj/PTe8VEKeAcQB+YBPpS
fxI042hwx9IUAcqza/dNrHXmUcTwANAbBL2J6YBJ/iSd+Ma6OmhR9ZZuVI5HJUBWPDBr1yOek7Af
8yuHEYd6048bZ0D0+PUgPQNqmkLUzn3OkO+RthPoY9x8dpNWmiiNejChbtgFroieWhjwsviCSzod
aavbXNQ0TSYww2lRG6rs5LuyS612xashd6fhncI9R1NhwRv6313t51pZuEpxqk/IjuxLLHaWasc2
7oTigmnIHNysfZUZ51jI6RRI9MHrAbLT09i6gYBX3zBK9pzvhWCKi86J1HdTccGejMoMdault3n+
ReErM6+gyuam0PliY9+ddu/QIfDMSUdSReKakPO6R94pcWk+ep0gd5CAMZbA1ftCy6tc8yl8DtRQ
FuFx9SZgAoukBwl3YLBEy6pLFSkLRV+XX/NW6I/opycC62pSvCcZU3sr5JFA+0g+V28LcyABJ1vn
mfO/EOAFv0XQStdn6BLTGdaktmJGVQhtZEjVC53PLB3nWa+eN5ebzco1TJaY3Ku5mocXElkhZDfa
vuAr4yZ/+j3iQYuYhcCZ6XrwehdbiDpus3mrcYlLiGZXS1iKPmGTzTNmJKr7+9+LMJQ5bxwIiR9C
Ox8487ABZOfipxezLRvRrSO6Zs7FTMTpRF/CRyDHlEkKe1XfR8J0XarZj2ZD5IUNaZqXP8uhACGb
eHerKxCAJ0LYyYCu0WWEiRLjsuj3BLYOQD3QUg4jFU1rLIexCs6X4YFLVZbgg8BbuF4NOE8HNIc7
VMM7d1nxBdYPK8F05pxs3rmPdTcVxtreX2lfmiuMybeg1EH2fNWAwhsdBQiydI55adjq6FM6Reio
zU5/8zhFI/AbKgETOx6vrnQKy+lVY09ooXI8PHxBhDIkomp6You76/YqJllV6OipfE15yu9jvKW1
uLt1vYvOKqdBTA5nS8+s0+WhfF8NeoE851w9aPYvGP5uKpZLBbSfC62Vlv+Qdm/0T5ZJyozPUQMM
27IXC6Jgr2Wpab/ia9+X84dq+QnsYovnFETZmYgt2GUdTjadUzjTUmMqm9cY6YPw8nkl7lX0oUjs
JgXqCPi/6mPUv/37T5cpiCWrfq+PCf7gZpcyhQX7TnzyLVw+zeuBuEwEH/VEF8Go+HrbVahS6cJT
VQS8Ft+wIq0XLIX8Hb3Iz5EQUf0GUwrjjjKJ2ScfEJfY3C1rvt6+4OLJPpbTnlHJRQOPXqguQ7a8
huPmWtCMM90ZSV/jAB2SlFAbQjMrIiu54s2X19lnQCOHLJdY3zhbi5uYYSk+sA0m+6n27hAdc+SD
7p9ljgX5nZnSqC9Lncve7TG3fDUW29aDVjV78Ic++UCBEka4tzSVQHDJZTDBK1yAVW714EK+i9Dc
+6zFIG0D8mVquygLi6+DMsFZICUMVx5Oe4wNefb1Gd5uS03M2wWBKwLNgnl3G0hTburS9jHIsXMQ
oS+IkK11G8V/CNHthYhYdYo3aYQNCPfjrRvQsHUlmQsttedCKvNSYFWz402qffPZKauCHwaQjzkt
lE89x600jLXoJmBQtYyIOTDDSPpXY13MuJGaEJuxwoMMBDilkcwOoYUl7jdVjfSnxkxV6G/VEqnh
yvzxuvURfrAnM+pkOjFGNfqx94NMV6b4/JD8YwJOxz47bXrJ1B8EQvNJAjfXZecxZmJMPLugmBIU
kpp5MhJbeQjNXDz0Q39m0Kbk89eXhWlPf+W6rspe14s4MCq/p2fl/Q3vgXgIKDs+tat6q1PQ2gpP
434SubHkBPRp1AS9yf8RUpaE1vjigRuhoJ74ihqHBstx9AKi0mw6xmT75nTzEGbMe7dQZofinpAN
gtxzAj9+LuKQe2ObFErZedtYQJR5GxRdN8MzUVmTbgHQNIaS3ejcLYAuS8XFAvWNe0OD7Piqj0vQ
wUPKIRBI1fqRE7FUGsc4D3N8DH9IS9yl/RWlxeOCNo2s9xfYmN1f3yh/Vt8BoMIjQr6YGTw187oD
kYP2YBUrJ3cGbvCQTL85K7jjv7vgptwuvTRDE5kS9btXWJWIZOmV+WkhMCuVHMoPKUOTCpoJrYop
MZNjqwYBHCN9wGEMYj5KYOfbNAROjvIgO8PyD7xoFv42BRqruOpJ2e6ekF2c0RgytYW5H2ezgYxj
4jnno3qWVC81+GcIk5aFb9ODBr8JQ8aU3+vBjRPbB6rssAU3C/c5aKhNtYkhj91jGDthvLvPco/D
zZeJMtpeE9b3loZxn1Hs7yIlFyPkLbzO9hLHv/82wKTA7lo6mixegZ+V1mEIAPSlP6urBP1AWvTD
Ky1XCdETSWkeIYTzdk/n99M2E0SCXq3rUoovhdikjBAYCQoRLMIdNvxgam9kDNv4U9TCzYTqGnFG
66b5fme5k6VRwpNg6u1WXedwdZay0Xm9WifjID45ljnSbK6VFLiP37tF1WL5/jiqKjcaZGeND6El
vkpFMjvJFsOlg78jTEPx4a2LCoina2PNgymQHZBvliDJLrwENJZqm0YUgy2ZEPqED4OleL5Z0OXg
UkDkYV3MJAwZWaQOPlsFgdx2/hdUAKWcIZYzPWMEwntZQi+LqdX+6Kc12IBHpr/BaB6cMJLUHG7+
8Yy0ir5XG2Shduht8sbNgBg/aN+sGqshhrWUyImMpxe7vRipPha4utDlfcJZB89vdL93eQqYa+pd
gYTvGlVb4a5gRN2y1Asfe0DoE0rn9bLf4YuS8awgWHnnhmqviPr67quqAtJOylID9EGfti+hPLcd
bRoL0fLhIB+d9OGEUxZtwLFRQYyQ2gm6zwSOz3qbnrrmQaZsmHH2m5CsmYSwDYd6IsOnAH7dfuyU
S16uNQ/seFoaafy6bDUXWD7ciS2oNxvTKPdNGs1hocRHP+y7/DCbnawxbP1AH4caezfDrgGCYkJU
RNah6IMIn/Mh5z6U4LHqN6KFj3sVQgyvhbSu1xBifeqGBqYHENTb8Z64aEAODMMGovzxphKYDjDK
X79AFjRi8UOgT34rNuq70V/e2DkM1LYH9w1oO2EsYdpQET6wIbra5wDihsKELOl33Rymy6mQSaC6
FHDlq2qPUyvCwFp3sotDhUe0tz2lpEvmuv52ESNnZNa8F8n9hxI9nLe9EIDlTtzzCk4L5GjDHOVR
lT7jJJ+3x4h2fsODwThaLh54fJAAIriMTMJses1Jcooa6FXo2j/mSAmdsnat5hYJAyibxaOykjZA
phgO06it+2gOHSV7J1LewmJgSrdH4IB7qiv4nHkXCBMxW632SOwEVZfCGnBrYoWfmH1+Rab84bly
Sk67mxUnWmk+ABbhPIK5vuYWj9REzjw2vczhGyTmFp/eRQC64E6ZCwMeauMbLI1fcWWqsYzRNiKX
BPKlsTV+/t9gm+fk+NWeEuVpJCKfO4fKqNfwJ5DpE9dXgGycFlc2KN4WZlTP9tDGsj6DVBvathof
+leUtxeoGNQ1PLh7mUO6FJrf9K0HEf6NH7wauDCxsFJyQaIZbr/1GH5cj6GvPPXqeBWfVGlNhIcJ
WrHnOVl+LBhVr8r1cfTNZ/NDYEqBocX7QVh4YtD+YPgMRRCIr6ZEuxFuXzmmfQzk2aVm1O7jD7RO
ZSS5vjmbeJndn5YFv0ZwWGQwJ0QJHBJAK7xbvhl0+wVjdcqwDoEVeq9Z9ZAGywm5XzoBLRlpDpXa
tppQVdwUPbitF8AsaxYfBsCbJ3UJ0faiz27xfyLtEbOWE4YAb01dQZ1XdWCQxZL3USPdpRQxwZqB
SitUrE6XHWT1yKYyYJZn64V2jNMme0SI1cgtWxLaVR5PnIOA5kcxKBzeUbJ6kr2tJ+RQQ9dEDmiO
/4KoMzNkMMOzoiSTue3tVQ1XlaETb5Ja1WdYKj7RbdjgTHF08oWTHyacraWosjdkxekkvQfyP5mJ
LZBJXoy5vs9+rTTYicqN8SBbppS0M50ZtLMM5XPOm5PHyrkQ2pgaJkn+JqcI6QXQW9AFMXQUjJrh
rIAzcr7t+VIUzCWTpbOuy/CaZf+mJp6iN0O0M1TrDXUY9R75JGRuDmCXwzkqcRd0VicQ9+k7Efei
Cd9/n3Xg1+IJy0uEnGvsUXdJsdo1jmBkFS0yzeSHUMFrcXxMmGVpqJo28A8fELyQ0dFro+A4+T28
RAQxvaOyiiCmAIkyctBUrb3ednmtdP2/1aJFhWsndP4lHqNhjYcrcosfUCYLtXPL/J/y3XWyGbWg
s1xEcxD8O0kSsdlBV1ZX0CkAHQHwssWFdMOEr6F0UKcRQirEjtnY1u3wUgFg/KK95rSJzRBBGFsT
i/pMlM1TO+sM6hANoVKvZsCL4ywc6EJpQIyobBGyxQoT7wBLFpj/SY8siq+x7tFMHINM2wGcjFTP
VIzt3OlIm0sPxxH+mM9zvAWXe8TpgIc7wOeXW7NWLulyNabXlx9s2Fcj/GUPnqtnmCcI8fV0lbIH
KXNF7huiJjD/1oITmklpia0HpZKlatJHfEYh2O+VYFEWZtc0Twwh0T96XI6P/bPx7vKkpocT6uj5
AE+Itkhn0vD8SGr2m1Zc9chancCO+vvORVrnC1Hdb/a1cLKKcew4L36oGmeK5ZiDLQ4EKifatC6R
sQdxyTcMEEzmPPgVVnL/cN/qmU4WF1hDJJ4zpBSW4382qCWIpxRNcF6ky+YL2tsWmM1txajMnkyw
cyZejlVl40qdSF6tVISv55O4WCdMVZrdNUKXNrFHgs+GkPxlGY99tkO/s4bwh66F1vOd30eUxdnC
0Z+LkUchAKQhiKWXQiexDWReXsq/+m9vVNe6qnnh5eFboNT0IXoN91hbEIAj5ri0eB4cwo8HsYl1
4s8Dfjud9EafEaWkHhjfZ280QaLz7sWDnCDTNt1LrPEA9WyFQ6jrdwrtuN2rPlPpTN9XX86U97tK
q2xGNOptUEIcy21UcVlO2gN9khgkH9xjE4C7mhNhBrPgk/qqeOtNt9p3pQ7K/JD0PuilYSnvedT4
qDc5IpN2oBabETKPsoci8cRgevMZ1xTra6X46IC1NKRjHdXv+XBaMefBppqnzARVIV8y5mGKUrrg
3ZJTK6ILWRC9n+Oq/ZcC8gh8WySOe6uHkhGMV6w+tOZgesF7VzUDprOM+ogJ16+vLkOqTR2H0p7/
cIAFtuDMgZKpA5zrCkI6700pLK++7DjuintVFr2B5Z/I9/Ml/eg6VwoAJ1yUG5qVJTXfCdqWnD0O
bbXLemfbQ36KCbcvnOUkg6oVeS+o4e5G5QYNBHyziBolb/U+mfsxS79p9V+XfDWFH82P6sq9WU0v
4HmPG2Tri1Co9SvNSO8e6dUmPbV3HB/zgwLtbXt3rUf3YRVC8hfVQ0Fwj+tQ4wTshUOVzfqXHkSq
Ldv0fEG1HRicy8HgC7Uz7zDA0OeRB1lekojjxEU6j8L1ImsjzR9XRpjk9WsYXYAV/xRzu/9xBO4C
t9zLgronKXco6Fq3ISG96iCGvnm9CdMCB3jk40pR+ZsIqZDGY/iqRrFE8Qf3nuuJFOU/Xs92w/Bz
b/dK/4PoqO+hczgMLd8mJLr0vr5x5fDAMxSO4Af5G82Cg86Afk66V4BU15h4S/QVhf/V6ESx4Egh
ZJcrokOwa3n5nfIGY8R3SJzF0EHctfighkg8Q35wOe8cTpVVrGuo+HitlwwKC5qYSrZh/Xw8PyGa
8DY1Pq7XlGLA+wjPi3AXNAhomr2VTb11QxjQYrx0xmvgD4C150LBy44W+mt9T955nif7Edz6fk1O
ZsnaAKihLChxM57oJSwZ/HciIGbm9+7I4tOvc2zgXV1cYnLcJSm5+x37GkKz0OMJy5Og5c+bXgPN
2gmIO44WcfprPgahoHocWXcd9l0LKkx+fubT/OK0V/olpJrj0FrblT+WJz1OdKYVvxPU+Uxg+3Xs
BiISFnRmwvn3t08d9+ggFBxrX+hIsOLbJTJx8ndR+nZXZ2RbUJR7lHa/404mne3L3MOxhiCqlB9t
oRKd2zKenjAdvFZOgZPzE4v359qLVOMZdBdaaiGmNVOaoZQFvY1T3KFzGDZdWW4ZXP1QLA0IwdqF
COeHwWmm/jFg5g/7Uk3OhfaMJGw6h5R1fTslB0GDML0VF75Km/rP5lg1iAeFyKZXtzEniRpYIu3w
ZdbT1dpRIfGyAIdTZzqTZyXpsOvc17CBKhv8Gz22wBmB9mgC26kZS0iO2D2FmUTTcnvSDmN8klVu
tl8LckPCD8BMORpgXVRsi6CZr6BGSF6pFBqnLax6b/K4o/3vsXejF3CD9I1FxC0vOmN8f8r5fDJP
nDk3IZ3HHgNxrtFa4aSVqHNdBlVN1f9ywJutj94I7Zez9jdDh2RV9avg19W6BkyPPz3rQkdtQHZN
g0QeNNZbItxFM53d1p2xXhP4Ci9djpAiwMvFJy6nMCWOxukIiC3JF9gBPMMj0neq8VSZQ/q/7Pa3
L9XL8cydN1NYXWRUqxbFWk1fW27DnwfWhX3SlxJ2AsZWE/aPySGOiEnVgDoOnFFTXyh5fZpg4WNv
eleu3GfwOXdAk8/BPRPL4xYQ9WITG6fTh6JbJPC3vJJFFOWu3CFDiwYYjc4NQlXqmvraXSGWu8iS
0nkAES9fs4U7XB2RELwFTpTcDruFjoxYpXz/ghKPrBAVO+Vukoltfm2DjX005ltTFYflWovRCsTF
1RVWx+24bBuuc9yz1grG4pDxoVQ/DEnmoUT380dUeah7RFK5xA1eAoBLjn6Dn06Px5rTvRYmac0g
CNvOmYQ3I3WT7okgltXeB7WoP5FFV1j0jKnh4z2Txp2D4+sdGMmJJY/0qZu69mCAWDFOMSH1nNJR
t7kyBjvMBKJBTcB5nY17qJp6BmeF+4jq534pujsoURWphCzfmnOyPAaY0ofGNR6uxg/GUfaUegRK
+AQYGgsNCrUUcjef5tXgJScy2/E73FAjSf2OEj2hLcLoXuUznVPiKp6VScjb+N2wLbHnMtHjebCE
fViv5x2MmqM6TZURs4pkMjzbGl8YTrNWep+5fr33QOl6bOR2Jgnzv4aSlginzAtbD5SWn8FpmRGZ
U4hTysHjw+C9cnKm8TJ22VPIi78B+RSvmH9dytHJPqRL8YUsJGypVf/uXESbdW4mFE5A6ooNRnKQ
KIrPeZD0BPpRQIuau+oxqjxd6qceh7KuuwfZDI6Zf9kEK3EzC2bksz/NUUbOmKCTTWW8lUtwXr/2
ED2k1HxUs6SurN328dt0W9UHN/JLmHJOFfQZJqs75QOVr5aS76seh5kqEW4G0KDX3CFaFn5b9Yt9
2DpKhVqEJWjKomQnuxM/ENXB4YRAc5CoLAzFxZMvjPLVNX2qvDGt03Vh//RqWUkoX0veO7a+CmkN
MflEy8dXCoTsHy+b9lmNkp2BPY5P9ZHXAQ97cDYe4a6YmK4azztz7N08Xp3MQ2v4XZqT8zCbcvBE
QVAiQRP6dWGw2Jq1+FzD3BgSbzCoPH9S5FrW8j6IJqvpKfXQptur41gfdlH2ZQllfyad4WT9s/0C
nkBrpfYmYnwgiFSSjDqxzGaVockDnAZ6/u6Vs/zYtruzzBRlmroSnqFY65NwvMstfrcggPvt/WzG
Q6kvc7suPolZd21e8JzNH36Ttcuu9F/sg52qwf8/Iz15rBxRnfEjSdvzW8V0RI5IDTWxpJFayVKu
6hH0CIyEHUoi04Aw7C6dsUaz/Jboyan2+XAY4eI94H4vTaB2gGEDqyyl6S9UCtqFtVusIOjz3zo3
Yqy4pQ7cvBiowXF8g7VL+wK1Wn61/yQVSQfVoVjNBd5OYZeGkRmA1RkCvACYRibD2A5Xekt2/L3U
9BJYJuv1Z618emxgMGJt0fiyeJTQMXKWQJUZI5X+xd4emsxhC/58Wa5210gOSFp3JhYP6P5/x9Yf
a4UPrCuF6ZVeXOYuqlgKhqMskrLbAL0e0gM5jWs69J34rgZBTY2ivIys+Zj0gl4/C22Miw/3O9WF
+6q63nm93WQR47M2rMLuFKEMOpmxhIKzzksvaWzV+X9tu7F5dWKovrW1/UBTpK5W5LzQuc87Tkon
EPtDq+74GXQiuuFh4GB4qcuzvl3V1i5kiJFSZU6uYGB5yWHh1XGJyD4JjptPAibQbBqyIH1SxWzr
1SIlfpNabDFns4ES/brUJtOTlEn7sfAaoghG5A3jWI+aSMxETfHXm6BwV4bcJy8I0W2xdY/phnmv
AJlveqP07LzGHhqfwXbvkW1j3GxomArSqtj2Jbtbl5doTZDN7a/HFYn8q8WsGHyUi0MbgCp4aDdE
iJvWBlsv4r9kuqvLUPfmTc37etjTUBKpMEkAEHwTv3KQL3B+FUUm78hAA62C2esk6Yw8eaAz2scH
oqPGp1opmIVHZbqLOcqo8sen/mD1+y8XN5SBSSOHjrzTLceZ3qQEPadb4loVwbxMdXic7v4ov+m8
7ZYnohcGue8fJrzEOx87noN4qSF4D+FomNrwPb+PUvVd7J59EbO3Xa2PmKn2matXVcapsrea7kla
yuVnAn0UIjY29TyfK+j/3XrSdhCKGI//6eMW/SysuRVP2JBw61ia9Fb5Y0vvVzf88T8yBV0oA4EP
iKGpyBccX4XM2OcdsnG0qh3MC6suR0snKLhZI07yJVFJP27f19HeFjJWoTF34ayahL2YLniLx5ff
18+t0NPhMWO7Q5w9LNlgLxf6JbOfcjaDT0YhacTLNWsD4u2ke3+gBGWVD/m1S3SLg/65kHZYn9CD
04FxBpW9mF6qjtciqGDKqCb8L0N3I0X0pL8SomnG3ScFXHlrWm5XrozKvADW7xlpCcPxIwtufti9
TSoeS+bacufynghhGl4eq4gueA9xI2/HCtnc7hGurEphbyvdrhMqOMpcP4MaXtbBPDR8C9E5xkEA
brkSBSawtQY3NJBDH9vIU4fAfmntuiJ0wunqfF8r7h0JcTE9RU7nKydQawdCqics/9LC3i3BDtwm
R9hHaWpSh+spLrDWsJrR7eTsvGKtFNfSGndwl51gsth38bS6tzHcqzDXq/3jXLJxVTmZnGB8wSAg
GqgWD71Gjx+tWFFTrRuCZ7gYdycM3cVlfu44otl9DBR1s5YWzgvRByPmVJD2vJ/Wu+befuLsrsKM
w4y6pnIJtcCqsamSCVAR1i7fNrzPFBEAgOr6fS4ZgoPAcXuN63kSpzneHalPZkN+Qua+p/kD/PEH
AAEAcwEv/il5v+DPagYZIGCC5G8qHKaUhZe0EO7iFfBI8904LZb5OjVOUF5KanKYw4V3xOZ/oNvD
1SEA02Xfg6vy+RTLKSPn7k1AQTqmTJK86RAYLxV/qEtB5MqIq7hon+lR7AjLRSrlttcO2pmcSpU0
rpbSwhqcgPuEefopBC7vbFLtW8RxMgB653Z+WJ2cfelJicT52IpwCgi6A8uWyQUv6VpGU9YbNkst
BFwLsgtWmCDU9aHJe3r+2REqz3shx3OGZBHDXRAsrgHo8fpST2qLeA7VrMOrlymiqwm21pk6v0SE
lbwiSMV42lXexOzSmFCRshqxkbhSAkITKayQJUTmlXTZevAegOlTgPM8lsO//BfJ6TnAufvFJYF8
Xbs7owt2vN0It/Jy9zkcNRVIFlUSNBVpJR0EU6BGVF5aQiaAt014tS6mHTmKGtqUvEN+DOr2ynrA
nT1Wine5qF90d5u8IOA1m0m1pNdZP5B58ukgPEsUTDyFxICaqYHE9sSaaaxfjF5Hcqw6J2TZo+LT
lYxFZpeprj+zwlpUPFbsPWERpbeeQ44hRFPCGqwoHvoGrr7c6SdI4GiKaqyOVQnRdRxoYDBGaQJi
KNK7jOpKZbRUS2huQOpkvx2Bzc014jvDgkEtyGHbZRh/Zj7wZTSSiak9i44SIBMBSrAXWhAhsIXI
2TiCO0OHADnAoAmoljX6IoNnBjYbhQDiJv6QZt92M/w2nIuTGW4udZidpAhC2zV/ZWoBzkD2gLVn
24RE1AUNneWE8c8k3HACNPzjVQauqoXAJPH//pfIkxfS2ajDH3Fd1np8b1z8ppyb+bUgUjM0dohD
YesHuJzmudA1/FTLRBojfQAArbIUzJ8LGgSJwaImkE02teB5ttGZlPGXVZa5R2z0BYOqsBVhZOUH
eZqKQ8xatb8bEOQWxHzpV34qfr5Gf7/AT5kpmb2B0/wSvvuXSRbg/yvrnCxPx+MgEmJ8v/a7HXYz
wM/nTHafElb4TmK1qRCNZPOkQ2g/GOpmtmQbsOsPziqS88QnLTqJX9BNV97xScT4kf36oJR8CCTd
7Lp8OP5K3m572TRq4lbfnEslEsh2dYiMVWIYmYuquNFbR79jjq8lsZLCS3iYrXDicmw0ySJKBJN4
3JvS6H4MHAD26PRNKhQvdo6GahdRHYXtfu3rfHRQvKFxeEa+y/0jzhDX79RBivJChpXQHf9TBYzO
M+sv99dmoprJ4vv/FYwVzdVHU/Qw5zuQ+twXW0n+Vb+wqrvV6r7CpJ70ilkM/Q/31XbbOHP3JtRR
8okVOtR5WKxnPNzEfnJR13K5P6AFcDG7Oq0DAjwz+E5G66YcFNlMcEiJ6OKC0KEbttxhRmDLK84j
9URgC6BsHzUaBTKrQQvGolCh8iX1bcQcFo2Y6Igr7ndft5T2nBWQ53IEyA9CiVs0EcfkbpS3R7s8
oWnJrzDhkpZdtVyfmo8AQQroePTopODHutbH8usVhnTz9Xh8R9appDWYKsQpJlOifSlM9g5KfuwG
HzlVzOMgN0tsBCpZQz0dbO+ngnt9ljsyIJoSSVg/8N27EOO3T3cY0AKG5slMAYY3NCrDgrdt0zeD
rIHNzbHWNLp0OTEFgJSYpl6KEAG3syRgE7gsMhvY6E1tXm0EWpSpcax9yDf3IldVVgXhL7V0CB06
vVfT+kjA6kSZYjbbfDROLZs/ibWjyI0WVS7rw4tmhGE270j8apLPiqmH6h1mwZ0oRsXf+E1bizuf
n47hO5AG97tLQVuWTSyV7ECVhIr1V9fVLIfeajlKjgeyuvQviVFtSb54PX1r7rhr9UutXKlYDX6V
wGziETW0egivw8LYJtdwIyxKXTbL7yDpnoopXkIW3rhFc6SRbNciuQvQagEAVovfG3vx71tjzw6O
6XyHJ5ZfGMmEGS3Tp3LycNvkUfEEx/O5B/fzLoHVJMSvXkeaTJoXOhskbbLNR9RQGkPuToF9Bc2h
YsAQUPbJqfoRKVGyxHx2GwyDvET6WkX+68SrFWInXg56JDIWD+ayiUaAF8yLwQc0uMbjYbcuKDLS
z1Uo+0mqxpdlFEv89gP1mORBzamn+tq8Wj1jcblwA4W+8WedRFQxpFgGfAeNd51oiirxf1iElKFT
Mfwg9vIeMR48MiCipUREix6QSI97f06M4ReptVheP5kl0z4zCPnxxdy5krgohgxt5Q7n5EzEgrjl
WBCZXnMsfZhAPzu3A6MQDOd3f+lGDYg7IfD8Dpsg6zxe2JNdmlcY3fWHvFCNeXaH+nrbr20P5vpB
zMkn9XSwAmT+WctjNVLLB67L8UFj0LcHgfxO0ya5aJHbE8JGMvE8kSZqQLPAm9yJ5siBv3YAwkxE
i1Lgr2zaqb0L130JR739XMC9PJhl6c4o9lWXGziUg7l8Pxe2ofaL/QTWQ9WP3RSbKgZx4oSqdSzi
5bJsiw8nCEmLu2bW4wTJSQSHqod71dE/74NnDqT0a+lNQncNRmvLlU82Exy9lMtp/5buj86m4CH3
7Gnybg8vPMy86aSGPvrrZBL9GB8EcrwO9tgfg6v5pjEioHCt27zjT+wJVjyiQKLbeOW605CnAMpL
pBabxTxC+0cze2GwWJ4rsIwZe27vuVFXPKXm/SDWO/Bm6AvOxN8M61FUnMSA6Z7XyEuhit7YbtKO
VnYdMPZJ8137qbO/7Izd9BValmT8QqoMHgopOYNVlFdG9xoJZex2txpQZHJU+bUjeDa6CtRDaCAi
lnGyCsLRcat+4xX0tI+c7xkQROk+czXIf4JyTfFJdGxcHOJeiqQIvBXTXE+s5mtv81YPqUJ6HzzV
gidnoTH8WMETm6ORaBBohz51QwDyH8C283xNOeqd4u1oAzcC4dAIG6sMDhs6cYw6TxHkIE33zmjN
XsNp/HPaOYf6WA6l5TM4ivDL2Fo5oKQ4fOud3Dwg4V3/QllPK3VevFCPSufmPJvL/eoW42t2mkJk
A08LJqjfJMkCKc1sGWyyPwUIZS3KL/kbl0lH2Y8JlMSennx8mfMUsH71/A2O5Kvua0J9UgW8jMk5
OYaHwECdXCN9DwApHv80ynBWmna5qNFFntwBwws72HQTKR2Zk/1nZyY/ffWm2+jxqtshe83VJ349
f9O20fgPe4lcqeteKKrK2Yl3hQwG8c4eJ3lHyBfK+yN+2uPDZBqGY91Fhse7WxXEwJBdrddy+/kG
DSA+kNJpw6Af0XToO6aaZGVq/bBZp65kP9xF2EEZm0goCDFFprur5+YD/8oZeb36YJp3dTn6B8Th
+G2YwI/JpkKmEQm/aym1b1fkwm60VGRlS6m4GryBAxbYxZOUkhSuiZgm2bDy0NEnxUJMTOLIhRa6
MdMwcoGCz+eELkEWocjuTUJYCN4IMngaTkmspf2QiohKPygGCCUegX2ShfcmyBhM7IAfaasuxtOo
priCWo1ESBlDt//1RWKp5QCuOzg5y8TQVAkooUjFEkDErN+tBnbVPUi8FJngZptQN0c0MivcHu3b
Uvnzkc0o9vrGP+0/LAbyEwNN0LSgn6GXw/RoCgcdls2Ij566nK2L+f9jUrAJrW9/J9VcUPdeExOi
9w5nnbeSoA9gDv4W5x/Etsw0Nix1QAJUCtkODK9mi1V32OzcUqF81dlbn/QOrH4VT02SpLhoINyA
9jT4iec384Ono7gZIZd5gWuVOKSFoOlGsU4m488w+nCPiW/ge654d/Y1Jw3wjsukbWn7qxf4wPys
dvIJqx2olo7d5Lj+tRBGv1YWReGvAI0WEH9IBw3UQDzfpYE0vixG4Wf3c6b33eesXapsYcZwLCYU
LMNy32FnTnDvOq7vpJII+dRjvDSYHuNpHfiJjlgKsnArqY6kN/ur16k5pN8Txgd3iSapJufg2Eu/
dd3Szn2EqKXoI/Dvuh3l6Q+1w7v8+08+68OVD1cSyCAG3UQcBxAfDmESjWfMOng89FCKQFU4vdj8
B2wIS5TwOUl3y635ExvjhmPgiCUdMzjqlfuNzi7pmp0tbz/ea6uBc1eBzwW6TOkWch/C3qRfgpBE
Uqo8Ta9fHevXwwzIPdJcIVkunI4xAoqaHRgRpYS4oB9X2ojFqAl7/Rk14vp+pnJX615n5tOCp3Wm
puBHlMBswJ89+wm2HzvO9cESi8X0TyHRRgtJTRljH1ST8KAdZMeEyxt/xTxW79dvpPLfrMW33B9+
5B2zp4gnRcwJKg4Jh/i9mbcQx4+RW+iq2uS9BvrqddndI9mfRCPyY8DMkrCYemCHM8VXodhE97XF
jZRYb9lgG2yFd99ZNQTOmyNaAi9xFDrbo6+tMJhZkrmcMZY7INM1m53VzUKeRxUZhMEZN5syHz7o
TkMYG2h5EeBpkec9BglxGBKpjyOt+1BBpc3HDSMNx5/quw3iqsp8Cq8TlK6NYhUT7iOcYrYIGfiy
jvTu8/mJwmUs0tDG8N47+wdq56RBtDpGEaVvjDCogZ0sj9DSWnhM68TOK7gJIeqy/zXMjmrRfCL+
WzL2foqzOT1zOdb4Y+aWuPi/9yPVKcoexSkcYSWXa1mq6qw72AG1JleRAwEdaAj6zvmNauAqOvmS
jAx8eeHXXNV0FAjYWnwOUGRlQd4iamd1mdoYN1N6+BGNySX9fm3DVNbSJ29HyfN+if7zABiw5lhG
/EMVrh406h3GMYKS/fUSE17dlT2U0NeoLRIu8emrZQLzTuKXNptVGOT4wvYDjpt9zvteDgR/ESOA
kAnaKdxjGSP3oZdZImX/IIxSpTBFCCOH6M3we40YqyMiL1sXRy+tqkEQCEItiXvz5fNiqvZOsQSb
tWFPR9beM84EOVgKvhl5XITzVZ93yKfusGw7IXslYTirC+7gqNScLPMYFCOaCyWLvs0t8al0T6ku
VZt481iShTWJ/BL5KIXgEPG75fjNljWnTDQ4M0MCXVAhgHlfx8IDxUFVditvVzoK+DX5SEm9u/H1
uZmrSnpof4qVqrwxBLMWHfIxRTTgoYPZFUCG2dYTTJaB5HOJ3zjlqQEEfzNVe6IHq4MCGEuG+DuE
E7zX2hb6FPvdXdLP7rU6THNdChhkAxNkNAjxHjtiFwCBDLptvqdYgB5YmGKR4j561AkB/x+PpeWB
o6AhHi3z9YcBiClcU+bJNbGPsF2xV+oZPgak/S4SFKlOix3f4YPcmZk7/jIgr6pbGfq1kbpsz+YW
99elPdhC9LzsMetNj+fWaPCsbpZJTHo4WZoGq6bjgnuaOCod5/xdQLQ2f64zqigOrPjxsmcia0i2
EPaWnVECxRM6UikWuLUAhGpT4JmdZTxhiyw+T1VgJkAqpt6yTODDdwvF3vVcTjx5xlX5mRSSNm05
3lKGqGTHTglNpIAS8EvWylJ9EkS/1teOGoGmkjnjo2XoSUYGGJfWp11Aljc84nDQsfz/59244fio
zZe917wF1t3HqpdominKnY7p6ByznWW9GIkf+Xe6HezTTzB5z35wztAGhSb2QAATwqiKSNs5JM6N
2eclg9M4n33zpNcTLRRKZUDs+LCLVH5U2IE/vZJ6C5IOx9dhnSXAOOp2dW0ouqWDuAP705UGWXax
W6H1nNnF7ODBlGzrG124IpC7ATTTIzkU4AdccfhV6Oq2+dCgtBvGSlmoU47iUDz0v6byytC+vGlE
1dEZi3a5nnM8kxo3EPxO+mYki+R/mbCCiiKwmID/UH17r/xYaptqUIFPIHDEPMQh7tIQNMR33cyu
iKQ/maf/qFHMtv/3DvMdFa24+rbk5kQsof72dyjejRaNLI3rX4DHank4BJCkWFibjE0dXhicaazh
zwfkmVbc9uVbO2+4hlKbPtFXfeQhyeYIk+Ht6i7wFP5X73IuZWY9C9lyBcG8IvuhQPa72xqr5AWK
OK4mglEh4HsfiKWvLXh0zywy9+ddWq0492cT4ie7DZ251I720kPy60TZ2d4cgIIOGn42bFrbIFee
31J6pmNUurhDyNPzPZWXcLru6NSCOUrkzBPiSkg8ZKhWm791WRFaoEqh/a5fgHhvZvt4G2dUwBgB
KjHK+ronGMnKytCcBCK6/vDouxWXbHclGiW9hFBHnpxLiObAfUbmX4ci0vhKtgEIlls6Xh5sVE1T
VtvdReBJffOxRkgsl2LkxDyF02o3OX260l5JZc2DBzW24iorP3iDbxtA2zznXkxgGPmHsDLNsV4t
LSlSLPzdiLjqrhaBtuQ/wRDMF2oCFnWmrQRQQRnaWoBi7TEpxKgKAl+q5HzzIa+TR7XClwimrboS
InuFeYy9RImP6I2rWZPubfTIk7GbfODhy4B09l8zOXvETgza5whqANpHGr7QWQGQMnsIW0z/zi+y
WbKuwjn0aycJGDT1hV0UsnaErsoqStfAX+J0Jks8ruLLATGOjC26ltcIolchiCXnauj3wNanGkP7
GLU1I0l6lkBNVz73ctKxZFGYqetPg6/AwbDwUu7jNM8e9wEoVHjyx4e3vQoxXMR9zvixgwhSjHxL
SjgrgaE/EJGxpklpPdrtD6G2rgFWnkuJ7mLqloN4TNbFN996hba9JvoiBXMk8OnCeAFSxIEceT2b
WLExTPmTNxd4fr0aLsIIQY5piS4gYYARUnCnB+y/BZwtXWqrvFtGiwC+EQx/tQpmwMUtqRBfwiOv
D6VcBcCcaXclWDYPXa5+MKKY+C+14K9Qz4wueeFrU3p/uwHmyc15x80yQL+KoPB5QrEof1bpgSrJ
e5sJQ2G0Y3RhvQTR+zsE36GXTaMguPHhYqYiZCAwR4z3jx/TmDVnRSf0Q3nkq8Eg+ICNEM0BcuIt
HCFRSZgo7t3PgL2qtQhcAXcYCaQ/WS+8DWhJkMwGYIG4dV89RwU/aqV9uZzeecOKXbQyWH+uSMcg
X+4UaU5H2ye74CJ2wYBtcqFCJGd5Eo88zKdPTvWMtvUWn1moVaWqveK/ZBr91NI5UZkb5zpe9BBJ
5OmzAsBq5cFA8WeVSFPdFjUNPL4g4886MjtNyB6HYXqLzc0ztBjzzYirXhskMtWB/F2N/n5vx+o4
1puAfttkf6asG9MRlmsVLkwhou2gI25ui55kQXA0xrs6yf/yoBKd+5Rj4OvxHWGMZH0DciB/twiF
/lpGpcPqJGZvtPdvpYczKZQ6L4ddYPXfcHE+7N/2+scobssAHLirdFu1T3k+179aEFioUQqelt4W
z0rgwV5UyQ+5tDreTvipjsdXw20+0laM0Xsg5U29zIEfTOtYWTEC/03cq2TUeLhAV4Ce9fL9qK19
HGtlkMHHzteqMiZ2w099onXh5anyn61+IsSqdxSqWygjuE9FCyVdEqg06qRDN/ysGridb3e1H9lA
ThFxLJKBCRjKHPHrHL9N1j9OTQiULO21NL+PSMc62Rv8ZXc0E1UeX0WM7Yl41KSJycWmfglnX+YK
MH0z6mNWUSTmHKJgBRgC7U/DeW/oaLIXeJiauj3sclyAEssXj81TSyrMvkFI9IhaZBlIpg1r7l3m
moXHzKvp4uIHNpitKbvLU5uTW0eB13dfBXwE8w4EFzcmp57gEjD72CSEUML4eUSwnzTvuAY/DGOe
RMHP/gVsxmff6o1BAFr18kgzIGhG0v+Jp9x8ObSkgRkHLqTpa75opmUIIJtwNcP0OMhk812EPOdo
gyMvwG+U7rh7IU96PYVQGfjZk1G+u/0GeYz7rajPowUGTZT42NJLV6LnOdGMGnlRFyOGIs5j5FVq
XUvyq2AI0SEZ0DDzloSIFTA8op9LZFzZT7Fyos6zqcudRhZEagR0xr4jjzS61uGLI2v1zbU4eNyy
DG3Bb2004goT3qurjnpikf5TUDVMX4xIINxVtvA0Rd1vM7OVXV9JpzbetAzfKwRxg6027xPgqizd
C44KfFbsYofJQ8zqcNGe1AL3bNgH9SVypiC8/5Iju5djYG5KrDskMq1qhrS1/WDNdOtTzbVrYLeZ
vyQIksLmZdER7/d6Hf78MGGShXL0ssoaTcwe62y3E5LsIedVbejQwf1Wzm3lUHK/Wg2EBMI5JuGY
6ir43LW9tRN4DvgMXrmwz8AzkNss7MACErcdUL+2P7Hqrmq1PpF6n61iMr1O23SWvl5Qb8zI9+WO
Fg+RrWTzRGzru5kDDapF/p/3bZUZf1enr9ZtX1WX/BJb9/2fCz8/8iZ4lVyxiVMQUvt3pAI6SOuo
4jU4C3wKmGblksVzBhBNrjroF3AG8g1Gj5mA3r3kqxn0i5DWHG1W6+ozlEOQmRSxrRwVx7lJDLOj
gtONIUOza8dZRSsnfSDnpMe9o11pB2zfUkFasuuGkR9fHefwZNN5ZIlfE08BTmcCzuQLulhJhr2T
3HSQT8CaOMdBxkO8OTTNtFhhhFjgdzElPHhupvyp4HcQDC347/ax6RqsvO9MDLH6/Ku6I8hdHd/V
C2yrQYOiendcSHN8VAbn+YaTuc3LFhQnwDu/2IZuLlS4QHIPPA9xLipDCytZDnmprWoR8wiROPjh
jIGIOaicYCJnVS/EOfbHjyQSy9Hix2oMgJT3lXYCGWoiVdNKqD47G9+iDmVTRHTz87TgGKvAzEVA
8imwajX5D9VdkcZdBIcdCqu1AlcTlPKzevcuJV7wq3H107KjEHjjgG8WZCTDDaXv7Emky6A03c5H
R8NGxAO0OBSzIeoKrKanuOri3PDhhMY9e6yUeU4rMR2b08SY9PXcOp7j/swit+LdGcUO+9r34aFb
+IZjvaMTBfa8CX079wk18Nln2bcdR4AtkEKVnMK2NseJEoZ8nddhJuOSS3+f4vj/PB+e0RmJckqD
wjNNY4xL3RVikFzJqOTn3wVGuu33MgWBYs+HjoaRrI81ugBKzeHVkAScBGliKM8dC8eoH8ag9qD9
lDip0tu+L1jDTbNc/ORmZemyyYbbN4GsUES+7Mym7an5SWlW6ZB+d+PphU1LtR7iACQhjTjKTdo1
IeL+em/vIWNGlY3tyZXa2PfXYl8H1xJfo8xSEIQaT+XXByFmhQhKHXg3IME0ZBh80dszLphQs+1F
1Abr5yGOekmktHN1lBusM9dLTntuIz69/4UX/j3NoIK7tvEpDE7cLtO0cMJ8/siK5oFykPSm6prF
KEuEcZR1/v9hJ4AJgIZ10FrrRBTd0H5oywyW9guI9q5Ghey2ewUhtagP/7nh4Y9ynNgPKO0U/Ij0
LoLfT9WQAyGRWF8T1GiB0s5VZe3yCr7/+YhkBIiuQL85pHk/wIjRuxfy4OxzPGxIorb+1jy/rHdV
FjLpRAnO9+D1+hP69W+Y4HINupNaQh2xZQPOWftcMIIBdt+aAuU8XIQPr3+fz2LyvNCqnPL533KC
rAAGyrItVeVxOCFHEOvQ+M+I8j/6ueITE60SfbUKr/lSKxpyDefi9udyx2lv7GFruQXE0tYFoWYx
sDV0JrpfdB+wJFsNalQ9X/TDfzBYfduTAN/YqNmd94eKNPH6RPZ5wFsFbghYyroG9JJ9w+2LgUyO
/Lb53bWZIUUDBE8DJRAylva5a3g1f6pxgj6TOqW+N7IMDqpsrDvIzvoZJwnae9sXWPfvtvqDwvDl
RziHv/fIitIbHLWL7YjwCBCIxob8q6OLRJYBks9mo1mgKQZgd9MdeVPv00RJnbHRgQr3cc1Jprre
awkvTNG1WlxKBYSfybUjjkyStspGgGEFsbsHiriG+b8vZSNH7PSwnNpE6Ildf7d/OmzCq4vMyXe0
/ClxYqy3NeggjDTkEQr0zI17iDloUVSvpz0WmXe1lL7wFl+9pF81otRAX1SX4mnyAaa0O3Um6mtn
m2fZz/8NVc+8NT/wsvwMWvuYfQSvwi1yFFekCFGJdqCYEyY1oEtu9oIvuT41eeuaU4u1haqdWUBc
VFsIz4GCbAmks3ncJzvaju1pdk7zyFFvYpyDAakGCDWDmIby8lmk8RXFUsensIcPquu+ci8D/oC4
E/Drw6UNhQ2VGuiZ9gmNQ/mPGDUexy9gXZQil5wVqEeqyAtRDeIAs7RtJFdwCd2TjNZ2zxH9Kaoc
uCYLG4lwS8qM25kQlK1wstZpvvizDkQ7K85/PK6YF7tPc6jW0fQcb0NGkMXBoYK/dbjcmAJ7tDxe
wxgyak2bqrGmn8TXGaXMlVdx7bZBbWkH2zqQm1QqeM9A/eHMG7I2RClsIvlJ5yCjXbB/zHHQAmAe
OD3KkLo5nLelXSFnN4/7/xOuMrtzEw9h31TKvMZiuOQryVsuP9nNzyRxhl3Qna40mZm8uDb2nZvm
l+pAhX+tdVXEOY2uTwZPPwkOXley9Eh+DMJ7nwjZYu16qYMHhqhO4ENiK4ugis1GQN1+++6VsgkW
ZvZtB3tRvxppUM7NEowrEDGyJkNB1dIvtgh9l0QtUNpo15PNU1zYKGEA6zHqXA6/5Rve8XCRZ47o
YuatKwbKvjAuE5euVUKYeWLs0Xp79b6Ff392SI1vK/KeXDqIJxT4HBQ4+2wS8johGY8HYl9ydc39
ACr9LTnQyrPO55MqsCC0beX/4UyuI52YEF1Fe7jekkt4EMrLLu0o1lcftiwliLy6Bx5J6i4I/Vsv
7pVUFYGoDFqPH6kXrAvQRXWLtMFjdNObqNCuEgmHELI9dORfALyquBz432oMgAOnEe4fhvo8psnj
MxHUTUA1IWF5O9Uyw/UEDOyhyGlDCIR52naPyeUoI+OD/RI8nnZqw5YtBYTEBdGFSP4ndi4K5ZhS
W/YE2GEZiAvBkCkcLw8p+5o1ab4749P31e5/Whe0agQVoYGNkLw21mPo4EVYCtWYncXF5OeCDqRX
hA5PHjbO1yPPDsYZ1AIaY0E0Tfqe+ws8vkzimUQwhEo26vn4uPrzzgFjXpTyXiWbZrqYwq6fatvk
03f+nF35m4+zk/B1Tvj7E1+4eLT0ebEBXu6JO+3lZYVP06a187GdvjClFjCcRfXl4hTjtSBXm147
sJDMkpFvK4oIzOidMtpQR+g4L0cLCiE6WkGrbibH+05yWUpyaYFVbZZvnTOVQhygxvbMeQBa8nAT
jHbCyj9XGdw4Y8FjhJ2xi9SN/V8Jcxl/qmMRnx+nCfgCGTEz0wp122AJs/lkSPHR1leqZijRJRHw
tzVimyqjkahi8jRLUum0/nxexsFZ0OXAgnmDrbsweROBOsavQ5c9KEcylA/MNgDEv7+ZYbzBI5v5
pRr8t4j1Krz5Y4ZNvFAuYxMjMPxV7725cvI3oXebIGBKr5m8yCEqYQYCQJZI+JXRg/+ZI/vWPYSl
pY6Q3nM4Zi/xLVhsjI2eXEyU4CXyB0pUJyqgtYyzmV02+qAdx3fGDXzXlmeWVJ0EnQUvhRJlZIza
zDJ17kWa7YpD9vTamLqDhC8tfAkT06RG3DqgkVPozsKx6nL5/DbES4Y/MqvmqOFuqogevygq7huG
oqOrhAfdu6IXNi1sz6CnhRCA2McBfSOyRPP2jK6TtYVxSZ22fROFuKpMd8AJ4IBx0R9ALyVuSElm
Y1DlRkzpNdOWpuCXD/xSRCbS7WX+STCMVovpWApRDpbNEqRXcFBsxhCj3Bsy/xyVcBc2eXobEy6+
vEuKAamFQ4Qolcj7IMBbtoAR8zHXNdaRG9N2+KuA+jOAqiFdJRoZdctom4alJeGWj6WbcOd71FwK
diOC3vk1KP+pLZM1jD0f/Qi4LK1vQsfTlzkCqmsgYwXFc8Dl81PB6o8PLJ/DkiqVOWBsG6PCg/+R
+vOGQTQinuU7GOlsxtb9zHQwDT5zGkWr4kFx907gAXpYQBK8OBVKYaHqr5j+DvzAcfwJomJjwTqt
nVYI28O5hZ5hgPlP0d3m4NEojIZ/Vkex55UrcKB7UD3CboYYufmPhfi7abU0Zov92RUyWjTitf3q
WI2KjZRrRAvgWAhVOPqs27zXEASNs+oPCMz0TThvgTPsvlTttxePXhg5OEfArmL0fIkS+mNU8i9Y
MsNZlsdoJVTiR1f1ofzWeUb1kmXMmFitbONIZPy2zyHEhLiXCVpAmmsOzmVNuvBqlH7HjC/BtkZJ
bClhAb1zj2tf65pJKOmOLYEMNbhy7nj4tOlUWgSZGa9Udgp6JnH73m0dKsP3UecTUe+eebEAQ9f9
JcSGP3IHCgnVCvbHE4qlS15rC9IbXjQdTSLr0iu7gL5kPNJfkvxqeRfNSSOFP2ByR0nKpF3Xus+E
FiJzEZw9j66eQda44OzOPqtii2QPYTq5pBqllDJ612iHe1jz+V++uRWCLdqRYPTipQ0EwO7SthJe
ReKBcDHceuQ9wiRFAAkPYruUpVcv0bgOcehDTmG+5l+IHj9RrTW7wjmq+WlZzVBis++hWIvYWsFC
1Z9Fi49NXMaXcS2eRFbpBFUbGEyrhIAejO5WL4NTachGoIWwN8ruZLST1IdE/VJ7i4e0wYH1TuYq
NdjnQdgBzi5wQqAAXw5cejVLcfNn0L36woT9jl/Bi55aVnX413RHL8y4AJbVEPW5nrf/JQz6YRSz
mZyfEKMspeMd55xFdHOR/foP1bVzANA/TcgDuG4JloZwDU+q7FwD8tRU1fXUaz7nE6UmQPtVndDR
3cBOgJJjTobPSAiFb8SODHhVwUNmnjm+wtWRUi54pmt4VNHbeyTOEXW8FZRURrw3nTwCOI1waC42
WSpEp60iUGY4ZtzjZIehgQd4Rstv/K79C4Zii8vjVl0kKLRyt+4MuabMTAVyMlJysdy997NY+C37
QzgihmveTZbLX98lhCntlpvRFc7Re+64l+3R3m7BN/4Cdw38BbU1Jy2YFtREpFzdH5acxAWcZVv1
Y1c7IUBeUi8I78G+mMtyIQyY913M/JepPZRg5MiWHhJuZ+GGui0jmwNfggZP6tfOGqu1nelg6f9g
Z1zRUYsp8vgj0HvvHkQKpiPW8cfs3pZPrUrRPnaq+Smb43dz/cc6E0WsPYCzVst2sM0OeFAcM2zk
DiNtYVQuWahuVd6JsgMD94oTjoJZh3/N2eesLHakE/xgDaH+/cjeS1vFQDXyznBYjMC8/lqh7S9F
/5aA86xeC+kJHrfU1Lk57UrFULPrh4ggQA8Y5oYN/lu2sySgW6JzEDZNBbojEKdJjNxDzE5PSJlM
AxZyhWfy2nQcTwaHTvB5XpTKKPrilkKqwObZ+Tn2hP4BAuHKeniUQKKrd14LC+4B6VaNH8Vq5HRK
/38cLosi9UII83G+zWpnIKb4Kuj0Mor8ViJALUy+WrMXV3Nc8F4gBKa4E6qc0rtJgaZ3V7INV6rQ
8gKWx2/daVpfpcEQD0T7pzwDdHB+XbnfJxsq3rPNzzvki/oRGrwWZFPFWqxxYS7GenJfaKJSK/aI
1YuNRoEah/VlMvC3YRLtLAecUm7fFkj2Bb9HfJrUPCGh9gMW1a6gqWTBC46rTyWI0+3aOskGtWqm
2ftk/o5+h0Z9fhuKTDeKZeCdjgcSBFMyisL/+cl1QMHLdkDp1I+eDUxNwcQj/OiQ1y9xlXgWDpvC
rkYYTQJJVo/wkqCeJMd4TaFBwkHuCB52BhunYThFQEtd4sFSWJG5F+nadANuNGffvS7MyV7V4Abu
rLJUhp///ezNPvf8wDT4cArK3GGyFMyHSgU75hyVZ6WIaAqQQB/d1rGJGi0+C/9vGyV7PAVM2hrz
cdSguiEcWWvVi8sngs/7YgqiRPIlzLHzUSqrHi2pHS/9OYe6TPOKr/QraBvINEqA2efDLdK52/0U
hfAhqNnbabQjFQ4yxfnRVPLDM0+z6mYIRLqqMGEu/iEr5Z0OZtcNTbXIyjUZ9m9WLQS/oEiC1lpP
vK+/TRzNfeehJ0DH10unv3mGNOgBGGzNgtiur6uxsOcnyr11hbOpdpTkFBbn1b9TfLcmQOZTv0qh
1vfc584u0v6p9w/QQlNjFxekiuDvEVtVe8es9qcXT5XQCrBdwV9lvXjYFvFPoKH5ps3LSi+m+sID
ueHy7PcfBa1Oq9rnLbt2zz6cuwEmWQQVjycgkV84ccTvL/jx4Ex79v0XT7RniqL6WhtnTUalYRvo
sYMOt86YAd43nfKQZobvDRVu94WQW0SSjOXH/Mslm0gC/mJ3jxNVgt/X3OhxjXcEaLP60D6vxM5+
GjEIBaRUXHlRHjpDmMNAioa6dSy/zQL4GbOrp3pT+amSP5Bd+9laghyhImA2a0EQtYmTadT2w0I2
MBJKrt3GRMi7uxtJjYTr22Gf2338eXSKoXPCEv42jCArt+wf7iBd7YYVzWvtgZRyl1dnAVYaupXy
YAzX2rzchN4y9QdjukvHqJyyHTaa2mqO9udgC6CcXgbAzELK5kmRMZVAObw1Xh4b+JaV8hO6Au1O
ceTL6Fc1YBQIHela+8SAGWDToOMaKnLzg3fCB3l3yFNgmV2UBPFJm2r6urlkIMHNQWTJEO8qJodO
96VZ9qxQ6O4GRo+mw7rLRwmQhgC5Em/FNSCFOByJQp29WdVuyhOonOm8NMQnqYQDZ3Z3nY16e9A7
qIUGNL52FjxSia9zCYehc2VnVRAfz/9OD3ue3SzixmKT8gj0d0/Ityt2+zqj0bacz8/Kn46JvN2u
3Xg/0Zf7ArzhxxnFSdTVAcJLSbIcnEEwYkJD9FnIGCsB4FgGnz4rvaqesg93/N52zV02AH63Ydt8
Un2Dt6pdz8AuoBiB1C5FMwo5YFa+dPoiqKw+OafgL0zTrKYtF6PH/0bYb5mKhLlu3T2/VLsrO4hE
I3sYNrEFsySh32vHi3AArkPgbNcqFK/yaW5F25TMG2dVTjqlu0IZLpuGq+MCfeBW7v9J+zG0aoQm
yys4vRl/afpvDfwN6OlybrD80IYsLAEhomiADqBAD/yv4wQQ6MFTc1LoeXMbOmUwOrjSeOoohIBp
OcSOTOWHZsskHmMXEGTOjAuqxk3aHwDTbJHYf8bdllvPQTMoVYJO+7Xp6P8cbBa+XiODT/n5rUv7
fKcAIgxQrpCq9enJspAT+BT9JU3wMu45/ocdMYmIyM6mKHySFwN8agMI88wDeBTdDF/8hyHWO5yU
lREv7P2c78gk+n+o2PqBX4x12RGhZBmf1x7UT80KFbat6F3kR+lnjLsRg95/pIrHy84bXqsn4Xr9
bPkGYmd4Mr09wnGasvyLCEl/gvHxkXWBqU2DmDVTxkGWTQl+O3opiX4zUlJM7r0Zap2mfsh8R390
h7hkzatzTVs97iyuPX60blzpRhJXNsuzMOqyuGxIi7QJoh7R/FmtiXnNl2Xce2xK+FwS98UIqmE6
Kbvbg/Tzivtr8SZLhq+Vg8JeQTvPLBxi4FWha9+YpckfRnyVUJebzgVv0GjlIspY8rz0iNgMua7V
+8RCp+AK9SgHFLw4r//bNcUVSJm37g0BaPtyGWOlOD6gMqFtQhdj5vOCXGReikcj52j8KSwAglqp
9fXlXsqKyYafXlGnozp8xMOprKH3P7dtbQu0r+2WHDrTQa1HoktoJy4caUWYOI5N0c4ngUflR3dR
8R9qjebojKQH7a6Pf2rSXyrh5XUx+a864vLl4H+5G76u/UJSZ8ZudRs2otzEaLRa2qbVcDOpHT91
ItWj+97yZYyWhfSMdszjgrGpn5U/fXr3u7Fnm2mMwUlBGF5kP0w5pss1BXaYtTAO7JCB8etc2/dH
frFoYc9CCLvo+oGK6bMDx84n7djPKr5fK7YSuTsYolnIQL9DpvQNv+tsjAxsvQEzN8qptzOoDyPV
aJC7ebviAs835LaZNE1BmKFtEPt0CxSzKWL8Z1U2ePRyxE6cvXst8T1fw4IqvX3iFSKiQQWzifvo
88mlPPEsrM0BS5397OvYdf6v/pZlj7LdPnR6v4fg5NGQiKVoixCoRsxyPCEysZieQdJu0A7jtQPV
fq8tX+I6jpFLL1UcLk/c/rbENIhbOdTvLe81KvvQ8NOyzoNq/L5N9bHyU2rWxGT4CFU66aNzEIUP
bcxgZLhjSrj6nnukCDcvidyS2HMFNABumx1PVqvCqGVsTVCWRV9gGvaE/4B68QWDuudx/UisoXV2
chwo+brXRR7wfrH2jYJ3SljThWdNb9fvaLh7Rksh3RLrxyidxzkgEFFiL5iqlkk+FFzBqlHtQ1PA
zE0Z/W77XZrrOK99chrBoprCvPGUuVPJlAzYYy8tanf9ybb9582CFyHLGmDd2nFtfDD4FwFTvYSI
TwzA6IBZeI4jVpiPEkyfy2E2a/fVCCDIgu15r1RDX/4CtU+SpnoCxkGdIGbfBT0db0eUY79GPNVL
XgZbtvJ0o1vDtOXSPC3/7Utc5yH21CEYoM3G2EVz1pzhMT9A4DkCFeFbc/z5KYWq7UWZdqeYVaeR
lNqdCLsbYdjt7v0a5Ib4tEcLf/qd+xrMbv5FGT+TCmsT7D+eR+yB7OMCEfu63kybNx7JOlcNBi4b
a+yqvcmahHJ7bu1Pv5Txq3jhauD1KB9VDoTJCIBzfDmq/w7nn/I9DjVeEP19zqKaGgZsk4HHhcnE
KcPfXxYlJuUicbVW9UF2MH98P0K9IqCtHs1XsuBZveK1ceIde2S4xB0RBYuS6lUfoiHwtmpY7EpV
a50rKhSNd1aRQj/Y3lwI9TCheWmrOvzXkxu9tgO2pHVpwgw5I9DLydGEBQLsqInfUuG3GVQBgQoq
iQljMLuYKjjDoaB4pShzOhviPf7WFjPJu4Ieph8BAJ1aSNnIj9NF2BtHW7oVsEXZGic8WnKDGO4c
qeyEGLr6cCITYdblAFnmPy0z8cOR/RvrC0CC4A5d2fM9BmnHhUHfvBSXip9tC3MCYwOQu8XH8KXt
g+2qWL7uXAmCfrZvLkJ/+OEjOof6v6+KvOM7aCrIDYiOmLUts5L2e+W2gnBR4qtaPqyQy0Hkv2pP
ou4uYldfLSPX/uNyZtzLuRLk/101URZyNEDAnvWwD5LwVMmX/fNvYyJhpY6gUU1WMcWn+9Tpra3l
wFTJ1ErtksQxwPcPfo3jMIFURQaLAE1y+zCSLbpojJ+arf3dSgxlsLIUpl4sHoY7lwYLNI/bBiUl
G0S+NdniMU80/LzrjaAlVkW8iAWdKlZipEXe4CKp0Bn2Bl+S01Lc4YWnbVqqozS2P3rjTGctJ1qT
U/5lFZa3ddK1KLOPDtoKqQpmFHG5nhvxvQW0u3WtknM56xlB2+YBsF4aQFTBBeEt92A8eJbltt2e
SVn4PCEQ1J3g/BDazhVlUs5DImVi8jbv91JVSgm1kH/u8zdJsyWGtyVRIeCJqUYGSEM50gJyvTs1
cthbMkJEoNcFaUyhaWXtqBeX6kHmVhkwKgk/VdshY1nOT8cCT75RZ4bRF9m63wIM5CvRo/Hxsbnr
VoRmUyX77NOSn8/aam3egD5J9v9l++jmPYnCwFNwTfluhYTD/VsB4+NHmjHCWxErUOKE7MjGUgg/
9cvu6pklkocxrYm3AHjSYIKyNn06l/LY6Iew7WGqwfEdcnXxCU6k/WXyYj4Dx27eU9KXTk+bm1ma
bUI0tDHxgf6s4a1zJ5Hfs5vThuB1C62xr7GrP4T/7X8Ob+ZDEeuGxslPEqkUGAYcipjRryuDPEk2
YSgjG+F8f3hAZ3l+3CWcq5klhyMyuzvq81S57FrxD8PMonT4lTTTYl/KiSqwf+2YS73l+sjjTnLL
k33uBECJEr+JO8tSFDj7xOpBM2spkVV19o3bnDtptGzayby6LCoT/dRybcpWKvdLeUMRcdLvAcaN
xnniKQ6+6dfylJgfNLo3H4HgalKkp+pUzKnPu5Bh29Q383aqwHxG3R2co+KsldgukyVXRKblsFJG
QKx8Ux6SQIv+72NYlCYtmWyceTFXARL5TjH5jWLl86Jp0Zi9oMFOd0JWAkyIPU/B2rAZu/2qZUzk
eNfXVnTaU5+Ms3fZ2w2tGnxkZqTNeDnX511OZrpge1VRgRidQt9gkk64fLqyMxt6b+ysloAY1EAV
uWXJ0rvM+VfosZQfuqjlKzn51x86h52r/Qw5zVse2sBAKq5hZpj8nj7eJ0o7f8bSoimErSUkqJGK
TCcrnEgwlNSwKDpyetov6kpaqPruCHptCY4oRfbgStfZLHpFJHZilvBuyoayWqr93lflYK2LQDg8
eQqCq59k0tmAuqtn+/gQsBGLyYs4VE53Rrp/QGCUs2qDyMHfO3RKoxQeh/0zKRwgmYdy8PBBDM4u
1qO0wdcaMV+4AyL/OsCEm5RYzuxtXd1z+Ek0XJSL94hk+YQfP439feNqyux1JfTuiEMMuHvHfHqz
cqVBl4PkVewTFU5++ki2/dpwu4NXRr0OjxeB2PXvbWtuYc8LFbCnFsoKTzsxaeYWeLAtE7riTHfG
ynv/q4upG3AO2aVZ2FPJs7cqO1S02eBYbOtANvCmDDjc35U4bR2JF0+JhOfOptVwwZVeMojlgKD5
V5GDVM+XEH1Kb1A0iQHteJyjR8lY48FNodosocbmiEt2u4LOG4WNMak73Un38dbuXQkjrPmgLM4q
TRMYYj3Bu86XVMiu6VUzAjQJunoAZVvCOS2jhmPHIg7bNVFDT6GNTwH1PyDmFcPwgpnfn5eyycfw
q9hVsGlBtj/Usm2ZC4tvsenuQXezt8/F97QZ79wjH6/gjME5dfyyPBHALQk1Hbu8osyXGKnnqhRd
mepUDch9PNx6GlAlY8Qegji2kWuGZRJ+E23Rzd/h+9/lhNWBqNrJ10afRGy/1OnEAJthZZ3KY1Pa
frUhJZqKWIKYTrOD88lsiiQz6+cFAGltSSgGhc9dMhIpizokzyMnEtYbJ9prwhF+x58w0DdhaO0l
cn2q1jA6Q04J9YvHByEiPAh/o55TndNegDqfYKsi3a6yUrPISTQQoOHl26voNQ1M0T3nzEdF1Azc
wrswGzmgWtLxUGJ5MiSdNJNGrAh2KIwpxo99C+jYcXf89VaBK18RqUFATy0MY2KiHwOFE82f0buA
CfQF2Zb7VRhKBOWG6Z3icdNu9Wp1BTIeEacvH8FJ0FPIS7Bqb+VQsOrY0+0vnYUrdQrNtNmwLAdY
x4V7eBFmgh86o7ylGBNUIA2gQ9h43H1mNvUmQa0d6EGQyUkR2XW+rZdi0lO2U+4tylEjt42cX17J
6YQQrAzH9A3E/mLZBBC9mCYNGGlPPGekL/qq5qrj9sTFoUQqBDIPPYHZt2jsJOp6od/qi86al1mf
k94u8B5YMvKfzYBYo9w11nEmts5cGb0Ql/Ngm2Og6n8ZjePNn+lgJizJ7LPQrKv1pBfAxGdfshSS
DDUDMKgP3Df8RHJWxbZ1yukhPQxphfM/xApUymZPLe/5N0P1dyyrYimye5Bob2x6+YUhI+RYYSim
E/adBdXpvQjcV3+ucvSHaYqZQripljOqDx9L9PBE/Jk0BnoV5AUiMBOu/deNoQt1HZ1O8bTKz4HE
jWTsLd9B1oLlFS+MDW/nwNtQC8ZV3Ogt6HWP0zH5hM24qRsB40YwvLKUWj6WRYIE8bIS6cXVKvSk
AryuaCrlEUq+911EaAVBEIEe0JfHwbR1DY6/EpeIcF/eHKz9S6Xos95rxI2K7svTqZGaGJcnX2ZE
k7ZB1wo0xGvdf3QXcsJPrb//XecLw+kjE+5tcVYTDY7G3D6qk61duTZbCUYzGq8ZWh6bBF3YBaxr
CvmgNVp0LEJ0ZJeZQJxK4RbfGXhh1HXzrKtJrA3SBY+b2Z1BYozh+qVP19rolJYwE46+KQRL6njG
kYFO8Q1Opq5oYWAW+ghH2kmo2KacjDYGAvYsuokaC2tE9CmgmgGwQYJWSivRgcWHJmJHCBIkoj3Q
WkZ1O5mcdhQ+eOd5lzGWjdjHjr6QI6Fh1HQIXN1Z1MKJQihCfdfGtoXyzMM7qp0hhOvCQpGe6mF2
LTW5k3pVqLgJy6OMWMfzQc7XnFe6/HvYlPh9lFNDr2JjOwARDXzvfeJXuPpZOM0TJzyyr/G1DyCh
H8BLbZ9NUK60xOPO3jgo7IEzH9ruuBZu/ZQy63i9IUMjuDX1+IFEybGYxhaYjsjEAW/Qhr//2GJz
9nbYVhDxlRBZuKM+DHBDVP3QmLM1uFy4hfC5xIAFp8qxGxE+ptKnBCjpIYTd01uGwPCGtCzrYpeN
N15hIc8+vrwkzJtdPIERt3IekuJI2Gqa1dyii2ziUuavDBLrslRyTyotL3vD9d2iIDgdNQpPwCsx
umDp+gHchjy58IIRU9TO+8evzM+L+MobKPLLNeq4ma8fz4MFKwA0wMVH1UN9KpXKx1+JxWq7SSUC
j0brlIIRXGlBNPwW8RBv1RdZy3hoCImVURJAY7EPnksHJCNI5/4lWM/Iqhk7fooJ0FAWoWS7K0Oy
4q01B1EJTUY5V90EX6m3n27jgN8yaOMM0MY5gpSsvUzMWWEDGV1bC2sooDgJDxWdoreoQW4M0GSz
aWTuILZtF9zzmtBOaz7iK9HO4KChKAVt7zBYjec7O91zW0a0935jKvSGCKP3pR8sACTGNYW5sj4m
D5ERJlWPE3LAvoQonvHPcxFBeG5XiJ2ZxZHlTnCIOfUXEhLc+QtNoOE0MJHTQrnEEILjTM4RXHXu
dQR1KGqQ1wT6trajTZjKgNPR2uD6YYQWveDI2uH/kDYsh19RBHm6OEKkmsipkR/X1Vd+yuLu4Bvt
XR82M6Sw41F3abuZiMxlVe5TxdQV1nil34W3wXlVxibGXT8GJ0SoT/uzrB8impgIgsQnRiTDgZiP
g3vZvSi1SwJAXz+wBkmvp736q+R8OBt752YDta3wL4dLFfIqsfcp6fFZQwgC0Jb3HO3ZZg0qpZHF
JEjDGFSNXFGocryMLZwoMR8U60VHbT1gnf4Mrl5SzjD7S1kBZ4KY+LaETRDLsKoJBdS9cEbDQ6lz
UG6ct5NXg4lUFj+riehY3UCDlcP7PSyuBFLBV1SJ3Mf1HhHOMhMvDBv7fqkS7XqbHagk8KrMjr4T
DNTqbq8i5DgoI1eHo29pyUGj3znIWQ0YJPal+1uO7Sd93tByuQkYC+ZXWxcy2uOiWs8Al1hfD4yV
vB+jCXTESL+oZHRTbEXd7rRzv3ZGJJ+LYWU3Szfd8QQt//pXqKYOpXlc2Dew9VFOC9v4a3Ydxzmo
Oq0tb+gV8zRSpOxolKJdXwEktnWC2ADVxkH5ZeOuRnAZgjZzhjP7SWSK59Oo24K347kNzpWxXkqI
09y70Uj1qJIMUL1sIK9qhiD2VaT+fbgBUBCIeDbGKp/vjhIiRwHNGDykIqJRMx+qUH2p/DdPC8v1
ttnY0p9NN45HOGvqz1bNnGTfQD22KswMfvgXE/GbOjthOoFn2aIPQRMBoqFnq1XXA5EMvRYLbLqQ
kMTuey3nyaRKRtm2G69VczZKyXHyCFV9rlIbwtino5P2CtByH786UkmGdH6/GP0m5pX+FJjgkEOn
XCP8rUnMuKr1ZiZk4ILJMTSMLYBOhjv3+S3pW2PvZ1fBBCbnkYYvRMo5V700CT8kghOpwxJOiT+m
GCGHufVrAerrxPIWXvUWdt1lYbnuwfuXCOBz+TXYaIlG8LsOkLclbXEg2KKFExeh7LBqYejqVgtr
NHGVj1bWk1bwx4tMrYa17DSDMMLYBHkRuVSiVEG1H/KZj9mwcmq/z/tLM+zQMz5MFmACvDRMd6xa
dKCaLsnsQ5rF10FoiERDFupDi57lMBYrVgET5gSEuhsfu7Jzo0YbUv0IqUPkzv1ECbUrNyTxYDWK
iQbyLgoAOKxcGJOTS95tH/fzXLu+lppzitAChUl0JTEUl1UwAPKAfPxa51myrH/RFZzVZuRrOhiQ
OAuIfTz5iSSdUfIDbzV/PSW5MsUwU+7301W3G0WgwB/qBvllYKQsxzt5Y2Wj9WvPtf8J3IjuirQz
A6yq4/xU1iI2N9caMIpk9P5+B+3niyhLJk+F9V6vbq01QmBLwrGDvJY/w88CxS2hq2qt5ypPoksP
gSQ9zwE6jjqVA0f/uCy+sCC1owi9ANPrt+2vuF0E0Afnx11q3rk4I7gSRCwtmbk+cEcdOw5HviOH
3SlwBDUqkhCO0UfNnaQuPA+93/qOn5aSalVvHT16qelhCx54O0amfo501qpLeEfFHChyMWiQL2KN
MnlwBQneB06JlQwqqTzv/wYR+GP9RiYK9/pOnC/XpAryfiEOV+3M+3X55wq06cXTCjoHHDHpT/LR
pX1IaU5sPGgsDfMputbbAK6zRYQRX4aFbIHAd18tWpnJSY0IX6hDjyBw3ywr9GsQQoBCeuM/x1kN
VGGc3kSnBm31yVQ9vjU9ZbdFukxRLwaTWNCt3W0NPm+bESTqdgYAk3dgQUA4slkvHwSfmihs9aXD
avRi8kBrvURc6JH6unUwielOHZKCYB180sP7PMvF0oYUFpOTN2AbTcUvXjBKxbNzMee0AXx8pibd
WCe6X+9WEr3L0DzZ68ZnZsUCMRBBDxZ0LP68vMDwTbgg/t9UDb1JMHkEQU+gElcnEFblvvgyDSgw
4a21d+KcViJIpTb44E9QkMjv7Z7xu1aP0yxBDRksQl3RvhvrS6jwka9FLbFiER+DBIijUzb0egTI
Tdvq7G0PHHxLPB9zbSgrXuZycRaAteQ+ETgbBgDPrnBaRsK8oY1A6wOfV9KvV/BhQbwPFZT39Rx0
1ooOyJ31zTCw3ju/VQhzV6xpjSop4fYvVNlkx8G3/b7UfHZjv8NYEn7ldVliR+KkMGoNfZyP+SLk
x39y63MZCuYJrWyksdc03BWMFFAToRXf9HRBhpt3BruV/ZS/gCplfc2ozDt72ZXOFnEg1AXIqTDg
8x1h3uX0rWXTDTA4woe5IFVYxnVXnAavQjIsgyJkjFnBrl3UDAgBkT4RetgG0ON+U8+5LBMgtebv
N3dMlVibN/91w3qVM5q3qxmwzyMCMGS4Qx6bh7i0Cg3kzhpsZkD6GxxTJJrrJGlqAimuleqSP4YK
dTi7yLcRhWzt257xnHFqNltlmhWMLyVSb6RhXRt4lWlz5c2TJo5l3RKMRWIcBE1wY2HuVoRM53WN
tCzW2PuXo9FMxMOIu3Y00tr7fKXM7WobRJnRvkFnn8xd9O6xunAbMJFkkD1mnAEPe9lKzsM/B6ch
8tRIt27pe3/VRdES/4Hg9Tc0HEAwjPjj6olV1ReXrpN1dDr47ZQ5AxyweLG4FYFY77kalJpWmEh/
BgE4DNBE0DhlaPI23WI5dIjsNSuan/NnRVrXyxlL6KQbtSrqGZoPCmrIXKcNovzj/iWH+bM3Gp2K
x8U/njjxGJ+CNbHtoKOKKB58VTefId+hrdfroy1BedRsBNDFSK09+yFy0wchV1QO9qZgDHxYdkGx
6kxZefDI4P0pasIaSlv5SYynXqysNmacOWP0IlTyZyRn5tFiKxtRYZzwHVdZG3fa9xIdxBY5pe9b
b4gI/ip2hyZUxZSm4Esu8TtnjrGDZpxPv5Gb0Ez9HxhT2SlIdNX9Q9oYY0sae/5BGaqm93Iatl5b
nrUIevj2KPPCFObGhIBSZJYomC8cWK9h0K0xNK2DonlOfjCJ+hhkUwQcfSwf1ydCyNYcp84Ta8yk
+0RXaRjXN0YzxC+Ld3KDYkH82mjZviO2wsmYNM+DRiQ0XxIdfaMTdDUYZnA1JGSyg7GlgR412AtR
S8wKy+izSXJV3mMfZiMElSI1svZydMen+8PkxeJbrNGYZu8UBeR8IP9Mn5CLe9U8IgHiaygufFlp
pVDfRalKUpJhG2v7LpxnAgGaMFva0bwT8ipaYEbdHE+HlYdEQfsUV57/Kb/wKEqcrClZoIeMN033
OUtdvs7bASaRY3ckq1DOwyosLEnAMeC7EDy2Y4owfxWx0tX2nJUapQETzne2n08+AWezJ6ZMOquy
YWRThkz6/Mie9RpFuqLuQ/NetfLZyF9RUNJ7U4hWXvmrwH4W5IxIqrpw4rx+g0REEqYznelsKXJS
fi7au5uZMi/55ZIyzHV9k4PywMRzTkMokCg+ena5aBIVU1ipYIVJ2PYlF41vNkuhLn/Aeljah9R3
zupdzLDiA171egnFSrcbWCSZr+GVSp9ulUM8HHesaFghQcqy5GA+Xky3uxMu/+NQQc5efrSew9G2
iYaecCjTLP8i3C068eUpvKMrzGsmck3e/wq9TNHxKhyg9ESdgxOdk4UFW/ylUiS9LGQoqF0ix95w
wPVmmS8KLRhO/3q7qwR1e53Z7ytuyuVCWeOGEsrdM5Rqs3aWGB3pRZFu71gwaYVjfOPdb7zSMnB9
MOsX7RZir+Kg4qW7DB9YvnlV8WA2hNRLDcbwwi/wRTpSO1O+O5FiDlGbpN+HHKPCmgWdBXkN3XNY
oMXUMO4GHdODbgcfZCK1qyaZEwWr5t0+vXmPzgbUDcRG6igs32oQYGtfrJp8ptSl8F8nnA6uo1OH
t7eZ1w0MjCO/spNjZhehDu2NLBu882MB9IIeRAi3a6R64SjhMlD6oSTq9+5uELGGtaVTt18ojxDR
h3KY49Y6hQhSfopGL3xOWIugju9dex20zPvJIBj7QGBJVfgb827rJH3fGihlcSqLB8qw/o01jtrb
8oRBMT0wmc4ZfyBx29jajW62tNdtAeUzxBE86/ZdE0XgxK+4WLCH8Uge2LvikTOUTIU/Fy9nZF/O
6FRCwcx28kSEls1xNacLFKkOsBrz+ymUSsffzjL2X+O/1zgq/efPNljB7rO9e/qIRY+0K0QTizDF
lxpxZ582qe/O3kQnpHcr2x6O5xGfVtkSFfr7XqEeN1FlF46YOitoq/bXfi+guAzYPv/1ZL68CpPA
xOmWd3utw56Hn0Q55iSN87Y0bFyvuDoK0pvH3wThyh1zj0QBlDQG4EEkZmgInYWQj6NpRbyIuQL2
8SLsQKACW2hH3cHLKgj20jSRQc4VbLVl3bjglvmt8FoowWHh3OVkmKqHQA86bKw6NbxVqEyT7U4n
y5jmrij55pywP7GLBlfy4zL18ZS9SY3kT6UaUYo5AF7dI2PKFNXbdEJwWNeX994GISz2uTObnjgO
EBKHck111qS9eoGLJVj9R6Vtw68A5liChCzDh80OQtiqaXSW/j6lB7Qo+zRvpZ4M06ZwJFwu/CwC
SHu9Yac3BY8jh5U5uV86MIp2dtCQN5oDdpmx0vSD4zp5Oav1MccpN0ST4woqq00Fv7FbQVOChCnw
7auT2JbRcddk8OqJV6pTIg1THnLT3gmhk4DFI+NFMyfDWUeu+atHyRIt9L/AOPK9EIk1yW2Y0zx6
ToszEu/SMvrFpc8u/RsKnS39rBqJilN5irmUCWqWWzInjEAD61Z5PW0KlrlQAF1HJ6k5i0C0zRn/
tuqt4UP4pujgNLh/bXOSo8jBivyq2WLnDIl8T30mAMutj8dNRGSAa/iCrQ+k0WHt0I3W8Tf3BGyY
g4aGSZcc1OTGgC8+B8Rcy3Rn/FPAax7aXi8M695cYLDxQEWLH4nNE8rbCw82T947fNoUZn5zCKLa
8oeFGVhqNGNNy1+VYPSLlQOY+ez172Jy+UOJPVfvw7rgK3FEmnQ3PN8yWqkRM+nd0KpD+RW/tWls
eM74rR4fsKj7w2Nxh4FtK1aO8lB9P8yx4tUQ8zT1dZcCuHRqL+AkOznVuBrpbM4Gl6r+0IvSmM3/
6OcGLCufBftiPV7DzOGQlX/W6O7dHPoEplbC5jvXqctTqpx/qJwy/UetC2m+46ssWEsqkKs7Nrji
iPIWr7bxkGIX3ewuAnFoGzqcS8PacWHDOxysK4K6gnmRRId3ysQmIoXv4LvRU48nHmPwWAtgxsOa
HdXCwgJo6qzksTfgtgkAkSO7uWIKlnzPyMxKHJ43gKSjS3sUW9VCJQQHo5M3XNxjvFUWgHNXyqBV
Hovbq3v/0T+RllgBjs8pgAJrfKt51JqEf00hkO0Jw3z/bKiHtS9pGZPBKAkSwfrcqvEPRllu49fY
+WnsoU92mznWE6HWGfMbc6kDRUwNODXw1UhrlZPvNJHlLG2R6Cul1OedP2CQtzMOIdqTNZpQzFeM
YzyY2JeOXsRevY1fTmsGHH5Jp86UPtAeYbQW36x4Z3P4LQtb0vwo30kjfps2IbdUViaM4C3HcBi6
E6Z7t1xinMH1Qnh3R1l+ILg1qKlKql9FqTpbgGbx5k9JFnzKTkjo4YGozvyfTMRRPvlnxvH8R1wO
7F0+PO/dikBL6kncWleqSTMSz25SucAKpsZn9G0tpCDPY4CroqmZeMB5QCpOuMEI4IKHVyemagkP
c5N4uARRnpeXjGN3yi1o5fQQXI8wgYNwUhIRNRoc/euf+sspO17T1vY0wIAUldIDmfUIJDan3StW
gxMnTYqioGJouxHV0QwRx0r/rLeVTI59y83nOtmP7VdvnKh5OYVvNjjqJswqg7hkgjhucD+u0PxK
1WC1uL85AGKy27QXluLn4b1efH7PciQYbUmO0YL2K9GHP58gtbfJY7c3FCXTCLSO7v0mS5afnGHX
7UOdI6aBJPAMnZMb//8Yz+JTEz+FIYL2iGSB1PorBb1VRtAjud/EUrTQmsdnlW7TFmyCP0WxZnec
SjL3rX0dEXEp0EL91HNkoX5Y+wPLs+Qq4ELkGE5YtBvEpcBgkDv/pyhEs+dy6+ljuG5ek75nzBMQ
Dv0dBa6lBAuiPpd8y8hz+aKa3Xn8TcrDavUik04/lV4PL3DBMQNsrTVya5t2oHqZzmpDQkmktqr0
kXg24OLq/NIKnTQBlsvjwbbjsDpV7+ESeLKtzLOimm/u1MO6vMOJmkDZ7erFdNp8oR04d12EvMDV
ZLlSRoJEF9L43zJHJoLGzezKjsqGuh79JC68IjWXZy3KmetPHy8jroAr89afv73XTq27no8LBvOz
SsmcVbfBbu9qLXVGOwyLSXQOh067q10V2MmYQ5jJp/2jOXxdBVkd7ZOwMOJkU1QS8oj+99GzlnJH
BK2pyUPHqpCBo/WM7J1xHR/pJudJ23J3pCqzVFWKAtNSlEInuuWCSzsW0oPYoq/uRBseAmX89g/Y
nBqt5QB6qJQs4po9ByUOwQriJYcOvrL66X6KLSaY2lo/Ej0f3d5YJpWVIbrsqlEbAqc96f8SigiX
VmnKUQYPaj+5mfz3sOPzeue+2TopfkIsTfP/joFuuyRLUCocErXWAQHuteVSLJ6zmuQBkM62KTWn
cnA8l6IMAeEFHFMR88ijo4ShnCZtj5tcTzQrGCQhv0C/HP9Ry1xMITVSyOKioTww43C5HJEFb94r
1kTXxt49uo/YSKaP6wPOLWWH+JD3XF5GytPvMUOYvAHYtHVuOryJDD4nns8389gN6cJwDhNeQUb0
AZtWJM2b2bsyagnHOK8ZuB0FBqXH7v6PDANlhFt2qev93f7sbU6wvZSQpaPdcOgIoGNswspemaP5
fn4l5bIS3Vns5S5ZwZnBVvZpyYLOnnfb01TAf8HcBST4XBHKScODkDjfe+t7+iofNZwA0rTU6iJS
hbYoTUHBNDFufJsEMVj3N1gOVutnWFQkjXMD3+uvZ8Z9uwBXN2jcx5wHDUkfQQ4E2ES3ar6DFL23
casIV91I9Tdvw44mO1eLbZOoEgaVY0c+yD8E1+4txO66LvZOrWvGy2M9srKpkhCvi6rgJ3Wcm+Tl
KyFlXR16fKz4FbDY4Bf+yeZpEsKTMDnBx0iEcUafOCPTs6tsCMAToRYgOC0T+ZYtKuG0za7z2gqS
hNnm1NKf1A3m2IyQcKjrq7bfuVUGytl10Yuvu1yH9BJf7HrTyRm8BCIc0Tou5NocLIj75PtDCS1A
hZ8sFOiIyjOJRlooyuWPhicHA21v9AoqGt/+d2GaqV5OeSjBN0dmYwxic5s71AGaFcxd/8xMz3Iq
pJxkIrix8wLUn4cxYtemRcZdbhnKGSnVOVyxijSCpr4JA5l/uMnPkaGMFpcJuYW20OHb9il8ww62
ewzlQirFGSgCiCUyjEft4sQThz7GTzfqy6eP+PIlxFCvUND3eRY4/N2mIfu8z0zRFEn0aZ5NmIVY
Twfm4zW/wJtrHowecC7SxZPhLP6qZ4IaQaE0359QJ2/W9IQBpS8oZi9tKGzxk9rhlOFC4HwftRYi
ru5a/0AVEfzJQCWacdTtypGJkM/scLSJ2tSZPqiRm7VdfH7nC0RcQNOryR1FFTCrU/ot5mg1JTYe
BZ1hUF8z9WV0CUYTTQDjT2VYB2HzLHTz+TLg+lLp1hXVMjmvw3zQa18vKuxCZi2RKTZvYX5yOdXd
6sS3HDz9w94Bh5etk+/KIuzKT98NlF83sCNNvCoRAGAOO99kiInCs5y87ipDymbHE6Y+v70jRfS6
KIki+5OugJPGGkriqfxqVcOx3E1b5am9xhQtnGF8VCaoml9uKYdN5W32bn4/IIU/4RkxF2AYPdd8
khE/SJFUUVK8xu7Ga9NOKk76IltqZJLuFJNnADgfD8FCbtoGA5RI1f+LBNoWUooxjWP9uD/9ie5d
vGmns9Yauk+pPMA/6OCcYM+bOyy2FXBNu7kopgatVzTsjfQfRbXV/uu1nUCG1T7JhhWhR1rbsmio
TdS55TdL9W6dWnAk5hQWT8O2ZWcNdiY62h1GVlMaacUi+Z4FKw6PrTS4jcDlcSQ4lo9kEW4eeLc2
4N2ysax3lWG6fLDd1bDNeEKSDXKOBQB53c/IVR+u9SB0ZJeDl/5Dr83SDzzq/6CLzJ21wnhaSOot
uNYY0fNEwI40QYHJX3bK+z9LzRGNmGoi8YLt9gkyqZ528GRPXZ3SjMEwBPHzEku8Fzyuc7kOVQUM
9k2FH33W2pBVavHygiTxTaD2PI0oRftGzOgtUTNcLuBrisaOk1wFzHkqwASuLoYWJSo3oAq66rp0
HkhwXlaedDz6p98nJ0M2XItGkNI/hJbuA3YK6zOkcby0hPCgHVx6+tqf4m2Nns0HyKlq0r8or6WY
D2tbgHY58IiK/ZMHJC5DiGdHqjQ5kgQR7Sy+z4r/ok3vHFUHZ1SzK63hMAFqzbiet2tf+UrNCCxw
ImLKuoo8i5tGpN43e54Hq9pMIMIm2wAycR5HZUr3Xhs8xdN9Yv33Uy5TbnqjaCmpo9l7CWT63BTR
YDd0/xL+u1TEsr8bSmzQsPwxHOuzj6L/VhOSR33aOFJCk5h8gD9fH4QCM6RrLvC1DjYxsgDX7IE8
C9fCzu0fNhxCquycqXioeUOB539kmHaN9XOcppBjH8Q6rVOumIyrzzpLThvNTnlbP/CaOLPJjAVA
snaiXX+tQJLacQYYzq0khLs9+Ysw0PUtILC3dPMTvkob61DxRAz8y03xUEFE8ZfLXPATW4uogo6U
kezvdQvKDX7B4ETiESMNlwWLUtRzv4Y5daRFpCyxELSYUlQllcM/fbq8QKckHZ2Xsdq0QJX1kd9K
KP+5DbMX4J6/hTrHZThePdne7FlkU6DgX6DmdBIxSyzLOU4R+tEi2altIZnMNRJUqWEMGYZG2xYT
aZSWCQ/g5uTwRMU6kJnHVhyIk9+qMf0ZQNp/5fBG/Z+4XDzOCkpmNupswkXTiUxXVY/D9dUICK7V
5lrFu2ei7D+hZALd/InyKTNU5EwiNRf0W6mpMJmiRrxdlV2KTh569tJH9aafPomvVlFCknPFCrtN
PN18t7HX61jCjl60nIijCXILogPFxjilebBbh5fcP769l4UQEWlOM96G/V01eI+JydOZaa8f0ph+
I/PZl9nMYnh3oqRzRThGxoEFR0u9kt1JqmzYttSQyZICrgLijHbrnLHUFrnmcJe1JlfzWyIP+gBL
f0ZviZOU7eZBpRNTkde/VQIXGHTS4f8AvGwqDnKw2ndr0azLvVv805rTkXR81n3VlJe+xEtl2lpY
vK1EenLtKk1UVSeYo8K0DnLYb8nPCVwEXxShKwBgAEuK92suOvalXlHJSngPpa1S3Os5k1DMlfLG
K6eBpQfsLp8yXkml1qg3bcuSnWlhQKkQGf+MCV2/DAn3nZ4+GrdqlyxdCYPRfRbkIVKxZGiFHRql
hbnACjoSFqlib61HMJpolTMRVCI8kv5+rEw5H1K5I95vQzZ62j/brqU8NK6NYcARzIi5t3OENGDc
1VJMTTDkgj9n3wEu74jCo4akayKOoudogFKdP67x7kNzeH9E73BARZ0Z8+t5jKOHCg7o+xVy9uxR
dyLLXfgtLkDMBmA6rj2qOn+7yy0CAKKp1juPQhPYAvJC/ImLMas5LjY56LfAtNU2/K2JHisCF8HR
HSUnd8B0OBKYxpnQ2w+qY7LiurY1hz4+94Z9RdpLpPiZm1602MV/7csKGx0c/Qh5iYlyvSe4VPwP
WImVVFpcX3UYm0X6DZeijDYM8QEyOLMzkGBdRfpbnHyQUL+TJdQFBgmlpjR+RdIiyPUzazcydGHQ
k0PzvbKOWkizwabC9cwhwsTWR+WOPO+3Pxg1d//SGgOn4YWCaXslu/h7sBuEXQsBksIwyIKKrRgW
305MxEcBQpDnO7I2G6dXrleG+lVTOBQoe4qwq3urCTS0/dt8pOSMUsU3VUNO6sdYGOahi15Qq93j
HMiozZu3R/uNwjG2avq619x0epH/MqtBocr1dAkfWTci7QzrcjMwvJvlvrHZIQPd3tD1LcBLJGFQ
JaeynK0Na4glH9Kv/GhWWdkNDIvYFaz8ejIPclLb0mq1O/OutdhlimaRBc7E0benMiIg7Dcbi8Po
M8hHv9z6fKiGj8+HO7RP44V8m/emMgAWVY7As4+4tg7/gE3UnMwnhH3FjhGuXmtZEqX+wne1yrJ9
IBn/qBKrJWBuGeH6SZT/wqqS60hxJW/CwuD2juEtKt7nXO7z5jvkrMhaLF12rlRLWriG4ycjAXJV
CXnlcBR2L3rmGS+30yxPeGlMaERWPFYIABpQTYR4sLOsdhIkWYUfOYAWk8n9qWTojK5Um+1ZgRvq
ZiI/XhYXkZGPSqF+rIoZtpMDOodXYtmNd0Wl/1aGAy5S4ww9I8hD61PNZ5E7QqnevHsQfP/aVXCf
vgoM+P+kBeHQOX8QbNdA2fu9rg4ypxon5NveHuO129CPYu62NbmvJxYZulxXK+pqYrabP05N1w8M
o/wdp/R3fXi/MaRA5z/hMJBGsL0VCY/GMws0eNYdHVvpDt6p01fu0y763tCVb4RGHX4OF1Fa9e8E
9n7d/6No2biTOU2LP8J1e5EDH3dwiNNP7RFfvQkdBBjmdBRsXjyGQd38JN02sB4p04q0/8txEeSt
LLbk1SNEdcy2NvugOWzSVHZ/sjvyQmvZTrSZnfC7UEjsEgrvzy6SqEk6YlS+M/ONIY19YlHE5BWm
gKzJokb+Fw6pWdIigbhJhSQI/OzODX0Qy7nvKqwyjnmbw7jDAFwIxPXtF5PKvqcLG3DYLajbIcqm
QwhlgluJfQOMnXd/MlE2tCnWEEZweeUSMVb2GhM33NhtyDDxs0BGFNCH8d8riXSCpIfxI6T6ntop
uutoNVnATNWc/5cBn9twgrw6hLaEB3eoCmYx8SXp2J7dILoza8UGZwtE7X1B/NHPdUOFtd3pyg1W
BRFGQ2L8XCD0m6XPjw3ZdACVSwQSQWI64DWVFsPy9e6GDFOdBJL1sx+I/RhWtfNkhZoLs45Sume+
u9CsSsNBIc2DuYCQRC0/xKonAiMDUIr1Ci4GrlzJDMy1bxzhpQn3x+DOPNBBfeDWogHGcxX04zic
yBAA7mlpunRJWPgL0+AXNKhWo2JKircIwWLrHdc41s8Eo9tO3ofvkGka5tIX15Ph3cl0TONampUh
FOSvbvFiqBDmnD2BPpFa1xsU802SQ/Rw5PeZHxENl7A+9lTZSRBwfCY2Wg7CzNq1o35VRBCmY+e3
pOAb0PUoYGd0LXfml5Vw2L0gStV50iWa0nVhrHBSmN2rwlEEsMjNhkCbPAkDZltD/cyWZHimTNoX
vfBiZRGO9l4+gam7DNAEHdygth37yMF9YiIVPBEBJHbTqythvv6DujgXmwTV2gw/UXpsD0XOLZji
LllmW9iO2wiqsOkSbYMNwL0zU+w5OJxcteEM8UxZ2Tzc8hWlVGcvIOJ47bu/2gCFA1kyEaCjPea3
oJuoDl7l8gOz1kqPu3HQ51tM11jxVGaothqHUiGbh8F1GcmRvH1jC8lismGcTNQ5K1Gx92n7g//N
DWL2Y8xHaZeSMyOyKNwtPrObxV+JSJAoMkEiHFc70TQOMQugfvfG6xb5xjjI048+9SyNRlmsGu58
YThUhm2Wvt8vSaOFay5VQjhyCitV/6977i0h75NPzBwbr2QGbnM5GaJ1PhJm1J2NuygUS57rOWhP
Q8qaz0gU0Qh6wXAWwwdvWcKh5kbEdxFhdLKNbNSR5H7PZIcqejV+0K3PdW0inpnj+LLQkgFufxW4
XgI3YRE9CrNSpJJ1hKv5/O1OvaXCKDs4JKakF9A8wyg61RjGRYkdtR9ZjLPQzzuSDsDmg0F/XbKT
TM8dU2EaY6F4oI8SlSh2KGJ5lnvlWpq0vSBTPR7HLr++xWg3UlFsEk1xSPGOCp+cYDfEQ+phWEF/
WGR21vlQrExe/mUDBFPIWFR00jVOBuS6czby1sN9JAVjeKf65ZpBPyNjNA8l8SNwz/Xh1z2rRAUA
IAU4UK3Nkiy7g6NROts0DnoErYuTtEniiUb0EjO/jOlbNXxsRiEEsK1VPTAsqqWTsT6FkgAMo2my
mPo9LXLll4Kc6nhFlaCIjj7LJoMylbzLFX9GkyZuRoF5FyDYp/gpqdUvbWNvf/JyzdalmRkmbKkB
npugOwsUKnSeSx4579zabmojIv7+XH5RJjut5cuLNMyWKmSy7BS1vIjzVdb29kxBHIS7xtIsa6WA
FkKDvntOrxbnQGltLpR3p3ZJNjy4hhkS3PgcssbiGWkR9Z8IjkaDD6kRHO0C3SgD8p1LnzdIKbTF
ybqU0kS26KB+etB8WmLo0IH43oStCuP+ZjFHY3PpyjV4jd1E+7mGboBmVSa/i4iuIe/VXWiOmsP0
s2kLURA41HO+xEfyX14eTk5yhnwmX0C/QlQNtHSFDqEuCgIHaBXmS/hIoVEKDJW7oGzKA6yHQhuc
je5F7PBWNSqA3ElfFXvsqOyD/VfQtbratHVdOisyg2bniiAUkhU6whcH9E151oJeUTViyRhwHFlm
5tQD0xK9f4wwL0cd1Ge+1DVmwjV42uDTzeLNoZSbDHMxVUSz/QAE7eSDXByoX6TmFQpvyQlvwTDk
+vOfKdYFUOJA2SvdHpinJds2Elr8ysPDMajb+cAStIHxaXGWHQj3/8p63VryhIrgk3lNncOZnxoD
5T4B5jVMUjGYnp91qUwpnZBhIejE/g7OXto1m+E6yDbjt6CeTK0hwlSAE7G7BKs/mv0dtknFURZH
zGjWNC9fAXfOVrQy5MULyPhLullCKIMiyo+3UC2+ATeEcD+WSbPzDzUOt+E8J1xy8S/Dr3jYioVg
u/tljtGaBksIjsv/9JHOY1udNAWtcpt+lx0PZHlWXLziqxDhZ28+GhI6Hbsmx7M6qdVcTBgWGJKd
pNRjF+LhyWj5P3DXNobx9thym74J4YHwJloL8Hn7rj0Wt7lUF505WAGjhmdE5YVzJx93qKCw4KfX
z11eVo1cJVVnY1sktOnvtxc4FW0Dovvb4jPmnU9XF+8qym0WqTuDbjabbjY2KTGFFWvHqWwcnBjg
PG2kdxZt7w/f8WeqTN1GfdP6LQdjlehA5UhJ+79tvde7tMNGakhZ1tn00+S5rWqAc1BZDlBkpNGW
OTypgA0TYtzvW/Josa4V0aWNQrn9OEnmhizlwrhRzRf6mamPzTF+YDTmNXjYPfAloRgZv8hLttjs
kWqWtUdKvG9jDe8muT0kOnMsdAELqu2F4W3g0kBlbmFC02DdbYy9hmW9Tp6BcSv9L8UX5A7mahjc
vlshJ1yDjc3a9lre5b1qdqqOH1ZthmkMT9qNSA0FXQ0Z/zxJsstKEGZVGO1XHJ13bucHJy9HBDSA
3uBu2jx6n2I4P+TPlCzadI6lRF2LqtsRLdHvjk3gOH4mlLC75ztIlZrgrsPQLvcUlCJXDS9wsGGo
z5rFVrcuC1W1ElnQq6z/tYgSoZAXGu1lr/kjiT08Yuyg8uiNMBbQ2+bJw0tcViypu68EserZpQ3g
OyrkQhlRr83HYP+KgXcLah5KNX/BmmDZdKxFimnz8+xHZMni4oJU3qLFHvdfq+FoM1KbufS6WsJ4
+1srgQhymjgtfcEFqQAZ1773qxOETXqciVh923Mgp3il1BeQhErcAsc67rGOqPDvgH/rdd5oyvPe
V6mjBkBZFBDKVm2nRsEisRRh7pncGG6ISfu6340GcOJbS577I3Vy3nX3VxLxTNhRlKFPaPxokZ3Y
hu2bdLCRi6xeR17XqV9KWtkswu+JxUBIpXv/8NiWH+iZTuVlBIdT/+0SsNoLRtCslfM2gak0KrN3
hBrqAvtiI9Y5WJmYQE/hcW8tbPceeyeQplVQAeMM/wJtVzV5sZKQ1/ZuJEPzNR2e8SvJgZkPI1pn
Gfq1zM+j2nbhzjx8/D+1AluWpsUXFpUWRLRcQzpUI3aKIcH7zsWUehkOLmWe8Y5LBqeGBuYp0g3H
sQUCB5PMswTATNsPKJ7NmzSmm40WrnhR3min4xX3xK2FIW6VnwtbBNrN0ZGiolgGu/dDpqMnuIXU
ipQd1TwFffJam+ZlV+/mGZHDWFldzEmYfQ9euoiBcwdtdT+OBjeuQTCDzLo4hGtK8vR15Sq0ofoD
vLVvWEZ11RQ3XjXNFE/zLzm6DuoMofR0NHTEsl8iljctVEJjpLlfkuO0BlC2WRuuVh/DClskAHN8
FX1kgbZ7VowwwlZGuGBmAtRlxf8nPF5y6IPA94RMLED2tjxI7cNZziUXTvEklAPgMV4cX4HBcSji
GzbWhtcyfnCGUOQahMQ6xiU0+wmGQl+LbTLHTMM4C0641bG09nBsLYvgBCLCxCwuvjrvF/QRJxea
VWnVuJxnFnNKdNFKegobflo72+3EfOL4Ymbh7FNCOslOKPZ38Fkmr0+QkiuBScaRCzj6cXlLFCBt
7m/uP2iFqEI/RDz39RWjBEIhCQI//JEnPBg1EE2vwMUU4M6lZdtXSbBivTLvOxeiL2SWQh27k4Pv
ufli+hZ28XK3YrGZ6KQF7q8ExYgGMzer3NDqNQkTIxVhZ4UhrnCGSUsYDkM8fw2KLSM51sD5XvyH
5Za5QKWbXuT78saeGsXbwhinVqWKyNdweW0Riw7lEnwDMmmWyuvyVXgIdjbgvSaB3uSyK1WU68jh
pkeL3XqhaaSKAMqyUaEX0a3z1iXbQzvPkN6lb6ku6XlZ6EqUuPvnDa2spXYKzZ5klM8IBPTU32O5
U5iHJFF2dRyX1sdA8TQWo/owh/jLLpQfAK4P85FM7LB2osBridfY5f9DzofK+0uTAenocBnrUCAs
q5PvUxn7dKlM8dWsbgWiK2D8BnGjJZxlcL1ldjF4io3Wy8hQKMtemiNKhdYdWfZKE9hO0NAiEGGv
XOQSsu4DQ6AIudS2MX483cDGLLJjVyeMZOw6XwMWzf5DmzFLcxVE8NGg4KbvHvb8kgcQMuF7HReh
Uo/lVlMWSZyuycaO/FJWnkiZkCa194ezHdcaMIddMeUudfBQ7BN4A1NG/2H/pwuw2o8/3yJ6wTBB
I7XPvfvpvzGHU9zfc6g3Nmpud48BIBxtT2g6H3/bR8DmgFAQu/Vz5Cdy2wXrnnvjqofaDbRVshTG
MwBPm6gdANto+Fx/jyhoEUG4EeWGcVP3pgGsk8DHXC92Q6WpIPVbZGSvHAKkhGDpD1U9lzMzwSWu
LyIiCqLF4R+E5QLO7unfFyZDPXKo4C8Z7NyGyDlGgNaBtO8Sl1YkEjc6ZF6QiyROXnmto2cJpW32
p8zmWOW/2PEudPpDMoZ6oQsgVgb1wbX9v+7MbKkUhJK4BldqNe4FLzPn+e0zVApOnxLObitTREzj
6dWCxtoktD/1s7/N72HqK1oZz5gXymhmqRNeqC4vBihgpocLLDOy+HUwpBctBr+CEbkzPiXCzxT8
u+LVntw6RwkfMIH8RwpytIaxhUivsJShVQ8D2Bw6bfZpe7yF2Z4b8PhbwozHk3XMvHJd1FW8ISVj
zM9nAuzhxfUtcBy2/1wymmhdwjwCswaKwBVubueKDL1xlX0LKcEeS3AXcoZ3f8UEb8IEkgVqJlTK
BVQiqFe80uFuZhwyrjLWASOGdtebpBR+1UCE8041iM7MuYVC1x0sP1t1GK3DldsFY988o/mc1t8J
1yXHfnn+6ISgH/+oXvYki7tFxm1nTyB7qvwBeRAn7KhdaZDT1xEORFOFyMGtGaGVYz99XX14JL9p
PgHlmI7BUKVTD09JBOHvC7LXPz51zcPuP3QAHZl1SC2873cTBkB7+THIhKvWITCWdS8AhY18dcF1
NBNe43nyYeskR+4MD6/mHL/fBmDJXBFpRmDz/5g+kGMmhccUey0KOc1Ua9U85mJJrWf08TJSxjcW
vM6PRpAC+5eaBcQ5oTcxLUDSQy5FUNsdbA04tCEP+CBJsi5mx06YLS3vtSpJw9zoWia1rW/orvvE
R5tiTHO7Nx9sKwf7ZvvvOzbyTu0cJAeg5fGmNSsTnekRjwI3BHdvNh2LzlbPSkO2FBoiERIEPted
9utUXwT5sU11g2QRwqAy83Z6ExrWGRlEtDcfx7YGlO8sS2AbFBJ+wpklWkNaoLDWv9I+Sze2seVs
RLHXYdAkcaRv+L3k8Ftb7PPx93Twus+Ztgf5rrHEo84I8a2X6/RJZIAPGgUKGdivDDYTcOKxFHrP
BUmFNWEP4NtG2m84HTyDNtxZLrC60Dg0NNPhJWtk8Njr/nz9uHqHqWSIVIg7VjDW5ezoDPmh4/cQ
oN9Q+sXwzw7OB7faNr4/z5DEiZSA+2Go5spAC77HMCGWATGjKgsY1BGuC5AfBqUx1iun5pNs19x8
ePKUdCniuxpOvCKJFYgLUvANbDiux5jjHEWF0JRoLJIOjYO3XAxVTDdMmX5yMbW7vBwjxSWLnlMP
KgNzDCKvzUSKzZTCkB2L5PDNmnsCq1RG0iVruq2zaIqmau0XkrESP9mTi2kIVS80bW2kIvUghbY0
C5h53efSLHHB/KRA6/kMZacYootSHyoR8gyYNdSTnYPJvphhhfBP9AMx5BiHIoat0oR0yR5AI5yw
9GuS4EKDNfqAzlteG3CDKGsvPezRuMoRKR1gLFOgFkkp+bdcZcCgzFT7uE3NfuzbdkJ2Iod9OdfV
7TTTL3lR66bakLLYoDGIY7mG/dbeXyCUCFgq+iWXSq0z6MJgkBgQMXGXrjIaU9oAvipm+wCK9NzS
27WvYZ5CHa4GXHPZO4hq1wxB4O4yCsqgiWqbI6HeHtNjtbYqe2v34zkXjDSSPk7lnpXiTTOH6GYf
ez5P/uRWSlUeUumB1UeXCtGXDsBfIRzcSwpExzI7IOLA4Hp26HUW6ZUbvAUIuq9a2slD6SWhlJao
wFgxcjrPEjTfhFe4hM5FWicUUR5K5Shfvb/YTB7gMa7C3ImHk77Er42vqxuKbdPkKsvk5i3Jgual
O4ZigTTksyDo0POe+Z6tkkc09nW+f3av7O+rLBmHdbgFHD1igrcPNQaV9rUqy7CGRDX36YuHAjed
rkyMIh4TkC1GdDBiKefoiHB1IbKDxZvQP4uiWoXzXvPc6K/eSLx7PTB2iYNV/UlRrl4YCMFJmE3I
tsUCDSfctJDs/6JCo7aR0vnK374Cj61Eajwz4CnrYPki794TeHfrdJ/Vw19bYi3eDk7tlusjteMv
CoLLfFLIGrZF3MI9jQySc8he0VknyChIROmMg7Qum90d7tqxLAEgG/vI7n20e38j/pvgdmU6snMb
voSfJybrKXN+V+SXT6bfEzpdHOPHUsBpZ4150b9WVgqCZeJWzkFEP+JV9jSTpV5yUuCBbC0j7pJ8
kGuZ4gg766mf0f9OyOJUzFvxqoa4gTRGQ1FDUA1Y0dBn1OdhGVJtHG6bG4WPC3jibkpmyuh1h9Dq
C89XKNsCTAxwIiJ3a9nCZzn+7/lZT5NqyQJPz8f1HH0bjab3iUPvw3f3sKVkCSqnIEH6WWgRgUwj
GMUicuBpf1ntain5A8+AVoia+sBgfoUNVlAClvnJ7WuJWXa3I2D1epEI2bnwIEVoe54xfANefqZD
H5Ybk99AcXdITE7PupU5EQ3XHKNfWtKFLRqY8GSmfY4pxKZGpVBflNfDRPKOU0cwEz7lJn/B+Ppy
FQPpQBNrBuSqeIZTWSBijwUlS8YInMhhn6yUxXKUM0Eq+I88s+5Ir6G2b2Swoa/7eBN4E+gGg6I+
oap34vzgB/aSnriF6+dlLvzFvV+ZpkOLBjX4lKw/gfH/nWByYCzgcRWEExQu8iQ6e87D+dFheIO5
2ak5+gktFIRySgTwsP5Jxl5Et4HkuxRKiL9eIIEGq8XsKYkUaae9I6nzJzr8rLHv1u8V+qTftIAv
Y1QYhEGb4uYBbtWdw/XMImbq+Nwz9J/Lsm0JaPwcwNjwMYq+m/Uw2bLR6lK1V1WZKNeVWH3MTkcj
EEYFXy5I9WhQgJ2mb1eQx5HMNk5faemg2MUmNo4+WN3Iu+o6XLbKIuNhG1L2fTmfn1e0MEXqqr23
8Vy3aXGN0YckLRlgod0jCjbG6u+Rt2xjSk5ad3IN9/QUtKb3vZLv85GsowT1xW0ohRDAt0/Wgy1M
fLeOPpysBLvxaaS0MxQReSrTlY5PScSngu3/+/bKnXYXVGo/irBvKzfwLg4wBln58zzZ7/aoqgJM
Bfssljub6lbxeKx6pNzuj5hMmaPFL6KC2yxhMlMraSUk0j7hghqx5nn4DUc5YikizQ7HcLJ4dk8o
YmY9uSh36Tmw5mX2IAevJKx/FlcXeeWSmnOHCngVPbOLemWPOWr0ne8yYxVu6LYtE5vDlwim75rR
B13MOha06BdW4z2CQb2wgYS2sR/edcvowUmJsReVd+XvMbUWSxd9MFPO/eEZN9V6NYPhNLkEpGXa
h2CZU2E7oaY42uq7tJ9u6nd4UAboMTttuMxYM+LAwPPBc8FahAjVgj0GSGzKDstI94jGOtwlwzLr
dmFCSdZdceskbxXUMqHM3L6J4y8UM5LlJULhQ/9LlsclV+cDQE2obn9TZ6Qzqear/K/ZbCwbkg6C
KS8yJfomJvqHVn3aWBPkyLOnUbwbAjvw+TfPDrUxGVjmqHEvS2iENIdNVEEjG/SsWwAKVvbBClmK
t3RiUQj8RDn4ASP6HyKDM2bEgSzpTcl5ss+dv79S+ylwOwbrvTS9wykSHKhQ+lh2WGtyUExsNqpv
6tyJs3y7rIVCZckAaqXUmx8Budz7ZBX5wWF4sIizfUamqKHzsB6mappCXtW5XVnfwxj+ydJxsKag
hNIDmeh7GRjm4QtwiBS+pwEj6vhE1ktksVuFPtj6M3RRnoPGN3T0LA1DjiEa+YhXBuVQnwmSp/tw
F5KB2VCRrIEhvJmOb2KjaSQ1HJLoidsItDGvCz65T4tCh7TgeNIWGkrXmK4yshA3vHPEGZvXKu9V
8me4TreVUWrQvgeNiVKtwEqLilUioUap5lqSXU5efAVdB3P78kxO2NMFc6uV92w3tABCf9d1DSt8
JyGrYQ1EL6V9hQCNor8AS51GgFN/b9fgP8EfrfhleWOmUFvLP4k3nT42S/OTfTQoaC3cQVSSoxLR
KZ2/oehTIcFpE89Ert4WDkqA3qmdSdWu29eZ1TAeuVqi6DgRxoRjSmYtGTcisAZR1s1uVwHSei6f
tBXnvAVEtA9STmI2M1QVFVDXHxvqneSFTNQdl5khPRDY9r6Fe7NY53Se8/m7X6AES2yDyQZSpF5p
+aYNX88lmKGIDaH2qKNLYqPrrhuwfsGVj5JdoJmOf9Qs8SPVbgoF1aWh5jNb7ICgVuXskclBHjep
Wf8lclSnLdvFNYT3cJSL5f6XyKH7KMPy60pwT+UotDLxn+dM8kQJI5dVU7sdCtlsGEaUbIncqqSD
s8Ob6dHDLue6kcG6zsPMXY9zfWl1OB/yBP1+2GuZsmoYC2ApfMfpZuprDEZFYMA8n8iGe80sKYsz
3Ej9X6I16fnXVMbKF3nz8SgwMLFNvIYij6Sq9bAnA46h85AlNwpsIjhOZmzVIeFh7PhijJhg//YB
K2vRDLd7A6r64uplpRbNj8o7x+V3AK5NqiLmLD/giKcTwKMp7mO9BbduBNFTg0TDUiDabBJwDKhJ
Fmyn5q8e822wQMEkN+NVaMnDbjTrvpSihHvTUYSk2qtu7URDh3a7qjbxhoMDaKA6ZCRek5m7z5Wy
7Tp6/nGgTnb2sP5muOS5KkNlhbpI42pkefbv/s4veg+1FbggrtVDoPQpU5l8bE7aY/qUiJzs2TxO
fR81c9oT9UJxJTsTE8OctqeEIpUqelMHFA9uEL3uySr/gtETEx5UXzTc/GhmlzqTql7mP7qm/XY9
7GlZkNI9xCxIcYVbkVvP8N1Al0bJILlci/bJu8lUe41QXLamhZ9Qd/ZWlReppCUbRY5HBS7HiHU+
lxAzX2u2y0zEL8K8Rq3bxptzd/p+EJO3Z5bFofMjxPKOLjoS1tqXzM/6W5RCtGCG+6P7zKv1M85P
xFqVNnfd6i64gw4JbrJDJXzspM9Vu9wj2GeL2LExV8znP52a6YSbtmHo+9NMeL9+7x01gLux7NMF
ZlBY41gVRcFZjDTAAG3I+3r0LO3cFpjpDKA3FbDKZ41NYIb6tzs8bINI0jF5zRo2+5mSJTo9p5Q9
V8EQzXuccNJJqCIWF+rhjnRURkytKSqDXeXtdksI+h0Oni7gpL53p2ENmRCrJk6P9bIJWBMk9Wxy
xXOATRIoSPuRpcyzID51cjn7gVIV4l3RuUnaRlu1FtUWAlWGm2JnaD00LeeWnW5iWouscc6k6SSc
ANhzypB8YyGbWW9kiCqg+ODOj4dn/64ZehssfrHagGbKFSwR9aXBJtB3VSRck1LqRhQ7NBDx0e6O
0WvbJaC1+b2I8GYA9R8M+TL4CKIOAZR/l40KFWDJcegVV6ODcD4mnxdVL+AJJ6AWJvBKHBiUBqgD
UX4d7CJu1UkIZjkcbYrEPqtxpfg4f02DWroDVkyRrekdHUyWfwNOdwiy3YKFQGWhL7XMq3ZqxUQf
RMsWckM++4FCTNtN16Zgg8Udmj/nQ9m5jQTtLTeWUQveY+JhiI0gR/55ojvYKIhA64JUtgBktY/e
BPfIV25nxSDUGqjzMDN17Zl9J8xc3truR4M4v54DVF5DFHqxOcojjRXcPHDp2JLaWasFKp6rtCHF
lSb8GesNet++CdJNd6bmQhXeUMn0m69QYQTfBZyQN8UiDAtNOIGlMq39hH+Ybth6iX5s5hhzeBXW
rq+MdaGFOPne5VVLrUuoz43eM1DbnpjIR7ZjTNeTkWB2i3JZ3Qz4IV6+Zko3Wrpe/xrIuRVrTEVZ
u9KYGvkKMGEjGgzZEJIwQMl5pJY5wJ7tOplfD7/mf2suKuKHBEDVTnXc47MKfnhwAiPp1y3mY/6o
+O/BUgUHxoGjL8AQXXbVBhRoZns/kGXyOjaEfgAzgTshgTexKhAOppFCtNMYc3nsei/m/HnMpV/a
GDJzy1xBCiZNV2aCWtexU910uBRBTtwCeXrKUtKSPvcK75BSCTI0f4UYM+rsHnr52BCHLy4s22bw
RgSoUz2AShCUzMwQLfin0sysutLUFdM0EnkAqdYXSLD+EqFwq1ayyyfPAfVDv9yoLL03Ic4Qd1se
IB9Svnzr2BkZxzLU/c8oTsRhoNRXoBsxOmALa5SL3uNa8irL/Bg2x9gIaGQ48JlLYx7KNw1AU521
Q3Qjj+aTFewEtvzk4aEeWFYue1LwyXiSEZaAIJkAJ6ghQYQvWbNZfgFDmvBLOgmeJSH0f4iX/06O
rXIzZrYj6rt//wutumq1SSMAm0YDQzNxm0i1DXEyhoerh4tkoEtGtrOWhTl5S/McVVPamREO1oxQ
u3U2UI20zun1ovl7Gpcb5af+DQo8ObReUxzsxEDbCKf08Yn4D6/eX7jvXC4HyyAqI/0WjxNhe6RM
sQr2CphXvRU2nwre+YaOPY+iPc1ZhuyDKWjiJp5mIKuKD4ViRJIsPfFceu06dPGFq8iRUAz8AyH0
nevGgvvGdPRMu24jiDszO5kGwUCSgw6xIoXhrThgwWOe3vKjinMKbzQRr7FWgFRWzKBrNZjSq1cE
JjVCkFlJErPwH4occ+qJDeBSVCdRWoc7Y+jG6u4OBZQlHUrFsGsGhi5Oq+W+grMb6bWTHzSqhXEz
RGQbix4BV5XwJ9qy638mw3rwPgD4PR8znvNgnpwAUi18IRjrpUKeysR7PXLiH1XMfvdp0hvHECg1
drl2V0Dpuhcbrd31pp8GVR6iGsyUIrjgEZvv+tpUruIFveiYfiw8k91Xxcd3ce/YBrFMB5CY+E1V
ZK/GHEynZl1kafc5Svhk1tEnMh4mjlUOfWh1ZGYMWv/3blR34WsGDMUn8sUHrgKtse7zId3ZRZO8
LA7YxS++Um678nrzLxFGLPcAS/JZj1A9qXc+vm0FrFj6G3yQTSQaY/Dq2nDhw/oMX6yx0qt7lRw7
+wvJ/JI1bjO42L0NvcnGRCdlcBxMOoKy3rls8UGt+ThYxXb6OcTAI2ISU3WkMCM/4gD4NohUlJBv
CeSDd7gqjnpsIzzNl2IkhPvoc7vrQMLLfv3zL9H9K6RAUP+SfFmvdSMS+0sJsjwFZ3E/vSETiEIk
tLyjbPWvP9ES2ixnBQyKQOjuyXRhTOlTVZUU5aybzDqSz1XSAlg/RS8E+i5mczhRSlS9yNi0Yz76
PrD7UaoelqHVpnc4aAxwhsYI+OQl4xIdVKV0oh/LBG1AEQrXvbkqCKsp3LI61wKQdfJNQKOw6wiQ
KXycRz0w4fmWGCvbR7MHL51R9i4n4iUIjuOlwqi1MbveThK1AOOQ9Vi5x08Kvqe2IaMMDDsWsAhm
LsoKVmwZAd1XkrQM0wZOPA9sGZ9GtxXGlh+WWrFWh7Yo4ZFp2VdTlPdtyY3JAc/vYVxkaPg7OgUi
O4bIseYhsvos0PlP4hs7fHyowBZBkmPXxs9px3RGml/SSLyEWP4AA+6db/DGenjYADwIGouiJrBD
Fc4WYhC8WY8zq4spBVGWYBjL/x+n1bQwtRDWeibVl/LFqtVouY6FAzgeqAYOXO3oSzd+bGZQPjFD
qQvEq9aYuqVHOwSxyCBS4YWK7IDFlxb4QHdI1CO3yUouhdS4+RAmlkax3OUzES4Wx5Znq0wXg2w8
GhqEZXFvlNgK+CiDuaBG9AkIghGO3wBbJLauPTdlGhSMM6wDL2LNwiTB+4lO+hY65nVQopaMMN/7
AWNJ78P+UxVGAWI321vYWseE27UNnw/JQyTVIiGHnpeqoTTfP2B59qImoOhdYZ0uCxTHELIKO8oL
2nnfOeeUa/0RqD6YT81M2lRQ5eo4N7sz1gESMyCbmyFFP5/wJNs5ez5yj4e2oJYmy98J+iRO9MuZ
tuArWm+CsdsGDJncx/dFLqBK9zhmh9MDTiZDZSkzpJSdrdf0b9DMCWjKNRU1B95ocpg5jm6vuqPQ
fOMQrT9TN4WptYF6IdN/hkHuP9OYhxBZYORYWTI5GAotcGTlc8shyGk8PGMlxvfa5ajobXr2oqM2
CfBS+V3xu3HIqkrblLTg/qCVLf23UofPm4MOtOyDenWhp400ZCnbcueSDAasbOZeYp5ZcnuZG0Hh
a1ECXAp49lTNB7gRfpi5aHRz0ZZ0pQVSpBQ3eUORGitDmnvgdiXu+8kVvX2lMDcnnGTJ73gwQIPW
V71EwozFcDMPrhvm6iEUkC2czYZfttflFZ9BemnQNWlBbl698D9ILoWYPtQXhI+ds84wb2Y4bSVl
2XJOmRf9UB8jWvOOqndp60/gZennUEbNrebKt3GUVFmAoae0c9PIF6Xea4ih6/McnToJgSf5n9IH
h3QdcLv0QEZzQDBryAnmBE7YHt6HWflIgibG8j68uS+7NA6BDS6LenCwBbFstSSlO8E42KfjG8+C
x6sFFyRDDoYi9CF/Om32gzjDSrkcfMF5GI6yQxJdbsF4jC+qRNrTIFRfuLjadcxgZY0pacntP9tB
b0t/Dw1Wm2Jw1Eo5vpI0ZsvPlD9Nq8s0TZGbnKiDwxtgv9rjvuRIguZMCCo5y439GhKiroJyz/gw
mPj7mRuqn9yjXMnYIEAp4o6ee7bHdEKklKpixUFfhGU2Q3Dgo99rfoxZvFdIVsGdxaXkU6WJ1aYe
EuoQXuWDbCGAHacc2lvwTBDC3gKWrTzGzrkn/wFk+l9hzx+AIoamXnANEpvnZhWjXqzbMGkwMAde
3NKi4mzu4TzimsxwVQKHBYkrW1Ew0OeUKZdpZsv1UhbpfO1kAegRRnUaf/FulEtFVxyQeX1eFQ7j
/r0tdmhlFb602bnpcMFRjdeFRtWQbD2ivrK8yW9RbhNOIex9ESsPxPm6iRgZ1VL9KqtREVBDWsJn
huHdlHk082EpIP6rGcwU56NPQBVnxGcNTUAz0phisfubBidIZZxOyix0Xxiv3ukUDNsDIoNDElYi
CPceqfIaamW+9MiERtB90WRJOcHw9PsnOh29RE7HwAbPNvzLjJJdscwTOk256pgARGwLmyPaNrsl
+/IJvhkzPKthDUn6717jhCJhUD7fcO8wruWovTxaAtArB757sHGN0Yp2QFKyZs53bnyIDcsiCY2D
eU+5rpQm//C/nrojZ2XXVFwS5heW4RRO3GqhbApTMJpA1YnrJbFVjBx4pUzLLNSmN3zk9QNoA1Cy
M1mIVzG8b/fmGgX03fZUAjAUE+stjcpvp/8wBzlzK/Q2PTosdaDD23j9FoOZjCy5pmeNtGMv5gvq
gdRwN61Zv7+B4R8jGAzMm2MgP8LZmoYKAyIlIlOQjdyZgbF4tlLfNsjCHLq2YwJocJNgL0YgC6NH
jR9sn6Luy8li23Igz7TZb1gJh9wzob5VR39S2WAL4l+vwAWNjnxJlbYG5tI7F12P3I4sdG4Oi2uN
0RnVQb7OMIKAZyg4Z2qe4Xz9DcJ8NmsOAN+KBaep1n/n5O0592SJ05xSsRDnRU7Xu3iApx3pDLaU
3pYTkDgp0JdkMcGNVWylwoNI+TAh/h8w9/Q55oXEbXg6viUAAGTNOYggY7XmQVMrA5iOTUmThFVQ
NcC26XddjkxtUL/6hminCx7CoGR7Y3CkUwITt8tMxm87qvADqbOuAjitumEndPaeNoAaHbbZF8P9
C9pHEs2x0U//RT18b8uIHWoBV1RMNJi5VUlNmPjhr2HdjW7xJvfHCd6v+gfuGfRHg8OVlWqZYSDg
BivvxJaDd0mUT+joVTcn5pIpP3yBLy9Kbe/hE7DwINvLwwiznFD+F2V/fidUsRa4jqTsOjvQxROJ
a4N9A2GkIHg5lm2krQCuYLd5sn0hKOe9ryi6SV2/hYuCNoKUWDzrOO1Rz/QCHBamU765JjDYJ+un
avAwRB51ScX5XAo7XgQS5f6YOe2EQ5Ph+yMZFOYLbtoYJdMQieBU+jwApiZbfg3FetZIxgwT3n70
jrVYVcsLVIzaryxwCcFLUv5WkGoep6ZEvDoM8/5T7sjRpHvncuFFou+T28Rt2vSbNaWAiz9+O1pj
U63wyVuGacjt9oomK7secGD539MKixiVQ1HnJNBSlXOCxIrGs1QcJP6V5YPOLM1gVTy0MWh5gDjB
lG1s9hgXqnvw9t4HTIaCdIG3pHz+U03QnQ3e7Mn7z37dQ3Ew1GpOO3hykqlP5whHD0J6RKi1Ucgu
RY/FicNzeIsVR6+a2iYMTjYalTS4+5Asl8MEwxyA/958bQN3wJFvkIxeQVKwx7s4jJwW9RmlLU72
ExBlZuXWYV3FizyYK9cUv35SQGbgZ+DeX/7LcQ+CLi8WFMxyg8imKKn92HI1d7V0DGaS3ywU4fhR
BPLX23cJNyORDBFdg9OO7zQqbBZa9EVg0LnnASLVLz47bJnfFl3aRD8Xa0sqYohvOG5Et0uOqbO2
dkjNzdOYxg8RG0gi0kUy1V/q4fcFON8XU5fob5S9rWaKN8IeERqAnZK+p2IzTDikBK57Z5Km6hAL
+HgvW6AOS+3ltyBA1+n/b9EcwxEIHpQVUYpGw2oqFc4CJoggacMWWiIfVxDf9GftURFfa8I+TGU+
dB8cMJCw4Rb6YcBv/VcBCbElbNXBAf+JP1iENIAawZZ/TXgP+tPrJb0Uhnw+m/8pGENlZEv3d8r6
beJHwb24zhMsk+RD3OCyx0r7O3wU6974sJsSHbHJy5J9YpyXbfsPB7ycOdnsUCxzegAAxtmZ9AQO
LgAmRA+WyXq+uhn0IF8S9ftxE4pJwm99CSFU/lsbMFoJmB4zmSTw5Vh+J16JXFkfQ00MhBBo8Dv4
XzWn+eeWA5h2vkupRr/RLZ1G5RKEeZD3DTfPBgiAyV4DamvpCETySIkCVoJOKNWkzMxRLrTQbr4i
wtk/YC6rTrZlsXPhMYk28jetDwPpA6lH/BMx+bF37HuQam0dGnI8NAureMTwuvZ0IG5NXgKJqKwC
bvJ1QY/3B6FIBGzCj8foAPD4FboejZQd34NcqFDoW/BdRm5Ak5R8uBC+HII4V6SBYjIj2bJaKnxl
pDt9CgnSOHJlaCXlxEIhXzRsaUe1kDjvINPmcagorNOikpjmqbknazsl5DM9oOTf2DlFcZiI1omQ
qmk55g1iL331BBt+xfJi8qQNj/lKozcKWPJZ6gliXqi9/Cn4HUb6kD1BAnQaCoyea1rgIlYzicd+
2fA48W7TS+rXvzWaEPBLWEyvjWXARYSU4PKigX+HWmUMkyRwhvQ6fcrkBTW5TTmFkdPYyTY5ZAaE
QDaOFFDsXcGFBQkrqY7xcaOJpyt+LYKCKStg82PGESOAYn4WUUTknqD21EoUHVFdWZMYvjhejRV9
vrmF7oizlEpG7DRzrAPB7nBujW5lCtHq/7/4br7+hyDWGnQpdKviCkf8cbh4mZkFjR1LLRYGhHSa
TMNOY3dCFrgcA0tCQ7zNIwIfJGxJxiODJ+n+f5bYM8olSU4ctGa/M7YJjm2ie1Q+1xrl933VhRz9
T21oeV1t2O6ERPJjC3HaSLLgAp6s/nGwjDHqEXHK3apfvjzvLNih+aWzAGBgjHwXtwLfZe/XOaVY
TVyXwHM0c8mdVL9lN48Zx11RPEVEiJB6Q9EmkHAiIs/sS9x/7er5XLOtW6FX4pIZ8tCk0qpZZQ9V
Eh3NwAJRP2Sre9+1zw3owVkqlGzYeQWNPzo6jJazfLGHTySWm8Y2Y8sBoNvv8vzkpK/dcpjLqJKH
E0iyYZFUC/FI/bHHUf7/w9Nk12q1VnTvKIEkvZDU9+Oxs+VhS01SUQzro9351i/PFaHu4xqUdv9E
qkbJ62TpgnWloJkkViGHF4XnxNlvOUTSstL+JYvj0Ys59ftF1HJIWNXVw6lR8s1iyQnOoSxq/MaM
UKVw+D16SZXFiShAqt3/UMX9DTsJwrZO/heUbHez511ilFieT7jPnYbzcCiHCUGDYtIQvPNvOe7z
YE2lEdFGVRpsx2trxKUD5ACZniOUPbc08eGUB2oGOwUVeqbpSmybFzPgIe0yvg/pD+Yn89IBCK5e
lTbf3NTh3OYwYCqvPIZarn9NllFtIpHxtJlt3RMViDNfbZw1GqhjLLGJSd0scpncfMi0a0fns3gm
T+HJbzRv9zM7bHR6oiDpxORxKUsrKpdpeQyP4nFFh5ZMBzYkIDmPykm6qZz7fh2hPubQI9L3Olyb
CwGWSKgY6G2FtetLBFRSvQ3xr7vniX5oEXqMkd7o2/w9SQK1eEY3cu+bCeLzlkq6PCa2u2e87URX
MoalETSg6n7TCfawxcjI9NKn7ouLYPpQ3Zt+h3QAVnGdq26VI6PmetUVK7DR9pCL0xwdbrKrLnmF
CbVuwuS0WJYGynMm1+fwo3s/wfd8jxZqDKQqzCM8eWOpofvhzer9+AMrOAPIr2RTUkQP21BcC6HP
1bxpERIIDCBmTx0IOOioOfLoeomqG4X3bzNULOUF3Y/5F+jjHBJX2zjdJMqbeCXlKm9OhwAiUd8Y
Itb/QqSvLVG3rNEn1D3nm+JMxESv+ys17h5c/pCBi9bY4HjKZYee1rly7riFOl+cvOEglvc6xhDy
dJDQ7myad8firjiwHzEQOgp5T8m/ObV1ntfwUFL4MR3SY9Dh2kX0LiA3HBQR2LDHut2xnZLF1WDg
Qi5LswfwVklrDNKwIk4pd8BHZswev7t6bmYpEn/a0cn3xfi4OKHRshTC1rGS48aYzhQGsE30JGOL
uQI8FRa6eHtb5HlGl3KPu3FJCm849a4FJQLJ9KIMSuag3lP3pszjfkkH3Ri45VWvyXrIcV9nJLhN
o5ojOxqfjW0eEw0TbPs5B/GdxVNF4Nuk7+dNcDiYnc8hRQKAJdm2dmXRdYlcoZs1+QQ8UqexYy+P
K1SbzCdeQiCcDQoLmk6SzNbp2Rikel1gHygWWHmlC4QNT5NQeqi113wGBbfJLS0cGVDLzbTAk7Yz
sKerI8Z6IJLF9N0yZR/o1mDUffiCCA5dEQ+Y9buCm7kI3PgXDArouLf8f7sV4dOqWaf0LgfPSlWm
Ua0fDTplILASfDAr8W9q5pz2xz4WeVANJ7U1U5/785orlBSPbHklPvWa/oCN4MagzfAeaxgCW7mi
jTK9TOLNqKsjrR0TViZEeWViBE5yi8mdJ8ODWCIgj+kzQoEAL7TcfVD+wzEeHt6ddJtHf9KtXT9E
Kgf79MdOfWPxqk2GOvwOfVhj6q+O82G1/tZqVwfXd8O7o1pdSmHZCXg5kQC/0u4gwKr/s+QUpb2l
Q9iGHk/C68X79RAda1LMWYKBoVUrVSwbZEnl3rsHPHD2rL01P87v6eJsUyyEw265SN72PUnwiR8M
JDPriSfYMjs0iinCQ6h6SuV7BFYyHY7D5Lc/tMv7bO+t2rjbZsVUzI5oQ1zSL6bcCL0y3UJqfeS0
yukOyav5EPsQDdbNcqCI1ROxm4O6UHxo7mwvKYjos7slNKSTtbRb4nxSuugkIjlwKDD9d3cLIQ0o
7gB5YcKMWnmImmGxVpRFcWTwdOqWhZIR+vJ7tiYJ40EBJm8z1AK+adRkE5ATYQZyJW9I3wigjx4r
9n4pEifD8z/RvakMBF1Yi5uZyciVgLfZ3pv+VMU48QXyY5JQea/MLSw7SQ8PvFlQ4+IpT02CQ91e
ImV3Iv89gOvik175h8kmwA/L7juNw9wHZ0n4J3Zq4ni1mLZ59ZxwjYTZeWvdNuSli4UwNbXFIv1+
5uncvFNh4cfp6Ju+VSmO+8K76fi/T864dEPyeM7OciKkrO8HZ7LKKIvXBa7pMLAb1rbe2kekwalf
JfiDR6SMGgtLMqImue/+SQuc9o2qyl7sK6VFbVRgl70gQ0TWRv/uwiJVvkXFRyM54NI4YP4jopn6
giLhs8xiFtiZImTt7tVCZd85TrANt3UKm8z2UOnMmOvkBOQbPALLMTdPSgtXTuzwMvymn5rasMZb
O61PH8X4dAxkDMGnKjECa093uan33609abzfHfs57nv7ZNaeV0n6TjwVhQLfv7EanMkFWlZT/jNw
o4vCd3ajDB675IcpLfzDdKQ5wpEfDkT4PZQJb/Z2/rnXntGzYrxLx/UakD9Lu7EGvj5Y5pi4I4O9
vMv/Tw3VxyE/bQWd1ff1m5mCfNVTkMAlSzs89SkZDbL6UPfMdbj5rzl44FQ1CttE/PIViqmgBdjj
v+dFa+eJnAt5ioI1nB1n+r7xEPIDshte78Z77Naj4thNNte+/ngQlXwIhLaJWLhqssv09d02ZA9H
Fz7QB271DIhUD4dE9mHjJhPTg3K1B23lZkIAz1izHDOI2lA+zME254as9lASfNI2NsEWcyyEUskL
x6pkEcq0Ljhiz2X/Pk0uQ8iTSvxzxR/63TVunVl4FuNxzH/K8L4RT/U2QFCjAAa+59BVeW8x8v8o
vqa2WOhdkfzDDPzh5u4ttAqhkA0Sy7O72EzNps0BfBt900vLkJEXkI29Cz8lcNUZgz5Q9TUmMIN2
fNxqzMRI9NRsMWUk5o5JpAStWMjPg6Qt816Km6LufXldgDzPCR2YjKM3zNkrmonKASmUV/Muqvj3
ImAi4AtO/p43BSlOAnvgLK7Oa754vP1opVtx1FzH2f7tXub1t/uJIycXhIJkMEqaQrbhQAMm7nmM
hcOtbT4DLgL2b5bAl1X6oooglIANC1v8MT3jKUezCVtZrba6Sv0kX5Y3RVqbEKZv1+yrNqFKETdZ
kk/pPKMaxIpH6/f98FJIl3FlJz8bFAVqLM4oNs/wmqUxFndxFrm63lb6QBdxI5lkgqMoY1thJzPU
LNP3HKMQwFBVW2C6gGQixz29MYNHRykGcGJ2K64bGVbADXpmpwcWboJRUOAQZaFmwtX3ykMuRARJ
5/5TzH7/mP7VXujR6Ipifpwe52RM2h0xEohH49KXH9yYHFIPCl5WQm1XSDXhOhj2m11mFJPHvJZj
adDJYVF7d2KTk6HBPpnj1DeQ3nRmXmlZ7q1Q2fl60jQ6m+fOE3oUWTrM75IpKUCFE95O9g9qvs1f
UcBQbEEJYA/NeCoa5CrgfSyPRoF2Kzbkzy865udRE1Jzp34YbwSe32fXAH1suTacmRLfVpY/oOuu
1RsFG9GB8JIHpF8sHfAQhTbL3vWrBXRVDb+gYoD1T8ubv4j/aXnQfwzPlFkwGXI3EBSgcc/dT8ia
AKPX/pPVstlf9cHhP/SMPis0nNlgc/JN3P03QxgKrH2VdTTZBlfvYpjCXA+SiglRXlMpWWz00pRX
8wz44+aLaQ2forset5aqORU15erXAeCUQUsNQKSffiVNngkhUrLYQfMMp7rdXgie6fAdPApTTWpS
lAhjUdUZUONxa9ZrnW6LwSgYGhiulCwUIdO6zyFvHS9LgL+Jz24PrN+oERFy+HdIFF1dNO4HMBdU
w1zdE9ozQTzfa77DBniBfLPm36HCM7tHor9eZceylbMaFO+FZNX9xr2QuHNXWOD8DiOJAbkQdT7l
D9xLsngp3/Qn7b/+HbyJZntC0Acb6JG6pw6CMEhB9XZ3Olbij/SgBro8j2gUmzCqsscEHGKSZf55
Re8aG/PdA4CvdpBmgld5xUDx+yNWTiw5GZhyZhTVIWEGCPny8EsXCm2emRITgXOPyIb+I03Etrgr
E5zOtB1G+hE6toAEFlz4uF7eTVFMfRNuDSmAh8Xi8Ru5RDbO9dfKDBm+RMBmJqkXDtXMB/xSEiic
n54Iu9o02G6xKpVnsDOmHzGDyg9JXrkNml4a4Me5353m72I3KjX8KJ7SFfS9ziO1DZ1rSiAmPz4x
c04S+L6xhba1FxvG/MJ1rKsD9x8WldLvPfGGD8LJ+yIT8bp33onExG0uQ4sQzKlGXp2LUwKsgyAm
HU1Gjccgua+DWNZJJys3NxMTINRE8LE4BsQ2KeAh9Se2c5QeSZfg1/s2+3NeK+iRSqlYwiMiUwjl
eL5BFBvRcqYWfKzMDs84r8JsDmC8+j1KJBmrbKXNZf3kmej7VHCrrSO8q+oLoWuEBumlTM5paFLd
spAY83GNmOXezlVUExYoGf6nZk12cOG/Vgpwh9kaS+Q35o4/x8ajJ8X5GvdP/zSA20Uc5t92YV7p
tW64s4xMmgLxF7bCzhCNST7drESS2EN+dIqc6iJ3ZtrLmb4maJ+CMViSNbXm00NQEqwyQJ2P+N7D
R7vzNCpSDbg+BocG0oaSBGhdxkP3mv8WTCU/WxOAQSD3iZgCtn1wE7J2PLiuAfaD5Ik1DpD/r6a5
wCjaqgjPaCU7ShQ6szeN5/z7xNCjnM5idHLRA4NHvW73rrx6fC9H2kdn7X3pMf/vDxGMFyiNxHda
L4fe6eR3N8vvwdQwsAITNsRnzKl4+sLSCzCHEOSrPmJuazO0f8BIF5Y++vJ7ymtZIEnx7XMSuRXL
2I6tpXyO2NuN2dOO08Fja8zP/of57oJwVBjWOpSQL0IlWfYDgcCV3n4cMGnzwV2PS77vX7hA/9pj
fzJRcpIlubb7s9UsoRaQ3LwG4BSm+YR7ljjX3eX4fGU2V5o4w4NbToLinR/wzyNIIuFAYlkfjlRu
7zAoQEMEkiircgG9sFYzmi2JhmXqVV3N1XLKVDmhujp3pb8LHyPQa+bfI/xWSd48cGS0TJfZTN/k
6QpGK8e5FtssDyPGGkHdwztvCewyE/Ac02VYKizMDXMn60rPdgkclITkANJwy60G4ZETCFkvjIgT
bAbC7Dp/83VpPdliL+Ph8q7CMepTiVPKaTG+7F8CmSYKTnm6gXpgJ5NktWjNlR8UVzzWAWJPCTz0
GglvwZre0IbsQZhsreJQLJhKC561yS4BBxsFzjAqOOwPZdyO3avdW4QdVJDEhArzed3gbRZL/5RP
f7ie/9JCF5XIczTamdkjfu6q3xRFxD42THRqAGRPnrh/uP8ta/KXzMyvg6HV4+OdvtbpymeDeSYM
KEckQpZiGOLOk1nQcM31zJYzk49WvBh9qEcgS2K1fb265ychzxsQL5rA+48mE2iknX2S8zrwbfn4
eAmuL3fWzKbooblzBhAtfIvI2ki2Os+DOfuNr4hgV6GbKtjItP2bBeOx8UXJAGfqPckgvgTUnsow
qmVgeMWQgwcHlVCFJVhKxaciWEdwABnlXsUa9lnG2I3trTwhlCy2r9p3/6OM1Oiujjt2p0MLvJYu
TdLbLkELJpsxZdfsdZsH5NURt3NVYJu8Cwhv1jlDyuncGQ+/ZFPIvuLzLrJLAszTr/Dcbn8UJcer
6vS4OeCU2s4xcnMlkd1a6JtgTcix2BkHagsTu506t+CH4dis6ToRpd+6VC2mmdxBhfRV675/dhde
kJLqOUU5j/Kyq07837t/hLRmmNlfFSp9H6cfZhJCbs+9XGdWbxZHaK6m6tHSlP9kq0vmXkpQ7Kc4
vTDJisObc0tbt1+m6TcPktj18d3bQ8o2Cn6/FOMzTumTCFHysgH56r7zoVssw+GJRy57XOgeYkPY
5ZTSqQQqLG+p8kcwLXWiIMeVYbYsooZFSE3A+E/SfT5CSpkAphdafC/cdN0DF/3PcgJF5A/brdm6
6C/hgD+UyqN6t4Hyg5F45WFF+WOqtklmergyVHDDsGLwhWFFxa99Hd80S9spQ5b+hqV1XpvrMwS3
InE6HTM5w29/bC2kxyFsjDQuDv6jegOcM7qRS/5KrESBO0hkndbSbea3dfAN5HCL8zk4tvyXwvB0
GsrKkL7YcB8ACDXBpMlE4TJsy/Jtqdwi1dhKnyZBC3ueDjjp3Pt2LjZBb1wGZ9YZCt69q9AgK8Kt
KFpDbB6DQEOO+h6YGw7c/S1R83XAjv4/Atk8frnH0YSo/7jRw6LpnlOSQP+aotHRvdT1iOFELTTD
qzh5lTJMofk8REXB3JgzLwSx2X5h/q89n6tJk5nOELWL/sDwCQfEGFpndKKAMgrBdx2hwVTQ4lms
wQ1Ef7HgNNJp2yEnBgFi+8pnNsRuNWn7g+w4jz7Q3uW1evyemeV03vWSoFC/vJWKZ5VqVzyYzbQn
Srm0S3VoFh52VBNoXbSWcznZEHR5bUUDi3+MERbcw2RJsyKOh05fjR1OQIuFEPI/E7TtgCa7zCTp
u4cwAOjWL9NA4TeoD8p9s5x6DqLpsGwPwIu7waLuKxGI5HmqovOvqcbFJupMn1QAnLan/bOgxRCF
G3oWKwghSCxylSYPbQR1sNLMN2U1RhjNmzW+CicnccCNG1o8EZP6q1ybs0BPhoc/NWUxUWBbsRXg
5iCdQTmn0hJuJVxthTpNQ39nQt6VITTYddIUqKtaXOZbp7FpcgQCmC7DfmbItTdYlNjtXou7B3FQ
9hmY2nUqeWPpto2nKLbF4JKMnVVfZt0xL1Vm08Jfs1i35ZPgRbBUQhTiT9LEm6SIiCSxl0pWRlik
6UdcdLSqR1kU0qkCQOcI5dpxaNci/2xkxlepM8pcIGGYqi4+e3Q87h16UqlEYAgtewM2dol9AqDA
rNZRACl/qv5mmpG5XPxVf0WF0Tg65LByw0puNlYuxlTfrU3duozCGF2JTURygosGWQdmK0LQybja
A22uIfezwKik9Rr0Ctimeh3SrUEJ8iT01PKup2Cw9Aok17+RjACcs6ojr29DuuK2MEcgM3tRE+1F
gWpnmkjXjC1jDv6Rq0f4PJHpmSsvkO5NOyIgze04eitebeUMmbtx7ZeanDA0frrSvMYbVEIffTkm
NE6byyIuVgRG13VuamMyMVgKg2vLejPcQ7KnDVL+IJk4OX769lSokHCB2qo0huseC2omwtJAVAD8
+ZZJMpkXHIT8gCPAc3EBclpUehMIHN2fxXyiCQnTdrhIltAcIg3uINEZH+ukn7WYYGZ8UwxSPgdU
ei6DaqTNmvg27qNq69/Ee9MPMNDuYxfHlCcx+tnyhZ1NYVQBv9EDi0bDXdJDqmac6aDcxLoQLdTC
bfvOKvUCVjfE2yLLWQe2psan7FhrhikpZdMrYy51RcHaFzif3TBF67FlZOLe/Q3Z8i45hwJKlzi4
2kcMqlOXBh7wHOh8TsMa1TuABkaw1A3gLEucfQOgfw03R3d1tNUrYcMYumoRdurUGMI08YF4igHj
H+s+cCc8yMEnzzUFzoAMtLjoZl4WrAcxLX1M4vDcT5GdJsZ65IScQR4uMc/avN45Vo4Cx+GE976R
kGXXZfxPwVFTb541fseY+CDm2d0fgoJI9WuoK+x3lVv3greE29fEALK7b9Ab0GoryqRuP+LXwGQA
at6xRwqSO/NnWKqFz8NxzcMmHG8+qscLZPtBEvSY7aPM60C6P8AyBWuy/bb//8pPstqTi2cO9Q31
U5FUjItZcxv5mNTgPMhm8Cy9EYLBWsgQxeJ20dPGV5n8pv6gZjX6sIg8omj5zsmyeXlJNta5Oyyi
1orANkUd/qL5nOBCQxw8tputbjmYlorDfVY485nUOZRZr6tNvi+fmhqqsMXc9ExMAR7+DKWCoFSs
gn9dRISwJVbJDRE4IQTwwHobWQZu2UtxIiSawH1qVd9nM7V4OmDcLzYjpDpW7n1SJoKa5/mbuqVW
83/85giEdfvoFWJSp+ou1LXBkX3hhqK4DA7dXMImaNguwCTwEWM/kVQt4FisrHRZiTPcgX0qDW8t
/jj0/t2eLZq2LD+fwhimQRjzhMEYE6Fx6pGH3V3nKr3XSVJjlwws42RXrTsvef2TY0gBe9hf/iJC
5yKJSID/KrPjq89AVwwPtVXXjbwhwrXuplYoxlGqBK8m20+g3CxEnC/17RhAvX5DgxeTnWWbCDBO
1ONAj9dw3F+LqO8QfU5b+iV9XYmBwAeSGdSHxGL/UTLF4IJ2WSY+VoeXJ8V9dhkUW4Bt1NNePnK9
8fMO9g1VJbFaRxR0HQ6HmcVEhwXUsZf1y9w2Lv+eeiCxDB3pY+0/pqiTFsLwd0HYEVPgcV2HmFRR
ftcIcFddVGBsb5UwHxBnR2IJxumHe05YzWPiCYaRrPqEBeUyftXx9hgpkGRsQk0FVo586g7pEWGr
Z0D/9nJf40bj4owyZs8v/JZFN60OxzWpysgGmk51x7rWktnOdRa2vkK9PjYueDkrQYECxLrgNX0/
yrD+2+gX5yPRs3NXv7pcZf76vpEjYT1uD0kw5s+K7CxmBvpFkAliXkO4E0NLtGTq1iZwikhhGjeR
fYma4dKV2NyUd9sukbUG/Jn1u2zpXx7TyGAqhVFjd0dXU2xGk5bOwKyMeXV6v1Aja4rcI9uX/7AX
h4pU3mqtwc6Qc2f85w+jyH0tCIbVclpeO2ExJCE+HX8CeX7yKxgubNazHGgH/dLh7sJ2Yb3ylOhF
nRvmvzFwyjWRWiZU3Pb81SrtcNUTyI7iulnE6uGT7xQidtctKe+5BLaXfFIstCxElMfZGR1es/ER
MYOoldQT6fG+FGldHSUnkR8ipT/STuXR4rICCVyvFBmAHL/WDbZ/hqNEnxDQbeV3Q/yZ/soLp8y9
gP0Wd4Qr6aYUMBpRPNRi6oIpfkvbGhBHG9Qol18UYo3jaR/7zH3DwpucoAU6MBqm7f7TDfoQLBDJ
TSrVwzdRVdQgSAPO8oz53sgvPvVQ8GwT7oVHvaQ3dljCydbAsCGPLbrXeVsjuLBwVQmfwLBuh0X1
W4aDDnY/78olZTJeUzAMShtR0TDNr5vbDc/QYiV7xuFO3usPUxhkaTW/hqnkDStwG4J9q7/8cUHg
rsH4IbnA58hxeR0cmyw99NvMjjyT0daCpfXtLIcin4rxqv/DLsqlNkdCEii6Oj4bvS+Nhne+rIUY
wlj/XLllSw/s8+dfUgYIM/Wi63AKU7Ow3KboBirlc2DAD1y1HmTO3BHpxJsqnAs1mhGqf5WTGf5c
+TI0s/aqskJO4uz2/CV+u9A91sM7QbI0/dMktq3mGwGO0bXV/torC/A/1ByCMZyA6BYYRiXc0fvV
aPBRvuwWAU7WGYYPMYt+kxnxGin1ZPYcQeuB7r2PZZE+1DylHgCkqGbofGxCYAODHAeyHpJ18NYo
r1T0t/NjjpvrG5taWee7hQsLDsGVl6OEy1pVUcJNjuNGg25G7zaYrB/8CUmoYB9FpzJ9536PQXDi
AngFO/paGKDFCfuHXD0OH0vn+cPk3xqa6e5zF5OS5eT4mu8tIhTuBudizcLgnzHZ/0AEj7AUmNZx
306ScnA+nNszjvotjfTj1F1wsICAjBsuLNoRTBKwJ5K4slN19u3s7AxYt0+umrclmOxw4YoF6u5h
TdJqOiShEb41/Yt6msIX7PW3TUqbQjTaMYEw/mD4gXl6tLzlTFpPWQR/oTS56wWHHG1QCKBgdzKS
pz/yCPDmOiXlummN3n8rzg25QBE2YagZUj0qLDoqW+s8pod+ZX57vgfExbROiE0PMsEdDKbrHkDE
Yf7uVJNepYef41XUDVGD7b3219iEvY8YkjIvOk95A/nTYAtAFzWZYg7GMwd2BqjWWU8uJNPlZr6K
XLxtwRugVdIMbFlhwBLkVlwzJ4cv++yqNL835Tyj5YEznQkFwvKmJfinJ9vLuPKrSnTUDn89WgUn
t+vg4OBrY8WK6YQSjYu5/0wC4vf7vzaUuigBk7wkIITq3VEinWdu1YCBy2RFIeo+se8SX6Zd8ewZ
+9F5liJDU6ICyLb7dXXPEq94ugWXUJyDIt0byXOMXInIbtfgAQnAbdNXoIByXeZbUcXZwhctJxZ7
U2/PCOC5TjAPMKLTSUzJR8ZAAApWfgW4FlSwRDl/Q+HtVz3ALvvON5AzxVITkERHNy5SXRIjonnQ
HB6HCm8P2PiWoRZ8lfxr1LLnXbVpWIXxx+JJZtu/45Tbsxsl8im5c8zHC4RtpW/Oax5R8ULSAgYb
EWnoj7mDu8MCPT96pEzFN9OR7sYpndeaDCOtfPAaRKH/qD+1pSWP60S7iqJlzrmZltYsJ+KgYHdG
8pY1XlasAL7qd8xRhSahzBfkEE0nNNorTKmhUSiXc9tdynvMONPkbjUx0JVb3+BxHZokMh96kA9W
mab3Gn3gKz2vCarfjwiTiPrNwxa3RxGHv5IFSyqGJTYq97oC84z+0sky794Ef9c362t097ttXPnh
tJ/Fw63srxztTgs8N6zt+ITnNUGJyA8gYwUKXZ7+IXJComVsXkyYOX7NUUaZwpOQ2FiBtsSr1nQq
wOxeNp5HKAzMOW518MCnTGiGDWbvNxLmTyBHYht0YSB1nL4pbVZcOqjgKpsHIHv2R76TTn1lx+Iu
XHXQ1pTqbmM/kxVmDTEzWvVK4S343xyQoY9c2Bivr0u2bLtYOuHF5xqst+p6RM5kmPsjv608etzK
V18BvWIfwrC9M+WxNY++NsCxWejeeTSExnOdZHHLYw7qCJXVU7NVj/MbgsEw3WuBPUK1W+viKenc
ZFfOhEaGpLqlE0K7ClC5iPDe0OwouR7zn+y4emJFRTRkKvDV/DlXRr+Qd2OLI5icr9ecNO4Gafcy
vZ8PjHWhF2fF7ahPFLRHDlBwns4Yd4TSpzCSgPqjR84w50TRjXzbIdHvxHqAb0sKls8JBgpIrkqs
AWQhL1JnX6b4tuqMxsXak38a/IlMO8D2QrOZ+dDp00yY88Mohw94Ak4yJT9UdGK1TyffoPH/Rgtr
8vXC6TlVtjYvMAwRYj+K9no0ihkyjv2GoUpYcRziGIl+hbTeo+leJ9quSA4nrk25x9OFslKyFneg
kIqpf9+cR8sG3KpjHSz8vjm8H6UnkfJB1HmNahiZymfve8+x+bPpjKDcAkCozE3A96m0Y/UoXpRe
dgdNL3ViFYelczmnEzIhRs1qrcbcxKA+T0dcgPy9J342VNaigThrpYf1uXD0YPrX3Mz9WcTbM8fo
J6Xb7sXlFxESxWnFbGvtUEtb4MWWA+lO8oA/jDlBpFvUS2jlHd9Ke86p66wgKmPuxXZuKDZD/1RQ
J+54bVtDIsGgn2fZDzIkKS2Cre1DSdOo7z28jnU78ZSbTRbvSWhQw2WbYAg5cgcmG24u8Y0yGfQO
nIjMBkiGc1nRbukFv8Ko+0AqBiLy34FkLonZl9Ff/eQD4bD65YOZrzG8/DqcjNhoaUYx3aV0PtZM
um/rT9X6Ahy4upDPco+XisyDiAXO/s370qy1Ctb4gVAbKYVncV0VpoQDSP2stPKDLOQEdZdKlFmE
srITJkkxuRTfpAQG4UgoRQ+u6oV5y5YPPFT+mcqCdf7MDairOKUWpqML9pjXCg0ewMQj7vRsdskt
ZrO7SRtt17goQoulGs65Cx93bpnXI9qzH1gf7npjB3q0UEyFRZCRvZHsUTD2kVUvm2CWsFEwP8Dk
CKq2zUGPf7FaDNQlE6+mCQpmbZsWmOKG1VY7nwnaNs5V28BGBjI9WVI3peAoh3u64+iLMDp7veE4
Qhm/oO9/k8KHXflSz5uic9vWRlpKB4NqpY270re6SESCxrjHc4IqIShJs0w9Vc1BoxUpOwOzhpXG
yPMBYUG9GP5syfJhk3R05VA+5FGn7uJ91HyZlwGZYJ7X5vMa/K0wa4keeCdjRc0x/SzkzciKvZ7S
Hu+t1vARN9FGElhucPBs6uneQAeO85oVmAS5aobwHcp5V4HkC9Kde49qHXxKsnm8oynY7T0anL1D
M2pLRsJiMBJ1ET1+b6tSNYKfZfD4UqWbpX5ZGUEXbbUOiKjd2yqFhihToDZuhH7G/izCqfLZ26wg
2nfnRwpR9z1wtQTpeH5wdKZNtkS2mAZHb62Kpt/RY5W94h/nD2+MqilmXxgj6sBBRw+VNqLEeX/U
gboofTN0/GsuDAwXK/7ZkkjfCIzgCEjZYCXe3kWx2FcmJV2gD0qAaugQ91PTbM3rXUSx8gArstvj
BUGdY1uy3wN4Yvg+fUie0JtC7vU1EpzURtdQVqZAgdnjIjLFQDy6llP77tS5TX+/xe4HaElB0g43
v1Ul512pWFbYoUY7NhoPHCCBaRkr66j9nslVgT2dD2XA8iAGg9DVjHKEZhNdpEozzS6UmvOc3yTt
JIvlpa22AzQrseUg8hWJgOXA5slZbLnqLJkhcAZ+o8aLQhaHBrKjg0ewtv8z6K4Yj44jUDd5TAy5
H7Tx3XZZcTxdI+PQeQnh34kplv90NRsFqj42aZzLx961QJh1hLFP4gH1T7mXkTWK56vaV+dRxgK3
y8sHa62tWZHIYtVPwNU5RZTN5Z9uVvrupj7g3eIVHyBInGLuWzF9eoAIR0cAunriX9Y4JZ/i5DuF
P2wM0e4Q/TKGP1LwtUGL4oSMn01u5ZGWCOdu8yls84xkdEzA5G4jz1VxgDt8YyAZQc+Fux4u7h4r
7Za6DBQ4+rzQoURlZSqr8zhyTGRhwP7sp1p+rVly9k5cUtsYWOT+ybzdOgUerQ5A0AEpt6V/Lv+G
VBGZpb0ioQDLHLA1ngcIZrYEeuo+D1UXTSHImtInbyDUwiTIGe/A+2H+YcVGYUb8Dky0xchOu2BJ
QB4e4P98rOBKCgcJOzeuExQDV+Lf4ClfGscoyzDf7z1cqKZ6r8tJwg1foArEyPJL488X1HGGlUgt
N13sodwc0fO4JwIhVR8uI/OBGoVVq09aFH8UU/NCh9OQ0UXKTehKEK9WQ7EqXfGF9pB9M6CWNtKM
igOIttJfeEdIQSx1FtmnWlpJ/7j2Z6xysGyT9N/LT6ta1+zIko+SQ7dOJoD6YP3o847mNmPGdHGw
S+FxlLacWYvG3dOJjdVOS7QrvtfF9RyPofMhdvTJdhT/tk7BFNwaMuVx3kSSkEZacj3g+b3yquAR
+bz5G/XzqDAv2jSYtyY8RG6JlmoUO23L9dkLQODM9IIAlw73F2yJ2VVPCroxaknDEzMjagwWjqa+
iWT539cO5tqxh4jYAgVzWZKFAk8HOZsYLlNm4oM4QB0QuIcgi3dGBHRPRSLEKrWoOXM49bI4aJiD
AvdX4AsNUbh9UgHc/slD8uXfSzmqGyBIMECEfaYQFFrt0awPVkxbmInsAf7a+UaKsE+OqpSiFwbT
CbnjPbaKCh4VPBSoWeDR3Ul64TXEZKmeRGK5JEj0Uhhu8J2rMXjbKI8ElHXkDKVk4qxmoBr4Ny7F
Svv+vZP5FEdhBnh+Yw79IeYjAkl/hr2Yqh0/xpZXw6fCzIZAQRmTb84uyHym2vDH0EKhsbQiYMhG
/Bvm+9koIJEtvEr6vEkwI8ioKK6aPoxxzyAdOIrNI/brIi40DvzcsVa9z/jsp+cndVb3x4raEhPe
GN82OZVcqLm/piCTZbQGXD/h+ALtUNE8G4X6omB/5N8UBNPzH10Jjxi7bH3uLP/zq+tCOpS/eJ2O
+HYh18hqMqwYHo85qIytIzt550jZovVpg9AH8L3RJxf/Kh7Q/lP2VReJa/+f2tTTIQhoLHgEQRTJ
OS6SZmkc+vp8iLTSorIFVN3UUKFiI3jvwLxo1E8Cq1LmPEIsiZiKhkLxVPktOW891zKmIVtoysCb
hTUtCNo7aJFXlGs+K/MdIuaMsX2Bkdpo8BCiRWBJCWsuG3bKSIxznrheAc9YKqUax9tncH3Q36kG
V+SWM5mh9vUk1gx6RMvHI2v6eKibGPAbds/qi5wA9R8jhA3BuuE4a5ANYNE77B0LgHEVn4h8++k3
obg9+fVChSrYIFXsBd1LOiBxL9nDT75Wa/8cPDP7fQlk6KyNL31/YG4mUBqNmUbW+tGGIuw+4gMB
FIfTzJYGIpsv/vGeZL+Q49Ktu9dJ5EUuhdW3BHnCqk5Ys5fgEOmEX2zqGjUfbuVJuvXHt7wSrPNh
jiXBrADFQABMits5E5Zs8BgDo93vck+GbVW69p/2Ds8ypuZOgERAH+0bm3GgdCYykRO7ZSjIeVHQ
ONEpO84QaujKWSiBpBdufT9RV2yK3XdHGQrhaOLpHG8iQ7bQ/rGD58SzSm49MwaoYqekBpmRJBds
5iEQicKPtbwGRUDW6BR1fxKEsSjLDFjuRRF3b/mboE2domCyACr79IxNe9V9uGCYwnaVGDRltgo3
x+qmuZqt24zvu+W19AgWh6/Tk97RaoJu5HnKZ33NG/q/cL7zSn6yx6ZFFPSAfrP/idP5pw+XknTy
Obo2vwWYLjNZN0jzeY5JIg9l8A6WGuD+O3XMiG0jVD4yJm70pfKEqP3V/XHxDY7serz43rubhpX5
VK9mdcYIE+NLboSYE9T1QcTeo6H1enW7gpyQygZ1n/VgKp45WHBtFIjVfMbtolQ0ZDGOc1l/0MQc
8/vuERBHd/6kuh1+krO0KCxgwi8OnwndRsOLvvjf2GXOB0VvGjFcjD3omETKRY8E9eOCBxDtzyh1
lmqS7wWOrfjvJyA27F+I50qIQBOkzJpubF15xsJvo5bGv4d9KafpgneetsHPNZVS/ZcIZyl0c+8X
Aj+y8NYJnYo8DiySiGaz9RX/YpNWhiiwnQ9cUie28xzT70Fvwa9lFaLyDUlyI7kcGPr0HDe/ckaB
8XtfUlpWBqElKhY4D6/fJzYd/+GU5oS+LAPRNC4FjlYpC40VnlRTAtsg19T7Faymj6Xf93oJiwaa
izU5QSw+fbEOyfIN+6o6hBTN30dYfCA1jrBIkbsjj3O3UNVWFmsLHjmxoG36rgwosyvoINbAu4k7
5QVRL1/wXmc85Tzt1Xrfi6oXp3tU+dwqt9Wd0CXhl/c1FmMhWxzhkHUDkXF4Dem7y+7Hf+v98+bj
WInCgynJX2fia4E08kpA1Kqu84ZwTK5b/amFF97fx1OKmozHN66EyFkYOyGRJPJdO+y9zWtQJRWn
t4qNwvMdRJ3KDsx/Z2WhcL5gQ4IaUMmEEio7SWjk29e7S9jb7BdvTe7ioLMwEOecoNaYny40tDYM
wAD4HHOVHF+jQMbrWP04GDEnk3Tr4ujLYGRTKkd+VbUWli0N4S88ujK0LjX7SNEx93E1pJF6cjsQ
qxG99McvocKxd+WhKxdCZQ8E9bIq1FC5yq88HMtcCf33+0/FEN0YA64M0RycgpERBwFnJAUndno0
6P+cKl7rmXaQVyHYmQgKe7hhyh3rtVUi0k7pbox/xB8HHWbnRFANWhJrKwJLTtG/i0kXm611t7z+
E7hLv8HJ55vEbxr5ll8erhOQ7DbhHojn328kLxhKNWIQ2Rj2JNXWIZ/msTzpAGuNwurnZFpRvMsa
NOFn/hViLiMfEEZbC696UPKyoN3ChKTxTJAMuhbhi1GAFJsrpqfJ5G3XDmppu8rLaA/DZsznszkS
FQwdRg8ijH9CKPpOT+3Vf7fDosxCQT7zeLeIGxdpotI/8ZOKo2eWY1IW96gBYME3FYCiVgP5IOUb
Q+eRJ9J9N5eMB5j93H86zYBCJXWkO6foPzMKbY6dSKFv5b2QZDxRLOVyyVhLulr54gNfIoqyJAY9
sSYLs8M0hC4G42zO5pNVof3aPSWu+gssasS5a/MQjO66H2rmA9SojnOjswmonJg6FOYGVQcvnsFx
bV7ee56O/rWsy+XMzN8HrJdmw8AFQiURwfXwDzo93S+aZxD9vUB805IJsZ9rnF5oUE1E43gOSJr7
rUd/hvbnYOYQ9TeaqhSRUSUqx1ETMRr84pLn/8MIjxRwp5YrHQTYF2FXlm48WVGISl7YEOCjNhQc
E7aGeuLNmsqI658Dv0psn5aqrxz/vLbDPFrjbliE9z5rwYJWW7xq+IjGbit9j0SGZXxT7X1CwzSM
jMH9MohOpg+t9za8JAnZppjDDrOBN8TWHlggNJctE7kP+xd2U9xIeO38P21VHvpZLrBDlbN4xVer
xhGv92xSupsCHEgTtU+5gTzDYfbMdmxaX6oOf7V6T52TIwxsSOX3G/guIiZBx8A6248V9dhKwsSK
hcyHLqzLAXZUsqmDLlzABqmDba5OtJOvNRV4C5pXxA2BIQFbqMPpv6xrTkFQRD00A1RxOHRUh6su
siEQX0dJufQ1zx5pGBObLVfbF0mHgx7PS702nzU8DtzhpEumoyM07f2A9uftCX81v+O+0hgI+I71
5Ip7ByP525iyzc4ZjhZAgU2/cyH5QAzzUafyjhdJhzCZskU4QOvcTc+FjYLfEh+oTKCGRG/KoNQO
/WJ7MKgtTiM/QB3TYrdlzjZ9zvoUKzkbJCCJlGBN5W5XFzMSKWt35Y3wVZ4r94zLsTjoKigFjcFT
7tUo7oIF/Pxc8De0AXrVI9tjyE4q2exQKc4MH32rO2Fvh4wVDfMClQNxWULmyQO3/BJs/C9HDKbc
KtRYgAu5kwBUyR2zVDH+/wk6BuSSWf1Dj+YkG/XgcMkXgf+9Y8yPvI8f3ar/m/Xo27koYnRUT5bj
yKcoLeB1M2efkmn4Bk3vpPJaVTkV3RzlbGsjAuMMrXLaDcaRYcxYCx3mQMcz+w0VdnYwG3cWyGBV
i3EL4jx4K0yaVl/wV4VfIvTG0XATSOzhyNnMFqRW/83PVhGV71xykXzNBNPKN5aToiybEBWguon6
uH0cEOJ9J1L+ICAHS1WcbPraq2Os9RfgWtlBUuOStGqitoqmxc1xFD2ixzLidnUejhNm4zmnuyEJ
5kq+xFcun1I9yWKIizAnDbxnkAneBlfU/Q7N4Pnh1KSdNarftsCRomgRbzUc1jm6cEeXZwcKPayT
+yvSxNqlLEVpGDoN/TxfMb8nnTM0kbZ2uz3pfMLKEwaVzpuCFhtaS8AVSXsqbmRX5KuCFU27501O
56VebhR9/cWYjoc3UuMd7T+OOiA9/y/DVucpzWPn2hPaiQ4a16EYOCGV2TaCFmrLf+hLXgushjE1
b2QSsPd1esSR6k5PraFhf3TgrwZD3ELfE7Hk/2R34gNYXfOl2ETLWeUym3HLjX5tlsM8KQpXLit1
Zcetwr8EJi0TMcnFPqx8xNRxNrZOLCFAKHDKLOC8VvFeFfLRvN6szChcE5cOe3SE5kjFAgJonmrY
3rVrW8ohxauVfs9jVM2Jr8FnKBEopEATkwK8P6kfb2+PBn/zQyVCjDMLFTcEPBI0D1X/AtDWk4VI
wN5bRhzfePq6W1/1/0YsPrTslVxpRFguQPhUcbVPalacMsrJxRIkIhgvMqpIfIYFCvvkJDctw4To
lnZGp+Ez68g/MomwqHku2wtg1Gh6ueZM2CEV9AVwQk7l6ejPCwsIYMxxYfTrncGCt5Zh1uwyAAU3
29qXDsW/Xt+HFM2htfZCA2qJUXrjBf4yIURRfLnw5UP8k3f0k76g9mgWPROpl9ebyIidyVmlE13Q
+v/Ed6mbbw+qd7q46eSVPAEBbzUBoTfgbFSnpYOwA8izPHbrkUCgrajhGSdieamzTCjZcvqYtEGZ
1HOjQ3ffiZECqF5yWw5vBViqufn04o+YFOytil/fi8h3ZBcQSahI0HrVxr1vDRistMo6g1v0EdX9
r9rjY/cPvMSfQbw+i+LhYr8FaTBTcdhBojqt5nWzDb277mzDtQOBxRt61Tp8rHFkf3/GHqfXCRAI
UaTZdhZ9GMxFq+OuOTp+UK+biRQk8S78+bcm0cK8TIuf66vT9aVZupSs9dE079o9+BQ0pM8lFC7x
ZujPXerlm3cvu0dQosmKGtZN0jhUd3DSVF07YYqdF/jViOKn/jTeikiJ4TAodkKKhkV+5uuS+Tho
5vv5SlRJG6iD2z1O1M3gAVxsPOlPnrWpXt9j3FTqXFBmech1x9OGynWpdWMFJag7zfrPiwHJRWDI
sVIactWmH0ZVeQr0SeKy3tDRhhSF0BqCNvpHy8QWanV/USS43nSynferob1hZet/ZU8Q1vJikZNP
+hBTVsPKPWmjak3NaIecM3Lwb7+yOzsXScoH6raruihprkO62WDb7wVL0WoPgs/VtfgvoW8Domq4
0UYTOnH7ITXY1emJb+KmsClKt0KRB6ZK0EqOTJ5nIZd51cCZ8bohZtULNTdbiQAESsMGVRWSZ6wj
8dZ8TxfBlcGp0sPe0PNM1tcFME8fAo1OkHr/kQzo/irryv+3SJ6tIIL167gb79XwNblPD+LlL5ZF
LbVeYneaGt/yxTwEKp+toTSQjSkIrKXI4Gcwq4kNp8Lhik/xBhYF2AuBbAG11eyatmA8BuAd0GPB
I7WIy1PzqcNh/XL5/lD3FxIa2c7Wgk+o9GzxHT+fXuRRGNaZ6Epk6XyBhc6Qb6dWob4FRNU1PXhw
9KX0yqUn6s5MXrIrEwmd9XaOgXm+TQufiRyNMFoau5R/s60MoKga1K7RVLeCEsFMdT8LAbW4aStc
mGrFLYmVFLzBKp169DDlFp0rmU8IHdMxpbA83e1M1Ybggj3aX5fNYBAwL/+gnvsMfztw8jLR3HjI
zQL0Xv2MmOu0xjuqpUQD0w8CpuO2wjI7Vu6l7hnQcudnT1VZEUj4Vqr6DY1eVFNxMflKA7bq7SZq
g9YiauIxN2E67iySjhcgzUw+pzPMi3HCFoSzC42TQpqpUb7CLhGo5Dn3Yxsbr7RDhK//gAEA8e47
rJEXEv7rwjrpuRO5tHOi2E6d39BFkAqnhuQbagah1rP9HVMepSLsUWDyHBUU+j81Cv7oduJ6csut
+RFEWvwTdApIxN9lxFdKqwoTI5mvTmtqsgjX7gVARwiAAy7MmJ6zY477HZ3Fz31PEAbBPY4ePg/j
jJEXe6y72NDjKEsuiA3vWVNooR/4A5TVAZo7eBCoipyWXcrBYSRXj/hkUvNhqwHFKMM9giF69czG
FiXCTArL7LnLE7k+1aCiwukSNXxdAS4JeEdGb8rXk4g5VhZhNDpKn38SKDssgI/uhDaBdD5c9m5W
cpTKNqWNcpRleVe4RtRdqctUA0ilAvCsaFGSrwEhIt+lCHKPZEf9mGCxlYxk3ClII1a7JZobEgcc
pBxlKlFvHUo8NRyRkcKXYtG40MugKm4OvIgZhqwCp43E3BmvQ0Dc9nOT8FjLr9tb/ChyhitzyhWA
5t1WyPDY3TTdLKbZLjh/Ybz6lSvqc1DY1BD/pWffNADVEt81zqgA2ALi4e69Xb8xuYIbOIdMq3Ii
xua9vZuCRM7+Y4YigPC+oQnR9hA4g6ChJV0XNxbzXi8vrY/+YiMhT+Ylz7dBxlhVfHELkrqlJyNP
QMuAHMJFWurUo+/YzpMx2zdC/+YENbbn5WyVrVLRR1kS+YlXrqRdpzhbFirqjCwkPiRNf5ZYv+bN
FKEp/YMfzQXuS4y89dvpl7mbPorSmG4eIiu0BkhVuQ2+sa3GJzO2d5owM7oli4a0h4xHpn3zR1WJ
fGwq39hzWr1Jn0CyCUqv6UA6wUnM6txZFr3fb+NRJt4RL1nhYKn6rVQZPLDNOsotBm5QLQIp0YgX
aeWwoCt3XVsWeJBNLtSb39dxSSPCDHxDSD0nF2TycL+Al0EsGbcax0miP3XUeR1r+ILbsAjfno+F
taE1Bh9QlAx1dIzuTSbQbYtI3k16bX+N5XmIxfD9SfALQEfEvcxk9sxPPs+z73dYphWgjx9oQEFj
QKBB+nMCmQ/289NRrfJ5BHBnRq9pXH8J9wbWJNNXM1xVB6RlK1YHeAzyGMKq+fb4pu3JfnFnS0FT
N1QiW34dKI0HXCrXxYwXBnC90uNSZWUstJqQvKPoqwpYOE8AYrVAwkJchBLL43Pu6tx6dPkpWTyF
FkBH3TQ1bE519OiD+IflsYMSUULQ/xfr+pC/tnR+uhDUvqQwCirV1xfA3Mp4OGy1KiL76xtFwExf
d14h5vlYBoOYe+FPafrYkcb1fdRl4sJVduJr9xsZwSsev5nGxHPBFXtR/6QpPjDPAUWrkn1lZkkI
DzlJJMirPkzihY2UbwqKtAwyfPLfvc0nHbdXVpyV+VWn4j52sGD42RvrHrwrdy+b4SJgHopTDato
0jCL6fl5gkTqyYIQ5bWoTEJPodvdopWOpLSqmAA0yTt7zWSdBjF/ICQcRBW7TXFJF+9O8/IQTYr6
/PbIY87fbarynAi2Ld/2K+8rlm/Cujj1hFDMhe98jOpalt6Ht6L1WMhyNkwQ4k05DgrG6dMVTVSI
5zs3P4WnTmgxI4KVFQlL0wXaj2TdOxLTOUQzP/cr/Hcf1SKnAsEEwwTbWEHEf9tm11FBxAPdYAvO
Q9ZuqyQOLm8MCKFIA5DG04I2uYymGIfhJ/njKrUsH4i9k+8OvXx0D3iTx1iOeF/lWtTr2OaJGsga
pMxVb6eSdiKzViDjN5nJuIntlxwoX+qWmBzxTG6SpK4w1d4PFR8dr0HGrff4PY3Gwez6xNgNFSjT
I36Fdgg5H9rKgaTbQSE33B7FMyLyjdQsAihO9JIMYYikXKL7NR9gB3Trf1Gp/wjkmIUrldyjk2nJ
NwzBFW3aUyM+6bORGoj83o66bf5K0D94phA6xtyFr1pkzMxqu1pBkpMjAjuQvv3KQnbhsWNB0uIa
su+smWgOOl7QpS8woYxpsrGMzZVzbk+8yKRF1PrdgacfCU0BnH75qw+ateQIy95R+o5IjPcRwaVW
Wftf9XeLHYwXe8HXJJoc72qsvBbFKIIJAlqaf95v2lnyuSuHEn4z5pf3u2cR41jLcnM0GLX45p3O
7YDeTk9RnztVzAGLCiQZcTxqyfG3joN/oXYegxZ0bjfuuOteFyBUq6lmN2EGhmgKH2Ql/Wqn28SO
xN6KpEUzF8BYMYt1gb7gDuFxP/ZAe+pYYTzotPEmfHkvcCn/bmgQ+qzBwPpmFs8unHvs4NXkjsag
DvuRJR/U7XTkYsaM5A9IU8pR3aXx6hPfjdVkmJwqeMK7BI2EgboUE1gm+n0WJ2SsMUq74WjIjo8l
guWnjH3QtV0fK8TLwSk4kgHfuppdsTgT/LaVsJFQzYYsmYnzwjmWDRE0y/PMBe2tMChP9oxEk80U
Z7WYkaPlWbNpYWxKL/om4twxXt0t3iD2vIuQJkHxgCNq70GvX7b5YvYJ/E9OTAJcVIHNbKUv4iT/
XrFn9IwoG5255eqBrsTCIUu/KpBMC/42AmlWEjle2osQmPLONc9/UZ4a+XaR6qx9xSQU9qDEgVTX
UOWFffLQAWy1+lu1BMukQBdtiFhLQsXSObLyBI+ENm/gJoa8eEZZuN7tDWNUmvz1FoJ0vg6OrNk/
TSQb/DU4sC+9Ca9ElhKMIQzCa5gKbg3db4En4AzP4eSEK37n/BFVnbaca5nPQkiS761SjzQZTwnj
0ICYVX4zRTQWkKfft/OhscXoXykCqbzVJwShbNtKszjqH8P+o7y7wJ7eyylbd+R5mOO3cN4gP0Lf
7lXgnmYA4otcEW5tXpsPTE8QTfh5cJerD92ROo0YVO6Wttp7thEnqCJeGup5r+QlZXhUkaFf/7fE
1DegP7kEllPe4QiFpXSUAicsm31RuL9BJQcoZvj5KqPFCoMFQPw+B79VRK4mctduHgv73/C4YZur
hAO2mobxp8aOOksC7ejvJn77xIlv2d1pswohpj2XCPCiSGf3HH2de0zFTYSJMMusq4wDuU5waZ/n
ATflo5yOJYkneo+HbRBr6iTVT5SHMfASD0AlDzQPmZWrfdmm2QVpCKe9PhMdyP4SrbFSG9xnrVWk
BxJfXxp6TSRNM8VqOrgM1dwCiRE+1rjdulEwdwzVwiXiXcqn/QEtjkAQXGaj/+ZCtwXYJasDvRIJ
E5qY9OtV+qLT1f3zMtR1iwGWMqV2HZLu5Y2omRWcMd8K7KwB9gFVKqTEL22tY9BjMu8fmKX0DNTN
hSIc8J2QG9Ldth+u0WrdAicrUnolQprVNrOB6T7rJUNcsOkrIu7rvfJ+wf2qyqj7YtdA287IX0DI
YIbMLDFxXkJbH2ixAQVD5odbND/NYqROGIMapKZafIMv+lZkxSp1meKfZI4eeYFNFR04fl81ISW5
FHw4wjSXaFvRkiuUYEJWPWVWj8DtLy5QyN+1f56F96xx5ZGGvjcTPoNfWJQ+O8qu8VfA9KlSTHzj
VGucnDq/8aTKKoTcrAgZDrA8yJdEUft/L9wWWKL6ym08nByJqt6qVoTY4D1zl7EtC8+84IDhN0t6
8aEDqW4sgWj+VerwY4xX0vngFy7UPJta3/Nohi9P+1UA85mlwNMnu9spKirKMGutmwxzoC5wwopu
OHaiTXwdHFbOcV0ZXcI0MZ15D29IT2n3g+j+UyMv+GqJP//MH7JnrAE1THktpydlQaTzeEp2RAP+
H6jlCy9qPB6m3y6oY3amOgt/DVId5MzG/ztW3gVLgYsfHZfZyaGxGcX2gbyUGT4V5Y+st57JMMM5
U1ve3uGm/qfrndpgNP3W7UrhE5kf01m8AcOWA1D8mkW/pN08//vWgCAN2Fi7zk96gzBqZcvzq+Go
Xm++wCxpRcGE7JGyRwQ7DcKM6cYa0O/LezyntKJVKe+4e5ysFtQDG247lJteVNPjPFmS2Bbcp1jI
F03kTK4X2ai4D1Qv5fjHU5DY6FfeZKs+La0i/6cxG7I7F2m5euGYXfIBuNLygmtixk710PLvNKd1
LcUZ+Zv6PCH5dI9XGFFYFuVd7pV0xWMl8LiIiwSHjpfsNZje4GS6vQ1pf8U3yQIv9Oie8SVxFTeL
JDkUUMwU1qGwdEHPfLSu9RBTxUvR5GW5Chls9DGt2aaJnS1FXnNiLE5qric/F9kWQKYEXS2V9Ie7
r9gi7vfRohnCnhfwHlIOQwORPzaqrKT//8gsI1hwmXUg51EaQrJhSnv2RD5q7Qteocb1BJugCM8f
NHSMDGsfrFdExamq+UMMn2pgdGjdGt0KZXXlEqz7Wxr88Lo8k9x1HA5CEiLaA6v1cfHVU2Zd2T5v
dPqOPftt9HbD31kqwfXtn2pCFGrhoZlj+UtDkLqOgD+wzL9Rjig3F6IK4nW9j0inTZhy0lZ93y3t
iSgKhZU6KV7OH+lvLNpt1kkGzlNc0mbEaL64yK/RNW2prwXSj6tmIKQIUm0anlANB/4mYpNhYpP+
xRAc1qhV8vc49N/OnLhrKaohCJhLM0P4mYAcj4VWff7/FR0rJFe/qUXiSeMYKXiiNLHRhm8sCENG
ZShOTp8SbU9He92bmv3dUW+w1/8mUuJl/dZZOA94+2CbEibwpr+NpZWxe0/4Y6jxpjM8TAK1S9UL
qsN6LE4yUpxxtHi3zAbDHT050+jVke9eiy6mkm8orjsN5f1guH5gRUvJ+DuFgGwXoceTwrACGIB/
EEyOfjl2KlwWKme6VtYfZ4R/d2J4i9dR6mt80rPVTxFJl4FHr/JkqCM0CDGycWtvr7lZBopGc9aH
2A3bkQwFnuaWCaokTCuCU6CUhpvguxk9j+7v/zxSGkYwoj0Ugbi6rgc9AKV0aW1HsCL/Aa74V5i4
X2Xye6KHZbx3pv2keskYsX32YqfVJOBZiPa+l8VqJRcna4KCtbkfcCPKPdRLFXC18r+XlHNFXect
Gvm/MYHG/ZlRGQ515nRyMSc7ecowfI0np7gQ03sN7qO/zt9LE80B9pgiake4Tjjs66SkcKBlsewS
e8R41UlaY/Tc4vNesXq7VxfWpXYKviXP6YnYC8M8tHkipc+2A4ebdJi5cRdlSWhF/EwclmsdiPwp
sD6x+Ii4TQvFz65Y/cWP1oxz70+buhHp37YyTqP7m9idMOswi9Toic6Dep82D7UJmAyJaqtrVZAO
p3HMuXCcPkVT5REIUPQpLqAi5WmOkiEDSX+wb2y9peLlzVLBcNHd95RvBoxan3d1IIVZcR4m4GAJ
kUL4PHEhj1KwBA3dKXD44+rccTS9GshZCU7dPL4DgZkdUrGCBBzmelG8yJ6Sn/+uQpF6K8AqDz8z
qSXjU5BG6tP4eJP/M1FJk9Pr8VxdBAbPgegOuhz6xxqviOs54pWDjGuI4LBDCoRubtkyRzHpsE9l
MAC96bVZFOVbP16WUn14aSwy+i5Twr4YQaAlVhfVaOIFRL6DJ73feeir7uQke6vGqRLJZ++zuBLR
89NkNhUT82CxW9ASJDfFctKUcyyGs73hQxI59xI1vGcf02u19Dd+frmlwgUVMiO4+UUXUp7A4Vfh
0pwEyWkRBnkU/NO6NJGcQVlxI+qr+/qh17gASjX1kWDYlwyLDKNfVqUDtgzqrwtExcJ48+0Jg6Zg
8XJnNFX6vMNS3nskp8/OVdhNczoYiWY/wfZZbe/u/PUbDPVS3rDOoQOx8wiSAgCDfxkUN1nmM8Lq
DmDx9sRxihcjeYwu+t22MGuQRZ31qcBG53bjC3FsDAYBgnmt96QMMFRPMMUzVuE8AfcQJ988oydg
hqfQ/UamaLXdZf3IKM2RrbVtXz5SM84XtQyf9V4Y5x04hb1N8wWF9UJjU+FgJCH3kD61W/I2ygW7
8iQGgNR5yBHbXOCXwz5p8FeOPgasU4wmG5TpN6Hhpqmh4O1IAwiPCdC6BPfsfZS3G+8VbSAK9fjR
rSbXwdkU/hJjKAbG/+r74P8pXUwDswBt/3zzlqjRDXQgxQAxLN0RCqf22eY3u3s0CvG+MRiMJy8m
zZXF5EhVbS0RRy5XhU37n5refrl+iERoboLdA7Gcxm29l6xglEkrsBHjo4FEt1iuQj7/nCvm/L6h
zwRKWqfs0qL2+U8JYlynpL4+Tz+TKCyArOCjfvbn2AWP4J5K75qZuH0DtiyhrvH1f+wAf1S26xP0
scohHoxU3QF3x+53+e/qTMc3RUIc3zH/DxFbBCPnSC7AQH+0RrxdhE+kB6IWvo5ZAj6LsDVtGESR
BMhrI9TybKlzvrn7vZCvx42hWXA4n8QQzlZPuy6e74gTtg1W/h6ZnuVTzc98HAlJm+GMyr4pLzu2
dv0RWq0KJ/3LmgxMFAf7m6tcy++AT5ZrybPTDViaRmN4Fe//VTP4SMaOS7v0xWt9jOYpsoZjl0s1
y/Aj3AwKPlARCNTepXyIjI4HZtD+ucnOpWXmVJQXIHAID/7wW0FAdg56sw5H98uEhgNgtAf01zL7
ARIn9scJFaFyctjTe5d9sJEiU+l8TjtIsOlKIgj4s+iM/RdrjPaJywDW0YxyS3FrfpGkMou/8ekq
k4Ay0EaQVtIwzHmRR7lBvDFMG3ONEm6Ec0QIiv0LDWs8KFoy1hFL/6v0aHS7/6D8GrL9r8/8eJZS
djlaOv5FzJIudRveVyiXmKPbcwZhUo5Ic7LDoPy6mV1nMfX4ljlJ4Jfddcm09RA/WsAKxoIiewzr
L7+M09S1UlHu+X5f+yw4nKXK8g3FD8+yC0iEVd0PXPmEuKrG0Plr7kmZSKdD2UNkfNaHc1dX4F52
ePXrOxstl+tDDuPinZlRpHRv//Q67FYwemMWbh+5FGGnJNM4wU70jTaeQ5k4bIl7+XhdNjiKPFrt
WpTzHQztaomGiSb+QXl/yz0X830fNVM/9tWinijpqYJ17OjHalzXr4rNA07k8lqV7Z/rMDQ37Q/o
V5qxM2Hqqw2mPRZYoadu9zWh1A1O4uX2UKwwDc4/SSZM40ZDnxjjYFKxoHmtkfY1u9Fp2G5TDH8D
NXUZulHPp8g1Id5bJebDT7aQa9D+XfIomDBJiCAUZBLGpRH+ZRptd9Z7IXoocGNhwV4YdsNJr73h
filQ1zJ75ZBFzuKQVSp+0QqXzdsOO27zW67nj0deNS3YuxJymsOTWNbOmK4IDdG8lp+4wgUvpGF5
kBLIKNs+Bkb7nJ5WAzzu+aeAnJvnu0Hv+4r3Uks/Ew5F2aise0TOVvM5peclK59Ivk9ZkKJr+c2S
7yLB0ytr6RFlRYwCtS8Ujat2THeKJSQ4/kzUQaHj6/YYRR0KDtavVT4aifnXWmoVh7YAs8C2QybV
UvYfLqpigunXAAwTB2Kn6JWRfDVDnPYNiIR9PGJg6YihQ2X0z6UXlrVwBaRdKh1vL/RbX1G1HDJ2
R4vf01WYRun1AujlUTPBWT8lJ8+b1yAQxNxaG7sp/KVBwM7BQAaZqr+47PZd0ooyHzwgT9oGb67d
uc/0U+DPRXgZnc4LmxThgrv37NuHIIs3dQ0DjzIYn1qUof8IQe5aURYJSdaeIB5Z/Ds7iizojqax
elhVMt+mTqds2dOF4N/HAV0aMT/rmr1gkSPKUXNylfEezrbgTxr1UrEbD/K48hVgNSnMBlcrBJ9Q
Ycr+e/Kfwio0QUINecvHrXfqZAPAC2yZ+67VzG+s78oMKPS7TR87GNZwjMjnBfN4QgDNEuc2Lt40
ZdJ8g8iOYUfelK++93avr6Vy3mJyYr+Yzt2/pljNWAkiVIUqa7/dLg0yA+PnZnuGUWeMkEKrFYR9
lGm0iK1oJZK48XJ+4O8M/oPMwlNos+TnLQJJttaHWY8oHRwEdzghY/pCA65x+IgaDHu9Nt67ijJC
e6HxFqU613YG3LZt9QPbYxmXW3JCZv32/cBQtOV6JFzzL7USNBsBjOx0vDE2nDIcbx/52hjFQP8x
nLUSdoryNHFiasg684s5abI6oYtMpg+0BhiBtu62Nqk939+NAfVpyeRRsgKg+hoXd8NlWMojljVk
IikKz/eXeTi89HxsaKTuRrmrdg6TrzELfGiaasMIcvqwIRZHboYctlRnHZIHNlFCz+Sow1EC48W2
FimZBh7gEmulcut8rKEEEjjggqgr7X3vPP5SvWg9bNyU50rCYOk9nN6rg+nSjzmLU79cMqPqHoV1
YWUqIe9lw6iiMrnY96wQ6sNyoS1W8g0EB+OY6lxnE1KG4QSwAHg1l6TguY5Ooz370rLgL2yE58Lo
i7dSG7kSS011uDCG7alD1bl3Gpl5k4B4wRe5Xl7vSdIdcxM6l6F4zhHhiPqgq+ifjC87zKtnFeQD
55epKKN/Ca2r8SE5LC2dJ0VVrY9FXLEBlHCFSlgmWBzn6CMDnuagN0Mvu+mSd7kL/e2LwsEx+KMg
Ny1rXaQVxq+RQpCIzvspWgnGFqqpuamJD2QPngNSUSO2mToLB6kMGAPogjmbIIQnLvl+FptlAXC2
pUI3607Ny284u2tAdmzTAUUq3/lb3a9LppaN2NFXAL+QhKrCZ0wbZRawdgZAo/Qes5lfgusYyP8/
B9nPsoshh7ftcuebl7eajQINHex/gQPU0FuMZVDlyLxJvqyouuR0BIbFk85ggahrapkyf+gvo0Cl
2NfCQooopxwVIFXs3CFJQWepg3rGGwA9Tj+Rllc6uz8BivT732zsakL68Tg7H1vmwxAR/UrZ/GlA
dJQj9MdQo9zzn8uu7s522YwIjoyLe0io+3J7DH5faCEt+VHtG3yctwJ8uM7DIFUSTEh+qiIAwMGW
lDqPSeaYC4XRbliqQer6GFpczpjONJ4QVspOPwbsxZFlRKC1CoIUGO6GHG5fLArTYqilax7llYdR
BjhezT/01fMkj3wyhwmSu6Q8f2Cw1Mlqlgq8N/xjLjoECzI56aO8NZwkWwSXgNMpTqi+K2GNvt5Y
u/4OceeDqZOc+9FxGFYmBYGXGNvYGHyEpT6Hb9IcoHsYXSCAo1Ja+urEw9BRLCWiLR/tSJRqumF0
3GJVtxKTrr1/tfWhazZXdrlgRJHDmKp/1ZeLrwvqoZP/YEeKevxGe71BHUkyv8ynCQipYQAnldq3
d9Na9flh4Qj30A+Oi2OYOLXUyORocwPLuKIYdn+CzxgjATxuYK5cG6UJJ8tBu1eXBR74HjcZ4xi8
P4bRArn7KvE9+YDU/fXfbxDXJF4Xpox5K5PkeHRLMsxpszCnodcsGovYVgqA6lvsKVCGkSrUeKi5
uftKEmTLoArHEoDCpaJYM/gX0gpGIKnJWf/QxrSNRcwjadrBWM8mJC785Yg0CbPThOSuUlCnjqD5
KyI70YeiiAQEpSts0KNMNSWNSzmUkDTjC4RFUx99jtqoOAX7NZHrbLjkB79Absg00q3qxQDHWs8H
HZWvReivX+bO6u+5fJGkYOqzbtQ/4ZZtByJsbKKhWUTcwpgE+Q8lD66kzuJJhwemmzPXTcoQAlgU
Y2OJbTnPwJ26h9GxPPplh3+AGgwGX/V9z9eY6JZaMpZ5ug6m85NbwCCzvFarYWOouWizaIcICB1x
GhI5V3vuuK4vbsku9MNrbGUTRT6HVOpL2zRWqwyLlVR6RniJTTk4kpWED0Z14lbAgtym5W7uT25T
3HDjYvoEiMxoP4NmqvwJNnKd4e8l8SZdDHlO5dXYqgVllMmsW40XK4Z4pD428ucdCrOBwpuodbPc
w7x6qtMxlYguE0Gf55zD/pa5IBsvo14wcCp32YJoGB0qce1lQwylycwBdiYBNZYh7P/LKgfyg0h4
FXHdS6Hc+SLhmD+E4UzGqF2CnPjWYyG7EV0tkCTkYmvwPGdCnXv/aEkDMbVTHWlZ6qi7Bn0jowAx
WAyU5ddr8nGiKEVnWr4mdTbZrBodrNJ4fADyizeGDykjhoSREEnL3ibH4ytWgOJhCISFuGGaGYjv
Scc4k3I2//0dzQnNOLrX3hq/CdwHibRdFeDtEy4UZazoP6Zd1HDEvxWQEO6qbbTcCC8Es40eoyC5
mJcpcFS8+mnGCCnEnnS2ofgx4z5j3RJqiXQgLEC/9p/R3XUaIhjkeyUbhI3ILNhqh0hTqs1MICnE
VgIj+kLlUDB/6Hym3TLMeaut0r0tZn+zylZBjPOBqru24qqu4nJKVqgD93bK4pLqi4J9Z5JuJS4m
eGHpos+WoWtxzCsOXQD8T+nOCslH0NEc21nkv3sAJgO2+A7tYimMrq4V8h3s+5ehe+O8aIjxGe6Z
ySuHd4+v+m54Ss6mR210AjAxLaTLwNrdOmmsxvhFkAa76y+F2Tyo1QUYf+r08onUpHVcBtZNMXVT
iDgjtvFkm9v6CzYMto1TBuj99ou60k6XaQ4lxpOiMeJKLmjJwDWpJla2ONkfuvbbrj9iDmFvEOYK
FmqibUwEJALOVjBb9OvbFKHgilflQ9dDbUa4sxlv9iIrNAALHMMyoKjjWc3r/ySxG90WLRQrpQzk
D/kId4/dwaK5t2bU2Wbey/8+yc5lY/7898fbBZL6EMpFuMhiRviZeTxICX9WKdUzt3/0ewwZ+ROW
Z83W48MwdCbzEIR3w9rZ3fEcE3Qx8FO0DS52p7dOj6fOqfsDFVpnDpSPWPz5bu6RPKCarfeQX00q
UGUXflOCKWoB3uoTzzwIBHHgID0yJIK41+exorczgYph37yVR/00D/czt20Tx5H4OETFh0es4I3j
GA3A1H2XJqPJQ91iL4zda9VOkDuGyPdA/8SPs0Iax6SCR/stts8zB6HTh6LQhhGiwwYW7K9ijMVn
H77KsU7OzpLOqCeD2XcMC1aPEgTdXB7b1/mxiMbD9q23KWrfnu8CfH+5Z2rba8ixrWrmkMZVG6TE
F0GZ8jmTIGEbwiDrx3Wnctg9ahK+MjIlQoumprTjTasKBfrE/ANFiYWaHXR9+4n1UNGBLzHc1yxF
3hWjfTeejwLgpWU6qS3jb6naNyTItm1Ucs0pJQYQfKDq+WaPoff0IxhPGK66F5VEGRefb3PPIo/D
mP63+ypaMO2Qcgnyc24RGefTMn6Sm3iaqe8J8rP9OY9y0aWApvL4+tBZd50QTKNffLx+0tPoDFfG
kpuqi4vrnvFKCV5Z30B+A0hQKd2xmhsyAOanDiHXvnZxxZ3iZQ2UEKQXj8VOntrN4Za4hu9GHbmc
LzgYSG6V3xTnK0DB91MDpWIqRJoMqIVV9JeatiKvXXcpPJCSfNE+6uOVXvuavTzW4xuHwm/zm5U9
cMwh3njLisu5hy/4rIE5PrGk6bbbr+7ByZVtcPcb9w3JxlsfLS3RNy/V06fKiMg3CosPE9lCq3QU
Gazg/qFvpmT9y4ake8EL57iHUw+kj5LxA6GCALAP734tqFWEVZffJAQnq8JqZx2x7kWfaH78oGaK
Imk8jLtNtqL8XLIRdDXClZ6RRpfJzH7Kb2fKVYEtU23lnFrq/K56pJAO8tnNvWS3aVwAFUtPmWd0
1RRZKio+ox++SM4sCiJVUvv5DwGumEMEoXjCoDjfQoT/KECtD98ckDXGjbanvdd/c+PQRPuefLec
g1uzS1mA9aFAMDC5niB+XkEfVOZnWw9Lt+dBDfEdX1c9nEFwf2H+zmHd+KHqeIgok+Pdhv5O+QvJ
vNmGbHE2NoJ/8ccKj48TZG+aqVSRTcwJX9+W/Vg88/uzLlBCwUhEJ9dSn4wLhEo09b9muY9eFOuY
NOsfjLfGmA0HQCex0wUlI/pXbGgOo7nxRD0R/JsSDC7sOK438zK0UdFRIsu2L0CbzWeHwbFgqHTi
BsfGVGfV7CcV+QcOkuIfsQOQ2mCJFmPIIpCZ+0cJGtzZiTsahY/C/Zyd/25aUchqmF0SshNBNIVM
L+hRWBNyJyc5Bv78iznqGA1zU67kO6BvbNoGZXQvoxUwyG9SZ2m2ztrTdIL3ugnjTlhO2NdLJI8g
d+7bK4g8rNST1RKmei15Z8lmETeXwWbeX7akV6gIcXD85WKq2STGFOs3h1evm91KPOKo1dRXh393
mgFQgeGnm/x1jlvzzxlgLjnhhHK2m1k+IHUbkLx89xRKTp7TMBa8y2HzZaFbMT/+MjT/tlBkqhDO
vGxMKSkmdDTiHUUrap0p+WP8w9rkr5Xw77gupDtIxG1yrd5OBi/tT6fLGmSspUlYBfaqoDY8Ak6N
CIqIzlJNv2246SDWFsvVXJ0sTRcrF0BHh0/ZnxlWyBAWWoosI9WFxB5TIJ9wPqPAdPHPfTwk/1Vs
NjmSZcEEhrUoejy42ZtC9v/kPAV2QeiPF17fOs4LWuH0q7te8a/RoZEZBJm6FFdYPhYontRVwdCI
wsPhBLvn3QAMIJ9ZwEUR/Bm8eZrjngv7x1ovakoMUECFVbeIJj6paASgpZ/wB62yTpzEhwMQF67h
ieQo0zBnrTdeq/QRM8KMIeRN7PhabzTlW2VW5aowPrCQyIIlmUN0iaEsI3lPUXgs6PZVN91nsCgo
2herGSP1s3tZIMp5SXVvRNzqIIFWkUDxMJMO2FKR56IZKQ0YHr96K0kN3NN0fG1KNn+i2whn4Ya6
M3h+L6qbuSrwtgpzfEpXoTu0YLWjRG/uMsJbMTvf1hPJ9wRXNg/xnFFqo/zfS/pDwjjRFStzeq9C
qlCFhQEhZ1ltr2FJj98YHAMUWFzxtI3t9XCDbuSWEgSdpwSJ5qpSDgNpMg0HJdWM+Ok0vUYXaKAu
hMG9EdTDnrHqFWhs9iPaclKYVIoL/BxENBCrUH9k7meKxUTCH393+0at0wSZCNM3iKXl5xEypMtJ
cfhyCgcEnjQwQmXDPm2ei99G3FPChJ9lN1Qf2DY2GB+FuqQ0CieK5GeN879nEKleRnA5oVkIKY9R
ZnQxmIvl5cAHFdqTg5OtK5ysElUnQo9fbUTMbfyBhNE0BkUznEu6sx3VnV0xWcezUe9OAaKbzs4U
JU1bORI3oN47q/XDJTrYLQc/2hzUttmK+Eu5CsuJ0QJPY4HleBrX2PpN3Ky8q9QlspEfUaC+Asd4
IzqhCYjW/rSoo4NyE8ST3JSp5mMTRtaQImXt+3wGLsK9XjeQ6voCbT4enC6aCIOsX8SGri/SRXoO
v5rghK2adwb8VNA9+3VzCjtWr2dnLFL3L/WWXvLr4j0VduEQrIfd3OXv0zH2B7rgjL5y+y4LKAY/
W9wVGK8jtdjbC5pK5YwSuuF93iXm05ACiiGWywHCP2XwFwWf8li74AeaW+akujdF8FUFhkBfmnhc
9PBHhpYucguIb0UncxO9c66zX+xIsfx+USV0RNoSCCYa1nW9tbBIOOuVAfIdyyV5o2ITsvC+spTp
qifozkKt0LpFUDQaFgO+aQoWPdAle/19nV91G6w4szs9pP77XdhJQp9mYBMqcjuv/6NE6Aanngxj
BlyxENuCB9xG7hC39k4JSriG34iyK6z04rT0RxImN02rgzOVQmqasQbVVmgf5AlkkBgaUlcY9LEW
gad1pvHW2mUcxKOPhzXM1E6lLbxiwRRvM/CmOqSDLw63l72jrZX5pEBVLck4Yh3nVlv2B52Mz24m
Y22W72h3vSb5RdLshmdUpulS6lrKFArg70crDt9Exw30uHBBzphwR9tAxHO1jSpgl/1kHSmkgjMT
NA3rmCLG7teJ16DKAUgLFBV5P5aqoquW6yYfRw2lj73fQwh1/KHORftJaFRDiemOWBqu5ldDqozM
YlNq4w7H7Bn07mqxkgXiOlMbR3+efy/c4S5/chBs09Llr3q9ygoX3r/I8FiUQ06EiyDAHxHl8FOV
vCzeahyJ1ITMIHIm2g16xYWpPmzE+COYbirETBpV5c53JQcViUoBuKwY+CEHJKj8L1aFBWsHO/QT
tkFyOYTQhLO73bz9MKr58RMyH8CfN/NHKP7i8AlXD+F2lqZ02mkI7u3leEe0JJ6pjoTy3zLkFNkV
FherjAcgIPrVf+p4i4P+eR4qidRGnh1qolr0W5uweApE0TUL2G5EjQ5IYavlzhlAbEmfAGtU6Phm
KSYKNxJABdnkb4kDr7fZUGqZheKJmiExAuD0R+Rk6+0qghBSc3qpNU/fiXYbzZlV4pLLA1WLi2tc
l5tt8KP9lxymKWDTIobn39SddkUxSCyt6kjVZT0q3cDy4myFPqV3xH9u97pc8rFK31MaYaarhafY
16AAb5o3NRUX1cDj4lhbRYMcSaMN5zWvAxh3BYwD8vEqcYUXAL3LASvQnoMARL4oUXf34YMLENyi
KDsXnccSfE678Umm+cnFXTr8d3m15Rf9fDsvtgHvuLFhrCRgz1M50yJnGL8fjfFHnyN6/4EDr4NY
/ZG8KbEdCExQIAiI0hwABdgElTh+l0qRO5W7D5YKW0uDFL/xMK2och+OZuEmo/sCeDys69Y4S4Xr
bCKZho6K1XSWKg8u2ye0oL/slSkMU6sd8h6aTQbbPyEQu58c1+LiNsu4Mv6C0LBO26vlozWIbWAI
6j60jLO7j0DnmaN7Ef5oAvW7UYp1QndiN5bVOpGZ3E5wcJuajweJWRWxiBzLvwJM4vyP43udFZHs
FttxnGS2/YgW0j/7ANITwGqXq5Ba3J5nh6u5a9pa/LFYkQM8iKNRWtxzUvnikBjJDBjfZqlqNm2M
aO+2VxMuhFSVVO5RX6dG85atVA0kxKzxWUZ1cTXzCscZ8NGmp6SxEwaa233M8K84lFLLXquUrezK
ykswnNnoJ5n8hgja807v7nOn/eTABwm3rk1wGXWle0BDOpRt6dXgiXUvWmUkA9n1W4AAxN108fKw
NOzICJeSH9hudDTqtptHyXMlgzQz/Th5nQfgRciCLi1Q1mOXWbO6RIKT1wI9D0yRhOtTMDFa7miz
dFgKSl5wna+HIPqNkUgErSS35b/ERl+6Tl3nTzbJVbL1vCiusTM6XPMBDmJK9PHIIH+g/CwqIy/V
De0BHX1MO1UOZO9a8MyK4RJU36tyaK4Uhrl5cS/TN4h/KZP+lwzGH7FFlBrz3ZaYOI8r9k+/pGLO
divDEFdEtQEHyHcsbs+taFSXB6L0N60d87VfDaHz5mJRSAnRGo6iXAq+ZcqG9Ix4A8obbKPObULn
1Ung805HiGtbgMdKDKpXcFfa346KZyunZNtdesRa7nS0cfpognae/TuRyKsUWEAKxUgzK0RAWhv4
nk2v1FKaNDlBzvk/oi99nWIzzBxcL6GfOzj3c3DBTvFlL0u7PyForRBw65rIi5FfAEJb0KPo/XUO
ijwDfjmQ+eWSjrVSSYvruixCFFEAL7Gf+GADh8ypWlTATaw5hxj/bXLKFqPA3vhMuw48CWQTMQSx
HLvITwStSUGhjrOaCuWK7eD03UKVvDpg0pEO0BiVQWei8Bp1twHW6R6wM4wycnI8yjiaLOCDtS3x
KHFNjlYir2KgU0+6GEzaDXTJRvcypfgUXirAcYAOzb/2YLbgZ6ZIzQ2GUyyZyYH+sWmfDGSuaud5
zoOPZ+3yNRMIlajBsUX2uspjAgiS/BXiNmzu2lCMEXWDrx9wBTDYXfgLx3Q1ahyBhUqXpbIj8CEO
Pjf1iYMsVtIHC7B0r6vmTt/d9A+N1aBOZ9KWT09yDXw5sHxuyQD3i6fT2R0y2buFmJSXTapK12lt
CqHfMOWZBn0LTNGpNqRLiBLUfh0HB3K/xfjFryoil3NdNRR7SNA/cq1MvwbCijCOmN8UCSWEMdLX
HnA6Dtq2bjCXLaaZ1sHRQ/y+VtOeqJMdrMpC1VW2AfP+jb/wJ016suRRLFaBJs4RVLsh3lvYMTSf
yGTWVZCMMwEis5S1dhpdyF6iMQ2O0841Qazbwts4nN82KjmbZpnTB/ykx9jNIl+AUZTT36zt4ubF
7ptBWI/puNmx9BOFaFeUlnhhHtvmvNNZrp/y5jW65V9PomhheJI6uCfBvPTZD4O878sCdTEo0Gom
LPqXsCsIvOUG8FLU2a5xcK6F+n8A1RqD0cySEK00by2AbEcjkSBS3E/niS+AFy4F1GYdnspSISPc
G4ojAGp3pMESeqgClWbbfVlT8Ot5N7jX8eaC1Ek/MZ7xXlLuXHQ9TnxlQwAiQLR7TMvmgR1iZcfL
vvesachAJ4A6fwtDBZ7bOFzO+lB3z+MxZB8yRpn1VjCkRVcMjw3JCUi9AxKlsVHwbg2aoOaqJMHp
3cBpKskfpD8nG6uie63eV2J9nDbh0K6s8sZCrH6dQs5W1Eh8AQFTPtLC5PfJiQ9g+qkleAahEVtR
sxfQMyw06uSFoKjo1S1YlLq+8H1x9jEyfTbmVuVtBg7T+E7D3PNxo+2Dyz/zxQQ9E0/Xyqqvy65V
SQQ84HvozJLs0S48HqQ3Jf8bNvf41SL8H8nYuYSSn3lKckjSjyN8r63yzjxpc3lLWCf2T2TODfFT
hzsbMis6yZh/uzs4VZrV19dLrZFgt0mT+67/1LJBsBVZQvOy/s7BQvmAy/01A/AniczBI/nWFhgd
ogGYQPGlW3VZo4sY1ZwCg89eT4bd+earm9Dw1U+vF16RVSzVVhrJRXk4jzjCjmAFYcIOdcWnnfyk
QokJxIOKQcTbT7T4XJGg0mW8NVdkHWlXOQRB/ZeTLF+rtFVLxlc+0Ym5qXS5uHCHCye4RNzGSBJg
tldvy0FXQAvd8X94gf2N+nVQ0sT4L14p4E/nXOtSWjlFwDG7uY/qtHkz8XGQ1ej1fkAfhZ3l4v4s
iugpB1MuuWWHxKebG38rSnKDIjqFAqGKhXzQETYmJiB+Cpd38duojEPaz07hsLzz2FWo1JA6dehN
aFrkSqnaG8Us74jaXi9tWsa9590tXpKgUnKJnqzj/HPUNIvVkrlKntMkXqaILfmiKRg08h+coDWv
HsKvN1SGH0Tnyd8ChdUxC7/3V+ULgFosFzNPMZJxfGGKY0azYeTdzdvHg0YB2mAp/65TzPByXQXY
vEtAWVMD/E+p9qcbAiQBcTxfTIfEjm6ILsmKhtLRTDRhd11RUaQBQTV8xOSNpamJzzgbVADtshsG
X7Kvv8ZgTbl92DcNoAmIgg9SwIHJi0ue8KzAcjdpumjwzhY+/twVKhkr5Im5YkwoIedAARWPEFgL
DLk5MH5KVmNNUFvYpn/YFUkrkBxIjQrrrLaB+t6BTEq206/HpAr/459+y/bfCkiNqEzWYNVbVhi2
+sZqSFc8VM0MFIwG6qBnJg1TifghKXzzLFwhYXm/kZNpAyhNG3UHd2MIKRqnMu5rTngXAHQeaHgj
3/OZeC599N3UDypTToSp2wwEpmI2Keu8lT2SoL9AWm7WnTob6QfrLnjZagFjzXjWoZkp08Jdn37K
F2isfVeppuzVamPR0Lal8mHIwtu6pBsyGfUwqKN+vVc4pIxbJ4cUycm5+LHRYW65Jwag7CC3JRlI
I3M8uiVOOdhCptu3QBlCAAXuFYMQiWoSYVMoMcah4/egXxsJwdnUuhjx2i4SXCxjWc+U4trQclmV
ErsmY+BXv4Iup+x7XpIQTW6JsA0BkzBngxTm7RjJCgGVBR/nJFeGiLxmlQrTBNEahZhcq5W2Cujc
dOkd4ypjnz9NasbvyBjZ9mOpE1IZ0p0Md7fV1TacbdxLkDNh9w0tpnJcaA6pwyR2/2h+lXYss5gY
fpxveo+AfZVishA71dD5sRXOAIPOALwNcNVOJH+D6XglBpZUh8cGQEY+xc3+je854AWr9pEe9Zz8
Y2bJx9gyk9HVQGLFatEZWhiJL8CcNMAJL3aXUeF+ZjRq5JRPirXBM2QA+vOUZAR7nYeyX6PCgPab
swqyNdrF4J7wrsm3ksjGxwoIbCjfn6Vkh/MrxEt/KRTFlV4oXSgULNJm6UR1oBeGkt0hze1XS2X5
nteXlH7mL/ye68FvIntzEaGc86mtlc4JVyg9lh13AOjfEDR7N2Pwic7pcnMMHU+EF94vbm8wqK10
atZRsJ8ko8u5n5yhUk1ahc7SllYYMsVFTZvEoAhP8jqYEM+WCLnXCutxWnsI/mNILcXD/M69/RRo
lXbFTTJR3mudbit57haOjR/90Zd/nZnhGn99/cVRfQM5BQFaBnv6HlLZSgWIM+ruH2dly98sx43q
2KDtnBCjw6cg0TZneyTU7wImG87eZvitphFATlPHIdDdUWamz9CzzUDkQ885LEFHjdrH4Qm30h6w
07JmrBHBc3/1BgQOZ9PWBdOB7HOTXr6xHafDlH+CkfqoEEyzc6fta7Wpaca9h1lSr2JZnr14bBDR
BXSx4ihBkDqLE8vd0NTQs/mlIZUiCF2qW9F0Z5kE4F78RCB3xyZ6Xf+EkEKDWLd7xxA/tJPFP6a5
6NBgpZrsKGV2Q9pTotrFEhvpLpz1svApGl7v7mtveYqNZYzbBxayfedT/3OTwSMSrQ5qZ4L3y4N4
2JmMFzUUpPvGDUFYKNfV2LOn8rhnFw99FNtHv54UooT05HAXN1BB5fO+SYtfIR0fovycmCjtFvWZ
KQjUbq12TdxxwOlQWjgs4l3xUQpfZvi9VAsUDJT3WDqc+q/5kMvYZGEl3y8t8Zhlx7Z34t3RDbc1
CK14FYRpNtBTwZ13azmQ/w3z6mwZfYw8Jk38astCwq7QSG9cP48h5inLUlE/xnnYtKgSoRWp6bWT
0AHiPXXHITH0rqciwtEK9WwApAHTvfTFFzlpvOaL8IYtmD40dPheYINe6xUGhXcaIb6XN0wP//qe
lQH2+qmsMxzTCoZyuu5cDNjxyoc/zLkV2xjfyZ/NK03NpMBR8gdcUV9vnsdcfeNp8qYlOBD6BonI
arhdp7CzFRAoUwBb9U/gBS/D8t0ZobEi7q1FYtCCP6nwKTl2mEVJ5m5/ZzIKyXQG9iHKXSUkpqSE
ZPKssFY/GBg0DDLniIvf+kHeUyclviD/o9IxYkzvJBzRk57Y3/ZpOxOfj66gE77XRZNJ3lTgyBK9
dSomtx81mpQmWoQ2tfHs6RtXydh5OTNW6rizszHedcwLw0Zz5pcizZNiIFnu6hTSPK8fKPJP1UP5
oTQ47PhZi323yaPtsmP/QUzNyXNtGTQTJ3tpnHM7sO2VwDydHo6oyAxvgbHuGfXJMuY2HGt7UNFs
ef3F7vPAdxbUA968JpAgVF8YRuJVCpuIsiH4aiHjqFkj3hXVagPKYr1+VclTiv9rsTi3P9IF/EOh
EvtUWnlcnw5pgwN+xidKdkD698muLHpNRgt0V7ldjmdZEr+C/efRZyBOpyBLPwR+XQDhCOGN3HTf
9ddvZ38RTqZfJcO7vpIOjYu0MPCRebDBxBGFeAM8vkkmlBmxsILkgTJKzsMJccA9fWKr/15fyj+O
aCH3RMRf5SbPMTd8Q4Mcg4TiiRMYaxHVtc62EilCO0S7vprofNHSG5w22ofKQsOaoIZS/8efqB/s
xIhEzgb8/rbfKf9gw1czoKD+Y0pNYrpm2rKzrYmDQGV8SsK3O8X1YWND/4894BQLRYwxAnJ5URSf
IjQKj8cWIYUKc1Y7I6ey2rx/wAqfgcpauDrX8vcrmJapubmBfFi4CKxebtKhChxKZsEUTJ+qGJ/g
Xh5Nc3J+RNgtBB1nGu/6LfAxCye2gTaAOyhsWQoksyXZ6LyxEAy6B6ZxMXP0bUrffzyvioys19c2
VQNn6MpdwIcPnrEHkJSLEYAsF+1aYH+RlVERoE1K5b2XpdoKSq/1VN03kCsiRYyu13/hekON3yGf
nd/hu+YYqnhKw/f+3KerFrRzlqymcrgiB6+UzHV2W7rd/1vmSHHqi6SLOF+a5+G8+YfxaRCtoihA
acnvIUPHqat4x0KBpzzSe0okPcEAnEahl2+UDv7gE+1RhVkDs28awXlBX3qtBCgMMBg54al2TfJO
cijJU2iCVstUevzGt7dy8azYapy97Z7dKw4E+sWnvMbt51YcqmQ8qPQLywEpuhzXeol2lQ1cm3fX
U9RzH9faKUB26k32632rEHdzJRyV5fO39ICT2m7b0FMLIT5IEul59VxxcXQcAsluqU+Yy+ggdrJi
1BvnQeEqic2vgTXh1Frk1dcjj7KbWKfRZHqxZ/mbeVgcq3q7+77b9d3ig0H6q2q7FSBOwR/Y6vi+
hnP7eZJNMdNoozkHz9BV2G1zzFfnLIEgWujxrRYOECe3FUqDvVvGsXlpYjQCT+Z15f6E23Cv75KL
OQZcYedMLdL/IR0Q+vBuCosKKIC20fV5ggLP6Q1HjmJy7aEGZy0Z96B20lGzImjjb2ZtnSYuNUVV
55lrA/yrAzejVwI0cTTTxFS/SmROChgI3w2690Mn1a+DG9QUyMSt6w8x23BTOyzw+7nCxMMEmPDf
52LHwCLJ3njSVTCjjTgEJzkrXz3Uo5MyA4JSWn7+hdXx+KCgRpDHmjRb1OSNxtgQfF9y13sWsflb
Kh88qI3ZaMV4QuZwnsqcm/t6McR4kLmBDKsJL9Rpi3af2Yk6jRKkERuMKpvD18ObCnCxHiZktjLK
Y0gBxPU5b3TxtYsyp24uxMyOZAKJDbLMLsS5Cb6bmZvP1rXR6kswht1xetTC/zB4EpeQS3EbjVmo
EtiiGzBKwdQxDR5Jp2gMOh5Kg3GfDFD8Jrnof8rIBnesfp65iEwn5RO8Hc7TcOvwF7BQ1ne51wHs
DNzHek5Xl5RkiQgVmP9zRdx6DH0hZROr8esA1e8owmDajme6mwGg8puzAXXnJAjEQgKaKITsvz5P
sQErshvgDwwV5CxPYvLy/rId1c4XL5f6TtSuj4btJSJ5ZxXY+GKFzDGHG9brZcXIXYyhRu9p+dYx
YcBeqiZMFjEzhh++uX1Nea5DTCQKR6SqachkzGRzFrwu86P64wSBBboFerua8VBfrk7SVvqLJhf/
wov8ec2bs7qApNGaqm/nic4osui9Z36R6pksd16CngPKUGT58CfHKYvM55E+eDLYB9f06BNpBzWd
Vwto3ne6kubJi+6AJHMyr1RxnGfDpxeBSoU/lUbmFwBb3g2xgRnBsU1+5sbmYqqaKfIttGOfGNsI
qMFEoe4sFl6vLE1m24ByPaGuePZ7BDpcL3RP0Vh7Dc8WjHZdNQ7uD0aXJ81RkRklAyxymAkO0/Q2
8c9WqpbWPHM/1XYc+eonNUukghiLU++4g2x00iMt5r6zQIIzhatA8jrYZ95kOCCqh5+qHi9CLf8d
YEgJiyrVuhbKG+mnkB1BvAr7C5Lre+vPVB0lk2VEyGLJR+FSpSUE2g0FmSdFjMASW0W2UpH5eDin
2aUosZtuDo6sK2qQrky/URgvKq8aa3aTwjmxrvw6+kweHYBwsDKaDYNpFGmW3v8BeJLvKTmNnwVO
JInu9Qn07WZh5EZ+tABrFSreQ1dYir2zDTlXxs9ap2xOhm9gaXbC1UbXeIv+dzBqpi6G1LSWSdoR
bJn6sOZ/FRZC031JpYzSf9dH6jwFQLQXaiLMPAEJf/5fM8YiSU07iyKZDvog8jdE6bY+XtYNlPuV
a6EBNfNzIuux0wN6kALFnXSPOAdvJv4ELdCpty2Jr50FLNTf3ZoBQaMrbAJOC96YWPkNOrXy7ct7
Hizt/aRrwJ40VNc6FInglCV2xogQHQMakHqUdrPEbOamMnQJ/CdpFRvmOe/xVA7Sry+JoWQz/WqG
HREdG68xAx8hRP/pe0QWspJs8+C7KQvGzcJqg4fOOiCSwUitWwMJBxeepMKJ/K3nSV1s9GpzhEV6
FPVm66Kw5z7agW8GOiIJPIprCyEMqRLmTUjx0q/IdMOfMDaTzIeagalWeMG+8jMJmB6+iwpx922r
ZFKue9IrkiqCQeLElQUgBh4n3xlp1NnBhJ8ga3ydPf2VrGS+0/zfjrHzZciXiFN4jjeyF3XBEak5
AkLTVBgICjnFwUiKSrwUUxH/Ch/PmXXyWQFriAbe8Kze9BkhYAj2vXHThNzFNIkPI3MvgoQ0+K2U
SbKrxogvx/c7ysv3h4W1/BZjaR0fBAPLfCCujFbzxoniIW36rjnDB+y+MWd+QViY7JihBbfI4oiV
IVUyWkEaDButsWsCFtaCETT3w5sGT6CVeEmMHgzeLm40b/DDgdf5sSp0r3cVPXsQ6j98Wl5MY5NM
HAiv9EAuJ0sxWvmbHWZr8h+BIl/X5rqLtKY2ztGA7wQF+qONmus7LK3uKIByC3de6hNtRCSZip2A
tttGwrqCo4b3AipGqTPo8gYOoEZJJ9+aw0AO1YPnEdVLVa90wMzWtTM+ve8rpsnk9Yui4Fbmsk+O
RJSB9VprRRY4Ku9x4bx/vu0hsmSRt/jDLZN/unkyFbAX6/IkOiEmZfuIkocsCruxZ5s5Wkdl1zji
TK6eb4gnq9wPvDWADu380c0wLw4XYjWTtHEe6idulKNHEHjO6VbjeA9E1eNfDeS7bqdWYhEyBa6r
neFVf01TQHstdlYL2VOla0O+6KeUO8xxF7nkKZKWY7fJWeaAvkFzzTi+uAgLdbD0Vyib7ZUkORR9
FTmbdVEwAlm8m2zxc1Jjnt5DGXHtgRVGQRoSBi/b8SpalCuNEbcfW/DP/wBUm6g2MrGgSs1CpLI/
sTpO436u1PGEPjLGTs6DufYHvsd74k98AtjqvQLLjr5u89IRmLC2dMCg90B5+73BHLA0m0ax9HID
CLRwgXc/43ZnYjtMC7fRRkkAWr3maE3efXsi5UgpreID4McKJTL+nFl5lG85ipfdY72TX7wb+YQw
cQlFICA1mea8XxA6onjTxhS7TPtS4JEzgxGQ7tR1LUlu7k8WT1g+ks5e1KjbH0Tb1zL5c4bdL5cF
/0+5G2XmW1m3Xibk5vhhgZO0o+A7VlKHaJ3XOgt5GXIITYTU0Z22nBX5BFDYASRktmV5J/eR4gcM
QwGw2Jhq69hv8l0NsH+zasyvQZaVNhBC9Aoi5/UpugxtFH7Dw5QaxhfEkq5PXTgcAOOa3TsKeczO
iIldweG9xW7keCX7azJFfsPXlJYXuLol6PICLABlPxmXmnxgycdzsVtRehojuMo3cmuD5XZTG9Zc
kDS3LiCYR7CUkpyW+Wcfrt4HfcIT81NsuLkNNZbQGNVFgsvBvllQCz1uzBro8JB1/EIqH1feczir
HqhU5HDbC8uAzP5jW1gGiNT5AMSxj3JC5LWKCfeNF5jZEls4QdK3ngK+AdQqvfp2Ajq/rTNrYMtR
ijJXVeX2EfTbngZM19iQCokL1e5Ijd7Gwre1Ex8WT5XeXp8lFstZXOwQbCoWtLPL81EuKZIWcOVk
YAeBSSMzUDVWrMzDPRvTB+ke9gKLZrFIOhh/ezISZN3zbtGC/wAQ6iQLjCDeUaXCbu+c4II6QErE
W3JOBb6CIVmAWQW3X80RffDMCiDPq5U4Kgm05jLzc4RTnXuM2ZDG3g8MyiprHBINbuUGJOe8DNGd
RmRbhvD19vm8bpnhDlZY+Zu8KywzwmNm75ztgGftfp0Z9M0Z1NI7uII4q3yPfBlNNJ/faFACmSFD
gDN5dCDJPuVlsi+JBTSvAFuOuPXXOmINcvj/42cpB765E9/WTSldTaC+4UBB81kL7RPY7tR9DL3p
/Plcu3t3dZU1y0mYufNSn/WSMAzAQlUDQe9dBDtmjstp/WSt2IGF3QYzN/mLxRTKsFHTtwcKxtdH
cItYLF2BCKT3EWCuj1q8A0KkhIyvdQ+JFxABwkbVe9bpnWAaOiEQURqXUN6XEFoNHwm2NN+MMs+c
QoacONTXb+5o62dZ+viBmPNvbZu6ubwgzleoS9XYhdt+1OD0+xGcRFEiZv1UgkS16O8iB0cA1juf
3X/tJQ+hl1JK/8K4Tc3hYW0T2DEYiYncgDDGUXZCIJsrx7kk1m5kDtKI4MtJv/P/Ct99LYS85tiJ
YTDNb3kdrbVnVDt2uOxzcRnmC2v7Em7LUmAU/W5fd9MJaTLDM/KMRB4DzZrUZjVD5QJ2iOQZTVUu
KxoCZjBocBB4S3owTh1MvnBqJQM1daNPypeKz3eirPbgMzjuH8RhHn1uWFbCSBdqDc0DLQt9eh5N
3ahMs3gUc5HTN3rNGQGEwrpTIPFdsDP5NEj5o7E8746jy43M7mKyWPaIlj/Fu4Xc77tax88wYQ/g
Ug9QGAoNFvCzDQ62QkMMY3nDqwqb46F5W/z/jbr+H7dQpV6w0xa3dWW58bNe014Unj9Gg5rk3udC
rtw/fEKSXicKhCbrG7zjkJ//x4wlq9i2pNlTCrJAKoA/j/LzmPy8+oInkLbeaSJ5XmmTJWDxxlWv
3pHFeCIwvAyhlUPba798N4ZgAgu2Qwc+TmAtFsAYXQ1r0Bdl+FwxiES1TlQYa1RDdb9bwB85pKhr
QPf4OP2IjdAn/0OQGPmKPwm4PSy7RkW+SkAkxfJL0QAp2vbC6Tp76sSCtrhsuMrNbSUsDb+HNvTE
Q2KN0g6TurfSxVnHISQVsYg26TXSBAL/CDnFZSinb8Y8H+eKDQ4Hl+FJIinbptGWUCXTHEq0T1o/
kz14PQNod2v+Uu7TwX0hIA/CYvrewEY3nqkrx11rawquWOt3QzecneFXh6YOlpYK7gzCnWhO7G2d
cdcJ5jr9dMa2VcdCDuDjcXQyRpng6+QhrBac4lm7cfOvwTkvlHKqhO+aOa5dCaf8gnYCYP2lsakX
lfYe+neO0dqJpO58ElpWkWf79SmQREB8+I5Pu6QMzClT1de/BdjyCTleGNgqn0+bGX1OF6hdvEpm
nJOYnu4uHxpv7jYQj2o95ja4N77frstUlnzsdZyIscVyZfa40Grenf2+a5nOQ2jrJv3vYuh1CCtX
5qo0HUUItdZk4ebPfosi7nRmnuPRog6s+rzE8yYF0kwCnH8QG5jL5qU43CldMwtubFUDnCN7+UfM
fDC3mMYhy+bGXxG7Y1hV1q/vtyHYUYP1M1sJftqyrBCR64E+PabLeeDXGummrsNEnwBwSAvIRUlg
hl44mXqDRphknFi62hvPAsaPOBvXcS1ObQiiBIFTll1nK1JOMVTA9IZgxB9MmnUPxTJ9xlHdCXde
fa97NkhK3Pj3DtGIbZa0OINwwvMOcc1eqkdywiTtRrcCzKTqtyg3ypYsuWrAqmjgYhbwbAOlpRPK
vP+gEvnUy+k8nMpP75zfEHiBajBoHuXPmI3pvwMCm3lz/mk+fmxSLbFum9IoUEuEs/voC2Z3kyzt
dVJlv+LQczF2Jy631ayDbavdfSiMjMOAUrfd09HGMUoOXLfSlHT8k5728FRjzyPLG2vkmUciwPwp
BgC16MEPWv0IQkELsUNm/ktViyBqNnCcjUj/ZiL556sMAXguQPV8izTwehg942qcSsmfmV2DY4oC
aSQ8umQJ8l3navutdMA5vRc0k2SZ8MVw7E9KpLDFNvF9HahjEZf1tQxJYG+E5FB8uK2e8eF2aLGo
rB+k4DYuUbQSC3/J3JUXZTSCUuE64YD08sPeco7w/rVuOG2MrqOa6dIZFrK7bqpubB31YfMvoKMf
HOyHGI+Pp6bEVKml8btIAYn513WsvFKwuOkpLEhQEgjG9JXkYZySwCQJtWpEChs6Ui8k7dTRCzzh
E7DJTKikQ4R2+sVhxwSgbDGcZuNL2GvrKyDvJ9HbVfjrBt2vvQMaC+JaZnpnVCywbz87GRxN16Gy
nQ1uGJEbuGujVncr4lyg667rExfNNkTWhUZ2PhJa2zr+WsYICnl1UbxAGsx/euTKoFFK7PoedoYx
FrkAFPq/4L5uBqlhuUWUYcVboRx9gOlp73GArpR+FTVB6jNrnnIOVbk63ntZA0UMsUL3i2v99gxV
SkNHeBFdI6AZoDtmnQSeCuJ4M+2mhzqPFqtbpAxLmD2wFw72IQFbIFxfaQ9CvyjrnK1a0oeeBRzI
tJh6IiRuPlw1d06KAlMcM9iab8mifZLyhYkMxs6VSFB3Av1ZLcVYJcxo9vQkWAUIsn0R9z6obViT
eSR/sSh+/h6cEAhsw1qodw5DMJ8kuslHDQrxhVcTWCbhNnj4x05ckPhwapMFQBIh1yUfAtOJsWNa
GIbNrSOp5fg2yjJEIy/2PQs6Kx9gsk0H7RHD0djAqLDxxxA5WT0Qhe2lxy5I4n7N7AGD5kZxbZzf
zmmVBE8Ak5NfLuGJqDIuPT7TgqoMteEPAwFkQworveoxbdcWMhtAqarSUz69nseisCSKb1LWIUIO
DyqR0BKydWsXJXm4ZUYEpBbcdXBTi2GnJdypDAmME4ampYp0/bKcs74f6d/eFCmWdhQxRplNcUyV
J60VcozKdL9bBqSBjs5NPaaF8IMwJyDvjQqYui0OZXpQYkXkzNECff0H9/HCddNICAYI/wduwaH2
PxMrtMO1e6KfNoL4A20fZ1mPYpHiAnJoVM+yl4+q+P/HYpR5EZXekXLD0TzWlAqLK4eB8hPy5tpb
phfU0Hc9LQQ+TZKfWjWwRGk/qH9HEJPEbRY9Wbvaeumky70WCk6ybR5thzMxHFujalVBSj7Kq+G1
H6WBfYfQC1cFAMBWjNDtlpT/Su7jeE7Icas+/pVaEPmxCmxHKUV87meCQ4H+i7uJpSYfk4I6rVm8
MU4WV8ogRWqYCOorDR1o2IUmLDOVnrddvWEKg5rw6P8L+m7qJ5fbHVcfGx6gZXUh30HiLr/kDnRw
NPxd86hu/AJJvxjqrL80nQEtA7WXgTkdKFLNnM2xKCX/0HjVjbVhjQrpT9SDfM4udWypWCBI4bZ1
QKp9u69fGAxocdZ/zV3/JrdMfn+2cVSOmpfmhb4uueBnC3JVn5FNfNwvTcpZoOU0SjRZrAAfua1H
Agqcr+7mn35b3Lntu3ZbzX8EIMdzNVawIUI6Tp9yL9GoP76Yhnoke/gd1vscQbRwxu84RLIBWJME
FvLuP4e1r/DLDHPww2SqZuloCMFzHo6XYHIs6HLd/rbEpePgg89xTg1GGUtyqtd8mT1hPToi8eg4
x7GYBoA+tvzNV2wEBScFbfNTmVItJ4tqNLbw4ENVEJG6Qq3190qvJ5DWFHUYbderXkZGfgrpICzz
gpuhWdA2fe65r1W9ncupKXE94sqa2vbKWe6y8xKBpSxQblj33XFocKFaMF32c8FGOpsmnE3pG8gs
8mtntUkgNSvGo2FxBDsCbB/R2X0HhJ115GJ0/MkRzQM0TYxaF5Jk8vRy1m+Dn/jjMbp8rz3ADQ77
pGJI/Z4cTrwLAz0YsiuVMIOaGg8nSxLysyV/47ZgL2iO0A0ulqUlaIDzFrnHYwGr55kq63F97ydI
wTUOL4rKbW3AGiK7bAxgoraT2/WhfDibEnYSahI+jO8dISUBcya5kzxfxyQ1Uv+xrBgFqN5hBW+Y
8TYboOosV3cmX4aGOuWC6vKcwrhmrPzGaeKrwhg7yExLmE2VKLTyFl5urLrEjo9WjmQa6wkhGtQT
XQMv/r/AGBxQrtHbxBtNBNLW9MqpAe1TmFG7tdD4lxVOy3bob3e1HTe4IYSW3a8vjZfA1u3995gr
sUKQ9nLSsXPfcbIQzl/JZ95PPwPbTuA5Z4/tXHZCZ0tqG3g1MRa7G+vcKrTjDa3MZxh3T7LIuBot
LzSLOQo3SD8+ASpWYMgjWYtHxfQPAYp1ZB1ZVEG1excIOlWK0HQYw2BPR/5da12LNhd2JFxa9EP1
nOh3L8OZYg9qZw/J3il05WS3riAfD9LcmBxK/lNeEwPGZ2XMrL37R/9R9Y3Y3KBGh/aOoRk+AJMP
Pjq0ps1l7Tr3gCqh47RXQ5llDZ7Aji+93ehAaMWhxxh1qjK52j42YDeLlfyjNDtgcNuHl7wDsSDr
vXD2JZ+f9ikQmUCQI1pmPCyvnEpPjKhKMR+n4yu+nH3T7Z4SF1OJXWriv/lKLMWVAi46yK3Z921t
JO4KHZ+nApzJ/go/8l1o8379xZ3parILsJrPdXZrJeD8Pi7o52BTvolAuFwgekQKAdAGbvF6oBVN
+eaF6u1u0NA4/hpQM8U/UhjRgJG6nlcwko8QZp/tn7hZDBjds0B9qcTdgCFlisNKjFwrG5uSBYAt
eZJ8W+FR8HycScHX/v9of3JYTJWc4fK6xrv7MLJ6v2l0R0UTYSZp/3Qjw1kut7sPDiI85tGWiC4w
im6EV5Gx/AnX+EFZClCEfYphjwIpO+1lk13rcUZOkzbutZvGGgVyyILk++960nb1oowzX0n4iP4V
pCD0oGGYupYF4cc/N/CU7KFr8z9h/6RnQMS/etN1DxgFOCN5zPXQlF1UfdwNxkJvieOcSugjEx4J
ws3P4tiy397g9xT6DuzeCbJ2mCssRllpW8SwZUdcWx0z/BjrbcQaPmWUK0jbrJ/ZiaodwKl9vNxU
amUtSqzrTiqzwApv5dy/Sob849XzV3NXW7bktd1RBxm1PBeHBQBv5Szf1/Bl101KqQYhutpyZo6c
Im1JVjQU9dFnhZTxitMRVsv5K8WDGadP3e7ztpkEz3ou0mnluL1lctS0wTzHcDGL/8MOG4HfO362
T0sa0Zy0yUvD4pj2/eP3ZBSfMoB6g7/WQ+lpbxZY4JawobealS0EGtA6yI85l3QoD526B7oNThvT
9yCnbAcJY+237FYyzJKJ4952voVdeAChywsQbDVat5sDfknbuZTZVspbyBxMu+O1723yQCr4W94E
1abMLfubGXZLV4f+JHibNni2qGu1KOCOTS6X5LltNew1S7Ngm8DGHeo42h97DIP2zEdi33rqO9Zl
83d8UR9KZJI6X1EkY5b2DC0UDZSS4awJyrq/TvNtJEVIadDSGmoc9RP+4SZ52SlM9gjhtbvhULjR
Xv0wD6CRUkzcIoLxQGxbFcm3VQOI7ghU/cUAaexfPvdYyWBe704/AE1N/2owR5vGrD5th1onNGWV
N3XIASX7FEMMGjuRBWh8emrgFS0/J7Q8z6Xk6CIuqgkhxtHWIJw6S3/pINK+oK0elJ7HLBf98MIy
uHfIi6CKq7/8xKwSoH/Uyfewkn98yc8HOFJ3WWWrsJXnndJBbecZhoxC18iXbrfZEqSh764D+vl5
eY8NBIK/9zyAIKK186c4AhAH0YWlZhvwlezCoLieUjPWZIVRCavfx+frMdH2ZqX5EcIZLMobxSoP
ylxLe6518rKnONmYe6D1oF/vSXgT2Wrvl4D8TQWAbcQKXyeCZX9ikiZMgUpkM0RcRRowkOipJ19y
9hO6lOcAz8djj72IgZy84Af0pC4f2kd9ck5AtsSIxqvamS2NTNOFE3f8xSBdQmrEjk/8v2jKobKQ
1x68XdhFot6PQmxSTOpUPhibvVBpkWGE8B1N/tNvaROryIvG7iqbpc7+PrZ+b+PgG8nn90h2NTAf
GCY/NVj/crkCnVCu5Kz71IKapYkxAQC7kFyc0Yb2brNcBQJuQ7QzuZ5SW3wVCmMopiF0l4LkHsoJ
Kxma3/tJIHPtZQlZGer5DJiaiuVVQXIR/dHodka/ra4O7prgRBT1RcBAF6cE/gpmwEA7R7voGVnu
DkjzDjwAd84LVLOxnMLdMEb6XfibvCVkLLwbcuX1S/G7ZHg77ZIYoXhgRCSz874fhnUgAmd5qG/U
CUdfEUe6JD0l4gDlXwFGdFwbkbBe9sb0mUxF8mQSzNEbpUGZs11hX08wArzFxNxvHt8AuPVuLm0F
Vkc0W3EUPMTH8WBwHB3mOKdlO16HuNLv49bxfHg3OQTyNHtLK0qeKMEUHrrqPHaqEWsSQruHp8gn
9Wlawq5NFDM7V/8Z3it/BSyu4RY/SoNXPO4gPw5oeJffJgrcumDFk/9DU76HJO7uREHKfigtq5tG
6NJFS1yW9oV3uhm0djkb5DcDQAhfANgwC4pd8DOjIklPmh2uKxf5qrJBkkHMilb44QWvKgJBQ0Ye
qnlZJIgskjaxEoOKYBrNsz1doG3IjebsdBg5QNUPzcG9O2u5x9z70u4QWaYb/D+W6DH4M9TGkwrB
x3ZsqrU2ix6mzpG9us5eiviGm2yd61EPYeP/PijRCPpW92DyDd1wIAfBUA2rLTcZSy8M/QMZCa+K
FNeRO/Uj/RjLXgHNZc0yXL3mWLvC1IiObq6Cwj1DhRStAc63NPJzul7VM3wmCu2dN7QSj390IaoA
OUvH0baDW0J0qKhxjSPaGcaXvlsWqghUfgOy89ITdD4Q8m0DDH+nlZSei9EiU8DATZ/Y9LoaXLZE
ue/JNY8FAi6T0Mmg5nLZvMkt6pEsQ6gxuLKUhXcdary6qVQnuY/qb02rT4PsYrjpDRe4Kcnb3bMC
23LcsjDV6S6C/9JCgV/MouBerX+CAOR1q0c7RCxO9Z0bsmUSxpvdlTxgiKqSiMbs/UWUpQH0qoV3
12idg2jCis5v4xYCasfPThn6TlElF9jPMpILl4Th5MQTV7Q3HvbaoK4ytjnSwEXLlNGmBKToJA52
j+1LS//TEUS6tzjiYilFexsGuTtzqAbFAvHPRZfrCgBthn37ltpOO8PweJb1PboMP6dOqyBQvkDE
Xt3sAoHEyvWgzy1Oml2kx9Fp4635dl3DjQIgr78K5Wy79F+3sBFlZ5r2GCzVyp2+97MzkSY0rban
D3nUHMeSM9anfuTa6Bf1BdeQ+hJdh58bPw68SesIr1TuWbkpY3CbBKbmURsA10lvdVf0+QkGZP0L
eNeCZDTFkImwFJDxxF1mv8mLC5iJ/6SI2VKPWpDU7yXqUN4Cv2qKavHnsol6qzSTUos+VjdGfS9W
jm7O7oMv159usvOgyTrc4kd8C7S4VytqqIhNNOGGZStpdL3J1hSGeFIPhjtOHvs6p/tlWwOYcWPI
Qmq/Sb+SjyOPBrkloD5VLs0ZL2hrE9aH1LVXVLsNGESO5ls9w9jyFmBWk7ajunFm/v3CNh1QbRRJ
LR4lcyEPkFklfb02zLTMGA/7z9O72ZANRNG7ggyb3QWV8wDyGlEHecuIma+ShVegcDlwLx7/NECF
EmZUl0Wm9aw6vzINlQogHeuQd3p7i3FuhzIwffRCSekOH+eStKKJ4SSU2jfwVPcLOYZyQoO34KQn
UYdpOBoVBmCrrzt8Rq5L9xqO7qKTngXNQdkUWqPDthuEEkgYkxh1sdLsjVOETVHokDUtxQDTZ65w
neg9Fv+R8jxzcIL0X7JTNswSHM8cmLyBcisFhA8hEXj1wJ6wZ+FUMbUQCWOSeHaKgJc/i4tCnAWd
HOARu7BOqDW8hJxxy2sE2UGc5xCbFVue4N7V2fFjgtyGT+wB2h3FbwZLfVbbxKWcIPep6d/+5M/o
fLF2o/FO9m8gKyMUUbkX85jUhBxI4JlNjDAvVJ+GggrRvMIMr8a999aS0JZtgYrRfR1uwO2SY6z9
89VhU9GC44koTBfAQYaItf7q4RsbPzv+QggyLUbCq30FEpX9tPLZNGA0rwRud0WuCYwf6h7hxCx8
kDSK3gBOjS/c+qPdIWUkzv9XNXvt++uz38ToFWN9lUDPuiU8gM9+iKryFsD7OGpLWmHi2dsSx8ZV
J/hdUSRFxLytdXlxnLSOojHrmIpwp6TuDkUYMJ26DmzfZrU0LGsIrLiaPPTXypRQddxe8lAxoWa1
EqaxwyJvntJ7PBHnze8iu4jQyCu/Jtqr4fsdtXhbyfasmhiV6pBj/Lta56PYBJZDCujH4Jqqebh4
mEt3CMV6sZnm74Lf6Z+Mpao+TFT2Mrat0lkk1S32xWbiuXi5y1MAuBDqbiSzOIP4mDlug7wysVIE
k7TNiRyrPZ82R2jDBO39O2gc+7DfeJQT28q+iL4OpgtOLqry4ycnZst4yd841CKf1wuPdPXz/tfI
eVlSOXdLXKTwzdqVs4M6HVsiFfuiX8IYk7nAfWn9k6Fxm+hQblEUM3AYNTRyXxrd8staljAZn2iv
EYLyOoUF1ENEIc+vnVMVYTiAeTiY8WD6ccRbhRiGDWpzMMLIJuA4xJwcGENIgO0AVOmxPnM2dzcb
QeYyNjIG3kPHogmQzW8iMu3jil+nHeFqkdAExRwlRhEkrRgYKsdj9jCryiWOlWWpREsZ0mO1Oiz8
KXMTLlDWKTCkBq1mofCbYk+kYorUBSjV5aVcPJhCBn9ts8j2Jh+GNPSoCYTUwDRdXXKVbiu8T+VZ
jVBJQE8dpsuMlHW1xa+9sNcU9dqypfiZwwusEWPSl0BzWbJh0sG3RbazgS86y2l9an0E4rclYfCh
OQ5gPe26gpYqkeQDx/6Hs52re5VoH4RrvtiDh8AlZd6PU0w83n4ahVBxxELdW/MnuiQ/ojX+YlDk
2godvxHOI6CNoEuV0ZEC0qsxhtqy3agjkbmlKNpA5wAI/4X/v+NBhAiwJ3RoX9Z9wbo509mCWij6
T3fMHV+5iPN/E+oAF5meY6Fs26X2s60YN+RC5t0W7AO0YydYbfS0otfx+xo2G8JDI0mupl/4IZkM
ond4jOcBfVilcVG/WH602EIzTDV6/n/AjzissJxNjlrWW8Nax6aUlF0Ki8O6Gox6dyMgy4b2Zpou
+RqUS+VmNzkuoclx1rgcLnoGlihfXYz+wU2crMSNU8VT8NnaxwFpqLsDyhGB5oaSVi1C1HdZksFU
86JdADZoTBVB2YxZBBoMq79ekBgF26tJqPjELd2eaG10o4IHej43ktV6JR9v1lVZne8kMRLL83FL
CaSehMk5ldEn8zcEjmlC5bLJHzg+gFm3z+Oab03PAPjPSIOz40SQaGzz/Vfo3QBWjWl2vYvm6r/X
hHwb3aBUyxFJpSr6m3CroMetkDwv8FbE9dkTQaGr9pN+pz0DdRE1TmYGC6sdlBJaqPb4PMtQebar
DqK++bzeTu+ZMq8lQYk23+LkbjBIv+Jz9YJM4qAqUrFrh32M1Mg7SI05fYQHlngXT/frtlygE3T7
Mbz+TEhY07Mwwz1P1SDpbL/MBS9n5Hm8R8umojiUMtMZ/HLKll9NJ2IuGzf4ashaPRq8dgiAvSZo
wPo4UjvkNluqY8jBBcoNhLtbcG1pm4C9qMib7u7aWHezVSu6z1ylW1vS7NRHceROcRAc6dAyqTCX
Z5bTLoJ1pAXqGWXlNFws4UkPSV276IW3wZhIOuzrTnl0P3QdLCxyaGyTl/br5QQhdMc4Y9TYOdHj
v/9UZuosOrhfufLx2kAi3DS26pYkRD8eBqo8ESc6ljPiE/NjinIDeI5F5pJpK+jGSw+ASxn79rcM
uCo/0fUCRcxvVPTs95FCBkBLMvW8xG6CA6F1r+fPwWR/JRNNgOvWi84OVqrOKsNXAlr0NAP6HLXp
BrgmDHweT4JWm11NBaDnwHBj1O/ij74nVQM+8+HRf+kNnHUMk9WfWnKI6G4u05wB7U6rP/FdlH7z
/OPfLTJyWKWCSK/uqfN3TOFiwwn//kPIbpnCTdiIqzVEasm8lnBltBTj6NqQa0Nxx1xxW5lwn26a
O3gRCPWIGovuFkr3KRjdkAVdUjG7Csm/LCob27diBK6mE5HkzF4mZTsR2H2clFXjgBCmIGcAE+r5
OoGPFDHbMdSYZ9JnWfyitg+8XqXNqxZHwS82mvq+41CEk0zRTXi+TIgrku6GVzvXKWd4PxTpe+3g
n+kNu6qhAdPTWh/OoQrRb7dsgKBBgzemjLIwxTKIOc2Rv6nX2KU6di+jSz+K/DNN4QYWHYm4YH2s
Qu930b3809MEZudiNXnwhcF9jVaRUEMaiVbMxhbRel5CeuIAKJLwosOdiT8NEaviVRlRhTeU85Zs
N5bsvj+2JwE327NioS/7NfbKkKo7Mk9FNWCq3B2bsmFs4Qw5tWrRG0Hk2qswljr0IM9UJo2hOCwP
KhaN77WBfsoPLkIpo2VZED+DEJ2l1ZFUnMEx7IzzEQM29CzQ7Jw5bjdFm9apc0rxVKD6WOIObv/s
zNd6KDT6cn4cZrtHtNxa247vc6w3h1s3WphJXtMt40b/lxQYGQ0o+H3qR0xtgnizTb4V+QXfitw8
bucVVVEUnCVCzX1AYoxnqO8EBIxBi7WOT3TuSgl1ARmYOBqZivhrikQ9sU0PTwXLY06NgyO7RQZn
GKkcIEKL+TgqeKvx0K/zpnHdW+X37PaAbU71WhUqQXAguv4jkmNBUg8S1DVL/IKv6p5QH+F3bCP+
/mQSpRTidy6EBGi3UeOh25YY88C15iyXm/DxJ616EDPIp67uba1LKvSJTKplVor4RdZV+qZIjQOm
88H8agAfs6bgIL5Bt1Vjit7xigCovNhbnAkU9S5RWhMqT20oe0lwqUl3/rSr9kkY9mVHcr6IQ0H3
FIL26bE17WtDZ7pM6xBHVk1a+Cor1ybYBcicZROUOyx7FWHsOqWElh4D/iDyy/ywjrGH0aw1mNZF
/arJYPj2eArd2ulG+w5zPKuM7d9ju9b1LikUqHw5TgjgPfPNzmayu3M/DN+fp2Yhv7TgTreGzPzn
U28KmqBaBLYrt5BqUej6drjgwHMb0f0Tau5TL0vp5fr9uHy2c7/G0QIBABp9l0KoowJ2c72i/tZX
N6wYcZ3nZDN9MCqoDYToPeBSQhUBKNJp+qcWlBbVHxN+bh+NJMrELeZ0Bzl7vUJsr1rPlbKEPcX0
FWKDIxb81a1f72dnLjSkfZUKojAQcz2Y+Q7oONabS8eQUKzRQXxpOWGvnKIJztTcqEplB6gqJHQT
t19xnvIAc35tuovNNbgN93DpiAxy7sKAzf3eeTe89+PtlptfvnrsL1Njfi//K3FKrHqaTi4zaBvj
U5gKBdIKgqvTDooBQgFpk6BDqz7bi7cL6p+l0fun8VHfmExerq3v1sW15J9bOxQ9H71Zk5Y+tYP0
tH0ZdD8CWCjI1Ha7EQCPMsMCf0JYuJM0iyeM/RqcgX0K9ICvEJCJZ4GZVH0ApZdbF8a/DdayEBvJ
MXgDZEgYEhjTAQjMhIthMWYefEsB5b8xMb8M7ti9pwI5CITUfJECKOZ2HrfF8JZxyf25U5ddBGBC
glj0sIbfkcHFd8fJd8c2Iv+Ljr5QgXevK9xweC0d6YgweYlzfdjERfOOfOJenzGEt1sPUzBVxEGV
fuZrEoTj4UlVGfCNQgdzrfHEj213ppwte7NumANXU4lleZHK+g8kDePAOd9lXpDfxnr1qEQz788g
U+/A7TgJPkcGXJYJ2f3qlRL3jn07hrNvjDysUq3Lmb08DhheRsYh0/epxj4IkPp9V9lt7ERjZw1Y
jE2Yv6xFdeuGqOHSzInQxnqFHGrG5NJIGVLTal296cwfbd+2JHSiLvAS9btumCcgmxTZwn8KbRRs
sG99H9W6W3EN1adwJ369/3uZDTPHnfDfD981/jttfnRjqMQKJo+Cgpk/BJJroDLKnBVecsWNYPB7
i49YJMTbtbUUuimLUbqfz2AVZEg7O73qbfOeyrCKgeIZcpQRSLBGOW+gR1a5kfjyox55whm/13vk
+MntpiVOh5gowBln2aiHnAVcldpKcPqZI9WGMX08yeQ2SGdI02wyOsXmcY+0EyHVxV6OXMkuTy4q
DhuuCnKM7syXgoAx7ZR79l2emsaCaIT7ltuTjcLwn5W9sfMFUKEZtXZoyU2QBQ93KVn89MgR/YaU
Q2lU6J6JaWMC1y0maG6bFuUBaf5NEnDQTwXn0BfBZrp8DQznu0a/g8owehfgohCRYfvKjxlzaLO+
ehLitCzPTtBPgZBWaDdT3ACf/jDSpEXBOkvurk3aOBVjlGtLnmHpt1/PugsGnl2Z4FPoNeqXoIdN
H+oa/+HooEO25o4ctMUIB5iH47YGA1zxsQkj6UTccg/+57XNLilFtbOQp+nIyOAu6XhkgtQOVK27
D4io0AC1HvALQy6omaFqU1ZJXABoGEd+kKyRoHNIGFQo42c3S/cvBD2f5XwrmFoOgo6G6ufyDfii
sqQBpINcM5CQNL1nnjf5FGeh9y1JLuJ5QFNJCN1hmUyD7kXR0poPs2aziEBZIikqIiw86S38DL0l
qa6rMWk1AfGaifgqwPxhZ+ooJfrZ3LuEGdR6avHaww5y9Qu0H8jx+MRYc6Y3wj8DOjGSaI9BYfkU
AvZZJ7VVCK1/YwT7YIw+QfBRhqSYW7jqleaW+e/OGzcCdtQ50cRcwMutesZ5yE4MD+XnSmhiBJEF
diWvjMyg8Jxzs4ZDWzjRB1RyIdjyNMJlz+Ic0ulBXdezYu8c8c75DuueSYVvK6PL4hKsblPdBT6S
K4+uWnyh6yymcPbiH16RtGSCx3WauZLP6R3qqipJ2g8Ynlm3OrHCCDICa8midh4+7F/2Udbw+jrr
CC5/bUWj7cPzKqr3dRPSXoF6+lPfS2p6EucOD3ma2zEtr1L/yJS/b20ZHMOsXoOscJywTaCOsraW
GsfB5LZqapGHEnz4ZZ/JztwWdkmd9YzCtp2UamM4uiT0gNb6L9uBrPIiauqLXZW2Dc8mYBD+KndV
nB9QD/Bg9UBStwwAFHV7nJ1T4n766u7UYzJhDXS9eX+xbGpKH3998In7VKay9M9anii+9J269/eh
+IKWTY6i94TOApwqQ4QHqDZ6rIS/yGthBk5beyvqM5ouPScZg1exeCIlg5p59qKHt0k6qtvnj7Z3
VN6yBno5KaCzKQS4S2xdSlKzhYYCfA1TC1wMDaowq++fP9cBao8HWyM9fNkW4eE4VXGI3MldRclb
FMdp+0SWRcJsLVzhu9wZDS3w0RVV4W2VGVJ4qlszq16nHFEJAhvv8Dhcj8inGSD+cO9PSbMYxUNc
1TMoy4IoAoUvyqHAPA57/5EhajCMNv48iMWh5pF006hI08p+qOJwn5gt21GZxPAdGAWjUBJaeuZP
zd9KMiTDfOITP0F4lB/7PElapUjbFYn5cPfMvrv6K+orK9Up736fVsTxka41+hP10uUj0oa/EQgF
NU5gIEvzIQ17rrGzkDbslAKFKmR9liI3ktY3aoYvUnkSyt24xjxDz1FkoWM2Gl0WdNmglcdcgHqu
v9RbkylydR013s/v5oZB/WifSQcISZTXFSDNoK4WqK6Z00sVYro2ysp11HTUJGWNuenhucpw5V18
DPeQe8+lPiqoTq/7V0MrSHsLdKResvi5SbJOaucpk3ALh/n+Db+TRLDRP44r/N9nrOl5Liyo8IWI
vLYckhybxMkNIrl4yDq3wJFTQiFytQRLwh6pP6YEG5LlwQJF+Tqy0gxt5IVlf00NYtaJCoFb3ZzF
V2ms+Bs/p5xftI7T4thQcYnHiEJW1OSwdyR3knpBbt3TyFV6gi8oyETfVQgFs2wwWypzDRCZmTMb
vTJV8O1O2HEBuodrhhXKW1+tl93/CWccD/QQHpvHaz5fiuBdI3O2Lk9r39rV8VQpsJaQhnMt6OC9
m6+7V/Yspd71eq2b0NBIuTWt2avJz9J8d8oeuEsTfBrp7nfZsrD83LRPEhCAUIcirNklRjxgBpUJ
upufil89aGEXYXtZgSwA07+M3rEp7UreY8Oqi3S3k53RHHK0z8r/xLIh3oBvo9rw9PwH6twFFsl5
duYM7r0QNYQ3CRuSjZYhms/K+pAKiDZ0UdgrM/awWFxAaIr/BBz4izSM2Q8j9XtN/RHzYRM+fQyu
JyxOI8yRk05FVKIDw63mwv3BI7ilg0peSdwf18EWSAAYarv0lG5AmWAKeMYcmrdwe/zhdngukJnC
n1jhbGZZQ8LUw+CkNNajekj1N+Cbk5ScCQYFRAS7t2uLM+XkGv35zMebzzDyUyWWmiTCw9xXyhGx
70/eSdrJY5XPKuqt7/2FZUMUzk/5B2UAP/HIuHFZmBstQ7KCh+6oHaiig+QRhT2yzSw+FjK5/iwa
TwRnBGULJ1lnrpy7okG5RiQkBWNChCkvEUBNXHRVd3ww0SykHdS9Gxl3zUQM0eObTq5a8LIkKgF6
8PILakrpQ+oRgEg6nov+qDxynYDwFEBctGx7t2tiKgkRNbXHRMw3YIZc1nMuxMc2+zSlvqBMIdq1
iMh9wglODGkUTrqwqqYWuZR8hma1m8Nav5enqwsuiWlrh4cYc9Ejo2yjxhULfrnZn18Ez4Oj5FgX
xuUnOK/gfz9s6/8KvJyuJPi3vIQfk0g/IzsTsLMFrCYU8iqpc2hhLIhSh6vfmUXFFlXK0SIPmyD3
8G9NvXdQChp8qbXwVjRCUiP8Jd+ovE50rI+0q5WFXJiWOkRcLhtU9ozgTBwKFbrKxv7+/jhL5GE3
/MuOBZN+TTSlOh9pFi9FasdXvLlACXpvBVeY7RoGhLi9bs7KGzel9bCmE2s099Y0ma0TRbyn0rCN
e3FO1yVpZjnSasuoGIUzFnbmguTrjBwcH0Gqijk+6IjDcJvkqVZd4Bxiqm752OFDmpNs2LWA38tp
71p/CKAwQV8WpQVcosFYUoKDhSl2pj/9LyB9PFZAXNHc9eVFOK/7hsABwLq20mfGS1xgZMgvvibc
HxvhpF65Jztw7VWXDNYF9/L9eQAuZCGmQxL0UXPmmdPPxEUgE9C/glbWj43E9TMBRURdF8i8a6xa
1Qqoa4kBZyOlbg4GYI/7Yz4SRB5sGBIJRcJjj/KPwM9jHaG81TK2s/6dPK4BSltxNXrACy+EPsDk
h1lxOm2pEeo4GaKIzqi/QOMXxEaHM1DSpqp5MLHGTC1yV1LhNZiz7N71Bd3CVjwvA3R60J0Ho/fk
k82k3bfxzTs3M8V9H+0+AQJasMUn9oWO3p/+Dz3GxCjA8CNuqJWqVzE3MFgE8qKJ1qOI1l8Raz8S
n3k9Npt0bzt+hXFZqj5H8kzeMKvygjxT7hyig4dAYwnvJvDmW2BhbDy3QVZ+kR9CHf7q8SSmUAqn
SvuttOQsgJuYzZNChm+BveSaCQ85YkctxcFdY8PcZvmhi3r4krjf0OPYWh396g37T457ogKStvxm
uxKYUILnrqBcTi4S5+w1KDW05IIVBGvq7cwFflPIkt9Bj2553ZMBdguq8ncK1ve1ZP/Twbr48BPq
Bws1+U00jgDYi7qM4WBrH3lK3PhQvy+DF9pVJ80l9HmwlKVY6dhLL0XooGY9cjXZpVEKGpf3MQZT
c9QbTHniGT1aRcvDogVy+RwE01kN0nIbmiPKqWVt6SgBOFkbyYPIleosAeOTCdxD0sYBg9s3w7Hn
jGpccGUv63KIWf40XNqU/5mVdN3ZB8L1xN2UXHig4OX9witYQr1e6w4rAtTs36L04A0Skn+sYdYV
kAHs3fzUAY6eDiBXQ9FE1wdP6zbMtLwfc7y6vkhXKq+RvBngyvivROo7VMPqTZmrjJEnz14JL+xO
VPRLHuOSZh6k6d4VTCAobODQeph2yBtU0kizGFGWibnVx2pwcKs2GRGi5MfnG2JdOqLBrJGKn2+s
MY4HywpTF5tHypMruW3KhUGf00EKRFjnVfBW6GtewDRsury3M6pnYIv7RkXyzscbxhw5eDWGoK7O
XIw4snX32eTPv5lo0yhomh5qMa0EW9wlJdGanpLG3yEJw9m/PSbExEEYQ/Z7x7JHBxlLfzcq95W/
gc0OwPso4G9dWsv6hLpkw1KZbUL7vMaXZPEwyQf8P8Hh2Kd1tgwSXH3uSnNx2xQLY2au67EKbgOy
aDMit3ohClRkyeypAjZf0gtMnCOt+1C05BCmknlUGV4jhSSiAdC5bcj9YhY90QWl1mX132trCCbB
vsQ00t8q6V6xn7qbu7B7x8/YNq72Os/trRNwDt29whQlKbPxa6zZ0cF6SomNhJbqTGqZATODwWhu
yORSCZ9txHm79xpDq4nEt7a2csltXgZDdLQl7USE99MRAob5JX2tp7nSNJMSRefTaYH04/JHtYiQ
iZVxxB8/Tda/a8qwh+/encscap4X5x7/NWsULxjPLDtMknD14//xOnZsaCNjKxXGBRKce9spxWny
pgPHD4KvNinY4Cm8YC/7sZBpn+ceN0O97QElWWYtqmdZxOaMK3E7wgRZIf3kglByS0nxDOm/a+dJ
ah1GwsxOZpj6N9DSxy7bQRmNblimnI+HWQ7jmcHVSNvZ+iPeO+PUbMDwunOHUOu60Ps8R25ywpLa
TWHw8A4irh8405UxuA4/kIISbYEYTLAGrVtfzK2UXz7IYBvV86GNGAGewAaYwUIF8o8O9yP/xD+3
A4rHeAJLlyPsMVwcHDhHNnR45Nu1PQ72wY2P6dVRGv+8XPPMPcvgF6iUbYkFx2xBSRJykkjXXmx6
5biuzVaNYgeBZlXtKD9J2VoA1AwMmMg/PFiJ8B4FKTxmbo+68olxcKARqjYCNuOj+wzimtTm35Y/
+4f8AsooyDZ7JG+WuF2yNURP2mVv9QtciibBtrwPllu2sDuEcoaOw2INQPlU3rxsgSZwgoBN0K8T
LxQe8zhI64LjlAgLlJMJU7qGLUaBgf+hZDOAo/QDAx+a3cmn3gOa+UQaKQu0ZuhcCGNzyrJ7eymn
CmfonBGvnzQsxnqXLlIrUTBe3F1QwvSa70ryBwlWBYEUUXd4Ath4RDUqrbG5k3cIplPJgxs4om/m
fw53wTSnJktzFmmSZh59Ssal1SZ9JQoVM2Gus1GwEqpio3eh1b2MGOhJAq05YZTUPiTvL+qUMym6
4Y7frq9HFnySYUXHn5Lh7EG3DhDuOYUkpXuR18t2vrFrD0aTg7OkHvW19Yr8NVsrPQPUKQp2Yu5/
PgjodyoXoY+orFyd4wi0KeE06eIltZg5ydjrv3dKywrrfZeoiGGr5uKfF5udjDaDGfTNz7KlvSKk
yk0NBptMqmTFlltAa66ZWMwGekSHelA4j2/yUWs2sCBnJGd8Dd7vS+c4GQw4EWulIQ90BWDJ4QhU
Hw8V54IO0RxjHi05IyF/TqIo4yIoIkstc1YUWVrJgWyivSBvkm3K5CXLa/t3pdpzMBI1IjSmLOn2
Q1iOdGbEk39G7yznIk9Ik8hlleNnQvlt3ZyqASH0NR0Z+ECI0INRajciQuN7JpdvyxCZVCOUoCwz
Hp3lAXVXHIm8S7bEbzfagLRqCuKNpX5s8UwjQmGZ+s0TdC4Q5adX3EVa0Ms0awCWnemOSgqvUBcK
cPHhIv51xDZpw/eTTKYMNIYogsTbKvxkMTIeI6Khdxun20NdKgPOmZcF0SkLynPwL8MGXb3DfyFU
tLh+jBrcDQUfQm6imUZA3tHWdxqKPV57UZALIj6gTNgRUIyD3k5z6X3l/fCQYA1ixwbyv54H+3gm
Hfm3pd4yNGZl3+6QJP+9hrRtxNamQ5ehun1v53qvJbEPwmwr29k3wh9F0uuYfWjf6+b9twb0xGse
DpIOFsLLR8GxFqYj2ZY/6UcqE5Vge49DqxKHBsCXoZqqM/EAPWveq+eEnDCia4VT+Rao9G7XSW8d
GcdW/T2Hkv0Q03VQbTcRbaTO7V7nuWge3+MNjC1Rj6EY7KVq6XF+YXVNdqvMNfbQQuWMGiAbcEbh
ukeRabPpFBoe7GiGVN+3Oj2IOQhRF6kL+BBX/2XfslLARTeLUScn93go+0YFsnxTyCCaTetls103
T0TsS3mAar29KzqFwNqlkDE6mG5QnMTP35erOdDzZ/poS/DrquZ4gTq1MsEd5Lm7iAYAXmuu5i8f
ifXlh9Q5cB3eHqmRme7Qi5qy3pClTU1sI18gvWSuA5WK/cuWnPtK4Dv4jq00Yp94goRQvneK4vXQ
Xgm22rFPJ/EKyp+RM0ixgh50nbUdM//2XZNmhEjbirdJ9XQF9pDnGqqe9ccXMcDVC62NhxxFvYnq
oDdsc72ycc/EyRDH01lPiJNn+wtQQWS/SrdAD7i5SNlprR0TY27j/Qb0YZQXHcSkfK6mPk4uw8Kc
j5CB9ycupb0Gj3JJSNI8Crdz2aFZH/F9Qf7DcWYmR6avVwJwPwIK6p4MhjG866dDorfGw1yLsrIf
v/7ZqcjtssT9OKg83pDtjzsWss6YoxTNjJCgRKewWdy/DQX8kkzUstW9wsCbeK+8e0P4IY1EN3+T
Q8E/fvoGH5bqIbitVXQCBSbOUjgDQh5mT6kyoSCl++21l7VHJp6PyLR2Spip/6y8jcyejD3+Wzbl
n9UCkNNQV64+aiYnyZuzkBEw70XXHqoD6sQ1Tvnv19wlmBz5ArO2scw8GfmviVIk8YHo1qKq0X/J
3hs9Qg1LO/Jf6jcYM5G14Cnl6Czw0fiWkPWu2HRZUysHGXIb9XN1Mn1pd+2uhyQ9euti65c4o5N1
M6QIpDbDPRuzFudB83DUNwipqQRdZyharrKhw7gcqQ8EGlmDB6berob6hJ34h6mL6dDOqB0JUtek
C7Dm7tdarW2NTWUL3g8LdE9WBLJpuvlxx3eRRChj7Wdh8p0zknZnj+LYkZPIlGOWx0GYks8E065A
VSWt5IaI4ZbWSTNPa4i8SO/FHLJv90bqxsIGC6WC3Q1Nyv2IwC3QAbGz+RYwK2CJdegvo1vNLBvz
d5aF4b563GH4M40eUWDhUm7rI6Q7M9tlFxwm+NYk/Omb0LzlXE17yyNO6ijFuk7Bzho+Q1Wj2HCm
OHtiW+Dmv4abhV+xRV6frJbyZxRoCH3PfalHZaSD73d0BsP7qZnHV0qKuouLtK1Whb0fRzjDqgCa
Ta1F3sADG/BoOxDRt5QvXGsTnJ/OpEU0Q+ttU+KRvmx/qP46CdTnin9Es+tacsSo/KLPoZth1UqC
LxGMpIKbxdYs3qQfevnkXF626AjBjyCN9FdF1d5B+yjhyphKJ9GOJMYzfgoIMQjSaYWrhm1aiTON
GkGomfJahLiWBXEuO80+lmLmVWj9JghzkMUl7BcRpOiPO9ZknDRt2mQ+ns34Q3zVs63sBaHM26qk
Pk9bkZx7cC+d65fajrLMJseShUB5eMaJsqOkCmX+iuEBsUUp9d8jyvAi8XoqaKkYW1qexz+/QY26
PPZ1ILmtgTNEYQQUiKmTB+Dx6e4UpkwoSvivzBNjyX7jC+6r2M5Xld/yl4xkoEEF5+9IvwhRp5+B
GGq6a+NKoVwJfpeGP7lgUAZJwia4e0LedXHcUMW9ZqT2enLHwX/3W85Qvdpl43CEpSsvPbn5tKtm
OJQmYvyr8PI7VglbJqzJcUxeYvCMpVu0oM7tjiHDNeGBzlxegPyI2b4b/RUOLulP4gl82NcjXrr5
9eYEloYOLnQzdeZTrVhQSOg1NsWs/tTxQeG8N7L03fHz9ncXzhk4f0Yw8Rd6kzlAaJDzx6BfVPp4
5pAb3DwHTY9IlKHq9Kv/qqwXl+0stfE/ZAet+LrNshUtJjFvFEqiRRSzq068XnbsyUhNUx9Hy1NP
yfrVb/dbVTbKf2Zi2IdA3T3M1cCWBALcx9uyhZBeUtw8M+P9o0DVbVUtc9rbvFtf3sBqvh7wI+8z
y9gtd8kLD3qPsojAJsNEWi6tzU9OxYwXybjYTlWQePQj1JfeyzHhaIu5sUKqcRwpstIuv1HGlvV6
qJEbUwbLhG2CBLnCQzHAeQtFcxDbjVYob2PdIClMYfUin6444uqqmC3McaGfugl4DEl6/mQ/ZMzM
xiDzZxpAFqV44PMvFbUuaL5UlA7tX4FqRoQ2bCaKMb4nasPLMLEAuSfEgWc1qYhJZyFOk/sNAUQl
3tSB7NzvsuJx/0OnACe+/q0qmHHgP8hnrUcrre9F91nq3eacRciaR20oMUjz2pXkWqWb8+W9vMG9
pfjbbhvPGVpDWUNoMaCiAUBS4ZzdxQgnohJ+7WH80LpRKWQ3WNnjOiYybGroi0UKsZnOek+to81a
EaV20S86h3tuzhNQRh6x5r6rEf7867nSjhY0RMKUXppMGedmLbpCPG/k9Q7J2YBAwYPqfT0tvqTV
sX8UcwUuMzuLoSbahhvR9AcBWl/MgDR7l7u+1Tpv/LMtWk8TXd6kmLx9UIqSj0YUR5g2yf9QfuwC
MCHaMDPeZSp4fHQaW7PPsU6cJHofY7lZKiPRdl3lQROWycEhqNWM5MG8n58JpMr3zBW5Y0wbAK+H
VqPnF3cQaVASFtkIdVgXbODaN+LUx+T5PEUgmsO4cp5i4kRumErRcvuAvfXd8oscMC5F9mKiju7R
Olasjl4dmWho7LcsmacAFTLKWfqDu1tN601R1taYMRiTvI41ED4GX6RS8g7mCsxEwT0zgR+dEEVZ
7M/4Dxy32qYolVxo5zxKZ0tgRlQy+HUwKGMoCIc9ydwno9yg4EbiHXe8wolJ8UsDJ9Ragdjnhp9v
QAUNfNzDTI/2MBvDSjdnc2CsnjHqedsy4lLn/wBlqpiB4yFkL0+RG0Qqgc4ZuBRxZeQKjXuhKFTL
XY+yNBmqF+UI9pS0kTaQ/qFsLWiz91zFvSHfEobEQ54i6nquHRxhQijVz34e4VTUcMWpj/2DW2KR
qNiq6nQid70wVG65wrIc1PqFCwo7xaI7rz9cl2Jz5nnTEfWqwB+/Dpqw2qK5USrUKOnQSIjGqVqD
XDpkIUw1nZvb1oJqwo9ls8aZ0zpjReyTAyVm3JImDL/mhC/VmLpS6j0CB5KKb2Kk+EkWB//qFFOr
WXK1zgWKQmdRRA7Y3zktcmR2EHIzYmPhfFaBCOLAe5ISnR846fD243lXirshmFa1R/1anmz61QDL
j7GxiDmJDjrSMTgOpeZ4AZEQdcPJ3aQEnTvwIKS2mMRrsE9WgNSyb2ANfApehD3FhbRmdst/ycVG
ZdvbCExl3iL9MGDGL+JLyHWpugPe0bOVQrqu2wcsi6Z1TE2JN4GrvaHJn/DdShdmca+xExgth/lE
HlxX2q2slYwOs67cFB0xwnqZg6FfBF40L7g3jHfFldNCWw+cpkTolDc/flZ+W41O48DtsLWe/WAP
o50fM3gPwH9PeGVga2PgjXlHmKtmmQf73F9yhlG97k4wEwdL+UgrUOd3ScWrMmzZ8R5uC8Y3RofO
uDj4dwnfPOPEeLvmmFzOYjRrVxhW2aNM95oo/ZKbaMH85bC5tv9Ak26rUN2SlPZMATIaQBApnqQc
2kFfbPdWMzo8nnFQ6SFfIFCRnW5ERDRq3YXVDHVMpfMW8MDpyIFmrLJLuRlP05THn/iMNEalblM2
jAPvyUGOQWgSIsELutD9KYuC9JFv+iAZ5mp9L8BKwmJkDEvJBr+FJnXNN46GtNiixc6aONMKELoZ
s+HcL677zSOf1SrSUQNxGUQ3U31HmC7X2ZoE8lG8OVT9iLucwxpjj43Fa5UQ7s03QlQ3cegUubRh
b0wCmahYwphy8a1s0NKTj95gCkOHx+C3my6rxPEz5jCsEZQ+/XJnPlgiJPbNyc96Qyr54qxNfOVk
YTy+blclDcjrToNMnP35+mppsGu03PF/ATNRescW6VZNfHJeGkQO40X/2z1/HkTjJhubj/SAe6jZ
+P+GfaaCFQ5KhzdQY2FyrKQLhF/Mg77iRxi+986eqG30Ue7Zm4yheO4RKkGkYCgPMGBsxScAUXrz
DbeXWShFF07N4OeA1gzzTSIIfekhtalJR4woU7ctpORaLdB0Mb9n0e9nrCn73FmqywSqC6OBffJ3
fofOST72lvujTcsk1xBCiBTG2YMSqiOJWrTnl1N2pDAubyTEQ7mqoOIxQvp0E60v6PVFAUHRuSHI
6PQjaD5TktD4nMh3qJbQPhX2DJKOXSoOyy47pIB28Qgb608ZUr4Zov5muiniqsplczUWAm7vqDfu
nndIhQPdm3lQ1Rd9SHtiDotE9N76ZbQutm4dEb2PKAu71XXt9omEylhupSZzT1s1LxjviF7Hfcr5
MEtXKtotb6n85xN2xMnw0Z/UzesRHbNU0QG0ImwNXsljOIDcifVQVkAfuhoYzUISLbjKAnc7h63J
dsmVVE6xB5rNnVyzxsFfOnyHCo7O7OjiVM8cjdnenGeTqzEzJW/iLnciIv0C9hVxiOGrY5jGE22c
iBLeqI2ldqzaJUlwZMirE64jkFfd+cKwDwXC1BLUAW56MReixQDnWRO+MjbbK7WoKzNqoJZnbB4l
2EQnoqEZvNlv+FrP/J1kQ78i1bUDdjF9Ow4b6YIPyIOs3SN4d+yd5kGiQjVhi2thNcNAwYcYkFUU
oqDHU7hc8S1jhMrorwisI1WYCd5rN9pRmen9CYFqfCHqjwC9i1QujTDm7UBupgt0FzHg89SSyK38
J7xbGSklCLzlUiQTdIJXWTVYJ7Q12L8xNuM+tzVaVd+5WEqXFjrQMW8aDkYBvCFaI/bZLJmd7iqy
kUCnIKBQi4DO0f46W3lGh5CX2ep4wcHz28ggFiduNkTd7pHt5oZGb3UeIP2ZKPKbT3KKwF/3Z/ep
i05kc4L31NqpbB/5kj47I6MP5v39B7lIG9+CRXz5fmwkZ2oz/8hfZyIFrMV78pXJq30RRUuwFEDi
Hg20rLNm4TuUQMnm5MDstBpNAqVUwRyUp8bYeJvAKSuQjBNxzSDyps2cpgNanHQ7H5YGlFNzXLjc
sOW8km5RE9qL6yKgtTbtkKomrX4JaMvuEM0zyl0z01jXeikYmtIAxuYujPiQVD7rgQqzuR925eTx
w++PkVHLGE41s875Fc5cF1Xdo/jH1Ln8bEO96IvS/HnwgeomghBHBP+Mc0+Xa4XnmwDBLofaeQik
CQbzVatBaCo8F40pN7JQdIWHB9a3503RpXpTiL/uTqi9bChKPgtDsMuXKFRFzwViT35dqJuL722O
kYNRiNSATA2Ko42z66+n2DaZrxD8legdybCvf6+QpY4Nlh7B8AnsbJMi4MYbxXovNdde7OQtgP4T
IFNj88rtD4bnykT2wHpRLKkKr5fgvNdLRT7IORXDaADyBRKKMtmrIj4oE+HlblgGKuA8PLaFocXF
jsoHIfIp4SszR6Br9MHmV1CgXR9hTvrT4phyeDMixNDguwayAeoBrW0I4MPtbv0E0WVcjYKUFI5c
O7E+Nx0xYmGoJq3zQ8U4mWXh8nQmqQZjTqBRMmXq22VnQDvr3TwA25Rxez33lPN0uIoVV5ZkkPSs
EpnFP/4TMCG9JR5QRPQEPliG0Z9OpwYgvu/RoHMQ1ucjn0ZuTv23uFWOzX9TNNtb9dUjK02EJTDp
AZRE6NKRB8/s1uql1MS/RxjVJfnTCs+7mpZh7gi47QloZ8IJVzwY2uCYlOkQRNveq2NQ+yqqPOQM
LXypnMH9nrHTwlASi5/cpbXWKaOHONXDgqqdwcpEkSg+3ja0a0v85VvMa88akol8AQ+kniJedHiT
+FV8YYFA6UuWVLvXrK/Ntj5eHln3C6mWtUzpXrvjijgGBed2McswvYkqH0m5wMmqXEMHXd9SFsQN
UdhZBOtphvLC4MoZjrb7UgvcFK83iMBV62StZwQsZiZttdFKP1mzx/jI0MhwA0I14N58/r5xpGvm
5uYS54afdywVFb8UcXTCSAcjup++SVX1gKcaUnc2ImF8hwn6lOEIhImJS2LjJE98i8JV2hbnSQ5I
FlFz+YpBXDfAzLdRnOo1JhWn+MKHhYGTNfAOnzs+Ke1H4orzZhKg/cdrPSHXRa285qLi1Sh+1/7k
oxAKNutnxHJFRkiPgEO7CceEC4uHRCggYvkGsuelu3tQ8PqsjAocYj1WI3fJYG2sAlxlwjkRejNL
52YUMQj9jreU7VG7mFaYgN9gKaEGzOUAZIxAyYcCrnsnDQn4OyBCUdWM4LVTvK3mgwgny8cIQxGf
Bfsmk8u9jmjblGcpqx0335AZ3abuRFYPsGfx05klI76wmYKW/Fg11zzGmOGaHNUQMpbW34Jxnvcy
OHRMDVfRznfsaxK/BGiFbjl3oSh7fnBh7ov0nc6v0htKDb2G/b9U7zIBU5c/ceiclSm3clboPGoB
9GZCAFE1dvwBaBdePB0I3m+L59syV7zUmuep4C4kkUU/gQirrB8qd9wfAnJcyF3wL7fCgaAbUPwE
+OXmB2pXAnafZwA8I+dK5u8H5wzHQU57EXaRh6YvvvhvIqfPXFB1yA3pHXEramESnj+4esSLNT/x
jJjP6j+9vdJe1XIBnrxYBR1T5rY0r1tlMdkLQ0mr5K6MGw+ldxEwqsMzqOTDdZNk8QLeQ/VBXqET
uOFbRmIEvWi4hNIrZXz5Y8HPG5SMo14z6O9EXFnE3o28NwF/g9aTZ3yy5kevQFXaoiXCxdfiS03Y
sIWRV21fcj6ZFr8qct3qu86yLNnNLHR2cpy8DJ1Sbjpz+svsr5WhVkaMAbok1Nu0Rwa51KsUsveU
0yV07w1tMstORKOilb/ONAzJc1MiEVhH2I0TCFTBRnTpD3ZDLx3bR5TP0g9fGLr9gV/ddlzXFXM/
5zy22KW8GMrsHGCHjCOMAqLT4RvCDPGE0CmOulOQ6bPVU1N2HLYyTwd0131xNJDvyr8vccwYpKe5
+eOMNEJPL5UlODTyAKC55x2xVvzodUW8NDD5B0p9ehFm/ZRKNc2qgzfMoaR5oIIML1ySQMePgXIF
nNzr4pS9VB9iMcAthCv/VKD2C/VaeCw7fKDPjOPGSOc1XvkReEoO8RP9oA/zjlbLH5fajEs8WV9F
Hot56LizdkDTz2jOy6t4qjT+mVdTsKaB/pxmB3RZSCxdC8kFF2wedQWaTEMVB55c6ZI2n18szGbV
wHLgANxl4Wz8TtHab923YyCEjZAc0Y+VJ/m7LjyV+YdIh+J7usUQKSxFjUF+UFDeGLIOzzYNv9+t
z+HM+BdndN/Vs13Yv1RB2QPlUlgYbBGTmqD1HX9+5CTwOczsZhitvOrXiUnlzoTPA5NPXy1AWvJh
9JDdMUUfQDbApjXrHJRvOw4ghuC1nPmWgCMqQC/OuaXr5FNVYyWJFK/8njSbXwteA6Lgqzemmuen
diR6IA+kGzUbBVCnwC1zSZzwNFKOjtlONHx7J2pSZMfRKOo9BUFXhihLxvPga4BxM/RZByORYXF3
U3uc6pSoK75vFbdpsbanAOLcpqCm1WL/BnFtCTWZpVrrbzHHnyc/VH1bQDw6SIGT0NbxEWXp11tb
c2coQbyNK78AauxXBWHEY+zO0mJ3eMvuE0c4BaswHCDPw8CUnGPhq9HnsB6Yg6MKvO6wc/sr95mk
IecenO8LgEj/8sZZcI+VlrL/cdDL8pjHLRzCe0gpO13bIqe+2zrBzcYjcY+mOqDgQ7S/2fqdThVa
RNvqrNXoeoyk94NRGAvMkB7+eFnN09J4REMz2rYbne1reyEtN/Wse281e7aqSC+oIo1MkJ2ftswc
QIRO9IVUDIucJyPDSchYg2r+GLvDbvH+/t6vDutDvV/ranpnerKWTRcD4FY3DmY5KpaJR2qVmjPD
qWtH0IZXh1Vu6uptwQoZmIyYSjUPOlxpJPfa6gXyLP1MV7+zHIFJ8bHJfEOhMapQxM2P9xkIc6r+
Cgd4P2VklVvLtIahWJvxk1acwr0ksnmlQHgBHMDTbQgPTc023BL5mEnlNnXurzd3IqbTBbG+IuYY
s2lVcslGkwJ8s8FbxkBCx9lDQxQOn+Sojeg0X0l0tJFSBo3p3Xn8H/zdc4BB/Oaigihs9KiQJ0Ln
CrGCOnL3ioPRNiOXygePidY4H18RmU1zwv+Q94TZQSkEETP4MAn5D36mh0rOscmJane8nTmYyyNi
H3wl/P/+/00DYU+ZxmEq1clPpjEEC9g4Ughpm8ZFMgOnePu9HRV8EUThoEaUwE4gP/sD5NLFWrRr
yHw/c298vy/BLevzAc1C7LRyQPWl1nn0jirNlIqc0BPJi2dxwPhAFOJ/btMahF4DWTdqJf1sRYDw
0+7uHcxGQn9iDp1z1uqbVgg7RX1J2QwTdWuUtVIMqV2fCIiZKQCz2ATLTnswthbJ9VuuioS0Q2Vs
dq0nHhJz92XGw61dqY2Io41cNlJqT83hQnjh3vLUK9+PL7QR+gTJgW1PidJ7n9pR99fpuasMNQg4
7xho56MG7zARkTSYyTnP27V0JGhsIzIlyJxYjXGfLn5BsFCGqjNQc/2xqVVpUqh9Qy+I4LUSA1W3
PJLjVMgT7LfdhTrCgTjboMVTDyah3sozA5X2bDalQaSSF8DKJYVn5xd5X0waJOFxVEA2jTBxaMKm
oB+C7HRsFukQIQkxf7KwPZHcmM9JV5HKRSQY1pTLJeTP51G5mHOhdPxbGhcf4nW5ypI8Mterx5aM
A/frPBOQr1bSXuuMvdA8XLDnALX2XgSssqDbjb8x78nV2aV9KWhTZsj8AZ8xNMbzqoyF74WaOALj
DjGtQaFhiQUEwts/GC81sbLaxZgFRY90jeBQZyINCAlwWTNmBVBYrk8G273Jee8pw+ViseHjJfIn
EZ4zxASeNF71XQfrU9Z1rBrw5OPxWS0hcHm/jM34v2f/Qv59VPGojcS60NVSNu4itZmFeimU0YLa
xQ3LoWltsX8iE386LHiAJ/vaInFvrjPgOgajnai7/0P9vQrYHb5+KgLpoBfCTtscghfX+zh58tjX
T4axMuA1HX+DCkyr6T1+1T9QIpcBuaF9Vig/Sf8AfcuFhp/qgs6G/SbklIFhajyrIUN52XktgmNf
ms9C5vYQiMBK8Er3lFr6wU52VC292SpsuTf9pMTAOOJ8efos6aMtoAdVugHOEl95ucSnU0rTpBL1
KCixu/zL1tyh0nUBkQEGcazTdmwXc998XPzCiyLr2J2INCfIB0QstADfI22YAGJPpK1mlhaxtym6
kUkR56MlMUPpK1cu4P1jLvpus2UfkOpmLXoBMqKQjR93cNbkEDp+jqVgYTufacq9ie2Z/TrCEPl+
MxqZF7MQG+gHbcsazBNeRAolX8juUVPXxBB2BWPcbL5PWQUj82eKWPFSlmS8nPFjGUo8StXIBIMr
njRh9EojGIHSUIQWomOxrtr0P62V2z2g58xfq57BNThMhxiU1Vh3WqUectLKyY7BXaSO8py1dhLv
NlfnAhn9yvj0uvRjkb+Wlo75WHQL5lZlaGzfeCwzY+UFqdF5rreB39h83hTmFWf5WmFCtL5VqO1F
43X6E49TzY2ujVe+sWjBXYohX1+xFw6flzVZ8LaDtpcWmKOUznHKrOG9nd9XhkBVUekGq/1BU8hr
zBO4feunRzEFgHGboeaTl0Eo6RSWvvyo32dG1ku267Pbq1mEod1PmlbTNPlbZ/ntcPqBskNFvD4b
tqqQvc5KBfS844uAl4H82hUCwtVnKQLFWH4EcVTztdc93buaAdk/PlufHL+AxNlvoW5FQtnNg7CR
HToekmZs6m5RjggtaysxDjzcOkqM7cJOAI37KlcIXj0+MQDA81GqkpFaFOfhMgbJSvt/4SvmtNBk
noGBewIIfL3XVg4rdffYvSM7MKn921JP8IIDqN/md8qMApvbUuDoA3XFAt1kc11LslaPhaYKTCkk
26kk49x0D0+Ro/8ScYAvGY1b2OiEGf8RCUvDgaT8RgddagfX+TSDTj2G83ViodRlgveKxyRe/dCR
vN/qsMLSpqgA8T1BiDfnrOT9Ub6xFqDIPcZBYzA9aflKYZg1oUll76+U4p9znPpOy5fGkzVJmWIv
/rzHnAMAo/+6N3FL99MyrJYRu4wS/kCbJ5jp4cHxjoNF9usR0ItY1+M5LM5lAfhq2gijuALXlbZ+
h73Wk8s4Vyi88G3HSuPKPRe9k5Af0xoVR2cotIlWiFgWDHsk2lRFGRde10/CNNN6hBkYRJVieWXX
VSjsyW4Qej6h9Oyv489BPrNKGZYhfV51coG7PQ14LPG3vN8Xh4Yd21zYYz5FMVrtsstYax24pc+Q
duOz+fiKkuh7254oLuVWbSkbg4reWyu7KM1MdSaypzq0DIFeznV24wIKgZdYs23YdKxoRBia+IRL
XrTo/AotBg4zm0wV3AjpGs7lVw3izWTQ95aNDzJRtST9KfUbElS4c8YlghJ8m9RmhhA4XlqubI5e
Z3T023+XWSNIdmZcY4mFw4s37FUKKAmmqpo/3Kt6o/e9NbLM8WQwAhlcu5b4c6DCQZMcgSJmj1xV
KfLYb75pX1fxMANbqDOyN/XZGE+uJwQmZZWmbuyq/O4XMsE/v3J5KuWQl/NJlSg/mU7QOC2OodW6
qcwPUQqh/14Ltjh/ILfgkkeHqQ5BYoVvgjvv2XvQi7hUMssPU2BjRau9ptwo4C0vrf059yi8ZbRk
dU/nFNXyJiGp8uoCBrNOM0WWsxeIe6t0mmQTa8A3/YnDU9u+ehmZRyQ7RRsZYQDup3PpYNVC9uxE
t8mC4M6BxMPmMBmiE0JcRihiTrWRYjKUA1M5oLkYk6cvAkhWKzXRYzA2wMOIciJvzLcNCwVK+0Cn
XfATfekz/5v8j7dZ8m0rGO3gN4SIflZ+/UZEuHNWn5nTIT1Tv0d/TRcp7+QmQZQMeMV21+iwpD7s
CPSw0Iyhxbz+UhAMUya9KTN6GQs1GZzsuba2hHxqN0wG+qTZ4hFW5mjcVe8xC5biAfuzGdJaekAT
dDnypVwxMsJqtp+jdZXrsWPUY3DiyA46ltiDcgJrl9XsrlsSxIJV/Rej5f6hGYOjXqN2svSNZiGv
GHLwjfwGpjaXzjfkyXmePIwMjjRnoheFR0+QBC+U8zzhqz+e4GeuYTfCGsNE87RbRSo1jLsiPjD5
ojs0pDPwmd49GB/6s7o+saZ3WnRVHWWZ67go6ipjKNXAbdXjf/Ja+Ua7S6Fv65baFnvZPXyNsVie
Q1NDiCaOzaRnJyICTJMAEXzEmdhUUAB/b/HbTb3/sdSyuDo9RYqIHknqduq7k58EJ2D88S1ZTdwX
XsPUcBEPO2cXY+t2A1RQnqIf2FJlVwm1Pz0j4tF+VLLMPeCJ8dXQyu85bKZm21cc9imXwpCjI/Sf
2gDMeV5NoWPcIJp03HgRJpwvE8ypd6/bPN2Tbda7P6xzNENdd16lJmO6BWqj+JEJ6vAeaVdEvUY5
/KTfMtKmYhlaWmKzW2A2b3NGifC8tLkbV/sQ4kiLfehea4HpKj0biyant7+jUhrEBmGiMlgyg4JN
1hFhY0xPpkCIbFUAbX1XA4jXp4bIfs70HVeiLoVwQI9qJBbWl1mdGkLvrEn3/KN35A4zj5WniUcH
Oam8lqN9TVPeKnr9UXciyUPrTbGuj36fO2hba9CFKUUiIwo7BRtrvMa9gcL4sNrQHwh+2gwkjTes
Dr8YxVWE8wzGU/pcGulDpDp5ceb1GExRRTq4XApjJ9jDTmDI0Gyl3QCoQiO6WF5M9T6jczjlhdR4
72P1slNHPIf5cYgHUBYl5Rzzzm+x0Ia+3KxGL6l/TVd8oWUbiFXkWAC71cb1pXJO9ibyJuYika/5
6DY16u1UX0F70COwLzP31TR1jj/de2uzCv7mXVO1bSBJKnm0Yb7S4zJOyzEH7I7NqK2QZeFayf5n
lAKFjWJLis62NW0gv+iqbub5JOw8mgTAtb/mTlcLxsiXjFGOMxtfK3zIVLyKeqrvR+vvxC6rWaGu
bW+KEiQftIfs5bYX+FPpZOmE0Frhla8VjqNtPkohOW0C2SntEM4GvHUEQQGJTfwDRB2QfM2VcHMb
QnJvw23Z0SWWalKMhRcOGwaFaxFrEwqD0hTktvYxp6TyfocrzKsVMVON3TMdNqQsdNGTLfGEZtxb
p64ulfcjgcdibOe0QmVwY3AZ2R10XjofnXWis44Ee/IP3V2U0bbGH+kM51ECuE5MO2tJjiYmp4MB
pVXK+UGZPsWKQsl7rG/FaNgxGXgROHbwfxSQzSr7IC+R6cKszI0V7TKQWTXvEE4rVBSpk7UD305g
qb2rthkBBZNvEbKHEGe3+l+t8QKs2nt8UCQlGP0wuEeSmkg6bZG602zZhSQiBBv/5EGGkMxtFW5p
pm7K4R0CtVQCQX8doMsrHTN97IddhtoqfJcN5WhmRXd6xWsLdmWZK9nmx8rI4004hTj5VBn9gK4f
WA3CulGtt/4TEcMKO5yak5oIp9uLcxu6Cn0bdydUelmi7ve7+MJoMUtksgeqT6b3kfV3sr/XubsF
JoqL13jGbYdxj/yMIGU0a8MrS+HBsSlL2VMxsUQvQ22rqnh7lWVWXbn/oOfy/MfRbVUurfkyQuRP
bdzbzJhnWL94/Wdvsk3JF5utGmjaXf3kKMcn1oZwt5Z8aYnpKI8zb8kHiqM/FPPzS+Fn3tJ+w7W6
uCXyue6dmeZ2kQHMxIDl1t0iTuJ80PXByQbSzoUEPb7vPsR6SBEsvmzkp00LTQkOwo+vEwyd4cz6
EuRWAcKggJNioIo1l2Hhh8/84fXMvXc61B2xhodqdV1zhTiw6NdAjuvsCB2okEXwmYuF5OXqzoci
cgrcL5YQEjlAu5DIWYAHR0V3c+s4c/ZTk3gph5SiWjwZgGQPfATzQqcjpKe5o1XkYS4xMlzoSk+e
KTHMqMiKIYOe+5QD1lBbXDYyMeOrs8t/Id/q7hZeHOYk+Ri9mqkM+gpXsAgAX16CrL+qBCoC+c2z
BczwWbAjZwDpuz8qaLZLklJhMZ70xq+wlpp36VpAJyTXp4c1tHFbTEvn5fPkXUAh710Wb4FI5Kos
aCNDKX8PXQo3hjnN5lzKArGfuuY7j+UrHnoR23AWX9dQajw1cwK+SykcZ7ajCjm+HxFMJBBlvjv7
UNl4bsR7xscNpowLnT8VWVHM86iBHC4eIOsTWE1J2sY7fGafz6/wZDnkdICBoaybsHqxRfhr/2Sx
+zHYJPdTykdFAcY1OZhjvhDgYcnSTBusyjoswftsGKVdGgMSSsybEppuN950B5GeUZ6xADOOZwN4
d2yECS8ZlHigmLTLso4+esF+CCZBUoyMeLOyVN0GL0dBCwQPkUC4k0mBM/E+tSjgDhZUn4YrGWbb
sYN1cc9jAtSyjn+FJodDVQb3eZkXC67T2PWUXzcCnKAOPBF8CQarQt6ZOr1PA18q9nHBxIo4zN/I
J7Oc+YC5kpJNqw9k+ubuP71zCi4fvWgxaduQ6evCwgA/LxmVSp6MclqQKzG7J5TXxtfMPnmPJx/h
WkvjkcmaL5EJHDAHdwC7pGAEhGyK6uj2CSdQtT5uDTQvtHqFr0cbbS5uWTMS9OG22MB2E/pJfcp5
8WEpLbEp+TnovJjPqnedwIz32FsnsrBc9rDJ0OSLewHuKp+8GILb7DrcKobYb5h8Ea/YnqZLrqVe
Gk/T0qKRDgqCC2CBThv+lTN50BUOv0NtUCOdxPniaQQB/Qo+rSt7xOspDYTCRuJAykcnQlbP6//f
f5EXM1of7do7dxe0HfQU3EobOaHD5qterHL5FZcQsnrv+3yhknE26tuLV26cVZe0NQkmU/hety4N
Lwdq8YMrgiCGgYag+k93KxXLCnByc5dwa9n6ozYCwpjhUWulBqfo0m7bAFQ2tCxkZGnlWsYPH1I8
L61QkZv8wr8jPqa2r75xEkWlC1cAkPXMdIF3qSL7vcgUz4CYec9hskZKCC9Y4XCLFR6DzmJlYzPp
OVW7f+YG0E3g0z6TOjieJa8p8lIScAx8oEGSyQq8wQxoOJxFHbYZEeWMfcMTY5/3msdIlHpOMQCe
gEoMZ3Rz4OGGR9xV4yXLkFQotZCQQiotJxtV3ez8YM4fldLhZwC0XLGg+f9fDruoCIV4pRnxbvzc
eM/uAtHbEYOcwOdLg+DaSDcgDlFA24i4hrD2DwAb9kzXeC7WvvMTmuKEoQVrY83gsrjIErRaSDAF
dtpRB7iSbOf21GfBZzwoPqzVsr5rngK/kVBtb+qVTHlmng3fnuDcqziZQQljeOBaxhFVkkoCQuME
p/MIJHJNLKq0I+aM6dxfrEUo2fso/3w20gqvQtfXYKmJFFoBBlXv77cts8m7iUbXFCw30o+NmgpS
gRtCCoZ3J4eoRAsGngRuiYR7LJFXgAYkPMnbFGj4icBI6uKQR6Xh0K2j+1Hwx9c0fI3SDtvGzbvz
P6ltgboZDh5ricRYQ1Tl5N3AVDP2/nSmcTnMLha/7UBB9IoUixjMuLXkfHdZKLRNEE4GJYMSIZBE
/qo+BDrs4xnPUT0xl9f9xMt0gYthfYHXZpBaV+1c1NIaQN9wNeRPbDJG/p0fSZEcO1W5FCNNUa9M
Jg0wxin2TmpL/RWG8DCPiMskZurXbND0HOOEXO1bbEJwOmW6yS9lT+GtCMXMzZn1wh4xlOFzhIdb
iHHkP/jEmXCFcb8iI3158iMd2icsswIuEQO6qiaxE6OLtN+cvyvdILOaIUJy5ytlWoVr3K3+3qYx
G5Gk06AGiCmKL+FYo8rQNokuJYldZG5No8cQoysgELXyYXnNUigXJpHaMpUeyx/MAzQGjCXpZl3H
FpjbQwBiFJRLX10WFBAVI5N0kP4cCeiGFfd+6W4sG25+js7Koqe2GQUADTAaJu8cUJTRnpE0iY3q
7sxvnFEjSwVi5Fkh22Jc/cKmPLJMy/vDfi9+KdTDsYdbG+Nc9VdNLRPvYptJpF/0Y9asTCj49Ahb
5ttbsSa9uXEdAkraTw1paaY4WGKbrmqAuE3JnXK1X2yi8gX7q8A2RT0fcNP0xFmKhqKinq3yd0hp
Bw1RloYtXemA5VxyS2oyl3FxmkL6Vn5ZEQSatg0FpLWmpb1d5ec47e6hoqTXYAKv9IH6s2jH7W2E
EbHvaxSxsKDOJ0jE1UpSbK1ME33s3NLD9E4Ut4kYTU7gJwgGvSDkWwfiJ0qjMUBZrWHiqJz0NeDG
rSGFPLah/MeRKgxKP6nVrYz61GZG/QaPpoiKFQGdhv9GwyIacI41OgazlCtSCaAC0T+nQ1PpkHzR
9hy7V9L1NxMKV72JwLEK3iRU674Ag7oooR0h7xWsmLy42lQMRoPTDYKATjrlhx5/J9ueSq799SUu
sRC5YgdRP0BaV2tzaTEouPT4ZSGdhnRpEz4b8HrPOccfzwCjFHJd+OZrWIF5SV4MHHDEIy/g3I7E
7M1aBX56gg5cWSjPGPfiPxJAiXfpb3mLS5ffdWITQLZWZDz++TmThFgmjbJ0/r8xMgWKsj4CA/0m
8udS6x8nX+j5Umnl8ZlrD53ITYR+oukoS8f1bz/1PkZ3y6ZgidX3Rlh553//hjFH7S0TXpVfa0SQ
tkctcxWqTyWLayl8+JpBF8u1X6364X1DIdTgO+dKOENK50VrIt98U5+dJq5KgGHBjFhO7tewDPAz
zlFJVs4p743zUFflfo9tFZ6FpIP0nCWfUaw8UkIHP/rgHKbOlyFRRmNiHLcMSFGhiQfHWD5R1oHR
/I2iKVlkEGTVtr0fS2qo7QCMsEdLZBMPkXsJwjCtCGYmEGcV0kW/rzqEpCEX/tX9Nf84MKxBp/zz
3yYQnwj9dQD5nA4uYq0X8BCArqIsGvD5t/m2FPZyAawBLIHZ4sQs/PywPJtRsdVXixcfV2cMR5UX
sJDsSJuRwSQucmUC35RUaor/xjbEcX/RCTDxNBYSiFm4gtgMEtX8MCu4JeD/M0rPK3yKesyA/l+i
dum9RLuoAWE+APbk2MilmHlGQFF0PZM2czx+u65LCzriqymrPVxMUPLw97BlFYdlpmvuVPYt+2F4
qk8o3JL8Fd5893M37FJtNUPZ2oPwlQBQg7No9F/vcu9EmKezQa5xg3Y5DJQ5rC30a3QQIW9YLBM0
Wuvw2KRbf9zOKHykqJbxCKk/befEnmztBTImnXGsVyIX5xciiY058gNZDvGCUYfrbyVhyXpkmquT
0EKJjOmXWClKK+vySfXE/IqHzTBtu++K1BRdgo8DurLZhLCmkhd3YIlRkb+8vHA8bHl+0Cu4Kuna
pNwnRxFVLUzhnB3YpjgjX2/33QQgrUHwXQ44DQkM5NWojH4N4o/Oh29NpA04oJ/+tl0qOf0hSsGs
W0+BtYhUwuDRUYd6GX6LTFWXIXrnANvhe2odMSLpLAEsumIsQppDZPYX4ynEV+Zq08/f+4mR5Ymi
NTKJeIdkzqoppe+ZjMqa1FrPfJ2Ew4Dohw9IVqZJCzctSypqJQ0/+S+inpdh0qUe5mjyqCSIjDTJ
It7tUrGaK+2xL1J67zoCrsRbL7VZ0wxNM9UduZAikdNPHhIwR4VWIPc/M7p8fGoPnFy8OR2RL0Ld
lc9AeAcS3ZSXPcpT2KBiSDP54xHkFM+YxONIrp7uWjiarzsiPotHViUHSZrTBSGVNSW00akmllHt
JpbxpYuE8CQMe6S8FRBKvf2e3nJGV+91gZwmrllg/u2HacRltdS6WO3+Y8KjZC1swt6w4rUfBBg8
bbrgaYqWJul29O8pZUf/IhWlFDcO023JyShkyhTKqZlwmUAYTFcrW5OMb3maUlAbGnYrRV/DfTQa
O0hhM2vn58KD0oD25XQwD3HjTnajuxjCUXeMkJvTJZaTNSvmRdFvjknYpSjiJhxiTRNbNB75suyd
IAN4G2F/+CeWZWTAUe6cty8UbUBEBcjGc3a0YgtSHtxuqjRCpe2Gi2/DK/pQFHm+IK+f56EcIm7+
mGQZHo/mcf3YJM5IxFh5cBYkX2tBsBLRtLGcLALI/bNHvgGYeMIwcWRJaS7RrzA/IVU5yylaqaXD
k6IA6m+Le2GDojErcCIb0IPoLbCq+NQZaRDXe4x9Yz2k5QDAVCOLuAwVsMi1tBcQS7Z8D9FBl/jP
rjJj4e9XaYPJot7W5EVv0B0YZlTh60HS4Q0j498RLmtHfmYFwNcpu1RS1dqE/IT5JB7Hpi/1I6Wz
zgQmHXf8pidK/F1cm9NdvR3oEzEyJCXxn6xDxgAdxgQlJ66QBGfT3yJVfOZa+V0GswbPnZM1lEpy
+mdclW1bZaLCm3t4KBsR6kuHpiHHok7TNHF3zCvLyBMr6vjwlBQgeKNuWspLshIkFhplDXpBROsz
6MkAeRBkLLSDPCRCj1irOBTjOAHOsFyHX0UoewQdtyOm+DHMWDDSS2EKNgfAnbDw5G9ygmhrc3L8
EWRILFHxfmY8AWwQYSXawQuAgL35H10Mi5bMAsMZdN+7+ZeImrnXIvzRsjtev5pKDvRzvXvYsJBz
4IktojQskAHS5UDKQPqiKAZp5s73uIM46OTqpYjFcOVNlnRaYPKlPtrMeV+Y58bYzOb+BsfvLyXR
oz6XBMrnrmuFz58AV6zIukNl0+1ebgl2d7bYUs5JXRbIQx/qzGiOsCLjB4ydwymaiFQKMaf+pDPu
XLkUCLuMrfKPVcDUAYqud6klqVRATXrzoRWOCqpvp8YdSvqXtuu4oZCpX2c3DNu8p6YeBc/jPoi/
tX72Si3wA8Ui2rPKlNaLRPzWM7iIMZzFLcnxbWsCGxtQXKkYUFnTC1oiyv+Y44Rxm7D51yfMD7pM
Yz7nvHEdsDAgizTK88mZ8VQeM+g0iOVCR7f5ifmx1B4BkL/c/UfrHsBfy69z5nxEa5NbJygURXwP
+Xm+UWYDZaH2qGXR/zM3AX7iMTJhL9w1J2zhdgWDdd0M/HhNkE9ZMxxzKXXwcik19ADreE3sLA5O
x4vyvY6M42toxB+Vwiy9553Cxks5pK2kSbFHf5tuzz4VpR8CvIShAXlx1qDy0zr24euS7ok/yHYK
1DMkvrSNADnDY6PnyVnYthk+8Mu5VLYIargnKFKVQYVveMLGIS+W+8xrMnOcA115dxiS5O6oRMiE
k/1PIRF5swSdzS/aubKmrpqet+EA9CRmWQMM6GsYAj6VhZTY4GnouoY54TpN7TJF02Ch2dgwFtxn
dVvhiJq5NTodTwAUmOpJaIQ2ALQju+EcEgi3NRlDT8/B56EpYjfJu9m97Bi/Hs3cX/sqdz2N1PON
L4I2qOTf96Zbwdq+PUSrgAFe69AqVzCNiR6QWZ8BpTOc/R1QSfkp4v+kgl4c+wminmu3O9Zm/Ahd
SqGNICaWzi4w7eFSLjcVFFdWUPaV+Wxfatn/VpRVMthDE+2oIUWZTvJFJW39vjntFcAC69qmRonO
1xddSMDmlu78lr1XmVLcrDMJvDPnBQXDqd7Xmt6ZlpMP7rNxXJH8eLjHCrzd7apYM/oaCn4DzmRI
oDR8I7nM2JKsR41C2eBy6B7vzAuA6pL5S0UNGm6IAR1finunbK0UQHL4PBceH+bW9YQzRfZM17Kj
h5CgZ68JcP5a575wK26EDrl+/H0IClKqipCT+8zXlFF/37TWtbd7EUkJeJrQB+w9AghuNlT7HzhL
dHNrDe6YD+mSFPeuhstfStU2dyS3zV26UtiRQtYNtHqdcY1JoIYfI95ZwfEHDqwLwr1dqFgGlvF7
+x/vfc2fNBPNRnTENms3uEoTSYxBR9LG1+s2kkE1pcAYmEYuUMJAxRHXlQ5uEtuWfoZk4P1osz4R
VRtVfieES0Ri2VnhB4VWnFenHzdIeHSk572EE6SjDItwkXwYN1RCA2sFKhUiAOMTtuxna1YV2aQ2
x0Lydof4QbhmPDS9Mpa4I9LUUsCwGTmkds+8sAmF/Vujqsc4VrX8AMW38vjryqDuonXThRxhF4O5
Ib0BRS111H38XIUxn5VixdxHVseiWATfSZl3kKD3rIeB11K37r6EkjKx+p6ruzz/OHZHMb2rkroj
cpzDN3zkL4YkSca2Bb/FI654Lk/s+EOrJO2aujCgPjlDokCb6SZACihquzG8zghpNffPbe9cbiWN
/v/WkbLbqtI36OtHmWxuPTivokc3I6T4jD/iYQp14PwOTFJ2vjlq7SCZ9EKwEYU4XQ4zdY/bZ8bu
xU4hJJVvE/D8+aRpuBzCzrY2JhnZodOw3eo0wgx+/Af4GOGg0ltlR4jSu7iTXO9tPzwQMoF0LnB9
7rYvp8fBvf4BJxt0JHMhEEiTAuLvC1IJC9MO3QNZbHNb9sGqYP8dZDdRyNhPub1O/iRj9eTqzH86
IzsaI3tvjxddDgR2+Mtn8P3HRzXDYllmG6I/Xv2H8nxKfz17afc+uG86UAbh1jzpA0eYGP3znARb
6ZTFHzAfOl3GCE7e86s7QyL2/5FleSQq2BFDE4QXi7aBDxIsEH9RZn/ncKT5+2glxE2MOLxOxRHH
U/M9Dc/3R/PII02uUAduj2vzjWutNG+Ix/gkdAXHjVWRFij4NDCYooUUb8Mn3IrnIrPOc0Mrkdtd
aCXzNpCg5tPJsfPj+ZFh4Y5px0bi0TAyFuFF1eDVCsSPQOMtVkmp//wXQa1bUZMubwNhJk7URRik
yc2ZbVoKFy8cTL1P/nRHzdD95pe3gLhtFiVbR22RVOYf1RhElZ/gQyNsgmf+dNYFmvLYuQO6l6hD
fmqVFs9x947tQeQfqt8mC+LPn9NpDcGTa0JLmc9FwCsJ7gxOJc+6cnEiahPsR7LDhnIWELsT8XLL
T880SLG04cQ6Qh8TQomvSWBdKGNMSfKQiaR4zce6ddqMX/9Iymv1k3djeVosTnfAHd9+8r9NLTwk
QWSCUA1s/5/Mu0VAXDot0OrOKSCSHtuFaRAWT0ZYtxlf18AJHpkpsNVlstONyBk0pH4acvxrdkBq
E9/eo6GFuoQzX45JE1xpzZNwvbmFFRWlguCoSxFmU5hHfBFSYR97B0ZnOTXQq9QvuQLz2Bozfo0I
oRe0KB2DvizAAvBVsYKxDydyA9+iECWB8Co1xJC3PD1NtieJfKrHoVneVfHeLIl4E+2R8+xutCKL
GgJdxHZKSu7NKMGURTcUDpzTy1w1t0rOJ0SdNzVvYtblDGMeTRhpk+ky+UI1EfwSxeG61vfOIkTe
3DV3Cq1TBzVCzytlZX0AvbxcergbWb8LG8mJ6wodQBbm7SVRP526TZKZBv54TXxwZcA1onrFC8fE
LEd4ZjjFKKjZLe4700PGy+hkyigyPX/dWcLtWuWpX/83oqCufa/8A/tilTPH5YKsyym5mPNYaDEP
VzIgdma3PFax7L2vnBLkgVjPUXrMPMiw/AzWUcn/IOIrV4MTTKhLrFLB7CDe9j1GFo4Rsz/CiVww
De1NCw4QVOS/f8xv1dEaJpj+9DBNlytwZop2x3whyos3ebOX8R0gJCB8KvH1VAHbXfCOv7qquWIk
cdJm+IfpYpZVStuFLx/4kF48dS3gTTnoopMqPgUvFe647smVRc3Rf6l40+g1KlsIyLcibLSBVveO
GVF/CYo2FRDTD9WIj+h6f1Q+TkGZwZtv3tA0G7ew2gLAzARnIwGVHa+pPH7gz5xdzEkRtEU656T8
EiurFZ7iZ3T454AGt4mo2TKknn4tPUN4WVIqPmN1HCHpZvAmD6n8yNgDymI/Y2pxGevqS5MwkS3p
nHYtlTiwvjG/xk30Z3zhwHZPdJtQKLcrcqUOq4BHXRVYPJ6pjjxHZmih+Zdr7zWxZHeb+aiz9Q+r
bH+SSgu5BH2V61Vf49m3rp/6IvU13lHPjlNZfHmTwzu+u3CESe6j/MURusQVlbJTPkOqEP8qs3k9
lnrvlsnoaTi5LcL5f4Rlo9Ma5N2lQ0Yn37Nq0sdUeVCChYDFTQq5r5x2iARL+GLPtm2cGfXR7xwe
Jqv0gQ5QNfqsJNA5TLB7jj7Zwp+Z4lUlXy1Xa6Y1/B+celJBuXB0f1RIK5hVb+cD5CGBwxnn2ag9
ysWdGLOYoTkgxmSHd4tQA2SO+MAiKVNC2Agf9ZgYoidOcICDvGEcXt0C7O/y2gSeTgG1Pg/OC4cY
+KGV4K5QL2kiVoIP0D2s8YoAjoXUd0kAdICpzn2aec6817mNZ0HDWW71+X01XbjhMsJwH5K5pOso
b7+0tMKnTG+q+QoL9JOZWJ9efnSa46sFGN+ux0J82YRrlITAlvoAgq40KV472LprEYcAb4xEy2CG
TKD2AcPFOsl6Kr5yGyHEG33XJ784mrPX2r/oPlvlogfMIrDHqA/VYCtV0GYaMl708CqyhAQ0AbJ/
Nks7BGxFm2M4FwNQtifb9fN7o4aB//2t29M4wGOG4ApXT/B+OwoitIHHP0D8BiYV63JkLv5p/0Ta
vjp+juKzd0+lCjpYI6w3v91OzqiWrN+nW1szC6IE+93VBXLQgz0W3Pv0b+bv/WmcHeJwblReEcJB
1oWgT6J9O4zzFVm5VypAqK7vyDzBPjy8Vuersw8EvKOdpkVM6nfPvH76zeKVjIfo5Z/5El64SIYV
IzQcEHsjettkMM5AcbOgLZYwS8KvgtTcJKAIZ6Ez2izQBVfW+3PU43DbcV7qBm3gogzp/uAzYiSN
yJumEBIEEFYxO0ol6Rf1LX9ER+pwFLdnT9SDDjopKr3Lk8m+qdezxv3Ok24v6LmnRH73e2y+8+tS
WugORNoycUwIp4Q5T6+qr4w/ZlZ3NUj455JjSWlf1aWp3EyakrahQ+ggnKGPH7MATxCp74T0ixrA
pASDv5U8aXB+rs4YmiBmXIlegYogcHpSszqypZxlld0j++9S0EA86CXXYrnJvOeZK6PEalQHnUZq
H8AzYyR7g5EIr77j29PUfuHq4O7s0ffMvZVOcMe0qSyrs60zVqe1CaluHPg02Wv5NFOjUcHQ5kYG
Fw9uGO3JZ1sRytbqokLf6LlrZXRQPkXQXBkD3doBNXwnR+fHB86hQFR9Ic++/lLnlBbfEXv6bjKu
nQGN9qav+1V1lKYxsCplK97JiJJx+RG6EJTQ1a933as5GsAyAxKM9Letz/DIdL8E549+YheQ6aua
x5LFqj7sgrRBtKblyqZan9Qmx5usiF+gSMsI6s62z3qH02IDQHOlRNlpiV5FUB0ztu40t3dTBi25
W/u6sSEy65oSWUddZliXI4cnYMT6OiMuowZr+6zK4niyAWGg1KA/MI7iv1ZksVZpwZMne+5q3cKp
EPt3CX7FZUDa1TxZBzoDDnCzIMi7owMqhpdeFvxbKorEFJfj2Igeh3muqW70eyIIym3vNVjo/5Qz
K9R+JLN5htcZPjpoXaQIjHwn8Y9JK5RMWrHqdHJXhfJPgJojg5BFHSaIQkTOat3mW859w2mWtZfG
HS0anQH7PgVxex9LeB7OnpyxSEc32nNWPFc3Hu43ylrOb5ofuUnHQ588zaOHYF+cb8LAPgUPjqbL
9vOnKO4TmpST3f8lTbcwWJf36gZupqe1PCNKqIatsX7fdToHbOwv1bi0gNSkuP3WUqPIuod5AC41
YJ6Cc0j5Hijxina5tOXLGF+BeVr8ogpPUzlJnqD/FShWW/pNLPbnsA/OPCDVQHf/WUdvm1UPVDPM
o2X0RDQZxLb/oT9iqYfi3rMPN2YX8qxZxf4mKQwQaRZ9PbRs9WV0rkcTsaQ5kp1GbCwL7Rh7Gk6j
mVILkcmcbew6zkAvcnxNdC1mkLEPtOM4QzcDgOfGemwMSngZGhEr3pn2cYLUHSEstf7X9JGrgh53
FvxzIRzbYGjUGa1zypfa68l96hmPikqM1z4Q4sFH+QN/NgDkAwvBmzgZ1+uamDysHGK+FwYZNo3l
HrQAF7rphDPX57DMWMLhjdEmFCeqrjkbWbH3LSfLq+WZxRnJsb+I7it73ojM2iV0AkmaP4+iwPjz
FL60YtcWRJfRmsdzF2ykYtcvlXjaV8KFIaoCl/dDSlbLGekeKXOefna/7d0NGALzSj2j9oUk2B89
RI4eLd639d0qwcXsDlQ0BB7e0drbPTUinDi0ZUWsbxaXzBU4sqaNpjDKWsjyz30G49xJzzv0opgO
EaSAqgKOW0R9ucNlY0eBJ9CjbT4hWGFRz4P3TlIpH0VnEoQN2C7Dt/fJvH0nkDSbsiKg5g0/r+2B
8sEhoe25N5QCUiH97C35b0ZeuQOiDbSOhStHAqJxubw9wKFRkCIfWaMJR1e5pFyCYht7in08530n
1JFj+LtUfobiFAlLs1cMRYbly15dCnDalApKrub63S2pdZxyxNDLhVwq9s1+E/yDTIXfvRfddmF+
J6LRlRHs7y+jK41N0EmPx++/Rx6KC0szDzpwWavzEKORsnAsGFJVuoTGt2gAtnHvn6TY/lK9JzjA
f2uVxdgPe/Eh/fkBbZ6cHuJ9jPGcpgAUk2zmmgWls1vNS8Ml/9CPhvhNDizf5Uqtvdp0R1HEhc70
lH7Bjql1P+rcf6MoFtZtTNKZJYQoIiNpeHhGiRp5iRKm3TYK8NSil5wcvLwn4BGgDyWyZuCSqUIc
+MoJrmN3mNkiSim8cUT7ZFju6J5wevlAbNUejsbqfBYd0Ed0Q+VjvVN2X2OyJRa1tSRBpeF2qheh
O5fLrffqQqb28oNjqhaYNjBlLWN+FGgPnKTmMsO15ITJbGov+7E9nF73nQXkrI8wmcPU5ieL3ubM
SckqhLG17IC8Z8oX76pIUGGMAd+AS9bRJxz0XyCjK6S96+IXWdNE49YTJEu3N5YROmwipBAT2yJF
OCBnazqNZqtdSJhVQs16x2FspVKhl3ZGM/uddz14EltI/27xUBkPt28haJbrOz1Y3Ccu/JmRbr2c
znOMzkF4LR8beS+l8iQrnyecWj2bg3rFacI9UFRe8MvyZv8TU8z6aQ6KQhi0+v+tZphs9YZNE6aA
X6kKWjqLLsITQkPJj4FlLLK28QAR98UW8+E1mJgbEm9UHEXZ9DdUgb3z8QDak/UkJjhDjipSiK7I
lxLZC9YFHXMUR25TN7W1OAfTyrQkH0JiwycnbufYs6/2UEDQzB8eX6o2b3odVizGr+0aw8i/5osE
cddln44grdmyreciMsFxYfav7039RLzHebKurIqoWk3FwNz5VcxxQMez0r2WZkC8d4T/abSdgL4G
xZErNulvyjiqqs39TVfHyUQMXWuv4mxbygzFz9UraU6Tt5sXQh9SHsHCkKikOCK+PjBoC9Sg91a+
KNLm8Y41CQ8aJRBJ2zm/L9ALeEHEN5Nr4tqVQefm4XYCX8lehVsJGCf/MjbCxZuqczSvD00I7dY1
VpeL7YZFpOSt4JSf3PzHGOJdlokiLnQ6pildshBAiV6rW8XQ+pSPxEARqaLP7Msd6WsGoJH7+9ky
o7olGRZdOQdXmZTJtHj/FQUYUl/uEllAyx8p5Iais0ddjSP2xMMmdX1dRvRYp238VwsoeGabhZlE
8Q7E2ei++36jRmiVdgjLRqONH8y5fjlZ7DmSqG9OnG2gKjiNPx4mNfPE84B+arHno5XYB23FwUJ1
831FeyFGj/MGEASLV8iYn2uJIC0nmOLc5gmhpPU+jWLUKW6IpamdT58lq6dJE6N2HFqGEaNbodJZ
CLOAEzK38YkqzfglAYGoHTq/R/i55sXGCmVaycZqMrIaPd0++kjkloTPmxYjYrR1QE/NqP/S6fUV
y1Boz2YoN0EI80N2EyvPpZCJNx6biEUtEOF4PYiEacWAX4V7Uit+3EaojaH1qDlb6GLikREgk+K/
Du66/wOlOGALdO5pM/NJ7VdqUW3KXcV7zmIlY3F1pPv/1hPelRhYxOwT7ggOedSPq4E7xfYTVVYq
Htgc04vzhaqPzduCXjZW2ErJ9Ial7tJQ7CrtkFDV0z5sBYUVHwhSjTXo7oQfz5/FH+ki4e0yxAI/
7rKxGMEXeqLbEHD+iRSC6qObViV6EPcclXCNkWkZxt4tXfG/aBvPIk7aJSWFIEpGatWykUfY5j+2
B9gC8UOrw7mNPE03szIbFq7XkjMZ+c2iDFRimEJAeOzAwnqliCFyWe9o/sRh9my8kY3OSblLPu6i
n9mxzp5uT9kK+U89yee3lvSVGvQOyJW0d6V9LLlO6LM56Fqe95HYhRQ5vTqoYHECGw/L8cY2uUoL
pMm6DyJLuAZvZK375IeC/kJRmhH+9hI+g+oFVmPKB4tjV65+kPKFGDrFMkza+Vmy1SgQZVDcTZ8s
7Zn5DckIBK0s8/DN447sNjUIs+ewK7k3rGeal0M6xlGByQW9Sz916s0cIOc+ux1ptXIHYZ/V6CqY
YjcvuBqjBUzcmp5EPg+j5ZwFWEAF5UpGR3O7TxTQaHjXf1oPKr7ExsNx3KWYiWjSv5k4x61x6eIR
h9al+Cx9uJqvzbIJCqhMDwB05zUrcDGNqo3uWr1WREb/U9cU8GCkxdzmsV+pZIEsoZP13ZvW9z2v
mcIozKuUVBV7uwRIXddiM9EDWrPkpYbTioDUzJpZZAXAxKN5yAJbPSi3SV+sDI/j0ipf3c1Y8hZ2
hUWKQrf/dMGSwpw28+Rax4oOT74omN3co1sxm+MQoZ5G6EX7BANaUEzN4PT3VyQK8vvWWi6DyP0W
ZTObyQWXGgON1zc+qCViF86QqUa49YmYFSqCMx3Zo6nBXV8rSHHLSIAhe2AGUVwi13vX2l2uOApJ
qdQWE0hOefOp2qqOjG18DVwIrPvK/PWNBqR7hw8fq/s7CgzkKlkG0BXg54luMcgLMoBGhsv4b4OT
xUT50hNpSOmajUnmm8YMF6xlh5wI5BoSiT3TJ08bOuhZ9ULEnAHz/oTXhR61R9bZxgGdcQ/rc9/S
g1CjsemCQC3JJ8vkSgX1UJMhsQ/VUbiJBSoD/62eHZAYNuUvh8jSDoa2YduOIlGWZNORkboOzrmX
2N0WOD64umxUYa0xXuBvER/NUWtxaSYB5gWNZ+JoXfSFdgyjHIfhPTpxocED5/VWJbv8Yf8glhqY
ENbwtcU7MK5EQMN9zqUdvkHqgHYApk6hkkIIouIg5gEVAEoBGDXTK46mX/ROkH/+uZQA1CVgaaUP
0hpfiTFi8wqHgeO12Zwft5c2mtf9JbRwiaNNY3lSnGzIy/7cefG5Hfn4JcGCauzWOGNfxedGO2wc
Iciw9jrVLId0NhqEQzE8lJoO4Bu95BnlC8yXT5hxE31PqZNcHPM3WGvrpgSGkjlNp26WSy4I3drx
HI4tbVc4HmSdGzqjWKHz4+03FwVsgx/ksos+nSs/5ni0zgn/odKI7TCvKz54g52uS0L1LO76OvZH
HWW9jXjPQ7yfHq4vbwIxRg+kiNroIVUYwDjwkkO/zGMzKtJlBoFJEwUW0HrMDg7aQXwIJnedK8qS
/S4E5zpN8AO95gESNZvWwZWuTTV9QmOGIH3ATiyNCfm3i2my42+wr+kdzQ9uOyuQYbgPKgSLpuuw
0xIf4kbBqS00pZRCDymMJNfbX4yiA2LC6h4Uv2q25SGzlzagXNspHfTPVtsTA50sjExAgJ6kUMXL
Apilf3atjO4sJQ5r6EzGfOBvZEgil79m0+CwtfpJhawbsX1+y3+vyyj6KWQNM7kwCE49LUPNR9E6
6u7LoFa4eHE+xQNhVkCC9CPMKd7HJ41E3SiF4l+c6fwDBRgjWFp1q9cyHDVm+mDSgNB7vF0JMau3
pFk9YM5S7jzowTTVv1P09Vlxzn+1vgiVph33knGM/IhP1cqgvSjc3AeytFhO6b0IJp0vEcngnCpz
NPTEyLNPA8kyUhWAfZDSD9/Pp/pOKnvnQXXxaYjmv/ytp9qp8vqlp7f6s+HEqkDu8sRIO2ayVkFs
K2odZAzOw9w+Qx5AFve9e5oWG7rqhNFTNlpqy6JyZcYS1L6JZtweksnFP4QPD9qGXKtTDAz99ts2
HO5vfJrv3L0Lx4vJNBKZ/dOUfmRBlAZNWfhEBplnTKsmVRyAdefJdDpzX2BHIUtJ2IMnuX8XaDov
h6lPLdY0R8ZvKpWbw0n/2bO7ZBcl8wwdmbjjGTN6yrD+7cOhjoasUqvXNYXhV8zUIb342JxPA5pp
BYXY9nbc2/qG0GfPzp/osVcAcliHXd1WTjDUb/EwCGhKuMJYU7fN/R8uPeey9VLUHrELvgqQpPQP
C/4wiJGyrnbiaJtA2nYiyX5P6OPQxdnG4PKLTEYQ0ZakOnhTh/4S2XBeVJFmuuK+TJXQKbt9UyWU
fh/rEKc2SxcBv3MaHH/lJuVyVe9mXsfEE1vgeZhXgGTXY74Ysxx0EETR4HDyjCcBXuIlWWnlqQGv
YPnZwWKhYTJ2NnIZ1dNNxqzRyO+08rqAXwQYB2KjRpAeemzlkYpSdsQYz8Gis9CKtDngmu3Bv62z
8Pb5VB8DyPH0hdTrQ7Veo/iHnRSHCkb4t6j1E7JOWf4VSkY+o43l0ulfxTWf2Bx1gJNxNcJf2bVL
VnOa+RPRefwIwoc8N0MxrHoXqse8HZGbQszQkfHDfKYqt26CipA3655ji6zzm+xTvDZJZBjmolgC
ZE9yVPLjSvq8sRz3LCHcW7AQJaF5b5B9B0Gyw3FWBJIgCUC8zDqnhR3lHvwfjnajk5MEQ3OMx1DU
+LR6Tz5yVlzIFQoIM3WXPI12a0Stw7C9dTN5w3H9L/XtXoZx2pxZ61KXRSfmPGLHeUq5/MqW1Cp9
eibtaCUznc9PZv3HBYWAPyB6mrBTvhYwrK46ZowP7pcES7SEKw/5dWCHd8ookYa1X8r5jvY7QF8c
SCqRXjThFqB/bzER+Dta50F4I3FPWpAdSuRgH6XQueHRfkl99FJC+CrHcA2sn+3SAlYnikAXiRW1
1qLXnyQkWMOFVmAD7CP7LBSVoO/y4w+QtII6F/sSttLsp+tqn8HdRuonjs6oal60uE1y0FzvEq2w
xq3r9Miv6GyccPSJyleQm+OVbvMombGFN16Kr0husN6dbHRU5SBTezZBMsbMAWRNX+Bz20BJqFpL
K30xvG4MNSyKBWm1m5+hmli4P4o0j56/cbTcxEowDNdq/AA5nziIPQOm0AvVnaCPd7o3pXEmvlYy
G0cFnHiUQIK70K2wapozYJt5yLkASeejbo/lBLAgpw+VVX9/350PQbfflYz+RORt7aQaTgNn4Cxh
eDafXsJclke/sv0sYH0vagVCGMuATXBkflTnSz+L45azf3+jFoQfwy8kyh8N51nFICwcxolKH3fQ
HMIs1EHGeVsXGcjSBzUYiCoutLwaRfT82xW9cea9/zIfwnK26doAlTDamgOk+jqKQnW45W1SuIdF
rxfNtZ2cDiTee3jGqz0PmVSnCgn3XMb4BoGCpgnwZubgN9R0PZYOyuHqH/i4bdofTiVGGmVEKTMv
vnc2CfbGBCkNM4rBadmxZ+yTV7LR/1UPsHlprf9hrnCbhCowa+OxyWwi7rLZvxtZkZs6sQv2VWUi
g/s2G/WY96yTS6GSo7xar1QrPQFVHNxpp5Q6ZfEeM3sPZhCgpK7lekUzYW6b4q091/a4MURGGfJk
EfZkkLSP3QUYMc+H05Tm3/Sa0JRFgWh6kCzN7Xw16ZQdF0fxLWnbLfdDgBiuEvyVzYG7D9tc0a+b
EEy5w6Cuzw4RvbdG1/UORyfgvoECz94cfS6qCp0/HaZEUUTpsKRykcpZcBY4kVDO/ElNgryAxZtx
PwDqvq09QpL5rR+Tqc3wKnrQ/fAZlE/OyGqs5jVxHT87YhlVWsdYmffnd48aQW0JdWmTwIdw8EKu
wOU/Qi9GDi6smnQlbAJG3Z4V3yMbkYQk6c1s+YuNWd01lagDh/zuR1RiPe/BD66TagTJKZUwHy9W
R9Xjd2UKA35MOq3tVtQ2qtYo6eWA5Fe17NROXaJ4XfnZskrytotaluTBtBEFGOocfMJEKhoslpcL
fFtDMd46TeXmbWJj37P16YVlvL5WdvkSKfqMpu/3wln8aVkCMlKAFTRPo8KLM+HWcXpadYtvPNzr
KDEyfwGvDUSHqk54qQ2vyYiN9h54Vtvsoj3fay9UW3KKvWWMs9KH04h5tZU+umW4l5oE6dZE6nBW
D58UYpA609ViAnypHvvfMtBfG930+AU2fZQOGxuJNO6g69nOsslnN924WgNzQta2BjYJE5gNgeJI
h079C/xgoX3coEOwt1Wh5ld2h1F0xkpRu8Uhn/9vLMp4hx5aXlTYITJ9+y2/yiHzUpTVAppgvF5Z
Z7I3Bmgc/I+qLRe0O+RvcmYvA905vidY725WZSrGU9s5f/JBvYNHDYJdOENAXDHQS0diOjOf2GfL
rv3K6Z4QSetuxnkRAg0wW4i01dm+90YYWc+TZdGuefL3U7HZruNZQKe6pB8PU06lRs5WYCuJmS54
eyVgf1grB2jsLlwea+8+U+2O1MRF18mtZ5Im6zV8SHVJjy7HR2ZhckDROZeqtHPJumdEx1+rkfq7
HYTaoqlvZJ4oBNhj5CdX1sEvtCyKB/Ragt9g+H+GwgCJaAsxbmkbaCMj/QN/3tgWs7SsKUp1SRB0
3iFsAgcOsjQ09/R8Zq4zGMqeqNc5v63Fr6SDyRRxI5Df0/uhXp4K0P8MZdw9tLhPwcKQBlwzFVJ0
Z3mRR8RtOix06fjIsXx8U0ta38Bm3hynnF84+x9dHugfXtTu/n+ZR0xgZmMPrsqkbLjq3j8eWZPK
+z5/RcZUmGSHKXNwRqZE+yhsbWahZVEAWKH8VoyTiUumO9nVHQfF1UN07n/xSyDybKwMheovFJ+Z
bVqqn1TGJ+4PWgtYMuQgiLKN5fzsof3IV9oshCZXv5sMbEqfetBFzMmqS9Jc5tK4t4243hKrG6kl
i6jCV3jWRFKlnbR0pSTLwaCeG+VB8RTTqcjPi2uSDiFJ2t/ebdrBBgxLS/oQYtaHsSeSJPoV677j
ft7rRgpxuyXSvpXGdlsinWtnhLcmVy3tsBTkqFY9PXu5T12m3RZkI/JvZuoWstFZw0j6QieC+uIL
VKIwFZP1o4Sdc+3HTKNS5DHYercYtQhkzrMqKBxEKhySQJVmABKj58AdWUnMCz1UCSfL4hwDyBL+
ldvXEGsfhlOXhu2W44Blxjt1Ms8tqEhzlj+GWePyLeYFyr6MfISVxFPgyqgPsswo/bKzYLDEwtyD
sFmNCfVkBWTYWHReibaBfety4SgvF84PWjgO4xp8hJf6EL7ro+QwzS0CqNK9OtiJtkzvroIUJpeD
twEVede8FsrSK55lYbFr47P+j01rgz1bA5pJ0TPN/dY5nL+mkwpC7KmzMAnTdJyUmmhiRrnwGveB
0beek5q65E4m6lLrtDb7K6R3i+vBspK6MIJ3tAYEOq1LZHrz59SLzFksUm9r68yRj2LCzzegTRNj
BhFJB4clU3zAYgiUc4uQbUBKJK6N42kZ/u9bKtmlV0OqfgYLFTVQEJ5y3B/cXGBqnF3u2DG8F0Er
GEIX2lOGUl46CbSaRqYw8JAxwXTG0SjBplvPN6Bx1eX6nNfnEQH+yYqn0/1f6pZlnBYqOYTCJPXb
seOeRQTHyDB6fLj69sJo77B1EslmFCRSckd760CfjpxOxw3EK+YVqxk9npMbp9j+spfpMQsuFGCF
Q1q0ahQ0/G4ASf7pxW5G2FlCvuXr+ssG2S/T3DYK5TJQZOqBhCRqzrkDvCT4OPlFjX/BwMJCAE3T
IvwYipozGPVtPOFmWrMAVeolv+UuEfrk8kQcPnctYfi5coi8eisg2WPblyZpwF+93lshXWOikcnr
BsWMEO6hL+adBk31uYPqbu+YW+jnGhcQP7VtCiSK5hgbbGooNqX4TcVudv6eHif5z/n88aotcDvF
l29x9WWRKin0tPJ+gRnl3DezEOs2ZlRF72VifMgOgwEYujsnhF5azWT/sOcwk/HLF9pvK9kpDJXV
Z71inCksAeNfAzlVs8FXdS6dcYckwrZ3jJlPt4ByWPZ0T7869ahbEtikvNJmIlQme+1AThzxMYS3
CoYcQPP4lrHnLlqPObqjPwXJriWDNEzL10o7gBikDIEFoFUPFP2geioPyXI5Q6JuwyLG8CbM2Uqb
/xsEDHPAsbzFbb3UgsyBXpCuk1E1o5W3J+5r2iiSvycooArLjUrUOvC0qe/pF+YalIWtM4wT2txI
C0+Yw82Rc2iNoF2C53SIfjKhSIeGYMK8gtdQiqRug3VYTIAU14aguEq4bMY93m6Bf3kKiJZyVzFF
zXDh1vcWfpq3Oxywr6uHF1hu0kkxfkco06h8eBwgO5Dy4Ikdvp77LuEgYHZiN+fuX4NV02rylo+M
yuRpMCdtznoYlLT5s8PgN/WfQazx8ZMR98jVWX4o5YNN9Dg6cYBPwf4Sz9K92SDFLGirR1ysX7K6
xqSLJEZKYH5q6dUlmRcNjiIjl5mJubMH3m8YYhBq4aGDmTMTVL3W5GYw7dkDZrXQBvduJIYz9uEU
yg/iHa8Gs5bsasLAKPKj8a0xP01e+zcA4+RHx4Ddohfv3VfYdjt++fJF1dErBe1G2hF0/ynQddJa
CEV8usKsjrRv83WvSkcDbMcM3TDe63PdKITaIiaM1ibDpjT7iPVINuuBANi+U2M7OfdCn4gJSmWS
LcuqK/6cgO+khzV/sQlHQMmF4jCiGAd+YibsxVnFiw23+CBEt3RO1h+wQ0+Jy0qFSp7vXJq2TiYm
CRTh5l18q9ctXugwKatrObhBssLfQsJyKNZFZ0uS42HUVPjd4N3WJvQ+QiwabI4GdidLk9C4abjB
tj6Agau6t+sG+Iw3XaAgNB0/+v21/s0hj2cqZMRUPS1yCB9zXfosqa9ll3EipRAdoSOANABaT2ko
QNo0q/Ybc5c7uVLFtQB2vk/E3dQHSaj2eoL83n9jRiscaNMKzliuPUcTLt9kBG5ysxzHXG1NpDLx
uSKx3+lQqlHEY6DrxInoz8low4B5sOH+yPsKNG9NU/IQUNm8boqsnZKKJ7bF22SBosRJkb1WEoDm
lMt+A56ZbYX6ZeINr4TIx0WN11vq4SNuT/yNGBlvCwj3qe9aNlGUrP3/Pf9ELC67e71tp5b5HoUC
F/lKQTkpExvnDnJNQtmWVfFa7XlgBN5nG1g7hhkOwJdN75Swfvb7f7V+lcNth40//nzG5k7EaMOQ
/tPDMryKvcOCg8chsqLYHTbsJbg7+JIJij+VPxRaQcCU1QKnS1CvABR/PvtafPojgrJOxHKAsNZ6
NGM2fH1Kv7I+1UzxlbKnNH885hBlkxT0rE5tuf8vQuMOz1wVpx31oyhZtGzxw49I8E+pM2tHlHQZ
8PokL4OZFCG54aeCPXVWIDJeWqasbgfQZ9SpdUPYA6UCsKN86CwX+BzLj84++k0Go9YPjiBUpnMC
WAmFoqTbVRd8j8HQQtgCFS8fvKHWXtkOTFxkByplCCfGymDtacoXM/ps+HvGYZTnVGWAbi1qmHMz
tC8IlMiPWSU28+jJ57gVmb93+XfoJIqKPCFv43RKr1VdLsFTtqH0NiIqnnYFZBZEvPUI+5uKO/Gt
xJ2loPxR8mE2GM1BGP4lAACg5MQop0Gq8aIfam8TGIcSvPfMfichNpr5Nlk+VLde/vidyxT35jPh
I+tLsC+c8mm7Ez+o3Bs0YEV50q+0ZlLpM/e0PYsSvQNJVsx6qb6zh6dgVaPHkPgiGcR0ApovfWSs
MjoRumgmEc3M0+HyKKXIFOsURuEaKiYWGPhG1S/aWJylK5q+vKue6HmfWxfSDX562qbir1eH8wSA
r7Ytvx4RgDfSL5LPCEBaXQtQbbkH5aJqVxiFCChwVpcoe0QW/w4tsTSbkg5hF4smi1+AofdylIEZ
/WqptkYdL+13N89xm+vt8PCLRpS6NFMDkuXAWSl3HA79AOfjnRUi9xPyEc/pnYdfvtKpHnjv7tt5
a1x4OiG9z+lwydYq5sDR8y3CHeTzA+2NDTQl2Fdk7WonbMyCsmfZfdl2hv+Xmop0YNjGJm2oPCy5
F2ghVbw2MF0Uui9F5JfrLyeuRrT49QVempBDNpHLwBqtXoPtCIbzp4FDLOHI6hv08YWgjsQNuHZD
Kw0VxsHPGfKKwVTWr6xirYrHQ+ZYqn4f/j9S8FU7tf+9h6tx+XOlOrkE4XBckiDaZc3Pcqm2qXHH
WLd2DJQzneenWbrplV1+05fQV8x+iifA5IeGJW2EuUCEmMrHbCmlB2URj1FIH35FVtQnj6sQ27wH
Ch1OR8MNNsCS7plpDUXZrOSHZNTpaDxJjcdy16N8QtRsUmNWZk+I1Lni+tn4nYbtJKScOLPCs1gn
gGaG5aTcn1oQMVF4b0M+lhrQ5t1Iak6oSXxeZ33pW0ZK+RyJBYNUWWl74boaMJKalYDovDTRaSNZ
wm+NmuVKDV1EPJ1759cw87Mkdu5vK+99bnSAYDfXLfmyquVafELB93Bg6pR7rIakzvL8eJXJoYup
8TTRuZArlsQyQVS6QCG/trXvOjXCT/NoZjul4Is8GdDdBtr7R8xZdg6yRFfdq2TMiu9uZvsbjIXX
shFNDVjFurLOmK6VKjOVemrDKOtGbHNEdKgSz0v1gP+jRLqTagrulS88wToL2bluo/+78ZXdgHQX
tUbFfZ74NqxfvsSMxl7xHIdE9UGoQYanwe8gHmjZzjCLnXTRTGH5kMvPLdne0zdTwp6Sg/nTtnFm
LZXnqBpmQ9Y5YLkMu870KcIr/spBSzIDR1vIHmNTEXvNxsHlL1opLL6Ri5uYCYFff7xWjcivzb15
HsKnnGNZ9hDqvZUL2zkkeJA9wx+mNMbc2LAymXT9yIJvpNp9q5grP/hfCg0vqS2rvfjpL2ZbHTMM
O/8BFUfIDAV1K+uAcNbPxMfB9/AK8uk6qJd/MmJJnYNx8+ND3R7fHTggoNO0XUNVTI01c2BvsKkP
GqI9FGN7PDzlSdCgpaEJtZDEOFuNq4DZXdU4JJx2bIcw4tK1n2ACeyYUxcCVZZwK6jzZdj1hjaQw
QJWb8hkXyU/tTLt0QiYjpGdOIfJuWvQ0izmcZ0dYKg4ZjNgFLdfUu9xhRjY6J5HJnMeDfFPadfbG
fEyoSdggLl2TXDy60o9VK3BwijkrwZX1bTyBUclzX0ZV/qRII9s4bA2QerJJ2gTGhI5Q5UpGzbPW
axtSlMJd39CreCUVCCRPOTOYqZ3FULeazXKwmOhIZdm4afBPNDAJqjt2QnOAx/PgFv/DxUhnjDQ6
mgGT7hCHxgsSyE/HIE87Ff2yTkY0rUlJ4Anoqotu719MgImoIxRLWJvliWJkm/TqRhn6uDZw1aS9
c4Rky+IDLBisY3WLRcYWqqs9rLON0uuA1VdR3yJqMlGmKlLwcFXEC6k5y344EJnv/VNxUDGstdtQ
armZDPs3vAA9J8ssBwKnoJU8543qKKE7iHZDkEfCwqe+pQJ/hPau+BohjC972J+08dAFRuQGfPDt
iMBP8EY9L4y1VDqTgcY269nmFig91jKaoMmxFwIXa3wxWVMcMN5IoVjv9tsFIXKVnSFPgbPIA6MX
xlhPSDluNbVj+07EDMn0QaIHuiN8AoTTCHe71IvcsWYnbmyq3ZjgLNsgLtV29htiJOSh4epJSY6S
utjCrJHtjmoz1KASvlIFm385nu5L5pJmDhAIkoXKzts+lI0BANBINAKKD9FWEx3OOYzN9kgwWXKp
IGrGFIDp1SWD3jNyFDvYJcuhSuxT1RKWB41HHz8QwfnKTO/4wbqC9r9f6FlEjqT1SFyA+LXtuwpe
wnrCBze7FdlLIhQZD2KCI0veagBopwiwqt+jjCGLmHLLgWMveKxFoMh4dL3O8VEL8YaABEL8J7Ce
bySQjB3tqGPSvSXctbQhV/ODbJD0xIzr6FlmGUrzeu5c6cO/jlHPKj9NNJLALf20j1Qtxq65wWdw
qC158Qqijjg0uurEsvvqmQisawcjamvBSccJGO17lfTyjwBnLw5u2bW4V9aAg2yM+vcYXT2Hf/NG
qSj41pCNbIdY92xonBxDq6VD0Fkp66pf2knpoyV90JBzRlyVRstsgZZKnttRpikIgYohj54rUBMu
JOMTXbr62WxxZhjdogXzgFuYHbfvXNtoHPeB7RjHTurN88/PYmhbYkb/1xNMLpzzoWmB0dmJZHfl
C7iFxkWBmB5b5flKWENDSsVKU9Ultr+syXdmUA3qvf/LovJxVh/l5wodPI4EqLDDqp5Eso+PnlLz
Lx7NIZhvMZ4frkosTpzalaOzNuVh+4DhXJVGilSrqyAZdxFWcAmHYoGhO3/5+QvPCEPV1/m+Jsta
+gKOqg6DWZyxqZ56sHIir8owEOJOpWuhtxNNqThzu5KlZsHqrSnTo1RukwCnBkRhzPHlsSC/Z6AR
CPrJHfVzJSy2Y/dYGSD0LmNgznaPVNSq3/FTAS1zitr2AJdPY1mvooNYlYYDUZQePlint+8ULuOP
Q4WLIDLrLfYsS/MyPZUu1XTExs2MtU/K3J39ewdbniXu0PLxVA2R4DPIuBo+Wa4Idt0dnY8xlzWK
NSNhOGXOUQLgM9q6Hbn4YkHDjoJRTjTTPsN0PvJPOUVN+cuD3CVtruYN0O/XAv9eL/LfErDBC3jA
YPppxH1E0xVMbX/H9X85j4PJGKx4Yngo9d8Xz2yqUq5ctUEYXO2VmMBGf79CpzpnLS0eaNGiKs4u
Dvqlffq/X9VySGWSoOIAPuyfPtLNxqS947ebQuTQZomJuWzPLEP2zbaRPB2DwQqeh7lexB4akipM
F1KPImEncZo5QuRtcORM+KVVcWrcxn/oiQhjDg/t00NncxGRI05lHKYvRI3YaLUe1+yF85OIaArF
JTns0Rg4yyzEBtdpZ/nRF/V04HQ8B/VzJuPgCjaWVPM40IEtWGKeB9PlJb571gOA5Pruq/Fd9gvp
179/kheyEVBpzdxknIzGWWv4oeLD44iVyWVDUWdSqqm4I9zpyPlH/ckiWbq320P+EG8CMZaRbdRb
iNdqkGVK1t12eLI8F3SuyowvBEm5LysGz9CoRuqpelrGxhnz+858j1r6hArOEUZmEHkrA8Sfj/Qf
NffDzP6xYdUt6PXcXT/TgQCy7a9/Qva+otLu64frQFcL9YvGcVRRU3T3FflBJmgPqGNVdz57DYBT
Zzs8g6igsgF/qwlt4wUN40Ty/IS3YoQbtXQXErXJ8dHOYJdVlRMFuUR/GstMtCeAv+RwcSsE3FQq
OIxsQbbToJY0/51fhDDpSrvK/agePssTO4Kjky4eW0TTX444D1TwmhEi0zPXa0mSeMOcWNSh+oJj
fg7ROJE4mCVlSBK0Ii+eUsmrx2vsIv9oO++j2TSCBJzykIUrFJB9U8P0ReDgQ2Nz/fhlBAuUayZE
kuIv2O105/a4gj5mKP2cwenMfz85wBfCjzqPEbmkPqWyjVETRBiiN4mHQU9FmObq4j8EV0WioHw5
hoEuYtbQ7ogCXMZkwSaKkQaGfO8d22ey42M/wJQcHhsjx+T6kjmcvyBRxnot1S764nbhmYjvVaJm
D05S/ElgRFgYgoJSvF3AyYuapZpC0BOZ3NO7fVJsRcalIdZCEivLG/dRXGehBTqnJSBp0S8kzjsH
OQZ1aWqRQbq7ZZ4h8V56CaQ+JsJtWu3l3SPFFSWfGz0b2uNJKqEFE1Es22P3tAeAVMdEwQNyyigl
jajT9EsoNXkB0rnjG3U9G3NOjYHlZ8g9894Wv6kTwo3toHqq5OMCOeQPXMrYHVhBmLLHfUh+eTEd
6EeNCQTFurr2xRhii2VRGyr9BGtdaaIJQq8kfz/5xBMWF+b5LkjiRsv+MiE1gq2rm+OebPoPS0q7
1FRaM6+sa12iBT1wPTnu5p5DuD3SdfCZjfKuE4ujHlRDF5cd4hQrMg41cMw0h/2Xs3+EmFCKjbdT
rbUHATVBm00EalLdV1lxFe/V1X+0TsOmg/QV1sztGUlNDw1vO5lFPzvmJ2y4Qo3zqYFlKtJyfmtt
O0BjD9ZXAtrlzL01K1JIq2QubtDoZhD9iUl+JmGc3mKd38RqFRsW4RqbQGgx0RYZXylc7M+U9DRb
7BUXdGXdO94aDt83+INWiB+f+MN7L1g/haekwSthiev1wr6ZafHIbC9M2bl13OUURySsq/UVeGKh
aFcByGrvFzgIXERmQpCeRhFCWDtzC6g7bMYP6gIN6uMUZQ1WqrnofrWnEZ3N4I/BRbm9N7zzCkiA
wRs4c4uy8r+41SkCG489Lb9lI38mBRyuk/tR4oTKvxv95Gy61Lu8J7xRKk+/3FchuSjDazVB2oKU
njfOuj2E1jKHkIlEL/ipc/CHSqPEVIOmwSuKSioahkGj3gnZ29VDt5HhVBIOQ+/pHhy/aT7JhbUG
V30F9O+aIJOCQ+qWdZ+2bYTKmHqxqUwIohka2Xl6kkXoDnScdd0QN0cLRSClZtPkPlDyzOGFQXJl
ByprOrX6L9aLZS286XksrFiNewI1Yvmjj1upcS703OwSOIXq7iwD64gRvIZx2fkG0qhlnb2HrKAd
DRQWIbfe3uX/aYQ1bGroAaaQItS2IveOZDfGhH7KRxLhJ9Q3QCgrTQ88oYc/68vNpHXZQU+qxzAX
E88JG58MdfZs6wvwrYX9rAeSrlHeVqw1B9siUf4UysnG+Q3G7mQyJnucODtFmcf0IPk9fC9NR+j9
6exuDekbY9HbYLgFzTsAd5qRpbNJdzLalI1EAHsWBhDUI+plF5snTVKXS79ifaUF70M1cTTlLPg/
D3ZYxNKlJkyuP59snJX00+88KHp3FYavC6XBRXRhESkOa3pWRpihCirCHTirs1wGEe/v2txl0eG0
xN3KOQaegrIvHLnaimv+zZiuAkL8RdjkfKnI3wEADV2wvl3olMcOnJZEUXXXLsGsdSXru87a81Tw
p/wRhXjiWxYjSwSgyxbwta7nzevKxIRnJ9F2z7fKA/4LrLL9J0aFcf/4lsasxJnxEdK58WQYUCW+
axgN9mI+qXAdPxrlIg+lHVZlpbZ2LmdxmNltTAmf7SE/8leWKlv9JDrNC8ifelvXaQ3Cuke7rPzt
Ejy0M36aI6Yuwmq3s5MpQqikpeNPuTUF5B4QSCeQTIpsuwfV8ThbWuqio32g/U89KeYWNrm9qAZS
5B75uWtdNhDfIT+5LYD+Dm2ct8l8tXgtclGx/X9qDv4nAnm220XItS6pPnopSw7kBAo9Degtp4x/
z8gDeNuDqDPM30BwTLuNb1aVOY5sF+FQwewUW7ARL2bhvfgXx7zTNEVLwRgSof1tuypv/pWChWGS
FzgqnoZqKMSBBs+F5MhMyJEpo84rDG/+ENTafk3pNf51zoA2Lg2aXs3RpsypYoCPdnTYiWb3Sguo
z+CRktEfSfLskOoseG2GkPTt3shX/ihOeRCk536KzruYXcsWd9vBrBZw8WwZX9JfPPBqAUzx3oIN
m0R+QmiWO3q3iDeHF1WnU7R2OunDd5+xHBCfpcYAnkmDQowOZxsKUUw88EHU5kXhXD+QNW0nPUoF
VjBPPHQkqJ8UpF5BdTkQb4qYUFMqEFP7+ixw8IC0xCYQ0KppjBckQWotMAnljiNH1jRvsu0FICp2
90lZXyzYx3E6OrxopkVs+ovCg+FPey+C3RuE1NRDHyVceVVReKlmlXwfk9hBxOqJfrAYtP/MS7tj
7jWi35en7GZ2t9cFMZusHeUu1ouXhLwXawvdsZrxfYKbaNA1eOg9MCMR09x96IH72HMCffSwUWpc
1kDXndvbkulNwNFx9fgYDIyvi0+ee2Ggl+3wbC29zWVfyeOHVtAsHs0HJLr4HmCPoxyZk/lTxRt3
ouddGQxWhKoeiJrSxT0wrThZtfksVttZMhVuPYyk92PW8POXhjwIa6KkeFxRx2KFTjEt2FJxmPRz
0M87LYH2I1LKJ1e+O0zB8vaGZK0IiOGbsEyFALcp3o3K9L5GZ1cUvb+GLkprROACW8B00iiHOvvU
bP4J9mA0zFDdJnswW3THH5t4jpxGBFL8FZsxNcpIZElbPvNMyCVG8Q6QdOy2rs/qOAlHnxmrLGeJ
smyVoYDZIPN2HGfsDrkM7y/mmhoQxp3ZjUbIrAP2SLgCbFx1XmjoctBQHrFfO8q5lCoah+Fhz1Zo
lxrhEiTBKb8GuOloxLqd/jf25PSCSamiXSVv8VHEk3KdSxA4dBP1nO6RkwlE5gpo0rhk7m/1roKf
6SXyx1sm5yezmcjz264q+9P9bEuV62UTnhJOmQPgT5CcstdseV45Gny3oa6LOIwSYZBA3iWXVfOm
XwixNJs82dK1nd8kn+EVhx9NJNQFsnwy8sEAmXfVDL99IPw3LoV4bZryFUK2+/N0UEwF0UsiHIpb
XTS3MLL6rVJOLsoOHyFW5980E9bH28yI8tzeoFb1QSyaZvhsm7WujbbYM+wDNW+A5XjmGRVQ2Sob
WdICNPDMJ2D9LmSypMdvDELWRJnJFNFa6S8feTlL8tX8K+ux6CYSvL69R9SyO4ZMa5fBFstClmGi
cpsFyAuqG2f+bccPIqm/01N5QbJ00yxhFExyJ+cdPu1yhI/6ONmNdIvoYIeH1GbSwRIdYoI87BB9
5yeuxx5U8Qb73z6/NEKiUfLNO0a7V0f+cw1ybZ6uZQr0CxWdP6bcVXBXbFH0ZONVuY2KFPaoC57I
En0AsJNr0udFdhlfJ61lMHcc+M6NHgGyG6QxuDoljyqKEI6cnTvv2OsK7YVtKQBLIMziJddpCa/R
bvRuUNG4c+UJflD9MSLC9suN+sCg1kdmuoRFOejAjvgNv2UuK4smD9M2FrhYsPXCukJTo41Hgdcx
Ol1eWDykGEx+CqW8H86Eu6swePUCIJYLPd0fS0aAwPKTX4VseShpQwLSByCUcotu6NAlREIVsISl
SoyrH5ZJa3WoJrfbyISkGtDqOWnH4jFKbNDJ/2bLBguBmaHv8SA8gjx5W8OPC8cRrRn6R7jDAmc5
3+rITb9cRK3HJDP2lBgkwIMjJNDK8LeHa+erpP78uyFvrkrakTspUeqip+YH39qw3xg3FdOZqlUZ
K6yrtG8D/7ghkfjwOr0G85cFcyfhZc3r51wx/PRykmQW8bwbkZQGUdjy2uAMMs5YgWaqFhtHhPX9
NkMcvl7Ud4vfVhcEpYkOITgBGF8MrNNZ5zEAAzrey+OywNjOsgL5bk88G8igR34vFAO5C1ThLoL4
zNC9ff0E8OfU5OEiu8W+ntxzm7BvnpQpmXUcHST5vJGzVMWRsRPz4SwKdsde0zhbyAg+9rrBA9eH
CY52TrtZDDuyMpbT0Wlh92J+kqgH3xkZNWHwME9du7s5PS4Q6F6Gt+i6/5rcTPxBclS7VG7hr9pp
uomjNDMbH0rMs24aF8CLAsx8vmcPZO2Vi6gtw8XpzVGkjmTV2hq+t6q3ycQ04ENW0bWpyUzMpREK
FE0cwfu3myjx6DlwB9xOX38VvCM9t2/IIkQLLSGTNz3tMmz/m8TXVJrPsKs24hqxXOLuCtNblr1j
fHYrr4pOUxyrgrwZfXZBIf05Ov1nr/3AJjuAHJJtv1fg8gGGGRY6wDmncucqLddYRiZNuzpABpeM
4oJSRyJgoXy8XYWvLK8LAMnvy2ISWMw5jrGMubp68rqSLGcjUQ7GlL12tHJDVb721ZL3H/pzdgBG
EhUGIMnTA8MxtwhQ2zcXdocPzYnIb0PyamOx9d8ytDGYcB6rFbRPvcPKU0EG9KqPrAnzcR5ztH26
xSOCyjIiqzsIWrcejays/FwW3cCEPNiFuC8UyIYsUkaeydvrCyJ9hPD5VB8ohHLyj+/lsLO+3l8Z
yEwvTQ0N9GXQDjs8DrfAswF+MwekkfjDXRWH5lrCaSdl1O+H6MnfJnF+riq3SVn+ej/clgzQAr5H
ATDx49ovcGzQV7jZ/h6fY20+lbAKvR3LnNdu0xiL7aGGQvx+CyL7FlhpragP2OY1wejw2JU25H7/
R+Rh3PvYrilUKnYjdNP17kPyEyyE4kZXJ5+Ep/HWOYtP9yDGjEeH3CK2RuS0azMjAk54hEmBARET
jHtqJI6K9ebIIEOybIHRP3Mx3iuYRgMGjKdBnIgvC5CcdBYdU07r990fvdvdHmXiJtBuFSIcvZKG
72uCpeP0BQ9GMOyMOQswBu9cgMBukBQ8r/4nps4iSQOja/q/+Auo/06cFwMI3p/GF0MnIPv7JYq3
HRmiyILkJlGoeslVr+sFYotTtbEMWnhnjVV/GizTLWx7NcBfscjtCKSquvv/MDDTsnDD7OvOfMbR
ts6Z+i/Oiceo9UrlRBHqkpGD6Qgqr5SA4VF8HWy2z5tQJD0BkTSNWdRR/x9ljNeJwuS1kw542g6X
Xfz40HWLdhTOiLxoBK3jRt+k8Tpd4DkRWJeWS2QyvqOvSOFHnuA+LfBCoK4iohbEL46XIJtE0t0S
gLeX+3e3IkfB8Jg3DIodxDKb876dLa2WFdfpmmijyuvbnkJ+Mdaf8s0+gSrNMfr3aEpNV7ovrVzf
J5SJrFU8rsUeIknDGT18i1hHDm9behSKda1IhwDmYPtUVqRBEOhWsHj2oInmmGkbeUrmoMmx36mq
CYf8p2RHqMXaTVo+QUai7F8JbRlbza0Ruk3lOKKnUw7BcBRO9m4C4vPosKGS5iNwXPSnyDGMxnr4
aSROFwQwY3rZoUx3w64M2Bxl4auWuCfaBCl+mlMga/AMTOJQGD60jFVlJtVCSjSyD+LZ/ZbMuqGX
HjMJSFOFDC0kC3/1oQYBnazvSKX93iFHPiXNcuy7ae+guky9U6Yys20aeqEV35OFAgv9GzOxBRYe
jJpysdHG/0T9QCuJzLGlROjuLf0QPFugIgKT+9c3oU5siLA3WBshxhE3bpl2duvByqojIbWyPLtq
f3KYnnNnECN5SxSkefUG2347ETE2qpJTIH0UmUUnE+mxy3C3qyD6LLxcPgo+ueVRdyKmdX/y8K7X
XhYEkXunDPEvVl0N8C9017FxQGAylgWL6R19AE0ckyk/gUH2369d7bYV1NOIS0tDU9Ox5mcPOcPa
S//Va9KS+21sj62TCoE6GwSCvrzQbo1TJLLTPlS7vv8aie9XVf0gnEivf5I4iyQbzAMFVn3dCbDg
Er/PbwNdI7ylSEexSUY9ldB4wso4BuzmPJm+oV/wBthpfIRl/RlJBCy6KEW5l5FMPb2txjjUd3Q8
R6ovQiyHzuoOQP1I06VFXCbzuWCGUUZN732+mTGiSxw2frr3oDV/QtfORpTMw0A9e8GzTqlK+zGE
2regxm7ibuUqRoabV2/rs3IR2YhJ/egGKspEslUehjJ66Fky2uMAi24x69UAeBrh1s1C0OYgBYI+
lWeUSO7XbkgyKv6M4H/XViM2gMnajnHfMjrSyhqWDyPwwOBLAWLs7hn+aJETMSkWLCovgE3YGPjD
yaxtDJ2+0KLNJNF6mYYzlz1ay2OacgQxzXaC5XGcCK3jSqK6NQJ5FnZLWiWEg6S2oVI9nZ157xtR
J2mERHpao2SSloINwVCD9Ja6scDWpXldE4+VuVCHaCHb3eSvjAMjU9B0VbRktC3RtPCINB5Z/6aj
3e/IbJ47SCTfeMlmM5tUey6XLQ8YC+WPQ6GdP+6pb60BhYUTUua/WTQNA06d7AElqq85AV8WjIgQ
NgwVjqFTYHCdbc1wwf4UshE9iWyCE21hYjnm8WV5SDt17hARsgXhp7uGXzfzCF3JlMimexpizqIQ
wnbf5cYDobHQlHzWDpUmKxWCWD07SLUS/aHBX0EmjOU2a53ap6pNYyK/e6gMwKJgV+IrbwLSUjzN
m9nsg/7iB+2XoNnjW+8EVPozGtyEjYQTcAR+bmJ7fKFsQsnZI2Q+IPk4zDDPJE2/8WvoOpcvKkH2
KnkKgVdLkDpNmZjTJn3VT5M42MJzpT/ES/Pg626nxcj9+dsrveYCRruOK4aqg6gQFd5AFsyHVHaI
unBYYa1iWNe8TeLlpBDF0OX6FoHLzUnvKs+DUmZXa20p6Tca7pShFvDttOyJo0QcA8qRxBSeABZm
nuWmA4dfr31x/JEGh7Ilxiw+cStluUFKp40Xk/YyRCtvUNMn922lN8iz7Iwyq1unAaN9qSlDBe2j
DBeRU59dZo5AAN03KDuOvqE0sg3ezlFhhGZAIAg9Iqu9RFo4gJChMsGSfmNxzSG21+E+6GTBFKF0
d3OFIIVKO05w1n8Sfh+IpVznFxR87LjdAO7mHnHGKEf2KiOp/q5Wijr/D5JNKhHwJh/FfK4NIFc8
WA8wGp6yqEiEQWaTUdKqmd/uajjjvPDwz6cfg/WtzH6Ob1m+fA7SNNvSzLSrDpNSiex5OWaKvofY
6BO1LqxqPIAtasArrwafspkHvaGC/UxwhFsqZEprO3C9UgeRAsy8v70yH+yo8mL4kvn2ylarEsfh
jK/jfwGm9m2Hg2w3t4Nxnz/DIT99TUn4COSb8M60Zc3ewfFodUsXJrNK4Jalz18ltLLcYvwx2Mlq
WNXuwamH+DeUhdndQAmX+4yzB/lMX+mrlvS9B1yKiQtJjUHo68o17oWRZR+MpJ+uOqwVTb8dXsiD
f2abtVNUN20B9+m7dZYI4jtQyuUnwkfH1TKFRUMUOiH3ymMs2TE86Giq7L501RxssNopIO4y3kDv
6CIh4HH/v8dYm6aRjXbSB6+jEv0SMf6sDat+rYxMMRSPi+FWFH4uHpXLivGFudlHeHfrg7bVx2hq
wx9rKgkesfH/Q5vYkRMb8eQf7v5I6KZgJAkX/uczq/7ngz/q84TbvgXVRBgZJaPuiWpeaLsj1toX
5diYpsAhaCdmwn5e/n6L9lnrufdGeaD5FRzi1hhXD6kB4tOhqMND7mJq9pvkRONOtRJ+gVoapW3V
g4rwvH2p62van8UcBEogleUokI6L2o6aHONSg9cW8cwI9oNxeM6cPgvd9+crnvQYw2iECx7OowVI
nrvZOzJFKFRD9XSgx9H5CI6+TMA5hB7uN3f6Mda5AtAHAVgPNhfYKUoKSDstTR2ah55per4y9h2/
pNfaCYFYWn9bxXeHQeGNGBk+Gv4M/wW23qRS9+jnwerbqA+DHTyNtihNVlZtrGXfZ6uqApbqnw9m
pCdNQOavgwmkQ/TORrEd2KmopXjz4BzyXbf9kPTU6lkbN6F0NGgsHAZBDN2IrG0/rmxVofbF69Kf
PpytPjVa279kxaMgFjfNi67k5iRWLePOoPn3qSWKVSSQ9gvBDqSIeqyKl6xzVOLM/S9h7S4bZa/8
Fm1nChPA3ZPCw3TbRw9p6aqO6wYMIidbc+qshExFVoO4K7tNQTULh9D9HtkbtdPZRXOSqN7J8mfS
dmObfzioUOpjrFB9vRKtgzmUdYx23MZr0xf7gEcfxBgNG6XAJdZYxzX3oeL3Mz9SXYVhD1gYWztp
z35/R+pCCiyl0iG/LAiTTnGmt9VRGTA1OHXWy01Ysys1f3Uz1/sBEoc8ZrqIeyuh9Gb5Kgoo6ltf
P7oPj5EWHT56+ymkU5Zfz/TNXbgGwXNRMyB6C3+Gw03Ma6PN+0cwV04JbCtD8fJ/y7YaO7ExSIpu
RsBMHNsv7CKSTV92OPZV6uMPgmFrF3+Y1GqhAzRsUTsiYabblNlhcCBqUmPOI6FYeK9oqnWKFyuU
P7C1t7EjfvK7gpAkGKkSOtalJoC6SJgPipqPuYHZaflXJGTWEMK/Dfd1nOUY/18eShBUILVfof6u
f+dzqVyuQTSnQs9ODscuf+xc37ojftAU1sKPSBDjb4VytdD60cOPYZYAtSAyO296XSNSDuRQ783G
VKkYmHozEmqrnjUv82aYZ29/lHRtISQsWwS63XBKgZbcp9kXBIDE6/gQAxi8Otp80xTHTvOUoAtL
8UKxEJU5L1O5QCJGj3dpC/59R5Yus/YyXAjt4sx3c2b+bzU8byRV4LelGrfqxFMPPdmTlCMhPKMn
VjCbw+ykIQ9hT11cAzNjN370wR+KKZE54HK8TUBK5N+ZKWPxnQkG1/4vben2JsBqur0rTbomPCef
K2JrveSB8lK5A7XsVzIlDaXGM2u/4qeANxRRFPub3mAdod/lmSNb7ZtAAIelKaRGfi8l/P/uHMzu
2DjKjpB2kkvcZ8YCZtRTcxPuzpeMDXVht10aNXFelNw+jcip5gJhiMjsMPgxNvAvLZB0KA9jkgJg
HOdrdHPjQ6cgHJiGvzdnEEF5Un8hVpuuKYNgWttjT7Ptp/JTG0UeyTI9RRGqMqafNbdt66a81+Kc
lBZmAw44f/23Rx7XKfpZmyR5MiWKqy8EzwXSOo0m9Km9jwxocL49/EtoMl8fYDBEKYbZM//mfFR0
4XoE9bfoG9CQc1T7c8Gesz70PmZ4toWTpoIsl5ObliqYTEwz8191e0CDTepSAgX1Vdb4Xee1NaIB
dUtTF399GMueXqrq9sbdcQirZTT/fT+RUEuJFxfHsydfSHGMwYUSD7LBIkFQ6SUN+CN5KuKkilwF
SwzpSaZLXo5MJRLJp8Ic37JCcRwRP4BXybNZkwB/sXv3zrYcasZC+ks2o63sROedQcnFb4dzOzmi
0nS0EYySgux7nUqoA28Pk3LdHyC/D6HyyAIxTcUl/E1avPRxwmoEi1ABZEstKy31C6M3U6TIV9sZ
7uuUbsQ+VGmDlrSniKpINgkGGmTg3whBChEVMpKZg2H+bTUmjiXmOu4A5lDPTTdkNLWxEF/R/7GB
gTHKhPtIprfuic6qTnZ2WEbqwD3gKEN5O1JX+PKlRbE1uhAStMYcglyxhb210KveZ+ql8/79/KZ4
5JmWe+uSvmCAfSjigSY+OHce0KgtPPslemQNTsZFmt5s43Y0DRsiDTBf8EhiD+NBSLumui7Fzuj0
jgr80ovvDZfJJKty55Axne2UeTe6rDPCAZm5t2P4AI+jyguSZzRkLOR12b7NCdFUY2mJD2ZCmNI9
Wy/NtTxYw25SE4c08FvaSj3CZvLs/CsLhdtfgToEY+N439HTcKdtPyCzGLhsVsAMpasnJKVoutLF
3V3K1h5kPR7rGqNxBM9dkEdRHnC5Y9fD5OtK18xHJ4+bxj3weAOwiMTXWWPB0XiZvmXP+yXPpZeI
Da6u0RQa65BxLM1Adtr6/z26ezglMt8NWANByxJ4OCi0S8fjo5LCZefquNy+q+ujW9tzwZ1sejop
oMjX7K3nqFrFaxn6pBfC1icFCuB24y4HQFdKSed2dEzjKeFxwaoc9WMMqZQq6lP+mKEahieirFeI
/N4ubZRfMBCqf8HxXEIy0QCj+Z/O44CiaoqQwemV8y4wHEaxz1qL0fQBGugYKmmDL1eIH9O01OT0
OkewXVAgruJJ7f6mL1IqrgR/HPJIhMCYdyhxMfNPfEwls8X/KP41xQpB9LHhAc2c+lqyXzrTCCdz
hnsdEelS0wzbzmBC+K+sOvtkQamE8e+Ch0kdqLpa6hZc9S68kv4dUMxJTy5pBjVWpRlKZNknFUAW
yzutkTH/8pOnwdIn2awUOIlLvpcCWAme1i+WvYPvOIzKna4oHYe+SgdmeK8R8mnOzlEBTWpB7bO8
1OkxVA/4A4DY1gFEk0CFejWl5sb0iRBI5wCBx+A5P/RgbCjFDRB1RW3lpMjfC4SY1fiKAPj81jX4
W5XndPaQIZx3zUCzP/3mj60FRCIRBpwIFzZaWksp2GI16U1JQC+MY58hVzTekhj16ZEeiMexexeL
QOSyylGiYDXzw17BHIonmjHKbsEMPi6DBX8kdZUfHqIX52Kk0dTV6hLnZMpgL272G22uwsAJr5nA
V73YiAbA8INuFl8I+hF2exRuZO6BuKmAPC8kkUhBe9pA8U7W8eouQvmZ49NVKXOZVDQTuVRoVOCe
/D+6bWWxce4MfpzrDp57pcEHvoiZs9ALfz3FPgWb8yqi/qf5yr32FMpSDXTAR5jdEcfApB6S6OKt
/PxpQfA4XSjoxF2/yg+1N/OfLWEK3FgPLdRAqYec+aktO34EpsZ7aE9vLiEn8CCdN3HKZpHrp33+
93tI//p7oOlilDWFilIxyypbBMUY8K7wYIqxwk+7Bg1vC9wkodUsWCLv1CeDPkpqFADjhqygfa7B
6U8gh1j3jK3u3iX/sAN1pRu+E6CxpFwRH49tOgoCQrjBTp3BzEV72dLRguWcyI7iXdo4OYZ8P9zj
ALLvs6k1RiMW6emv7lCIV/bn/yt7ugozuvraxTUe3ysfyyZ1VeJg/dvCtPZo3ptXmILkB3qhLuxV
M/eSnKGavHDI20RyAqPTNYrorIzJzEV69uTrDsnvJqnnxYZO062IG0zniA+4Zm7XIF7Z2w48dQPO
u0KkBfQTNcZLhS0glbjrrpWqmAnyZ0BOLVpn6ForxL4xtAc/lB+DQHFBEqVicP2uDdsFaBBXrg3F
XlUEIexRAPS35k2UUL7725Qa9Gblt1GSIdZwNrPzJGfP6PnieBGdZ6+QgsstIQj58ZkgOeqi0cWU
A/6KqnzTOtoktdk0RBiyybuS7mda2nPN3a9ziFgQNck4OzX84dHaD8DtBG1KFjYVyUfXkfXvVOae
v8IJ93c/88pYMRobd3s7lFiJ1KdQqF2Zsp4Iof7f0ZQqCxy2OiIJY1EBOLOE9a8HC6gct+sIwYbY
1LIBwS/nLAJhuKlgH8ukUmHOO0ZEyHRVdmqsxObHLFOyFlsUBc6oIcS6sfppNUAVqLN27olC+dD1
Xdtd2cqPW1enxSZcRTA1xzxsqOj6RWcfQh2ljmrwLp2iI2uU2EsAeptRuNH3b5PImdD+yzJG+cFF
h44VpQrxR0cnmPT6VlvuqiyKZT9JEPIgAqgo7t58TaUvjn02icGQuWT9cEKXvX/W5ZpnoqSvw9P+
AW6q9w8qBHsed+CIzlROIxuYrgvHvSjf5CYL5hI0nWmBR+GadOqhR5V2YYm1/9MCLyW6azKoQ/ex
coFU3SgPEfS0bhZ7mrB6cND9rOalFx2zzxJhHEiTRGO5aTVR0lXe5NE1ZPxHrg9gs9ClmcWIj7R5
HXf5c2VLqUJQPkqesuFRP2QbArkMlneHLzPsUs6XbliKFQ+WJcQJPhTWjecuRRsTTy+Cw11PsLh7
WIANLwj69qucrRULbTyFqJtuc/ftkLugMeRtGyHKHLXqJmKQ810zIy1WPfznbPfRnwUkyxo3RyoX
qofVPveBhSCiTJebUaLoAu4jhvb22pgs8YkQFp0byQPZ0/Xlgy/tUTY8gIRkOWzbtUHTMWK68W+I
/nIMaVDzSOF8PBLA+fTp1YEJzdSZdYotFdp/b3pB3rLgeK2cOjtWJhF6lphu+lDErcB4fm/MN513
kXAD5vnxyQbmcPSg55mER15nAmepChxA6pTOt58kI0K+lawLspzjZ6O4EfNlcFD4mMCAT8EBHeJd
jCIzAH3KiqPCjzZLyoyXjYOHCdJOPhBDpCqQagAaScoxd/sRKUbfqHnHDFqZX+DwgvWxb2BcCP4m
kf/3GmiEhdzJdeWhdA3f5J74Ltv5oFuu0KfUvKRbnpcH+qN7/qjlsF5KhR0cFSfzIHR95UhzgXxJ
zKr5zRwJXPeY69kEdMBs+G6JvhHCgljr6a0sdjA8Hw5sx/ZfkpsuPCy3bBHRvDoKBgwjC5x0NPHP
8OsRT/ZbT97LFBLu0oFPIMG+bwbmjvS9lWat3CZubZb4gHdEHlp5tpOZpnjIHB6lBiqqI4ivKgND
EYeBwlxlEj9IHU3f7mc4wC3jTqeTJ7fSsV4c9Elcyhj6ZTRT0Cu30LZJWAFX7fuubKP2iFVy2Ah+
Nq9mBxqO61hUxR3PimdHWqvP4HfSv9xLAcke2+leBDR6Pfr0tsZoZOAzFdwr6fahXd0l3ykw4suy
+JWuC2S3S6ZEnCqRAoFlV17gABC79ynt0Qpy3Rgo97Hb36vitcZmVBJrUqFlLg7/rQYZuzflbF6u
9S/whTAoKwH+xlgrDb0wnZ8tLkIPMpiCMtlPkUHipElLkALr7xUnjtYQtnaLGfascZVUIuwnHGqh
RRI9F9X7ikOmpY/CqGywnOXz9/h11vbtazLbXQW9NZ9antgazrMpEwgyqTFv5kNAgQ8ieFvZBFY0
slIiJgylsLkbSgXSJS1d9t4KJiptOdnfqdTNQCWuCc0eDkkEEqjUf58pggb4G+D7x5uLDfZDsfaZ
e/BoBCC8M3QvEWm7N73SnvKEq90p8reA17hA1amiqeVHYh3QpuC/iIVCv7m5Llg41pXgRcd2sdqY
U4SL4k1QbCOuyDn9jjgq+PJ3uGSBWjL7MHyaqDjEKgSNaoRKLVNNTNrYOoXWaOCgp6uZEaQiYXnz
h3JI7OJjvD8MCDdgXQKGn12MwKQqSYM8s+/yWVXpNowLBcGUb6Z3+gdJiJO/KReZen9w+BP1rxwo
QqKTNbZxICJA80W5tqU69Z+VrXyUvr1gbdPuIFnl5Uq4xwunwrTGtvNh0tWCJ8ua7DmFd6PCr86H
ngucbRfp9jKh4iJYd1brPFpWtiFfYy0P3CVETndqAAsuU77baObB7zLHbVXXLKeXx6GbuFvbZi5e
j4EZsvsjVn12Fp3WAps+HcSPExxhg7HhyfBJyusQLhH1Dn7xyaMYBL6KFx0N1v4MN++QW+N6hlmu
WatGXPruvzF+K2nF27YSUOYZmxV0dx2Qmi/o/IvB7NgOyazvO6D8wRCtOuCVbdHKen/1ATAe79Fb
Pxe5MZjI6eMI7i5mt96dEMtB7UzFmO4aRs7i0INsLtXjvQkvjbw4kBlxitRv9ldcqoPA5mvg6T2n
SgrBbYnGWWBv79FRuH6yhOfpDEV6weuQboQNPgZNOvQhE6+19f/m9rD4VPt5Bf/hAnAWFZWl/6tX
EnKqGo/cr8YNJxKXROCd1V4nkWj+oQaEH1gdJJwnKQYonylsUGRHtDCVG3aCpKQv9HSagFk3+6je
IPgeUWt97Y8byh0rpx+PDRUbZ5DrPohlLP+lNmtu9dvSX+jJEDua/ImSgmh86RobktF1fcRjo46l
igS1cxTJ9booL+0v/4/WG3HGzTeNniKwRGXoycUuQYwIA2QybP0j7W9gcq3g1tuY/evnyYBGj0vB
AopWRi1e1bLeB7YfOXzL3Og+Fo8Nr1fl3Qs/Hk1qNof7yZevo7KxWJ4CPUXkM6ubMBJWHyeo6mah
esQwAsJnFogmjVeGcbgrNXV3YM7RJroB31YHlNgIDoKyN7ymmzq85tFV4Wam1FW2XDSJ5wM1Uuw5
UO8biYoEE5Rz1vOHqFMtloqiwGAEjdwnrMKXABmH2O8vg+E4nK/GTlQ8iJTjeIaCs/XqcLVdriTo
RXEUPWCAFqvUEd4uTJnvpYaiNyxpFKrZgKkGIfyyacWyNmEle/e8vXeLcrYP1Qofo66sQjbsSlcm
bQzpxpHUq1PbjIIAYuD3RjPEmWYs9MleyQogUXAdrwtwLUyY6cZZHpnxWPbbKj96/upXAX9vU9NI
zPp8dF6eu5NqRbbA8X6wswZ+7lBe2JqG5zOy0rysGPawfR8UO3CnVtVPArI3JiqduRw0f0VUMrwz
MBfIAur/YIkYW+Qs6OvfIKI9L3iYIuYfFtou0PD/7amvsSphPvsYB/IIjl8dCa6yJBC6OlX18yeM
41Ubrxnm975yAI9WEIHjSWSXWpjnv98zlwW5KUFfbc6bgI3yUt/2fT/knxnDL6MopYLjdIPGTkZY
liyh7h8SxzrkNlfYiiMq7PETADf6ssybq0wcaJaez5H7maMey9F08iTmbiGfD1jXhc0pVXGHNqcT
Rj3Di2Yx+frCcH6+wWGaROnD7cZgefEduUfp392r/15Mdb3c35mGhLV0AbsDWDEwfxgXRB2RNMr+
0+M0yFgv/hRvyYx7fswb4lceD5bW+8yZdWQeCSpAMhBnPK/robEC8t/HW9yDsbbqvGQRyKDJchJw
aBuYKsCu8qnXKGUbZdDjgd+56UUqHpXzTb+S867ak7NRVP/co0Pw8nXWCOYwmItLgEA6Wy6gnWy4
FODcb77leMOubBTdEUkjaH2wnx5Trx3gIHyJdVABiqXtKpgAgxBuvX6jSXpZPlpwFwSyCXP195AR
WR1B/tiiATKqPdWEXBAtcsd/YkgoJXtJkY7cFGYRLqoYQZDaoggRopuHpsJtZVMhMD2MVZ/cuyto
lClPB6O5y1d6nC33dZAqjdR4n+Zm4XwJMckTsWfblZFzNYtA78UFd1U36pp28e3zYF0KwSXsAPje
bgGJ6spwO3NBcxtIHO88u4WAkTLsjiUswsG42/sWMdF0FQIcPW2s9CiNlX1xax+XnIZEMRe9JCCL
HYU6JXv1fTWq6AkDjy/EmKjJ7mqa+PrxDRgJV++BiQRz9bCujjBlczqxDqmxPaQ95XEVS+XvT0jq
k1OC/DoEIIKXENv1u5Z43UqkmFhhHTsEmEcF6aavh1gTxBZnEXcMc6fI/UYuauU10RATEgo4hhP9
ZcgBXomVYns/asqpuLBdCkW7iyou+SBeY3EYfQLUizu3uE4YB1KSO6FdrWvHhoAzBDXMUzyqropA
DGUAkEC8OKyZnqflWgF7hpZKgXiQ15OvyNag8Uxz20Ob/Xxxno+TLly08ecXznMuxxaQdFvAiKXp
/tsG72z6mGvqhKf+nK1pSoWTwk7F2/cWcwkw2JTdCX9UEDIJbiiFUfZJ0eEBLjcj2OxtCUzkZ/+C
Zls8kKEtKFj5kvDMEy6bpokGULLTyaulnmJRdRRR/D4n1kY+0fN075t6Tt8LqOs26+RZ82oWVCTL
mlOeaCEjBEt8ULy42AfYmWVCwDJMqsMGNCUKrTsduRtXYYBWwXyeW8ZQy+XeQG3QflnC9IXIWyZc
floH1Tei4nrmDnLpTb1plSTzlwDEP4T8SfF25sqHddyBOCgQC5mF/ZbHotqB6NQAsiLi0dFtCsHG
u+uBfEAN3bM8pO8Hn893jarDq5yLcmfW5Y+XBDoxdanrcIRGBXSkYRf3H3R5i+TgR6mndUBAh58K
fw6ZCA117F2C3Kihgzqv/ZGpPvSXwGBnk4knaqcw6yfhUiqNcLS7J3SomI0e8jBDHKo6Imm7r4pU
xnWZ44/TgU9HDJFqZt+tAH/w97aMzvrDqxqsXBO4zxscG6orY5tsx4v+9ndLqYvchwRjOvB8xfK9
x4EdA8WQ5qMmCcXwttU265hjqI/Xm1UKFYy7rtykZRviZZrpujOe3oTCxioSPv3Oqst/7brZu5j0
CoS3tCfuM2ItlVOUQ6XRS+Jv2UObdeLi7fx7uNfJ4tOnYV0YcPdnlGtadnTSaM2mPdx69RjIRRp8
AvxJ+fyIYC8LrFyVQnRbjtX720JEZhi6s6I420a4u8rvgc+i1jTcGt7zieAr6vD4tlUqf20zQ6bV
6x3KPeDc0yzuTIKgIf9S3pJht5+TtvvjuZKcO1DyLOFGYBosRQ2/DQp0q5fNala/bOlJ46/qP8di
VqgqFFy3dbc/IUDY+7VoqqY/6LlWGF9KT5Ur0ufizrELck4Ne0EJvNSiRc1ZG12S8GfkHU/2UTGs
c3DoN6Y9/WCJSqsGXxJtEn+VIEMkbnuYkIyl8WOlzgmnZN8ZmdiXP/BAmNXliTXQZoMZWQdG6R0Q
n99FXfleI7P0soBVAC9VFRWzCAX/yHYygWf7jCYbX1PRoyR0DEHkp1kRCegHYBWXIpO5eH4B89QJ
vjrt5rRfnwB+LZY0XGLk1rQTv/ptI4OIORdoH1D9Aud28Hhu+WS7l28DqzlMuRw++qdVnxLoMKVt
TCwV+Af+nNB8ov31e7O2RcYYjFtr2ET5qeqFFru+vy8KCnLB2tBZGl8kvTwjYTYgeevgEB9YL9NT
hsMblhkxAPRJEskD7VyRbsMdmmKN9RDS0xDESFLGNe347540VJEVLmgtJSuj9F9O42Jr1Z6CI4Gj
uokziD1xK2NaPX/G29cSc5mn53h+AnyRyG2HogbKvia4ASZogsmnLF/kQQ0+jMfDehl7f3ZTCrIh
hmefzM2vQ8Oxg9nuFQaKKL9lLZ3xUl6QndSUDCWkfmRVOVCUIj4l1sCPH6woorCfLmWOF0SuMKhl
liIsNlBUczivzhp0JSMKU1uFUfV/LeaFmYD+1+NxGz0yd8VwaOiB1ELOjHEkPhzc4VLNzANGTCQs
HS8BKLzYsOiyzYYbxTFJ1zMI3CK4KA/KfeLZ5jKNBv/6fmymnBgt/dcNIGBPyo50W8cnNuzY6WSD
pojauApHvBDxsUPvMq9nVkhbdz2ZOg87aLIRpsyJ9Ze72BUF3Rl0Bc+x5yKRiHB2iY6V3Cts8WBj
qHG9/9ev0YiDMBeFGvkaUmLfydtSDrZK2oWWSW6NAcwKHWKnROlnhaGVe2BR0vcPMUS2ny/oJb+Y
Fqsu2WSJhwq+H7XTaiW6E9jk8m0WMB3nYkvJrYtGbcZOisKWMxSFnlt/8SepxWPwJi9VqMlBKqnV
YpM25N2+9k+EGFQKHrT8W8FiKQAWrbNf24mIeFwS2gL46wEh9i7J7VMKJd03Dl39akevAytbLcKc
KTaVHdLkxh7D903efkPOh0kbsJgh+SEzX8y6JefemUoQoGye/a4KO5P6zpHlFDrOOHaoWhwZrNv5
rGZGTbQF8QsgF9OlfGqmFWWYll6KzWd5SceFEeO+tMqAmS0eNWYl20X4WWViTjjBSRfNS0oOrZ/K
UEXiq8OgLe+wBdxYcZ1Mu+iHldevzeL/A91zRqo1t8wSusOctPMeUAm9N8b8aIi4UzPfm6vM+Ytv
asSFeqTRbkVi3IBMNKzgi/w26FsIf8OU0lnbeTwfNcbtRuGBp2HnrdXpXC34gP2qFWomD3c40IeA
hOICxPSfrAQ6voyqk5H4YuyqWZpdrkMKNB0A2XBwqSeNNYmZRNRXiTONQqU5ThzJkI6Dt+qySXud
dRS58vAKR7y+eHvyUx8wQX6ERhf7Ym5UkLLSnIgnL3/MXcUFTGrtNZ6ZAameqZc1hHOl1BkBtJU/
K3pVYjaRw0Pwfy+Be8Xc0RHyT/jIHO7Ay0DeCtx8xCITrQjwG0ja9RdpQUIubjGIKC1KJ07IKdbd
iwBna5Z0aJ6HiicAQIin9gViOd6O9/8w1U7I0cXGkgpYzBH3YYe+NTOv7+QXJLLvK7v4UCh73CV1
NRi7TKHfj8h6D09/6Unm1Kncc1UWqWSZrZ2pA2v4/lfnEgt48WmTrOs4EHgL3vDA6XkpHns98PGo
22n9YCDR0Qc3MABablwVse2AV3utN8h0t1tenIi84uWz2rLT7irQMVhjf6WmvRPAyFoHuyhgwcl5
CYoJw9QCavb+gkacsTBYCwI8OFx+S6xJlra2HzhleZFnNpxGOD3wvCNGIArcgCYXETi7WEAjk7T4
qBO8WjPHfayNMWs7AduDmPikKAeRzQSBp7ZtEcl2d5FwQR6m2D3Q8gqhFAODMell9S/wNn2dO86o
YYvV+RBj2EC+3ybNhg60dFL9dIQG9z5xH0LIMjvBFqI3jz99ig3m7sVGD42z2zH5lwa3FmWMUZ8t
rHPg0HpQ/s8kDzOuGkzCzKla+Cv7wHWdQCOOFP86D5b9PzDvZuDL/W8BOLP46MNwKDlEJJAW5WM1
0QUI4+ikZqcexRIrLFL7l2+2Nx1/SEkqC/ss0VNC6Mqo5VcpobNsvzVkDmKEqtdUQoOfYV9xFm6D
RlLfgtfzQBfXdwuC/SVKmvt4sazNTW5qF1siKQn7MkEfD9tUeHace16kHiI20Dok/8luJZPp1oVj
EOqfovmv3MgPwZczJZaGQithDRXeXPHPqBWL+30pOBf4XpM8uh6Xuozj122ZQ0mfOl89arXdoETz
ujcz1Scd9EvZ+H1f5QeHhctYRyczQt3pYAUlbykXUO8GQP2WBES/QqByXEEtZ21kND+7YIf0xORj
EShyo2CkuYHctmSDyZT92JT/BhBap2cHmnJ0AXQs4BnfN1m8yj/XTi9xoBOvl23F4E0LCGXf4Lnx
hZhu96TuVyldU0r2AufxxEjQ+3Ky74X1PteXJk5nCAECb/Jaij/bEj7JpOfsGwsmaHpQA/zmvYJY
rdRckBEfsnaXZaX8BShIzv+2ToF98Aw/TwgEHIG+NjAdashLMJHxNSdUm8xkYwepmSZ8c0Q1b+YL
PGeePT+7LJ1m2tk+lcxgT0Tt1CfsPsYo2HlogqyI9jwLtZhwqBTgCR9pn1eioauIOzRku2cRPPoT
v7XshZgUUZnUe1sbJtF3gAMOBVc6LrAKltzU00dsnS/0b7UABoYywWXOZpIeqd3wt0OOWYyvQ1tr
l7LmHjz51+Vzdvl8Zes+BDqPYc22jaT0Pc9D6O/UTmY2dn/6cEYJBy1B02b+i/ak7trZ1itV2Gaa
4z6s+4xb3o1qjUBPCz9z79j32vm53QXRWj2RVtQTuSo/yYlp+c0WFo2Ptl091boAt793kTQsPSZi
wTBAD38Am4QjvHFtnBEtqmQCi/kI3kjs83l8jtj7nX5oezcMikM8odxGm2gotmvdnKvM/PJN2Fp5
dFi9HvAYo22rkIiMmM4e5OdyA2JIaARPGMvuPbPjXjCtnqVTA63DDWQkZM7YOl8XVvqEFkgj2O45
VgXIbbzNstpIHcgKlk/Yr/tIlg5e8imo/fh/I2IRUN91X9wHtFRiRtUVsnvLuubdBqt4dj16El2N
sC5nsp08mvnZZJM7eXko9J7/GgabmaknfL7zSEcFGXO7hWsUDVINsBS5jJNm79Y6/Xw8S/nzOpWH
1IQ/YMQDwgFWwIbRzS2v0NbODfWbUYh5UTIdOhjAgvmrBoYmnys8oal3/yKxCnwJyh8cMiXYbywJ
NGSzjcEgtrcOtaJOnJ+oJ9/AcH/QY55xSCUAsFFe/6j4thRp9zo5dW9N8kYai61LWDmSIx60aA6x
WjuLwzEleUbGEvlVyOQoXH/P6pIYurO0xqPcW4M/K8k7XVjP466aP6Lq7wA2iWay6VZNWkFd45KY
dlLo8R4IBjN3OLEyb6+yp78s7L3e9JXkdCDiytFA1LZZfWM0PjVemajAViRdltnHduYYGU/daZVE
itjE3yzSK6akuWF98MJOCjgbsWUnSWJndDft7gUP97PBVp8bcFS3QTrZBIZGmsOToBQxpkMsRodh
K5QcbyrDm+LZYYRi01UeUQDzJiOaZrXcQ5f460HIq/76kfEErA8vcmvuJO/FQSeg7m6OpVnsZU/5
j8ghSfGV+87Wxl7I2QgOPxuF19C45k9NZhdDq2/e2hrVqSi50xnF3i/7IVF5YLqsNLEzmIbPb7Ut
m0XnVDzIHtZmPSMtZZEcokkYSpdBzlQInEZnY6XOLLgveKFDRWfrg94w0pysOGxsCzukZ6qBwAOT
h7oXjuutY331AzSr1ygyV/GFMdrY9qWbYmCsS3gcUw/W39w+H+wgPnAQlgCMYvllATTx+zKpiep9
6nImv2aKi8w6/t7ZjQz/uzisNYmsCnfXn11UdtaHfQnjSws+cXNHcIZfYSccNvGOF0td7B5Hwe6a
RaG0ejwzRUBXNZtQUyrr9nQcgZPfERWE3iQDlN2GFJNs6SItl8KpvIAVHxqBp5G1RL3x+Saxmfq2
wEdPM756TdVPKGAfWqgjBN4lLFfSFS4Vq6YhAwFQtV+cyvySUS9zKegbWRXbp54FP51AUwkU2wzW
ZwAf4/lPYQzkuZpLV4PL5GJR0MpvkWzUXDak1UYvEqvMv+AWiu5vySg3hkM1Q2QQ5hWsdd/7jYLm
0GE9kyeWf89OHup0f79Of0J5SbpPrMQIsMxEIW74inZiqPpgwkwD4xgRtms1h1RdDKktQNgGR4gH
eM/Gcv6x4KdAQW5YiQ/oc4Nej3ntCQPWv0++SWM5wi6b7jau6QSt/Osl0yQZrvxInxAMi2TR/lPf
stzWeB3bA2CHQ9Sg266yIcGUBXuY+4xcr2CLTxA1ez/xLTUkzfxcH2Y+3jzgIeSkZYFlzuF+Gnn4
QoFg0vm8Fj/8y7rDVEaCeMe9cXJe/hzEuZgsCRn8/dZuwn2ttcjIwQ5s8gWq9B/RadFbC9s8TKYu
53WNEZl8wM2n7MQn2RQ3ei+0Vjn9u2D6dB2o5alLmAQfE00RpABrMOFgyNmCX8i1gHILjFQR+Oz9
ZVT0S+F89k709LtNGB7YfMxTXCytxDiH4rUD2LsTF5W3EXBhkhSjb5I86c4sOv5Kwk9Uz1HokIQ6
ETXTgLCOJvVjAYX5ULxMzfSu3iKr3yihlrODb7Ql8Xi/J7w/oiODGG6ak/mV5Cb+sy4jd3Z1yWce
yA2k+SdcZiJqMxmBn53JGjkh1dT9a96aFIllRhU/FE8W4xWMIs7Ut7zGrhgRAdmB7PseKx8iwDV6
UaF135qu+qiX/6SXjQRctn4n9FAfVh1LWdxYmXjv9OO19jUZZdEaTPUOZi6xSmdAXtT5yNGLEz9u
s5cMougIzZk0Nmuj66zmIbjyzK66+EFU+ob0ZdlEKw5pl6mjWQp6OGvKiA7+X6+6rhCEfvIRHwSH
H5LiDmrj4KX6DqSHN3haUX+GgxgraOxi1mQuyRGnuNaBmtZyQ3mxmdz5s9xXBsXhmlBH/QgGYemt
vbPQap5BwRaR5WM7O273tAkci9OiE7AETzN0cKyIwY2g0vFYMRkUMuHtkDAJE/+Qw0PkcelLabXt
xvA3rWnnJKa/esM2cBleIbqbIq6acL9XbXgV+XKFYUQLx1++AyVdtnAjs4Lx5CeBWKeSb63BuJ/k
kutvIDHWOgi/GdKaDLHFAu4isJbDey99kOyqFacyow/CWDxOnS8xrWTQD2W8NfHTY1pwpRwF9scK
m4X0w59ElQx6aa20IjswB7vITlkH7CnXGFjCiKBkqvotjNB4+LhAzExCK4VNRpQyArbebJEZhucF
g/kpJaSEBDb5a93r/l7tXBmtbMqHLtuuOERVrHNSdHD1dam1PX5+xPn9IL9RT901IGdMHSfL8Xf1
uFaBBoj7XClmzrp/XlMwu1/tRuVXkx5Jv4ZrE7lIK7/ga30a2+zW4npgsRcgYtON7JbJfUZOQjsC
JJ3V81Mp7GGWHXP9DBKEm2qay6EXorm0wX8bIG8knQer2vcWwXGXeve19G1MXdLOjqJhT1ywv24t
AXX3up2hXnTpICpTnvgQvua8yaOhSRMDahczAQaw1hDCudPmQoOktgtIwLU6exCPzS5zs2/hjZHW
kZfUY5VQGU7NmE35Q+mXTo5R9EllDDNtuwLyl28BmFKPIIx0PnwurBItcbKkbfZpk+vJXJgwI3Kh
togpMOMzJy/S0O8FFHjS4rEpa+ef0Hew9dSOGDxETPuU/tS1PMS9t3hfV+vOTVr+Ecc+bQJGdVlK
rMuFL6JF2e9wP/H+dqz67TdR4Ajrm+GBYvNQ8EeKTbL4as0AsL6Y7KKwQ2y+aOenys+YKnzXx74K
yJ4ExDsqy8cVfTySeIYJRE0okbvawcz0NVpZvYG0qvjQ6uY9b74XRQTlwdlHxB0x5nNPLpsVplov
81HdEgl+F0RSHZqZ5BYU1u60b4rOvMH5jAAzkfaMDbdPHoGRSziKnPsy2kDayn7EWNNa/gDmkTI2
MWyxdHkH3bHjHK/HeOdGNYKyFMTnAWY/fssrtDXwSQUtmgoxkly/PTVHqo9nnHE8FL7WjmsdvNmm
4w1QAwm5uh/ySdj6slfOC9NCWekCCuBcpefltxtg2/VshntsEBGmX4qugg+OR29WocxCMeiD/QYy
lhuHry7RrRrTglQlby8OmSNpM/WoTeD4C1r3kk1kFNbT3aZjOhprHEbwGZk6V7IGbjeN9P3qGaSd
yeEDP8FQWefLKU9LAv4DDyPFKCMkupMxhbxRmuUT0lm/tardm67UtKrmP11f3cRHX2x5WM1+6i5N
LDmcNFutrg2f7T6i3fOBuseUfBYIV27Rq4qEQAyjIf0tvkJnl5z1eIaaimUv578e03t1yR83eH8v
+zO6whYfXvuSlgBfx3AIUH22K4O2ZWlCbJL1LDOR7FVHha3o8qYNYq2SpU+QEX47SymDBDHpB00h
NSRK3mMCvWsQhJXxJghV7kAn+kxk29P6XnJcSQwF+UIS4lSqaQiu0PYqIHGw2DJGcwBMw2acu+iJ
0xiJE+SzBHAzndSjIJH7EGNYBw81PUYxB4DBdPFGFvBQQfS+7A1kMTDL+9OdAZajfadAKV37P6Sr
5AIYWllRAKNHVaEQByr6cdIUj6SmgBG6aYj6gm/Z+CPntb/UAbEBfkM7c3t+Y8Q2D2mBURmXsU7Z
cuefugPTWg1zXZiO2QE4Y7n6YQ0fs9yPwxH8BxUVzrPquSP4zd3uHdiPdFrebUnFF1CqAUI43UUU
Uat5xDwLwsgwKCma3AFWWFJzS1xWXoRiqubhnGN2Qcnqj6lvAKLgpnXCflgdBm0/6JpjWx7rWG5+
YRrNHBGhq4Ttsiczihp6nxym5zrR34RlRA4uVV7E67CSPl0buk8euMCKZ37mwAHqjkQLGyHQE75o
Jn9q1AlPKWyf5V+E91wi42amULKGtHY7C8nLyaeHEitxK/kwOtCaxS/V8CQJ/oYMQIZk+E/j/R1G
bkOBknn3GWTLywmZ7A1pCsPLdf2GQekW7sfoxvD5+h3n+l6s6z1ImGUlswo6ZeYfYtS0d8CyQ2Xy
ndy1owrSA3B0g0ViJlUSBFVGVp9nBxI2usBxTFP8rdc8t0LBo2aJd/4qTYQSYQeLRgzyGcRymdaG
AHOwRBtfyNVbTmqLWzGWfpr0936ewZ5gddz9Josw3D3bErjDXThGPABV9FJ8M5TP2yj7M9H95n3y
bvi9z1/OpYU1PaAgwOgxAoCJTNNfBzbkCFntILVJZ14r4kKLoK7NqVU2EPfQdhIbeNezL0iKKMWK
amL1Sf1RqTHF79wnarbutTYc0yzyKPzvEQyQ8+boxWBy4d/GBQwYorspbGpC5eGclNJYLwoKlzgk
i0sdmtgWgjot1sF82kf88tIt0P0QT/QtmX8k4RQGYGC24u0k+ny1WG7xPhG5GHE+kkMuGfHiPhNg
AUox+SdL4UuQB43Cehbu/c16BvX++i5z/fOuUleaw1j7c7FoCNxY7CN3nunOQNQX7HPOIXlcgzHq
J3/fuitXtlKpuEV6MscKtkwjugRX6xLjYn6AhT2moDHXZ9/TN3ZZQSDg6+/F/OzV71s9YSmcl1ZI
PdmjZAh4JGlWyQxXb7QMrNTfzxZbK/y8ebKL3ZM4gJl1lYPFdc9rmi5R50zMBHKdoLa5Q1KQRSIV
njf24lgAA2MfLr42I1bd0pAHdg9hofCkdkCd/mR6yOAk9ESMsGUgxg7oKwtgpBZz3UivZvkR2ZFJ
50gJqSI8tjmdVXAZyzqUwd2Ldru6SpXTuRJb/HtLVZfik3IaDOWJhLoDEbbFF3vVtCwG06AroIRc
bY0t8l+o6TyeyheAAYFtxO9ItLKO6vNKwBwxNxTeA+fwALPVv/g2TnMEkKuBFKsdhrSBmAQa2ROF
Q4B04dLYA0QS4KbS+9tf8L8TWx/NACxvpHD7jU/1s6XTt3pyr0/oiCYi+ZB3PHJaUITulEdgqWhY
YmDROKtvUKTZGnu9xcwIf1WWerPAknpwjF/zTen05o8scUHQPMOE4iRMuhSpKBxC6aPxrOtQITRx
MhhmSIJJmjexL5ozeiQqADXTGWYhRjyocXyt4ZvZ+8/FjjV2jYWuVU3kdxs7WuJdrtGWWmwkyR/y
o0TEngManoZcfwcAgB7H3Hpn3224DCEM8/+xhpWr4r6UNoqTopw0RtzvMUun/g9DfI9t+u9F+gya
yc7R85fIRLPyJFdoByXTracJiT88yh5YroUDRTkDv1QI6HFzvf9nnRsJE18nNI7BoUv6G6rXcD8F
mZ9w86sZwgdjtahbQa/1oAiiJbAo6G7+B3Gy3C5JPkme6vDPY9bZmBGT7n1mhDSdHBOsp23QVucc
flSf5/p6ePWcO+unO5G3bj+seogCuQMzVeQLcVoDFu+GQ70cH2EpFR6lcrFZb7mWn2sVq+yqhSaj
EG2HmX/jGNOXhreIyri20j8CUr7NvOQ/iVLePt9xsBK5ly3sNHicrvtZCmOTVu49lN+9iL/aQsW9
UAihzl2uYzUeHj92YEu92W7hfLZDJuERDrf5u2Vv64aHpeMvEE86DBLo6UC1CxwNSGJCcJzd/Snr
RWsPsuR0H8KghkTmtCwFBZKcRN91/w23SqIvtjfknPXDJiZGneciaJQjI+i0mPkx+G7I/XEheykc
KO3CPAWaizvCR1Xs5Js6kmeH31Ny3UgKN0oA09d++xPCeo4Bm2ML6YBsSO0gmjFEGpE96ZZTTrxI
OQMxhcZkrPY65GX2D66wWY0PpjtmV4QivMuTjCp+yqPnfQ8Bo9+wPepBxVZqc8gyW7iDwPwd7ASG
YTPn7Z4pOaGhPgsNdsNHAZQYZjD7Kd9Fn2Z2wZekIOSfnRt6BKOX1mKgbDSTrRYJHGWi4BfkdrCb
jR3LZoq0nWL3sOnvvrPxccN4VhUs/m4lgRsPtmKfrjoPkunTPCAlrjT7PucjKz2VajoBPE2aZxK8
nhpO3RPZSd69Gg2DeJZnCesdaVX+BNDFHV9Jcqz7Qq3eCIk8mhisP2NHilU/g8T8Kvg67XyA3WtS
gzbeDRr6uMdhH3UquhF9M+dCHdmN+ITqrUI1jpb7fMo1c4oy7a0piwdLkTnJENe7xxk4n42mnrYt
1pdxwnHZwzF2p16Nbj4VlFppv1NzE/zf5E4uJ4tWwGIxPBobokAF4KnDCVpfqOXm4I6wJizdxKZc
LZ1irTdWTe9qoQpfgLuYv1N4FHbNeZshEirQE2XCwomjqSFf1gtUHq9fMeSb/i3SFxO05UBHu942
IB65sTkd8rNSLQ85cZAtIKbXHcU+WCnLmqKhfnUIbk3YQ9qDA8i2xE8i7gZfytm36vwfN+7tgBwO
OHd6vqyv7rpbG3lRRFw4WeLsGzUM1MO8TjQFHujZQIy6Q/638EslEbl1HlHNPR4E81iVaY/vRj0a
WnZcu5Linxph0QXRfVR/JZYHv1sSjqB2IR1lxlX9SLp8MnTZ+MedwF2pDZeD7NLYbVrLLd7gjCpR
nQ5amY40bL8ccVhwr7xcRRgaZ1NZRRrb+mucqvupVbOLXzx6MIVkefMeeLVJM5g2Ghk3CbQzREua
p7sZTzGWdHfgubOQz5+lIR8ZJZ0U/84OApVwnRvAt8tsOMtI5PKITKrx71Y8k8g3sy+L1wyfX/UJ
MuGyFewK6273rnMfLse4bRqKXKa9KeP/Jk0fQHXC+Uf4YC9/XQEI4kWG3pfJaZNF5o7NBysKkbsL
2npKWcs8XLikWpcUQAjnQU2XxBZbT16PuB16wXnmxEpvXR8NizJZgDzrtjVVd5cihuJ/Bc01jmNP
fA7ZJgv85Q/4oYxbOGmeWPSl1QbUsT/21q9tJ9LFPOHF38xbPW/2sDLcP5GHs2P1ham+08LRgr86
Ss4NnwrVAEaHDKy4YP7iGZERuMuFADjNnvug3SkVtdIBs0InwEnuCumEmnzb3b/c2QYuJzjjQHoC
/BnaQjFXJ74nXFCTN1AyvNThH04RY0egFhuKftdIY0vUwCLhLudPg0sa3BAH6iLcg+R0tEi9M3X9
+k/nmoLhAyCd/WJEG8zdck3v20kYHVMPA//AOFfLV0QEK3ya8tMQdCqXU+rOWeYM/AkmXNgvs2VT
owoJDJ4UaHddgiB29Hp7Wy52OmbwnKHSn15Cus5Zlz3oMsHaX7jA6HNkYlJyJMBezchR6XSmpELS
jluDNgBx0IUqNIuPEdo9zfamXSb1pcSmzoeyiuY6/T0BLAX9+GFKEbYuioAKj+pNU1up1dGhaiie
hRrHMDZx9snWPkj6uFc54+f/bflPEtxSFcQYEQn/pzv8mIXtzKJ1uT0x85ZTv1CojxDiI+vyEidB
0Bcvq3XfmTh4lZcLWPrpEcQnJCF5DlTRbE3PKWT1tjpz3kpDpR57SYP9UeP+3FfVKKOv16Oi84dc
1Euela2qdaEn9ijo2vXCAy5OitqFYOcOW9n3sNo6xj/E84xuc7SqkwHJxXUtmhAOXBQRzOfTVo4j
qWnq/FeJU/e02CXbwbnA/A2vXEVsF+6KLmALXwXEXdRtgg9JYq8F+tB6RAOn0dkEBXs8w0Tn+8B1
09IyrRkQ7kl0+9UO6JZsRCBvBW9WAwAVpxUPDFnq6YnHHpxcZ/3lyxgSIkzfJrS79GmD5QYndD1X
TF56RC5sq3NRHPkikoJ8Wx4WKHLy4ozNq+KMlfdB9yr2j1kt8m/t420KxwK+hxJof9ZozDqBoF1K
OI5b3mSkmJ3sD9uZVxdf/4RMKKc+lZdszVxdSASv3H1zwwkqZdGR7qEdna5Up7F4o2lbELR9n0TT
hiJcPVac2bLSzL9MWnNQ0ImPcNxkU2BkGiER/kdjfsTOUvxMvNlpJw/KGA4EsBe6JkN1x3rm5syd
tQ1DSKfULL69EimXLgzTp1twXTE4RvQx1ouyxJ6egh7ScRUjqmyQ74aBPnJowC3LBBcM1wfPdEPx
TvVVz5hTeHB015TdT4K4D8Q/d8vF4mMDNk8cG70c9T7uUugCcowiBUqE1N9VPPmL37f0MDBlfWXA
L5GKzf4p44p6qI1v+DjhdcKy80wJBlINkOYNJRGELDpmViJlip/+hu3cZLwbprkuRPTuUP/IUEMI
5MM+uyocDfhp5rBRVBD1f1q0igj6trwastDPmcEkYceIpyLU5Lo8WTjmE6qeduAAzHxwCDQ5lAoo
HzOKS5+Ftw78QxC6A2/clqtAJMSm6ZoI/we6BlVNnpz5OCwEnCgGH/xsJj+N7L/ElsWWlIgV9gRE
hqXWQX+z7NT0WngH+ClyVzyrw6kKsA5IWuaehoN3gujyQH2ESyx82d+qj+8uatMmwQ+D4XswRqe1
1yXgFKT6w+XNv14lBhDACECElfh9wxTzKGkirciiMpgVqAuEYK3w9v5tHLSvCVdVdTVGpXJMkw+f
ynXC8RQygSlay7QgtMUqet2NalVnYbC28woOA49Bq6qfnvfkCS0nLVYy4RtBdOCsCT/9yiaWNByN
+Wc62cnuXVHyIk2JdcrYOHTCD37/5I0k5baAAB0wTcFPQeEW32NHAAoRbmwIEs7tUmDd4YIZJ+l4
eq66bk+yh7Mvj4jU9T2RRpSeraI4Kq0m7+CSs6Cw2dySciEqRXWiHytaHqeTIhbcw7uIljMdyZa/
hRTVAMPu491n9N44DGlOeHt8RRTdJSdouULBR5e3+ScGTGXp+FvnCSl8h733sGCcUu7q48MYl4k/
SYMDRJYCOgN9YWiXDp6zxFDLKcL8X4qG+kyjIIwrU3xb1drlZUU4QXqP1YMBlG590pYtBPemo4ok
GVZD7rlalc5Uz1SLNUqoEQ5rKLHjnAIWY6zlb26s26XfioMKB5tx5l+DxIq+t5cfFqQiRlp+y9Op
bT1Ia2X5JMxZqe2s7wEOSOajHszFI9cNYroNQlbr/3nf6ZJ+7FrfJBI1FYGVm/IQA13d2K0Syg8x
zXt0vJ0qDABR8FwRqb6QPyBYGMl0tx4uPREJ5C7Ju2kBwdCcmhV3VvWWcQM0b7rdwnN5d3koMdfE
3E1wdAQ6xhjjRKdwkOb27+dDWkQM/J8yZPVWIKI7hS6SFX3GNeovTk8o2o4U3jbtJJczNNTDPKUt
zkSVtOYmqA22RRjd6hdVLcnT+1nDEiS9WShoxHs0Ckg/GE5qz4y4nO7Dxm7ZNlFU/mt3KhFR+DUe
y8z3LVkKtCpsNaGIpbHIg+P1+TPg8zMtLAUR8OFxAngVPOxaSeQaTSRoqGPXTBlxbjOEH2n2p/vC
Vwh8e3u0z4RJYHTH02kYtOkHRtwhi0TnC7UHH1MXvoGq11ApTU8UmDnL0krNGwfnyKEAWvpHGQJY
TJnrgHH/ATSPrd4akQiWdGveqHa1CwzUl/CpIbJlCoIfFJXLE9tx69+mguCBrlINV8oCKlqkDcst
bzE52qA/1PZrFspp8n3Ql6bVUAWkPXRrxLrroGOP9c2iXfDdpgDp2lEb/7b5YNO6Vj7TlgdH+7wy
wOp1pwL/GUPygb83wDgIIxcc4PSjfhabVf+MkWqMOSo+OivC568ejIBoPcC+Q8GGLenU0Eyyo0h5
NKYKwAJKh7D9UpiYPigE2qZs9EU5nkIi5CgTuO7ZcycdlLCLfSPC/UKTFDo+k83DQA7tngM0pa7L
oghN2YB2GYppVExgwmRvPSCStzQeDtIyNdrYOCIvdKNrkofoiV6DJB22hwAdnWJOkE216VDfVFdN
Br/2OLV1hEMafCUO7yIY2aytSpNPVPXpBZrbDrX3+022hVGGovqYlyVFLAg6ZkAq7laTZyzyPabL
qYcXjfNBccsBg09zkjL6ovWzXGRBa1edpkIPnb59R/lP5Ip2eRk5/B9K3552HL2ZGjnBNq8hjxG3
xLtlQJxLZ6s2tR5H0QoJVyUoVXIuZ/SUES1avlkzjMWD04WOwyf6yxb4/Po4x2E/MK5yr37IJEXU
cRlyjxy00Jb2YIPoY3BngOWzybsJywtdvCkUf2m9A1hslfsph8b0bz70l6Q0jkOPplg+y/C2hrTX
oguJRCaHaTTYefOtu35XsZioK3lPUfRh1hY14hM2YZAquVRgk9cI8nVidZMp7exduh9lxLaKFyPi
QvjwbSlsEwfyeghN/BvakI4x+jqxVz7SA6CYCA44CxO0gWXXvce13K5mKE+6RdPytKFOUzO9ggRV
zhz6J8ofapfVBPkk0n6gyOuUqydw5KHkFXlKM++zPW6IHf+7FQitKz7qhbI3MWFKUjaokePviqGN
dXgZNmetboLa5WXWWg1uYVQXq9VqyUB/+8ZXt9o0GCtySXBz0THZW+RGMuiIJ7UE0CqQsRobtZ5B
2TGLo99NTfjhVkxi8wD2+rSNBBP6lxrjzRxKav0tcOVnXHZGu1/pVHiPZ8dyA7rTtaxQCPCK7fZM
STTHA6DbHqAzEMrUOMtI//zJzks19kK9T8wer8u7X5LthMc2AyOeH20eTKlTPiVU4fEpJyB34M5x
zE76j65FhdEEsCLGe5GtVH9DcjU9P5RZdK4dTkGR4Sav0pBRXONC04aWkhqTa3RGTa0iCs+Ly21r
heTkOu8Gwdpf9WFiDt1E/kspFLPbx/4pLIJrbWfzTzQ/qi+gjisI8NVJgsc/o95xLMdQwj+uikUl
LIfWcIQm6hr4zrpbINvooFDfNwPDHWLO3GUAjjMOfs50hh7FuhMbjbGJxXWIqtT51jE7wjmnTPDK
nKFFzwa/Sb82kUmsESYXeGZKJR+X+fuKgqL18ICZjz74CtXtVYO49ER8uZtCHM9ED8YfOtWm5OBe
48rZXDRwTQo/F2I6JXXqALuo1a+0ecV8Kg3ZxMmTd88YCx8s1kEJkwfmWBmBaU4EOijc8iHfL8dl
hiRCEqFLFp6DjfYyk3omr2gLfNaN6BsUrEFS2evmIrqxdsftpz/IuOGd4koLOVu4LICpcc7seTik
SwUkmljuv7eRatlz1IL7AKOb6U0rZ2OWpJyIrSPcWPXB4SvDPjQShlQ0R8dw0AhXogFmhTJmWGy2
eT2m2LdU9FlyL3NufwkKAZJ33Tg/UyrYKBYMFchbt3CrGgk0E/mGGr1OJb7R1LEEvE2db4xZEeK6
a4gAyv/C8rdeFoEZEIUSbugA6iBaq0d/46T5GFJcha+V7+SONFmS3G5jqATVZUIF4X56+4/C8k1H
BkbPMOSYs+fTtl9qlTVunFaWZw6VayBOJ3UUQY97zwJZe/R32m+gLMPuDjwyk4MBWQpCfvBZ8gKL
GFdgEfHoHrcgb0CbrKcQaa6K2Nm+ItcvVGnT9xvw/lbzTXwMBFMHWxEPRQzWtwuiynrCXP7e9YiJ
NWSOx9qSunjn3li0PsiOqHjA8uJ/Jmdmvq5GyR6Uw67441aVxh0kA5Ktu0VTgLJvcAA2Ws306P7h
fNf2pZJZUO5VDx+vQ7/mx+0QDKyPJqtla3OqQHN0nDJJu8qexodEjAbZ2ha3cSngqY4NMLV7zz8C
oiotsDW4gZkttfTd4K+sDCUlw9rnHp0dOFCfu6rLH1+YkYonArdT0kKmQtBkfKxYarokbVWGzyQG
qF3EC2RuASHvpCi2rrKtSO8EhMkpD22jo8KMyN6GmEcBkgGx6jyk+SUYY65HZ9FzJJ+CFdrOGyt7
Llr/2ruMcb006fayp7aJ77uPBam7oJnJvsb0C6yZNQO0G5FvlqTZ9essfDPcyONztzeHrCdk+Kl0
tmdIqjToZKXe0FMJZVz0iYZguCKkV2Jn/1p7IBmfBR5c52sPDLAHj74mQyDemvuL391BfvBUMklb
4gNGm2UUxAUepVUf3jtbdYEXeynEAy/avOu/qmmEaUq2iGNgp6l3ItOHdOwvWcLFuoLpEc2P4Iin
NPl0Xc51jGi6RZlpPbofC37ApH49j74/rFN+DFFkXDTDHvQe5r57hJxpk/LpSJZJ8Z1NO8ynlL11
6Jnpce1E9PXYbGetKT6tUtL2SEleaovVNOhKdV557PsBNiqc5MkEjuvl0e62+05NDG8Xk9CI9elF
sUjaWObsFPIuEl6I1VHVhCaDV+7FowxJspyN+RytsYnSL31IlKzZQD7zk2LNHj5gMQ5SIv/uWnfQ
UGFNCPtRkdUU+TgDyfrF8tTYAdaERM3u4r3EPwFI7d1sDsW4qns/BfffBuDOuCU1O0dlMQg0l84Q
jIpyH0rp015ZLPdj4laq7yrTAqrtMfh7Ay6yq/jLNtDUFOuRvaWouucoRfREfodH4+UwPZZS9qXy
x9raqai/BawxaoH+D5tkpSv+EgX0w6sJXkbGrFlSey04lOzAcXsVOJMAe2zpjuDdvUt9EF99uiUz
LYxP5XcqpeG38w/ooe/9w1MP1NbvTwh3PwOFpbLrhtea5BcyZjHtFA7dcmyMtTgGqGM4oJ2JncmZ
uOTKTduOsscZimEn7H857HFf8dz0OIVXhu316mIQKohvweXv63IcXwmUGPmVWPjSkBZ+TqQAA3Fo
pybidy4+tu+31Z+QlL4WZbVM6e1n95pnjDphSYJjUgcLhtjtiLsc15LcrBb/ogi9Co+gu1AECe4k
xNJMEvAOfDJsJ6No0VKrUvmFoTHQ3nZETxhM4PVgm/Fq08kEAjIh5IPO97CtlpRdbIBAU7Ugd6N/
iYlyVuLlzoBo8KWXBgmGkZBPfrlje3E9hTjtA7e8izpAPPWiZJJjWoQ3eYmOmq0E3BTa7vQj0AlQ
SNhgvabhm2uE3M++oq7EN5JqYfrVL+Sk/gJDjw9Hse14zAUsVxLmM7MCFypoE+fzmNsVFTgaWTNd
oJrb3K3rTy+f99UqSCJ44I/djfs5V9h/6XCPZnjPe6cAlfIJ4xLUx/oP+ra2RGV8KIYHtyMveFwR
Fe4DHSPL+5jowV8685gpxCs4dwapUrWx4PKBbXACbriLRtZSXwTCgbutxpuMFYSJs1ioakmCTYsh
UwP0DJPLluNHkMaX/jbmcWch2pY/XNDaN61RK3bmBULzRho9hYaukNvVGtO9AjIezz1zc/gfXBUP
K2QBVUwg+sbwTPj3MYz22OfNbehhqOlr+ourecOQpJJel4cmNY9gkLgJD8PzK2SolSDTQvOZ/5b0
oWJQKpuFRhSXTEd7UpMw85RkRjFWKfhovtpaMZpWIye8y5GviqXQHTpCGXDa1bPvOFrPM3RomA7Y
FZNhT1TAGRH8X49UbUVmb+q/SFs03S8k4/MyuPY0VkS3Ser7Kz6R7IZLRLP3xGMnf93yxVG0TeKQ
rg1Qww4PYsK9Ls7hBzVZcfOYeVs4nwTWs2wW+G4Z7Uo+4MrnWZvT+z5NradEUqCckHoRLXZ1knfV
pOvXOZH1g1GBHUJj0qDhTkcdxOA0cGXNP+tnw859IVCNXGrk/9U5ZkjAvlrbi8xbqDLXkypGGkJX
LDtI4U/yizY8niHxjdpOCewSKA0Z69z5xAEjnEk2o5gaeVpjynAEu0pff+2SKxxoltqN1L/+SL/B
7sa1jD95o+0+wifjYqT3dwG/9N92MziUwdH6ZwsA2LzlfA4mzFtsUocyftB9fj4ZpNy9EDmuttiA
tEiRQB53dH6QT28sgRyVoSa6YR9DGbgUyy6waejIVvTnGHzsmE+APXPLSQjMfiGcHELWLis9AC19
9Tc8ZZTeii/uGNxHx/6cPP+j3Zy9vn7WYt62dpSjyTqmzVvET6qDyd+bnjdyu4jwh+eOxDR7Q/Cq
VgKiAwGSxQxZrWR8zHYcJZx2uF/kfqUwSGFsMK2ql2IVdT6y7lVbpFUMeD4tC91wPRGT3rQc3pyy
IspyRF6to4Bo//+YrPme0vdJ5S3D2zNjiS11vwaakfzbef+jYFAI+EQae/WnpbwqnftgjZdshaEQ
OKefU65+BjdPwvcEjRm0CMr07M5F1RloBA10Em3fsR8v6l1E3ir3V05CJSDsk8H8ruDX6s7xWj59
WqCeNwfWwnpLc7v7LUAXw4ToQMf98tfcutEInJ9kdoLbRb4ERfy1bSQP3uYCKC6KnYSOFuBRK6YB
Kf3oLa6qgSIM174/e8L5UiBvj6DrCi61RjqY5SRSzC0xWUIxe2OcaS5BfShqsw3isrYkVjCtBd/w
m1AMsP8VnfJ4UAVuLk7SpWTlh2D3MDxImhYPP9mbw8Wn3LXtLZbLhIVr1yw4E2/Y0iHXeEIxh3Ai
Sjc1QyrGUWNVvMvIZqR27HgnL75XFqiL0FsrN7r5PGNeXkpzHo3npPB0y+LAGrE78vOf4xGTUWeS
3QZDMNvrvfhEGS/AIJxRbXTcEDdrB4O9yZIzVSIsigBhFVJRIbu0grlwwE9N5udI9AkoVBqyGdTa
Qaos6G7j4t4F/o8npFh+VHrq6iQygugTSQlY2VHlyq67DYNQyHETB+TzIBGDcwCCqozcgvA8CrHB
DvL52lbiu+Mtr2fGwTFZrWL8u6h/HwEcPhPzBIdiJrCU+yKxBdxtbPrXH9SbVoGEeYSh25c8c+nw
si8n9vatH+bDMmmK1syrDA5TttY1+/AELsJ5Il7ZrHQ7jlUyWmfEl60TcuWTt8fp8KCfiCUQsqV4
viqX/cNXQlTR4/amNXrlBfUw9yv18tN+aW0rr0Y15sAynQkxAWGBWotBgEASMdyVUxMWL2Q0QxDq
l2JZiZZ6RK/nU9eBOGu6FpOdt2YoH8iQKifW/sng2aKNV+EgSBdAv3bi9Opgb3Nhqtc2DghtGQ3N
CxqBrjzI1th9p8UeESmgJq2LkZM+31ene/K9/6yBRqDomGq2jdKdql1lZy3SJeelhTl+CtdxsiZW
17ofM1kmd7OcDnz48khSDezfNaGSMYStgBx6bYRJNtYefcDtdNm4Oa15zIHlTkSQQt6W6w2uqg6Z
FWW/Ct1owMtBjkSezzZaFKklvxLz0+lkto6Ui0zCSoV5JeGH9ipedx0FVqc/KbwbDok+DlAp//TM
hA1C00oRMbRJBc1pTN/slysq8h9MbmD0yaJGSbmtq5x57WTyMuM991lppWxUlMQlW816omLtlaHM
pfvRjEe64Xg1MShTGLa+Tqa3fY5MGm0m1hMZGqdovQZGKvQKZZOwjBL/Un7dJAdR7J900iUMoS+Q
pMrXb+8DWAe5KjdQaJ5kPeNB9+8zovIsMsgENgQ3xLnsOTesnxIXyLPKyOwGDtRl+vnsHXLG+0bw
xBlyeNkW/j2UiF7uZpDnqGH8CAhIhddZVFdPM+xqVgWXwPvqnuVtLceihpHgoK+h8/cSRUJmU5a+
Di3NpS0r+rgO14R40Qy7Hun0LmYSQrtvbavGW3XRnSRf5QJ8NED3a0aOQkfGaM5qEcLbOxFjViZM
cY3Ig4de2qtw4pqLpp5G0hQakCa+zo4to8fF3Yzdn75IFk30dde5JeoGBWeIU7SxvNoGe49cHw+4
AGEHnL5hXOZ2xRSLamBL56b16Otcp5iFCBhNdHjVDGHxPkkRMAnJ647UacteJ6F7PmCfy5AWk6vq
uWLybQlzw2voaz28elok/F1JKD006gAdrIgWLLLGa61n0jddSmwSqUOjPV2YONk/pePQzX5yOzUh
vr7DKrapqQ3UGwWPDohm+r3HjykZA64L1Op/RKGSoQ06BEDRzJ7QOrvrD++otMolRMyEE+QvvsLL
uDdQ1NcO8QOqrOSt6uFgscJSpnc6WrzQ+eV7Xdrw8omANixmB9XA03n66oAnvxnFFmtjFDD7L3LJ
rVDsmH5uK1V0Qg+NPDACtL3UOoSN+crhYIXYkr8hHqr9FkgBDSQB0ASGq7qFLZnXsARUtzmzHKI/
CviRc15KuGy5fIcapRCyMKSVGU0+CLF48QIqO3DYOhTTiY48iUfVlZijS6B98S1akhzt59ErbVDX
BBw8XuMUYRWtuyAGwthLyWj/pzStHHdliyke+cz7+RpvzRUsD1Pcvx3l661XPSY3BMzV1c2g3LOj
T6IdAdtpb5O0IlV4Wp5fOjdiHSngoznzs166Vfdd9KWrD83PJI/17juC7Mn0kAgfhp1bBwvoYE4y
+PYMJ9/T4ePUwQIyYGk67A3Ra3QpIh/OYykGtm+mjUOXJDqfWhtaBIrtul2f2mhCSm3E9/HzzVw2
cOH1YVh2M8ZsuwOkhmQjMqkeRsdzGdLLnzZB9OsWd7BkDZtw9ui3yiUg7+F9jQ01T27i9nXfSsmF
JqOhdlwsU3M8kDZOklFEenmjhwamtN/7rDnkIINdje2w5JnANca+7OTnxyPVy3YJO6DF/NZGBsK/
5j5lpcGltrCa/q7HiJJIdaDAAhpLZ9Sq9mzi1eQO1JMmvHixx3Ft49XX5eoCi22KZVbhxe8l6ONU
VCf3fRVhnIbFYZY20ZeqTH/brRfDp3aMsRL8dAX9nEW3WEdFL5BaqUOM4yDWdEGuG3lhe2x1Fkqj
HwwiwoJe6agYvAPqzmyLKIhy6td2r3Jpv140SuFshes+Z3AsjwyAixzktxeVBFn60tsPhXKVRbHG
5vE2JBWSzqC0laKsWVBkQOjscKvynhGcje0mRYClc5KWYLHNAH2fhp/J+Ug1ux/5aCkMzefshsvc
LUBHkBCJl4lg5H7YAJ6FiCZ70BFD2zbNpqxm9Ch9TAlPSYNrwqj6jRn/VI6kRmP8cOLLwCDB32JM
jcG7mCybXpqys37fseelyZaciUBVMn+Mh1yA3wuVL5JdSyIpr23AbS99RMI1IONyyQlRFLSwuxid
d6ERySzjYvhb+iyHCtOrSCQuKuXk6I9KoO1DN6KrkTMDzkP7sJlzVbkne5ipFoo0vzpWFJ1GO052
R/hB4isTY0tKTt9tKlAJFvSgzs4PX7iqgeY83SBcFC5feN9Z5AmdHnqZbq/dwaIn1+7xxg1mrMv6
DmWLPrELjet1IEr/k23JG7S+HHA5imVbpS+Zh0SUjlqNl3JBWatyLyM9TW137oPJLWOYmlPnqxkD
tv0AA3IY9/GxmsSG6xSLmssAYyDNlkMDgZc7R/NrXimvqEOsIlc4USTn9lmgzw9TmbXY9t7IAsGS
sKup/AhFaC3EklqKwyL+T8jcY6kk8xZ8XZ/Xdj3p+X6Jo1KYZHtZYpYBejvrZzjoKa/cZCK/M4Mb
89BDoQulJcPQ7/BJgeFpu2LkX6/HwB5l/UCzsVcQFigbDUJgD2nI2tAwWXTaQ3H7y0VJl6FgTeTv
F/W8+oUn4bykJjhpqXkAKL3sFT1vy/iHTaRZEZ/JkhEm69sn2ynSzfFBbo812PGcxQbRJ84nvIlr
U/+usCgV6l4pvLnuOhVTd8ibVyuqZYtWNqZIRI6nsW5rb8GtlLCSsH7/IkxPn4Ox1PFOBwn6Tx+9
BOUBVoLw/uSSNpeiy/Lhfb+KAXXJy9eTmDnXCNkizLWSDdL3d6gXUcaY6e7c5b1UlrYkZVzgEwfF
Uh+w2wv9DMGiz20yvQM4wjhfOQKv5G5eR+qFwfNOA5v2E2L6NYh1496qAwq4q+rX7bN7UM0o0XpW
oDYv1bbFzs4nLmVFcb9K8FTIxbC+awWrG7qt9Hjifg761v4OB0yqKFpZQMBYhB561GwIlUOd9++9
7EWQEmcH1cA5xnHco8ICDxsYzZTzQhlIahEXjt0dw+i5sGYl+9lHF1iwI+qu3mplQFmr3USrxTID
gGEMi9tZGZNcP8xVWqMYKKbu0+zRJxY19mcRrjgr6KNvSFMwgkSfFpu5edfsH4S3yA0kXewTaZ2i
c6C+bAET43H49SqFl4+IFGAPQQZ6rX+yIkapTovdjtJOuEE5ZFBmf6xs9AbRnsHzg1E8jeOJoaOK
nkqJcxhUV4Iuf01hPZddr9nK9fIlLAhnN7y7s/N/YIXelwucwllj+gN9m9rE5tf/87Dpg3Sd0PMx
FKUGWmAPhB3Fvwbewr0L1txE+lou8iPUwI4DRzLElosatC80aeou/lUroohke/9ZFOYN1wGCmriS
obMmm21m1NguVKJNrR+/9RwkSotlMEDikjMccmGE/yxh4A2Oz4ZjsmQU3jD3mxH2YjUwxhj3gMDi
BBXVEWdHCJHIf15hX0jXXLnlvHhEM8cCbKaf6oz+YVg5ObSKzaSFs+qr5OfLB9MtWigSDn2TkpXS
XeJBmzn6fqaVK8af6Xx08sNDkWt2J4oK3X07OpwA5u0r6M89bIHRUtB6j3NXvaiB8iYWmXZ5AHFv
0837W5SpxZ+bPxZqtLJNw6m8+F0PL6OBAsRJg0vq3iVaGjPWjhmH8tRh6JA8IDqKbsyAbZhYp0qo
nV6WPSf0xx3Ot16Ai1F5VDTtTLGLCHGnmkjZk7rPsx7DRBZCJ+hsVHv5HQIPXTq8Bhoo3O54gZqa
3gKp5iTU0EOkddtSsNI1YdskGQJ6q8S8VFggvu5J/C9dZy/fZ2UVzqZeYrLxoMW1fHUgoq9nsyx4
yK8Ot9jFx+Ylyn0DM/y4/O9+32naeAneYo52XN4ncBmpblmORoTzhWNqAwvgM+9ExA52BomV6SsL
DorsVCOSbSeTYq8uA2bwQCuLxB0eQ1WEaIjNmWE5To/4+FMdTM1abrSlX+Lianfc9YDEvtG4fZ5V
Jrpt/ukYqjKNc7lBqDD/C6WFaXJCZmqmHxefI0otS3z7E/pGENIKjRSDHtlX0Oj6CtnvbDDoZick
TNtlp+kMkeZBwkdnrqjOiu9ZaKqHDjnMgzkTWkoHE1izhEa2Gtp6vvyIomLCXkNs/rRBhDANVG5W
i5HypbJtYK5VECLgf42ZH+Q5Su3weghyCHjgVLUSlG6OBE8irkQM2BKioN49t3MVc5wx71Cb+AsU
N5esB7Jyg7SQxiUgp6V1LqTUEAcEQ9XSbfEmUbtr2PaTw4jM5hg5qXaYxHMDRPG6hyxZGgv2ghdO
AgDuaRfhM7gETLuEdU+fmjo+Xz3BYY/XuaoD1mvggg36lGOsAjyUr3J7xmb2Wu81MSjW/3v/Q8BP
1OeK+7o9ynshQCll8OFpjBYf7Bmp/89dMJFq0hUuFxa0TI4nax/laiPasxSg6CHmCCULi6JNTNdD
woIQ6wh9aDHlxA0p2489WQDBwVn+oiSp1G4uS/km6b6mM97AHmSmhKzSBuvXhMD4wXnt/uU1IRu0
hQWtW00FfYksU7neMRyz8EuClGOm4E8WlD2jYf8IHrEnKgE6qLHNjMndqP2MPdjSiooLnfe1CfnA
1euETUXGavwjDhtF5ybmYQkyAEeiUyD9QJ+wGhbqKxOk1MONfKd1+BdFnlt4+FyKZAAJv6P/oBgr
O0AELqcbrkGSKTmn7pmNkgaq95IeEuAfI99CXQuBKN2sV/GbOrAzqZPbbEWPQ9PpSIfmMj7JV/6B
44CqFjd/hP8RKKMDXCd7I2i0LTjrnoZgxLVLqlNggpv0daS39mx3PBarW9VzaoneIVfsEmhFwJnF
EyP1+BjHgfLzmV3MCmHOKIn774tDy0S8QyrklZxFlN+QNo2v/QuXcS22iv3eSz4pl79qVjnBo7w6
YWeLzszTmoEt9POYFIEC1UOXEO7Z7VyiQWHa2ps8vsDb3Uvaq1OoTOf0pnG9uXVm4bdQOzkdnUm0
TnIX254vvbgKqRDT8nUEEQ2voVVplcRRSd+jxKz1TUmHteCAw9yujH/muCspZ/M+z+4pyTut1trt
fVTcKvu6LqPfdQ0CEjzoZbhAHKUvP8o3DLbcVygnmgRvfs0dXZeFyEIv+mX8rggyY9QIRV4tFW1M
ZbM68HMNOHt2WJLMDdb7FjxaVPUvolpeAEl/FNZHpMf99Vi55oI7v1sT6wby6EE3hRu0gWXCcxGN
EN1tPYwc0wl5jSUMsY5AJL8ZrvZsCkgqTaEYG6Ln/863eMn2xPp24XnECOdDiFOoIS0clCsUYEp5
Bu+2RXpNdXACBraesWaaaVZY1ikmGCCESmUeOHDE5gCnuVm4Q50+s+SWfQOb7GHYVLA+k02+M9gj
TFYSZkjBvkDQwXBurrg5JwEjyCDYGLzS8LyI5hcOyPRXEqG+UdUfRY4MrxprUOYxtZ0wIr+OIBwy
NRWYoI98a0zUo2vrHLbxfuIxCiVGMLUhFdpwWcUujVDWlznOizoE/wHILXJSW6ddYMNytZeIcsDW
A23tb0mL3VSfa7lwLXJKmnIfI6CrVhLlmrb7UllgAklqvArYKANgKEos7JQA/r3U2HTX9WZJ6Euz
SiYUvyzLLV0qD06SCQhmI0iLdP6M5mfm/RpkgAo2Me622jOBQK4n1RRY1bfnRVrKQx8KQyJfUMel
M6Ju8nzlL5xjb2FL+UiXO9pF12RVXFPVq/CnYxNDZnsRA2PZYf3BYCs0LpHcUjYSAFalZZ9bIw1d
979kx658368UkpSfI2vSU5iqYqZB6mp5t6gZjAisURj2S1HBJYqs2K4vQ+P5VVjItRmG/GIXMya5
kE0u5ph+hOvWSpp6UgZTNb4wSfczV/sE4ZFzwCyu8nLoeqVj6zDOnSmy85D2r2SCvbwYLb+TNwgi
TPURSLkExAYZQHBoXCefi0yWodVo/8wdEIW/9/4JZ7SNcwBtHhRjhp7GRZlEL1qq2OgEYWBIfPzr
yssDan0JPlwzK5Xc5BP36o3u3HL9cmd8Iq44TgVJ4Sg44LYSLxQpipWueL6MBF9C0H5K4RTF12f0
fE/TfgsUVNtmBd0v4bNJSLRqtNau0EAJ3xWwM0ichEmqP0yMZd162q/UCbYj7Ghj2dxTflKG1gMM
83sbfA9yuGRM+11WZsF1wL8Qd8wdqqYEozWtKFcS9PU5eyaat+sSE+3sehkEdDSMp7kQWAr1MYCU
3r6FaBJJUL/AKGV9DR/L17TCXG4ukW6wzXYEqoA4siibzRdggT+fYFd2x2XcV2yih+r9KZQAEw7a
jTiaptQ8DhRM0zjyfaTJI43+9Tgez9atgn52lHL6VLmmytrokZacumzwE28rymrB1gKvBaWgJYGz
mRO5OIOk0dR8MgZ1MSdM5Q7q878iXZRpPzSBdWssYfJxcYPHi1LaP3JB37idZuEcEdEd9axongeV
h2A9fArcDYnuJD125LhS9C/gFyQzT68zvrrHB16wtKxO695KaAbqhapIvQ840HFZcCneyvcxRDA4
OkE7uzGwAEueGqkJrsR2ZzsDSvDp095XRkesFAIk+cso1DMVNgmtzrReo1Slc1s2s1QeTsOrSnBK
eh0rPyePzl/x1+8NbxZvzFqT7RKL3EkmNdyylztULhZFxCzj8zfmlq1KtwdH1vZu2Ma4gt7SKO2C
Nw+UpARGTzhJM2UYDORicIEnQ8+6PBe9+Y4bR42UgizAo73Oq93YAY59cMaQUVNIfZi2CqqOVSKU
7fTpWHasNhUWFX91u1tpbifgmiO3PMCq0iLOXf2Ykl7NBHT8HxnmsxF1C1dMgGkWZCsNVzoOy3Cd
+M0bP84Lv3jryqPbfJfYZ94ml0b2Iwgjc7e8qs+qLo9aulFUreNcx8TpjArokNdILkNltm/Rb3GM
Gm0evrezmMVAo7lmT60lA4unOeZ64/dm5ahWai6OT3xGlJief97i4lLwe3bxbqJNCvaaXipZRMS8
03/FojmZeOP9TNmkSRqMDnAdm4vaAw5oQRdbudPDe37T0wNLDLCn/OYavjMfMFNWa7+y6jDjuvn8
MvtFA0kDOCzQyW1AopD5MJ41mbtMmxUSmy8RyXug7ZeFLfNZ7CPzB+Pz3do5bc8CFYSBxrRSf1wn
ozy9YVdStr2hUDaacOlFshKXBFiqRZP+jje2sS3aG5ltNFSbAYoaIemJGN2u+/EU1Nv0pVWWCppZ
MPQyACbl6f6CPRDKrPUch/ygKSkXGrBNN0XBnjU3a75d7CqCJAp0kwcJ0jkhxpOKmV0ARkKo5XtH
nUgu/RDyQChZQ+CkgL7taE7G+LcqT5tMNNJFqJbnXbS4GAN3Da8N1mXpb4XW0r2XJ+WDOTLqR8tc
WTIdIK/xubVbe11gbja7oyMd/RpCEvC6m75rLnG1k3O+rNLx3X9Y/7BHm9JwUGF1hnkYuMNYh7qs
fTazJgKIrBs/HBWjo1qxPsmsYsIKpdhu8EvudcJ0pKechBK2hVLkZ+u8Dqekcy5KVvTwHZnbxVEe
E9Q9C3Mwv0lAAekd5XFo2O1e4vWDjhLyXyB2utyCkMRdDLC3w7fBjKcUtI8v2WD/d7Ws2QM3SrBg
ojFpVULeWsX63vX7ZJMellT2eTueBpT3cmNV2Vz+x7jV8kHcPlC6b4KHv0NHCMfrUn14hf7UkbjQ
1M/WPVnI1QduVZXzWwOThEwS8b6dUABahu84lm/X13b3BWZyNwVH7abakiBDmuiRLjobrIyCqqCg
1vBzb5DFuybk/hNYCGKAPdeYaEhnS/JnO3bDkuXT0XS7P/oJdrWH17gWro4sk/kkHDnKbD6TKja8
6tnOgm56SDKXmJ6hM42Je5TttiRKy4CMG/nWOQSECFBongnip24KuhRmvHmf2h6rIfTfvJbkIn3G
m91+5xmTpJlZYzKQ4jg1g/vdFa8623mUsvTDqE7uBcqUpXx+vh3k+B5G5wceyNmZifeBy7qtgLss
qruLv8ynU+FvlBTD9CCAOFFHrPMv5p4JU67ZV4/6S1G7Dux73SeVYlYF4o1V4Qcfu4Qj2bsdqE+q
sCPtJzgjb1SxCwcCpT581V3zdRu8MqFwKXLDM5TbWKtOlxfss8hJYwcIl4YK1algLw+T0ZacF0Ml
wQwMZ9SpgDuvxW8OJhOIoO5G0ZvKJ6N6xHRbMU5Xuq69yEA3GAz2lLjCNhlcSqJG8pg4h0MjtVoO
cxNyoj+1HyZP58kpXKdzurURD1B47A9Cv3o1qWPASuF+dZeJILV8EwG/Lg0yPXMv77Iyr0T7JPwm
CGCFc/I4E6RY5iXWx0dc/XEk1h4rynJUFF/q0kqcAacnSy+YN7ykw4bYPW10/33YUPInzu9Zg67q
z/htO4XkOWeiSv6I66EAUS3EVo81Nj37i0dDwx+Ih65Hiw+EuhWkDQ4/fGZmkuQhMkAO/L/ZJHFa
EKZbvVX+2F7O5p5htJWaermdBlBi5p6D7sCxyp7SZqGxusyGbHpJebTTQzz8lrR62XTeuE7L6hWs
I4Vma4rLfOAd2sHaXexkMxxFZUgLK8pt+rZvY02CMr5trMOJ+gWxTsk+kxBejgmR4Qg3pmj6FvNL
VlKKyo0Mp/z5pLRXM1bQNeLodxCpnAWjXPhNy26ZMl+MjPnJK9sA7xFfn6VjkeARUvfnMeSo/ftn
UEBkxMfAfXL3dGAfY/8smRHAfVWsqkn2xdpELtcAixhHnYTaXoLYIcivy/tipnQzt/NCg3F+goNf
tKKo1P29yQMoZKezUmeLQXdoNNpSS0ApLAW6/w/hMdbg/fNnffMMCtnAGKKrD71emepjwZkce4ZI
/4tBVGQpLfHjWd9xAK8lNX78Nhdv5RTzQrjDnoyhpvWPgtQe5qT+Hq36VjwfbKnHjqYRzCI8lkph
nzRD4XMPS4NuGDW6AIdr9uGCFC22XVvRiKV9SC7yTotUvWMG7ZnDUg52Djzrfts6rum+jEc3JnCk
uhWYJGFDcBzGPPRsv7GKsGNpuvgbUGHSmodIwr+da8hymXhN5DWUxUVyqlyxaPBML7avwA0dz+no
nFlOo1O/CUz7REYKjchGeIm7NWV2dZYp3Gk4Dt0t9XnZhLmOhpd8/m/HugPbR5wJV/7TGHNRGiG3
6F/IMewhKRi3iux8kOBfiB4Ua3WdoqIGhgsm3DMXV34AxJyJZ43AgvkEmo6ou4iY8xgXh5Z3VrCP
vETRGOI3pZdbisy0SnJn7aK3Ed2vkUxlIozynb72MQHuXASEmj7bk/Mka/XOCZrMp/mvVcbfx/L7
PNP+7ybJFvnjgn+asC+wLoR08sAjwZpxjySgfq0mn/HDK3fmF3wr5XsRb8+tDA+HnWZIHV/W0E9J
JeYB2NTZU8Ie1nGVeCv1vhCJDTa1A5kHi9BkYLoohNXJZaPzuNZxoL8DOhro5obSNZmOLVcGXGeT
OE0+hMpBxp7o/g6fDZZflXtNsRuR71cOiiIO3nCErVcr7isPXPiTgSIgyQjNWCBg7h0wGfVMNWQK
/L1EaZ0c2EY+ExfHoLxnfx8yAj1X+I3RNjxXGwI2ojiOSTqLqmwo/gFkLwcErHP3y9V8vu+pMo3o
g0aEQ04RtjcabC6WrUD9uv3DxvGOKIdqxoIp2Kj4OatqcRKIQ/z8TDr0prgB2BUGvXgSDxbwWCLO
Sh3v5TJa6BOFJ79f6P47d0l3hDye8ypT+hMMYxQ4j2it6bhTb0yss9Bz3kv1Mp3gzl38Zq00U4j0
SJc+Wzton4EiKFF+iFXj3akhFwjP7fXEv7FC+ttel/GduECZ/uja5x/ifF6tOTNKx6ltfu/d64pK
sg2nraDazx5bqqgrmtSurj+gwJ51AbrNUY48lqaVWufzZNOia+MPrDWxfNoooFsCuqtmerq1vchY
6geurg0/RNaAt1/Q8VzDofygfCQ5pzcht7umPMyFlTS6TuiTnCdjeaVMnHr4ZFcYXK+bI4+NX5HO
QcWyWWokCM9YjyAVxowx9jeQxt1tWScBuTeQZHnSQa2Eb3k3FFd3wS+XrdI4nO4DGTAe8QaRp+9a
f7FtmeDljo44HJ1cQafUIw4lGCyokRmh5zosSPB/6iU1oVazKkqRILyzgqezAmBVpAnxXiFjMnu7
zQ2nSbfbJDSTKY+fa0a1adrqRpQweily4MmcCKXIQBQPtiie1W48RL7AJuAtwL076/5DphO7qak4
GLlW/mAKgq2ILZny4XHMzvt1Kegc9eHwv/qcNlcfH4Ak+zO24cbelrUxFNPZxMQ3OMiE1M3/5sBD
CYn8ywZ8aQt62X8+W1KBa9i6OfshoMUec/1EvCMzVu0wNUgsQ67JZ4wm4c5GyXu+47nST/gEAp2D
H7K/DiyCXORKxxEv1JcTtoHMUwv6WM/mhHgR9HPNeigwqV4RCHPDnTeOUb1DQhEJKnfpQX5gYM1r
B9g9/hpUGryh6WGPY/NCM4e1vYN2usVfo9YK3nf+bKWYRvkm5yTvvE/uq7KoyPcnxjKWnn3ZnyEf
DH7Watou9pChjsiLdgPRtSJMSxr4cwCO0Spf1Z5jsmuDciJgVkY4yWAU64bNsjXhUMZJHs6gwbKb
OmyFWK7vqN24T+MQy378alSjd98JGhIZ6wBH03FcPESs1VsPWdmv7uzk4t2Ctnbt18hGZvbb5fJR
IHdKdTuPqcwLx7G3jzenH24adR24yxUJ4os4wWN9J0Wt4QGWJhiddLVBr3MrE0WYNVfN9PzZ5S80
pwFlNPNByufrD4JvsoJqG5mrCkgDMEyrT1J/9pACGMGsgfna6iZXwl1BSGQ5QOoddeHtrhxPPw09
MScQmub+v6f1QaOmRj/tB0hAsCQvnXZAFUcdNzp+HTVnaepQFPha21zN1fZofPmvdogHjQyYFL7a
+jPW1KZvG9UjAav/9yEAbjstKC92wScObmjJXgcNlTXU7t6l1OIx6lFTBp29HYy/lQk4ZVdIBW4O
hjglVh2o6I9d69ntP05opk9ncScRTikAZELkRi/VFoxr0lTpYvKkwULSNZJtnZkshb9e38C0kgxU
mq+ccGlS5jKqihq1BZ0179ICC/Fn0OnJ0Nj32u0DszPVJkqMR2Rop/7X9I04UR0QAgTdnoDZueAk
FNIXizPJxOX7cXtSqYR4+/MnSzYo7/Jrllbxz/bEnBfFx+RbwReNmcW+MPOO2ezlSTQ5Oinmgdaf
PH6WCAA3Q5LOy79jmtYHpSpEsoellCmJLelgPJvdAkvG2+lpBdKShK9QKtq0yZHzOLEHQlfKNERL
yNiIqM81KszFpSxs96VouopFkUZbUWVv5A+C+Tyr18alsc3LrMGhlg2X9qXTEj2RMGgfXoPMheU4
uhYW34L1kYixMkUOl1VxWSVw5qq5xOu4JqwS2r5nVdCex76t366xwQ+DNdxkd9r5WgzFEapPxQ1z
nxtIvmpIoYnMRffMhMdRxbF42G3XjqjXplVGzZDC7ulg3w6DaoqG5GGfNVSasYDUFLdMe0YmtO1y
cz2+Qf5uYKnm1eKPd6HHhgUszNfuZjwvLiXf/8EMwAYawuVxQG/sgVd/9PUTFHFPgzVASQ+xi4S+
3/KQzlAW2ILYVdF+pre0JCB3+5Yj9JlGtJak6/OH05bY7fjeham/QaP0tfOV6iULHOtaqykgiXx3
nEhSO1gSI1jOUh1pYb5JOkNwglRbfXqXe495eSdTDaolFkEytCkJfTkRrpM01ivIfLKmrEHp6K4y
zRs2Q1mkVL7uaOAkwup7NDQASSWofzBC3aYPo5uj0cR5C4tUdM7TbLOUge29mp9zAdzdKWthFVh9
2EPTecWF3qwlUIrzp4mTGO1b5h/cF9S2vgH1V5VMSd8+SIJWdbmSzCHu2pp74gMRbP2okufxK3N9
KJyFh2DD80bmlIuGAMw7aEciuqMyaoBnDoSEdmehdz8GmkWAg+AYYIEXCAjQIQFQxu0h6EuKiYoJ
NGccU7HLsXOLVEUsGw7sMLlm+5nNxzdU2+Jev4GWj5NYV/vbbajA4wiDvRYWiIMhh2UYNETuTorJ
syBk1T4J8PFN7dgfkRd8RkQwlsl73rBl+0y4C/kKai8An1cOO/vZWmTwQiIBsxHWyisap58SA+pH
hWp//jMcFnMCYovJXjwu85u3TNS+FGjfH01k3PKzEAL/FsnB6kpBOTPJixKHWVq5ppJJGEy8Iptb
WqMyUFkSudZW6fxA32q6NjkoE1TlLXumyGHAP0NROji2HqR6uDR3fXRB585OHZb/fTImQdIyTw+N
h8OyEXaN+Yv29Z106ujjgYO21LPWeQ+juknOZBdG1mR2drnfwYxRr24i9XGrtvg2uveGw57AGG2d
w4deq+WVij+9hZ5ra3suvcGQgLuSWd3VVOTSuYPPW9QmZUI2fR6a8v4ZHEgFDXw89oTELllVdICM
Jfm96/DOKr4SvUnguL714xNx8yD9yhFpN/l3lx9X0GnYgtgtvdM+9LU+gME3NgLTrO8pCDCWOWay
HaXxIlUrI8rs/QQBz+pIlDPzxxBnOQ3O3m6I7JCkmGbehacuvCc9yoBwMC1PxSvtg40tUopTLjWD
x7uE93D4wNOhgedOFdwGbA0gJJS31mmC95461h4V6m7Pzr9xxqgKkmIQHF9ezbSMVhzPnHnzNr0t
kuwnZGaOug/Kc6UvkGmZjAMJwxrjkBvmRK4pbfLvn+Esp/YlhqFHsiWYqNMoyAi6nDhKWlMI6C1S
MYj9POmp/PmsXKU2dZ1BFtTeQxDIJvT48N7tvgVq0e/1728fjB6CNZF6XgR/XrqLIsxXlm8DK0Ld
43JS99ybXbzB4CyXXKOI9Z7v56pCmNoUX31d9MsJh2rWv/ctmJZwPS70WrrrQXoz0gXsjkC5r2JD
brFG0x/CVEukXAEuPKeTREvetylXu3IPgs42KPd+3bNSWvlRu7ZT9PIr1JkCiywzLVo3iG6d3KLu
TtBeAIeQVPOdnYZJJYrxfKU0D4/9ZWiYEaANJ8FWQHQ4dOlM6F4qdWs/dTRZvqTlDec+EoGqtSTz
yISZgH0axv0TfwlfOWan3ffsh38eA3RLSVGRtqUKSJDhJuylmAILXDlDgvqlEzuT72QBFxlbKYd1
ZMxQFBfn0FORNmRS4wJS8pdamrIopmaLsQxniXQFhY4cd+dVINkY0m0Pd0ghydoEaxXBFOoFvGcS
Ov88pKhI1z7e90s5Q8KVdjRwK4fxlFQLtYYV4O+9qsHrAp/fdfyUAuJaNO0hy59W8W/Yz2nRAY3H
vwV7e0JmRMQYkn/Y2DE1aXuAHj6aaqTZj8mPnAMK0mJSZFrUQkE90JJ3GLjrUx+Tbo2mgPeMnHXK
kLpE0hjnW/Ij+qUwkBKpmI2tU/YAybr7QygzgHkggR6gpu4exYAEqXz1Ipwyyr9YqXh7sFfouONl
5qP+nPTUcmIe6NnbPYKZc/LlaHlz16tW8V5G29UqqHXSNXbESHmRjYfVEkiy4tmz14T1xzd9g0rs
qx5eBG2XCv94yeAKrwKEs1HmwWkrggVy0TPT8oe2V+1wiDF+IQsmzkmiFwvEit/PikHULR37Sgo0
PLJbBpmsEgwE4kVjgdhJJeJ6P2jU07Srw3JuwI3CBhab7hoJXTZuwFg7BnpRpPzmt388VKbdd/pC
e4FKrEHfXBObEV3zCIJxZ/MzKmTQet57J+aEgrLqHdZkhTpn3Fl3UZ4XiKeZne5V9RtavaH89At9
iuQzUT3Q5L3bDaBSPPIUUDUjkjJk2P70MV87TMJJZ9Ki6/mKwfQn8coOKptngXSs2K1K9iV/WM5B
xXLqitm6vkjrH+JIu7feAECyXDd1YrhG+gJDUqvsVcXt9xVIeuJQrL4JJzV2+c8mPeh1dvTiVFfU
ZyIO+hbF+SkaQuW+4eyvWpm4H2yFqpX2Ke279itIIaCHWkXNGqHgz2Fj30UoOUwYeQiAQ2TzAWHZ
jzpSM2ZzGoPXP7/Jf221dGxdfjmKQdEA8Oy+s47KMi6n/JwcaPBeMyfvjanUaYW9kqNWjdEv+qjP
ePfiY7C0DQ+6ETEnj19zqOXE9ub+FG8WlwYnvtFc8fA3v0sxsCprLU3lUGUTQ2owi4Cq1AA8SNKP
f/STDS/GufYaYejAP/X6APjPCnuBsZIL2B7SpocSK+OND5JKSAGxbPH2U1gwSCTkMgBi7I2qNXWI
wZYoEBNwOAei3kpfbVQTS0ZdIW4KokUUfE8ZnI+WHXp6gqKeFTE0O1biqRnyNPfGTGK9N2CptxyM
XBceVSv/5l3HnqW6Y1Sk/hnOrbuIZVy136ZCVmCoqiWL52AQI+dV+iaRhUu03JFBBVTmAb+aikno
YMj9RPrk/aHCrIsXzs+x74lw3DKVNoWIho7AsV7m3Mq03etL2m3daDZio+0oVrMNC1R4CRty7qBV
LmemYkqq/quKRG3SE76NagrfqMeWfm8jNqDQArxPwvnQ8Sj6wGLNoV93Jaxv+LiAnfmbnHyRYvDB
3FD76RTfXypIZrIztRVx60B1rVuPFr66on7bvOtru4QWbk8uzcGRslu006A5+W7hO3jTPfmdTccm
a4yFMV5fE+pdqHYzxVJrray6lEZOXg4G9RJW400kRnc1EF6zamz4sVsYG83SzNQGzAjjq0Kwe/0K
dW/Ugzw1p/C9rDD0Wu2kZ5ejic0j4Tw7H8KCXAjAPxuhvely/dIBX5pGZ02MurPt4j5+zQzIcXHr
aJdqVfaTtPLU7nI9yEDs2j3q8Iid4hgx5unb0JqNvt/AGY3jyqD8XSB6fltGR/w+BJ8oelE3pTV7
3ayA3VgGJSl3viTe8jniEr4DCv3fO1zdVJP1tCTiW8g3tw1Q9Xm7fbLycutuc6o4HSjOYVzMwMwr
RztMr5hsTU6KEjmuXAzKXTA/fOBxTy/b0WhJ8ewpA9W4dKzZ2wmro89WHVGWKAEWWtijaHB6IaFI
2UXEmjdhkjmRqph2j9D3mDMxCeAyVtAxCnd1ke0yX1vXISo2qhQCUU3vktYPdjh5RcRXqNO9xO3d
PlG6KlNBKRM9Z5H+qxzYnW1PcfoG+f7J1mTS61knpHEjo+1+ZAAKQ97MO/tyuzoYSXD0RjQmjgCR
ZTwhYpPRuYaQwKjlJz7Ti9Rn1mI0u7wd0q/NyLvGIOHPcAxjX9ToQMRblkC0AAcwEE0VMc6nopXr
6fgT7LBI3RZsWeGltFI9DsdkmCzGa1luQ6P7OEYh+qX2PGOgaBXK3aC2Z4VJPLsKU4UOimvt7fzh
HyRoV1usisXgTzUjzJl94XdjlnBUuB3bNcPygHK9iUn9eH7o3L9Zl17JPfwngm9C0P8CKgWOFX20
kgpgN7iRWgGPwuqEzumgWjK3ZzWbfVvIgbBbUxfwqIJtInBW9eWOgZZ5x/QB4L0gAjWNRat/jjc8
WWw/wFN0rH9O51cMuOi/iTToM83R+6Qrgj5SmsUoFAr4zFiwMdpqUnIxWHLHYcf6Puu+Ex86rDyO
0EcFInWqSBDWMhPDyZ40ql1iTTUo5eAJvoqUQUALrPI3RwL5QzXqBCdkntzmtp191JbwjMURmtRT
5m3keh4+6iKRw3HT1FeC+IwBnJHnJPR5iK/K/fFKfTfqo0FkJHwQZCdQOlkgWJV4oqTaYt/MsoSB
0N8DIas6RETm0X3njV4MXW+fq2JbSZQomw7QyqLTozcPNw1OkCZHhg/hanhiZRLi6za8eKJ3WWmF
jsn2wX2Qw26nP+x9YzdT1CQhjODT0sKNuuPrpUEXxvxthPvmbnxiVJzkTWuhTLNxn4i12YD5i+fw
DCDkmYV3+be9mDCtrxThvEZhAqwE/46k8CEdUCy8gifXUSGJA/5GT1kC8CFCoMg14SlhiZcWTEy1
NcZY6DNDhW4/ili1lf1bIGE92Zpap33ib730J53eD3MzH95K/gj2N+KcePGiEwYfJmFVsIOaRiAW
Leh9NT1mqd7DKyzxKYsBsw2YnngxsGkYjJekxrLj9uVN2eyAZ2x27VfQpIv8ZlPrcDMEq/saAsgS
HxvSTM1fIeX2baNdRVU4naqyJbbsV+eVd3LfibkptcQX6V9UAgs7hLTvQzip7JONzPCPalFNBSMC
oze4qCCZ6qnWo/IFLduFxZa+kN+2oa/k1PgYjDeCkbwvbVBdmVaRG5QyfIwvF0MzDPq7TPjqw7Qq
LTyPokE1UumE0UNigVe4VFrw2PSWibaMwCsA7dW7FDB5fuayK+M6+/GGszcZnfhzNAE1GW2bXEHn
dFBjwjbAxM1s3OhuPbkfoIL0rwQaWahKNjpG2l8clLIkyjm0QbQQFXmGvxQ03+EvY/7VD8SnG7Gt
Hq+jMW45MbyxZ+2OKUa4AbPvILR7DkVwMsFCDQiu7HpCaiGj2c66hm1UPlZ5mUfFt0iSxCYnuKV4
LBdUFCU8iGO9tzBFXkpTY2CS3nF4ON9NgM/iRc2rDR6otxdCBNia7TJgJD3eHm/2wNLxfNMfCQEE
aYu74BZjpDliCPdqXWpdr+kq6DzpPbiXMSBNQdmAI4Zh0em/VU/DPUeBoAHtZSa/gJ1IRDPqs10l
61YhbLJH/bZg9FiLuVVChXzmhT4IzTltH4HbJ9a4WDcYsvMgf3+qhWwmmczEviY4nZtNLiwNrf3v
bZnTryYBqsI3qGl2NWQz8M1D/KvM6cpOB+wm7J9sOXGE7GTYoHT7dKTLwjH2RsX5fllTDvVz6T4M
6tqq1KkD9KWrvAVQ0sVynj4SkwPliuh0cAmNHZtmibX1EgCUn225rnYXfjqFFmVhQlQpdOq7SzMp
OOe2sNlNBxF2rQutLZzWJpVBA1Xan3vL/34fSmpzSPMLvgZPWJ63OuQBqdip2SppNdji9SPL1shZ
V0Ey+MQZlSup71nQTCSZyplai86sKkS7OqrpMYtB6W2V67JCyIEfjrLRz4lFQVQj7nKiNho60B7K
srU4xuZr/hDiQBSGUFL49ijw4VUFlVARLPXLg/CRj834uyQ42rn1/HizXHAj4r3wM4X10uGDW1d7
2K3jd1tpY95+zqYIFTX+7sX7uFtwk+a5UibPhRO9AaBg+gpJ8BXz9CD79BMhL8PsLS5/YPcrAMVX
uplqJT79xCDq21C3HHsSUZUcRMMO+akKBbIKcYsbbcL9u3CS9nCnne0mGlGmWf0B+WMUInzW80Kq
jtg0eL6CzoKT7iasbOWhOpLGNrzsgwQgIgIHti+eqn5fD6iei+R9THXeZ6iu+2UxLPZYh6JqzGLC
bhJ1ywD+gdig9xd/JZenNZGXWAgbjWmTr7mrK6FTTqUr8/KX5JiFIzXi4uBuaCYIOAhkkswOPYSw
gouAq6VUN0iy0QTB4NrYDYj2cneHns/6LICdFld02ESVh8FewJ7InGomfEZkSHBqQWXbSEKq1nuN
9701rnz30fqfeefL+iIl0JjH1o3E53et+gKbpYrBHb2J3nffMuDbXFQNriNo0DRL1Un28BoxA2eD
5SMx9wb66jVXFQTFLg5YEcvjPU/zpKz5Ggq0lyDq1GwHUPmQJkSPeZ11SnxTlQhmn2A/8JOtUupO
R02i0w0+S9SAL2A/uyWvb1veRftV1ZgMIpQeOlVofrhQp1JsnVQR70q1C+hA2uwghkBiuoiHKyNm
R3V6erBACXUpM+RrVDXrR6MNIMOIXO8/8la2ZYeClTGbOnwBRd00e2/Wnk6Mdlv+y2nJWjhrnMSB
h5WIQfruIFRDu4SwpveGI/y4edq3cNaN3TkaokiVvUlx0EdFkjOCZXw8w5+wV2h4dK66ttZLyzD4
TknuJq53oinxguQCinvo+8eb2WSnltarFUESV7DHVHTmRdnQ8CnAZePNaFSXYMph/PC7YvqS5u3Q
dok79JZ7RIYvS3xSDqtmZqfM00mQDogUctU+FFkhcK7GaT3DdbkQoP3QMaZ4Ybyh4vfESKItixcb
AUFmbRaQvD4q+lNyFz7gbMi0rplcMPYo+phbxqBfusmMZfccsT/p7eskH7BhoBe0/2OSZLCRfQCv
b7SWyHPW++peOy+ZB98+uHyDR+WUVwD+hGPNRVRJQqw94cT8PZHivGDREFvR1j9TtzvKHAo5naH5
fLYiKbRJhEFOUoW0437Rdh7UKX8GkR+iJqqIbk8vXKn5Hs92HnSLUT1QjnaYl+uiyFfvRpOEtNoe
aD5ZZ5XZ6gSiYFGGrISVnsAplg8tE+zjhD4v1jHWNgnWs1DOf2/Hjn1TI8iZR/p+tF2ctQUPadM6
nG2qQRE9BGRBklybYxzOrTYxXtXg+kiiNZ6swMhzOa2l9Si64vaeIh55RugN0vEfMagZEQtOZBHN
NL4gudZHVZetdFDssWGmNtD3CJ+o3WL0gR+Bm/ukROAnfQGtJI+QD2tbqev6ktd/SFQYQ2kpjgIJ
MIWZOISUwWMkuMM83mX0D13nx4rggYGl4yk421Arng7H4iwDceb24A9F5OLHJQgiksbmWeX4XFGk
GFCYiaVA/Ah+KA+hvNv6zkRB3Ms+Lvga1GJWPZ/kx2Sm6eb9x/2nfNidewDWvkXkZNgN7QGASZBh
GhwwGHPk90iudfnmLuEnfwwLQO/8Pk3cOObL/qYfmBz4jvnAxNG5SvIYpBSfLnfLbF/vZHUUd/R9
zxjdPgwIm/BNk+2i/4MKowMrGFcDwZExghgGSg/mivjpENZwDa0E4C1RrLLzEMq0zr9TKLUC8Qwk
46HOi05Vzpimr7b7EjIdwHNVzXsvbWTK9lpR3rZm3ndFgFIRbhafX4eSgE/ODKQeD45MJsXoub3A
AA3aeYI6jsRfUKCQhMBofdyvp69Dx3jBG+/AB7DXVrZyG95FnTVjyDg4XhcibnUViBfrdBeJTFIi
rlB6h9UtWUfwcABA3cEy8Yo6zvFp8BVk/UuME4lfOpuwWHxj2Ck0TPE2m8p/m2YNaMbzXvLIUUBe
FfJABBRhffEiYioOr5nvnicUuqFQWsyuEiYP4Eq4Uiu18E2rRaAqbjDZjHc0n8JI5LF8QugNLCXO
2YMQFmxnU4ydpeHYJw6uQX2CXTxH2yj5Lgb1iIAvoHD5zqaP1cHdBbuOt2Bsdj0e7y/mxJSlhpEO
7boBWu4LZC3C0A3z7vH7tng+SHLHBaTLerk9GgfYiSOdVWRKNauhWreVVDnPa8P/PkvQA/S3HyPG
kL0Z0+v//kWDlvnndS4pGbCeTS8Wkk4Yjp09jOnbGM0NekNVIAhSTRHGxcfgJ3/mAukcVtgk4Cps
kjHRmK2qwa4TdsPYH6XyT5TlHHT1VCXleCFjg8RCFGW9F+H0lYx1wnfJoyxZH5rIwI9cPH0s+Enh
d1GiLEm09Bba4ydQ5Vb82c5ePccWJ5vY/4NYnXjOstVSrRDiMFutwaDmKp2JKDvxbrL4fW5CLXKa
A1+4iRwo1CoJ1wfy1dmwR8n2xv2t7/53OVTg/cZrgW4SNY2cTDJCd3I0PmdkaotxyFoLpefPSi3B
QQ7ZVFoLLktrLyedAPr/UHN9/EXMlIDAH5jl5OKHE8iUiO+MHfOqWtWpM1cCx0zj/wd94wOPP926
cxqdZSEWMCHUToYVOb1CgmAYEbOYyD0E7hQcsd4n0Bg6tCtNPPfdxUqzaup2m1pFdk1wc0u3BTFa
MLJ8VOK1hYsnIgIs1l8rZKovtws8ynjyVOzhgqHp0p84llp6CvHF5D1I1WvmRNr7fVX3vDqFI7Pl
7vXSdqrV0IR4i5KMPrFtSEQA5nVgNF0AeJrUwncaH5yamynQZmc941mb+YuU3AEzWCJCUrtEC6qt
c35uvEznCInLDmLLPLIf0BrjxWQSY99BXA4UPfdm2vsetRGOYI77Gm9dFMc7AUYwKoawHRw9BrID
+Lun6BsjWOKufZ+o8y3XKgfY31TNmUgKRRZZnR2IyNhgormw7yu7D2B1alSp1K13ERk0flhBYLm7
lYEsgypi+koGt733HhATkEg40ODcjLhNL7vT1X1qnlsLQ55KFXfClKthO+0X+dk/7Od09p5Phy6D
2Ar95r02D+wJcNVWHj0GXZ2YAvL86bfFBmeiPmXTYUn2hzJB9nwRZpfu9HZH3Niz+YcoG5sXcQk4
ke9tNPOwd2mpMjtZfLvQP1bM4M7uFk3D/3myXSKqyLEiWbWgPEnDNEVb4uGiV/zdZiTfObYMMo5G
/CVABOvyNgMw5q3zDcR4+SN+Ci1eBgdv4x1UuDK2WBg3nKEASb/rfR2dAn9CHiI1eR96Pbd2cTXw
iLXvM5K00r4L0V2/voOZaZ8ANBb+TXn8i7a+hl5MuPbCEZy29dYp0kXisQeEwkTg0v82FDG6j4x+
4cXWNtgXEv1DbCQdkKWHPnWIXetUwON9ftYr3MPI3Xeylmv9/oVUUZuNmeVFrcrLUciK5+8Ekm1X
yTU0mOKuOvUI9B2tbD6tCBrjMTtv3kMBviMysho/1W1AwIGNjbYT00JSNgDbrnyJFJ5uML3pjwR+
1tILC30YASaUapaA+LYzqUO9bCY0FeHglYd6RTWilvWauK9Hsi/GAfeBpd9lVu3BWkhMrNm8wnpb
g8q2BUANb/6Woyn1YD+f038YzIaxEByj3NwkmGPDcULBc2dEQHQLfi80L3C+LuPH4nq9iBB5mZMw
4D57BSN1kCVUfFjDgFX9uEEfA0qtLOnNIWzKvLjV6M5l1+iDgPrTiMaMkZwwFwRa/W/kvtmuploq
1ntxlCsgP6DLAXjJx6Q+JzdENNxXm4SVl6YbY3IlKuGKqswb2+1TtFYwxZSNX5kUCdt8NbM0DJdR
NdtjYYy8nE/iRVhQFhst6BNL9YYFboG1/H4wIK5S77j+YmPV592M4cKpa8xk9JJ3pADXak7n3WhR
/BGwGqWQazpGhjJI0t8sTVyq1Yvp3GWypkvUbh2bBwU0tR1AAaR8/lPjRxdUVvEWUjaBjPXHWA8D
WqRTCtOBHN+YIhuV4iC6btBuHgDhbPSAdZbqcPngrA65ySBua2Xn8ynPGsHl2/u905xr/OKN49vL
yeOp3AzbknAcb18KnHT6sFsh0KoEf09CQXnJDCjRHDJ49PWVIEpxj5lbE3YjMHufKnVJXrGQxdTl
ePkYoaRJXlGUCop+hwiTCNdTg9dw4TsDIsDS7fCOsGJWGSLyhNJV0memdO1eVEdPZOcvtIkfzKCg
3eNDqlfjpIePmDce6gqTv5Qa4nV7vifjD+FD5UyEj6j+VCVqhrdNF8qhbZ1z8tsiORvpgLfnRA/5
pdspx6jSHQUcqedrnDVXwVELsNMvw49bsIiT6eK8gYr2y56wwBa6kCC6mtEziJq2qpLG5+oPfBPg
rrnFMzxBtyhDPr164E31QGVkXXfYqwPoHMrh5prJqXfzRmoA58LjsyviTvj/mkSeU4ozrDLPego3
QJcfKjGwX0NZc9nrktkI61ZZ64yM8v1P4gCkrBo6rcVo68KSzX3vflLxlrRdsCYBYg91zJManNdq
iPAj4HrpSDCX5mwCCA6nrbZdA+vEepRhY+9WulK61SABa968z85xzgAtsgCacUXq1HL5S0QAL/yZ
Ie+JfgizlZJLhLK4WC2aKMoV9wyEnn0BaZTOKmmQP4EbzQwgxNPdZ2V6oi0xF8R/YgL+RRMfoVFB
Q9UYpKltTBd8X1QnGy/Njo0a29/Rb5JDqfIq+DWEjjuoDSC4pXzA0w2juvASSb8s2p08H5Tq7uDu
cAsk1uW/fHddXlhjlIT82RwNFv6C7AA0zh1yuaP94RRYZFAKowJX181tov2my6OpZ8X6tv5VvwrW
p+ONkIxamTSePB6DAnJt2tNlCFxiQaMEcQnq70nvggkARvX6vPxc4v5WXzB/YuX8gcMQRGjNpVDY
oF7MTwMrHe7SqYTxKFhgrgWt33sWdLrQ/AzQztXo3ElYR1ku6/PN6v6vIDbJ/QkkK76dYdO1/3Sc
EH6eR78wjUuQdcS/BsuJdL1qUYikHAAJ/+x+3y9iNe4VKhAlHX7/vBpygjueawvS7n6BHaZxleNa
SlcjET25brbFWB8okjUcgPTCUPH4P8iBQpT39HNaB7uFjWuS3rfnzkqQHEys+NgFCkk8WX0YKEYo
1cg4C36MxhNFN/7P1VrwV7QKC5XJ8ij3/dTMmYtjfnvSSubhAS+9M35LTPrrX/iTjc0HzmqjhfcI
+/H0eBT5cM3VivI7GpkvQR2Hc5MT59Jpmud70QCT7o6kblUOjIJzqRj+Axwmu1/Lg6A742cCq+X8
2UiTNCiEcNlUMZE4uUaG/FKLPGmMBaDgiCndX4fl2hj+KJ19+zAh7qpi1YcR9XgR/JDL0HkLk9vq
drHGBxH7d4LzPNGc5iB4vqTyT0fE1XdTx2dZKKfAd36bCsv81KEcNO2vRRtWVpxsI3OUdz+7ITzp
lVCtq9lA04bic+SrduG06JNcKJzxdCrzk87QM5QLMEbtYp4JgNgte6hqoVm6j6L22aWytzCnN4It
XBnuUBoxSEKVfFMgLQ2ttgKwKYsAoVbEah1qTEuNFmjejsAB47ga4oOqm/uJbv0uG2oKrgeoanD9
wNwgcM44RWWx+M2HelPnDrfCMioNZxElbsHspP2nm8Oo5nedPCqFxzGl4/0kwNUmXON5fpbgUEMo
OK5txur9/68XhIWIvQlDjI++yLDZXISMeujUJKWPxtNGq3ErQ5LPYyVMX93aN1GcrOzPBIyWTVZn
7pk9ieuys3ZZlorNeglSci9JvYEOwqQCEaFENeyO71FnTxQNfs98o9TBQlppAyEVRdE+sbC8r/x8
DZCCUDCPowTGexGCvfRNWoqBzB3itklGEej7o9irSQVRHWEwlZLfJR+xn5VkqAnnbcuy5M2K+mXX
ulVZQZQ46RFJ5JoPGkyKF1NG9VrKub0KkCDzn4FTEK9Qpg5U/IkVZ8lhf6c0YKewSN3hgWBbW58R
t+PTDgFEjQB0x9vcDRsF1IIPU9ZVxHnxc1m+h72/ONEApIbxudh54wSQu0QmsoPQIswHfNxLbQNn
+IKWkZ8LB6fByIVq/vtpAVdptzc+rlXCMZDdSZLqo0/vCuUJO8oTuGF4TqqryZCZI3Ad/WHmHxyU
OA3nBhsv6mQnQm8zjDi0PjQPLv6RhhFCQXImaMGzkP3XDmIjlaPYGngdwqB8z1xiPykEu1GkLF8S
yqryu0Fx3SJZPAGbBIlOZX15ivf1ahsoyuCAyYAOEClI+gBfmuCgaGFL9+Tm+XvpErHwzEOly+LD
b4xD/6kaxMZKhP+YJARF2tzYlwiaR9x7JtX4d3ko5BWIHOcEiKQ13UkmjiZGj2M6TbOABfTjmAsF
6tFernYyFTWfv2a+RbltxdXuNcvtsSX+rbAGrHTPSElSobX4EV5vP0EqCxMt7zmXfT2c4KUtFSWL
orICPFAR/hFKtehY5ABLrFaT+91C3bzxWLTIqsg1yxpOyUQkSFWnHRuWKk3fn/6blVgPowIxJ3+E
Az1gXvooKUBooGNJXwUsHuqKjJHDwWoGNkFWsM7bzp+qVJeooVIcbCvFK8wUKLy5oNhz8e07BKvU
GWoKYLBLp56BoBIGRjrvI2aK5wipsUFhPqzwr4UnmTLZgX5j+T/GtW1Xb78FhrjHDv0ROwKzuNR5
H+Ha5UC/GKOmaIlffhrUVNygXDzAvzS7hvQzRhE1SF7ZPTxS7SCCOzVdly34j5rpyGVXdhx3tZf+
jIkCB/8NrzDYnYw0EB45PqiI4jjsW5VA6nu271igGijOXeDfaFkl1yBcILXV830WGm8x+HA1BH/f
3M8orlHXxuUShMZSxjPodG/4ZRDHnwHpRfU8fDcc7zI5kN08Iw9QuWeSSIUBO2ur3OCSBxBNhEiB
bktpXwODRN3ZqJGOh1W/N5WN9vTsvDcfU9i5+enHCdk6S8HiKpSf49LvKGSWiUGho40hLh+PphHZ
mct84H32SBAH2FAy6sH5++j0RJ6AAOgva4wJlXPcsuHosPU0Y4uIuRZhlN32v1a/T+3CZ7Bz6FAF
N/9aLpAQIAXHH7pX+ALMKvFPxDEUKZFwME123suvOlyHg3vOBJZ7tDPkeqvvIGGxK2dQlc2NQOoy
xckarS537Ihy3rDTeTOFw6yvOOa0dPyDUR42GnmQm/Ex5G9IrzIdrMwSpgEzhmbHSB6osBsl1CGk
mipEmPUaLKZdPMo0fcGbO5hXtYrmhGZRXInCP9CPlUi/pmYiOVb9XPE2OpP2oVwozHbc7d9n2dQk
ed+SW2dV/hyzwA80rwbx3lgJc6Uem83Jzrg9aSTEaFWempp9/cD5lXXnX++LyE7jkRdDBmeryYM+
jd3Tc3YmXoGWW6dY+MdLSE24AcXa1tmgN5hAtOsIU9PkRGQT1DMRB9EODTh8qdx/fD59uExJ/+Bu
wpM8fO/sSO9Mg1SQZLoOW5aqmPraN3NW56ZU36ZfXMBCiSGhwm/yA3FTcjvIFQYiHnBkHOhzRUKY
3p5WKrC5eyYDzrCMFBRpFTl+wQnTWW4G9eYAVkUx+riPCzMo8n2zg3IWrnYmParrCRsbnhu9FETe
HlEhKpEokqUc9qMxzk8R/GIPnnRW4DavXB0RX+1Qj5PoryYsHpGpOw17AEqhdY8htWLeUbxW1gIz
OwbHzp7UnpHcrI+666n7B67OieQlBH3uzxuo4Obx0GNGZyGxEHbxYaSfXWmBtoZeFexUS086lIZK
iRmuGHJM6/JL8CCG3lPlJ5n83dJjXzctUnKXCj6/AaCrJHdDENtajhuEfvY5s3eeaO5VXe5Y9wVW
w1jTJ4ZL8/5l3NQScryx2/dPOKLGOyzH0wCyHzgMgf7PcmqquMTh6mIPO4RY4t2GnQGbGF8be9j8
EA1fqjjRUWu7T9RbetoGGT66FHi6ZX6fnDS8Z0E3bS8+fPVYOROIRnNYT7u8eEHU5n5gN0A0deE+
sXC8xF7CLJk8/AEnXwpjHe8P8ShglHnadfFGRyOPBdb8/MdPuMak5lYI/hkztGjihpEKmY7JafqW
9EB65fbTDx/9U9bD2aMFfO6hR8d5uBGqq7ffVwm/hncCg2cZqVrgnJiRVTligJ4tJyygDdmlns1M
qxAgPFonD7FVuf/u+wUO7jMKjJnfz8NcWTFyEEgA5wVo/Tye3DPCWdoWOgfvmQDOHPi0DFFlRoW/
csA0gTD6fA1QbhiZNJTHKRfJsbdr0FyZQNwOtp17tI+MENtoTLj4iRkPKkjhR5+Mj6uld40nyukS
ldTOKultZXxjx/hK/YeNaPebkF4/mxjar6XF1popPDrkjs6FrXY6TZoTC1gjrOJdZ9t0Q3zbhRBl
Q2hHICNX08X71oyCoTm/bT4ROYoJPTWfRLIdJGEOgbqYICSXalYtpWJ2E0BWdcRkrGhjEA+urXqp
2Nh9LMH1pWe2/Fv1MiQJASnlxKMbNm5IdfIbZnzVv6HyKl30J/qY9sPYf209GBGCmp+BbYckH3dI
pYV6aca6pvBIwK2DGNYF4keUTI175KscxTncJ8xyEW4HyIiGCDEBuZVjXj0xPUf+sTO2iu9HvzlQ
iD0iHynqldwhz1W1BXr17DzEVy47AIXHQHudSnBHL6y/LLKcMesBShsfj0DfSH2V7vpUTaubpFCc
4D8T1DBfDv/9cznjBy5ZJaqpyw6NXtUfiQmeUYZ6v+gQrj7fAHPU0zCcqtVaFi9LhU2R+2x8mm5t
YsPWArI8VUljF219pzJeC/Hintt8MykO2LCjsLMxiOSMbS+hXUfMzAeBPqSdXcZODaNy/IJJvoRb
ARqSpfAbr+Gcd99PQPvLZO7JruUwbL7MIqvbnoBkIMBVpa1g0N/0P7dtw2pWE2+DJN0Ws7Cxdiem
/TU4/kulsfK7djg0INMHaYF+wbvXe4Z7y70HYV2stMo/mouiICNG++nukw3C/eiJdHQ01WCmJS5Z
uEo2bGwpafTpzwuY2qmpUDMo6UEyqmU1iHngumK8yg37Ds1h/saP6Wkij6tbmtgvkhqEX6nhMUAm
AEk8GL0ZGezAPjqXF/jIekVOk3/MwYsYlf/CE97Wf+zxQ32Mmf9rywiUxjXw0wPBmskP+PYMyX4y
XSDptlDiUuoyDMN91RV8odVKbYLeMz8JMYUbP53DySZWCeEKzrKBnFn4kksF1j4ZipzG9VRfws6h
r5Lo1zZiBw0u5xHzVQsGz8vEBMiNuzUc1n+rR3O5aYUMGXPux/X8wrZIdzpKemnXK1bCxoyFCc9L
RvUNo/yQCxFJf3tnvioSmi3gQdaoE7fGuxGQUYQdZTBKQYPUFdjSdunwUMt3fXmTPwi0O7fGquII
qgFIfUyKUknVSBivvz+3cU+LAT3p7fuCMbfnk+/Gb7RlFN4U9HrTf6wEEtubEAZzOSQ4YdrOW8ua
VT04gJutw9wLsgmP8ojW1ltmg4U/h3tP9NqBIG8nLMhCVRYxXy1d2Ma9u95wUS/OtVunGbRLYam4
qdGgj5L2URWOl9hEyQo5m/E8ZkBvduTe//xy/70/nKgh9+ODI5wY3FCXfqvYz1dlPpIMrbHE/skR
aR2DXK2EhX6QXKmPpegn9p5t1d/TtJzl+mjU/PEIfC6xCTrcyaqX31bm767/RXk80GjFiUYIsndc
ZbZlDugpKpoxia+4yH8AbQxpZz9WLgc47vkEQUZy5jtUfQcDi1zYGpGdqv5FP6jLPs00Ve20Cl7O
8EyvXNtsWt9RrDWEjh6a3FMD2cGr3SwOH8qshH5t3loCfPya1rJmjw8/whHdWjhU2pqquAGnLyil
wXKtcIKi5EwjT2xz/9BKJVDbQbFD3ViW/f8AbXNrTnFruUBCDw1g26cIslJcx3KfxJOJViju7sbt
CnVNId5+mu32lw+mfqH6HdHDlQTZKIIPXNXvEL8TlFqRDS0KT81kv/YkWDij1EGHpUVrMSmykwN9
ntcaw0RT0vmXQ559Dp3nLADPxQmVKwB0Z+43TxRk4vUUCfvAxHweoMLAtuRc2mpS95f5c0vDMs0y
Ll06LcD0BeOnrvlgNRCKvA6WWgWc8w8UuLaEKQvyl29bzEgF+ALP3zvsB1n1/dW0CaKTjJGkZMCc
c4yGvX25Fmv1rplhJlC6uMOWldYeedmi+QrY5L8HWRZDoNi6SdT7HQFkKaD9dwZ+ja0hn6FTtuPh
Yll+Mu2K52f5s4WEjNC1ZTYc2HLthrcWWd+TAvqxmME9pJ8FK7lHOg8FdJbs2oQK7yqk7c4gADFr
p+lQJgE0QSWkBD3fWbcaEkaU3HY2kB35Q2rX3FICHB1SCEM7V1CzarMp6zsc5YCt24QriJxHA4OW
cARCuSG/zJFTX6lW91R/DMB4GGMzrsttSLxVOrv4tKrTK4+BIIC9DbcJf8og9eTlfrNSFcw+tyYm
J6CNuVedc/27V8kXrAwI8lSVQydF2nvDIwCevZFLLB5eA+BdA8wl55qoP2tMXj29dPTPHKFvR4ee
8IUce0yK0fFGSx5zf1DVXFtwnpxvX2dfuhD8gBeQOAu5X0qdjpvUxJL8YG8XcPkcTXYLxDy3WrOu
IQVBtD6IbUwpcxVFcUUFLKaD2gZUtPu9Fqnr0KNHkm8gPn8j6Li8mMvTUIk8kZId30wT2/sM1s9e
8Mj1D4JsJlYqVMyB55MgSSQDWfgbL2ea0d1mZ6AN8yfp1l0P4F5BTzy2m/0Mqxq/dOGSKtUno3BT
RSHThTsiB4kYeQLXK/yPeFf1V9u7nfHmrtSBITdhxuFajcNNND31Z8Rdfazas8Yf7+7xptcaxmYY
IyYmTFKa8u/ipWhbqo2yv7lRVhlrYFgoCUKprkiGGV52LCFwKUSFzN1UMlotrq6hb/DBFpGqwZNA
m3Arb7PVF5gr/nngSfUbbOStfgsr/tfNymBvOHKF287eAMsw2TO0IdP46+BEEi5C/4v14RAqXViX
hFYwKL7hfyQQMo/bchW6qDQeP65jPmrmbMyNO04p5EOz5JQKo1BSyKZt7rXMphzc8Ef9VFqbsZHc
XszrRWC9ub++LwNm0LgLrrH5C6YAbXaK3PyDadH8FX49qsZU3mYU/Pd7Q1mEkMhc5cs9WquFkdOb
tjKaranP+vFAyHpInvxIRkvXo8Nl0mzveQx4IJ0EZqMetkdha0WH70iDu/EpKsZHICvtftBDArSv
5ju0EDLFU7O+DvOi+sCryj9Y/kbfkvuni4H28gcLg3NzhOdL59K9/YOlxzDRzEGK3CyqZlS14E8q
IxMGBa/36LtXIkV6695f+kuuBdzIKPkZZ2iriTFXdAKPKUcsYewa4BAhLv7dCz86hxaOn3nj4U7M
wHBrt1WzuB7/NfXgEXcv1OER7P8hWxur5J+8fQ8i1V5yMdXG3i0wgWqoJ0TWBMRck5UXkjTC7bIx
JXFpsiQ/d2xtxVHuvBKhuf01JBHiejAj7gbl45JnPoy6FTWx3Exy+6qAycKaiRC6WpbTEcj1cVJU
TvC8sosO89Nw0OcPapC1mFKXF+96Y6rjptCmNX/mCY6MCdJJHsEGWi9bfieshAr4nEo9kxVCafzk
1Cl3+gZ52GtYPHbDYZwqeTY0NOiDbpz+pHK28okSvPg4i9QCIjOBf0xK1wLpXRQ6abk7CS5ZCn3H
8BENq3V9cgKSuM1+dFzZ1ZqdNrqypOaieOKbY+b8QoEWPtxAHCeI4eehZzZt8tjL9716y+KMhrFK
LcsoM2RENsGEHWdutlFo2Tz5aJdq2JNa3iS7HfcGjmX5K4wDlxLcJg04HzuU21wjSXMTOZTFy0S2
VTXld+3amYxmwvHtIALbU2+ysF6burbRptG+KxQjo6QcxmvQLjoXOB2ijslWzn/6qJKgXxT/Myma
ZVsIpyli7KVaUh84OiR+qiit0IPHpAthu9PasNyR3iQqGaq99biYOEwUNrMpMZchYbHxw831TqHp
ex22IbEoU2Z1/ju0k2jmzCOlj+kFNzcK55a/09Tvs9CMBSipIY/Tar8sPR/+ECNCQADu2yln2hCg
j3AMZCfuyvOsP5HfPJDxONQV520XqI+y5kcv7qaQykM1wHMHJOCNyP8A8HpqZG5fP+2K/Duvhw5W
CiOpHio/lnnIhMzbAqC5wibZCDUcVWidvr3cg6BfJWjuKGbVpcP/QfuFPvBWDr5KfaXcAWh8gVvi
VC3rYdal7nm9YvCe0/XnfJ1uPgxtTzkxTFmFjowpbbNjlL/EZNyb+DS8uXSQO6sd2+sz0tLeg3oQ
NZ1ZU89RMKBkHBOmitA8VP2vma1MMUsqRDCf50aM+kKVigXwikfzj56gSzElk+4PRgG/uIGrBIie
/P4Ytd17niycckCtsm/7LH/El9vl1SNUe61OFOHcS4KrLbZ4iwHxQZUF0xsd6ALZcwX2CY3qDkxV
NL81BJBxO/Vubyfxmv13PlKgoWM/dnSU0/MflDteOVLoIu2Bhjb8uzN6zeyX7LyY3G0lnLVzqsMN
AcPbuGhxFuokFYxaWr0sxQjRT611WEXRKwwxPsoHzBIbEhvTgv8yaUi1SYxr+y2h/xvNFk/TZJls
+AX+nOqQTRKpfJpkGyjrIoenk7ujbEiAxDzg+QyG+Z33Rh7L7PfKE8LeE5rSe/u7oG5CO711yM1Q
PNAw0lERAVUBK4xWz29l/olBIxPP8omCdxclnnYCJW/6d56eiGZTSuDBj+7RRqIzo1mphp9tSYMX
+PM6N3HTdfmvnolXEb380JpTqkrkdWv0EWlESCNrsjlbEn7QExQ/ZdSRSxz7PP5wmYWPSuORJkAd
JVixmzHhnf1cAFso1SeVs48kRQS7izNVmkMWRA+gwp29kHj05Dgye6vUG/eNrvct/WCW4nvnZwPq
mEzDL5GHxzDL6Y6jgxUD1w765T7cxP8xLr0yfCYMfMuPAd1y8y5welloG1dGHky8shoSDdb2Zq/9
A9gbdhZDYA7yDUSTmsGvXkCkpxtRoWZ/khrXAQbU0/zM3tBlCqOFAXUgPF0rn0D4U6pygiUujEJ4
qGC0qHiBAoY4iKndc+gkgcvJGqI2zjuhPdK3//eywEOOBXQ5F/WxLj+04O5QnQS00SnwNp7ftJyP
d1t/2ik33wXc3pOss46wNoYhRREvDaVzjfPcOVQ5nTmdlPLqgwdnbmU3UOizRRyuOq94stTgywQD
PC02sSP4yV7dSFev5h0sodXoxxrQhfJNHHFL2LHDdNyVTs2ffD/M/YhYg6/CqZ+oS8nRsaA7Cp8I
eoBLBABu9eY9Sy+7RvVcroTqbQDqgBynV1Ib2+tZFsbDhslKWGwDx6t5Zoj005Bs/E4qc24ZdL01
OJLheDMQw4HoOLUo6qHr3mTKP2Qea8pqMw0t+/mZl2z8B8lNjRf/gxZqnM+F9i9bPQ7m6RpGGyIh
kdbqfXui0pbvYnDBYkmep1aYXHO9ZOFk+2pDAhQPMv1lDCSAqAcnB91N9tLhuneYs/HV1wJ5Pz8Z
DNTbrM0LXVtNaJmAtD5/zRL+UhO0ft/GNXQlfpSwmnJqnagmou+Md6pXW6HVuL0UgXHOv840hz6O
5oDg6zOboQ1ZAu6qamJRLYgJsYHm0QelO0Skt+8iHGXtldODqG+sXGS8kqAgf9qCmS4vO2qTYEWy
WBrQmRwQBeuQJ8JaH21KccXntKVNh4wuljrWCrdkPqKVN3atfDmhYbzWTB60oMaROq/SNCn6eW4A
lxQWZCFiCfZJHm7qTJtloJ49rzqD2MFiC7T6L2fiC1qMMZzeRESYO4YX7p2+RJq0JprByDhTj2zj
/+LLAMjUwpsAT3HzFm5wcwkNfjqGQSOlPqg1F1sdhUU2c/UMZ9t4q07WIh8TSqWGLcInCuqZHL52
hv9ZWDtDgm7odQcomZa5n5oJGezEHruJALCmWkVsQxNDVc5J/UTx4Ushc4HGQe90Rc/+a2D83Njz
vF4F3RuJJjibwwjiphydaUvPdVZrKlOId8+B8RV2ur4T8Xs3TczUFPO0xUQ8Ltntq18vzp9/GySz
OvH8JpFPc450iQfMC5n3f/qoDB/bGYPwXoOcJ6kiNjG5OrDf8RCxJwrmvinWJ2aJebmC4PbeeTGz
K2jnmDwkUzme8GV/KKUiZl5hNYhXxlgiK7Wrf0IM6Yz4T3LvvcoN9z+iJR2MIg4fWiDYMrIreWb+
BtI03WK2srF289zqcGUp9rZJrGqXMr4kXay+VrrkJQffnpmkQU6qynL0gGt+mFKzvLZxJEc8vgsi
Om5oDLvaviQNQ0smnCosGoHQzDVEIFLVvJAho0R0QpKo9cEEFh2ejVsF78X0B2fMYWaXTtUBvEvq
U9iLY29yk9J7myoSxlqqkaKZaU1zVYgRI2HlBzi8mWFBjzLlR/RRWRByhW3SrFoANZJwrCST39v8
aA0R2uHpM8txd6gXSDpsfVjfhrkZ+ipbYqZbZF9HUS95j5WSu3WeLbAlQL39MiqUVkuq7nkW9A4G
upZoF6wXoEk8j0STvAo9AgVrboGxMgpsaXe2a9XEzc6u2OIcb0CO960uX7NpQyBnN4VP5jGLFicy
eHhOTfDqMFh16k4VhcAB4JwNuFQd8QPqGp4BQVlAP2K5yCPi0bzaS8md0kfGkN/GRae1kuz+e//Y
MNnOwEbCmDwrvJjqyvJYOJZXK6DaIH+4bOzTfnvzpb+BqwdFuMTBF9cGuYpBgHCTkjqXIQ7lBr+k
9VnoQNmFj4sWHfh4IrxHjRCuV4d73hD2iYMg5tSLgAOjTJkXmRRIrY8HG9aKTB20DSl5SPYzT50a
mKKAf9KNP92vyj6+F9hwbpd1IpR/kX2gB2wvKPzeucCSr7GLKGr8C2viPzTiDREH5L4WiALczL9B
tpkUar2JW9FZtaor33QTEsI6Q4xnpDjz3fX4yT7oTaIPL5LlutnQxnyfinAxNNrSAzSUzUddjQKc
1ujYmUepGyLkauPxwPHPLpklKIu8yrnZZO0ZFrPr479mQo5z6N+vfFTy4xf1+1kbPvu0kX/hfiqH
lIUFP4wuap7eSOQEbkZany5OBxh9oi4DitJXBf4s56pBJi77yDA8LmRl7PSEm1QYRh0TA8UpVtfj
zmVAphaOHYCb6Dt1tERRo/iqrP72rDYxlGDPhkKpGMXta2pSpefy7HMCB92X5AWp9eeqYa3S3ABT
8SMg5WhnZD/hgY4uZhXjpVh2L+wyTa66QppG6pEtPOuw9wwTzQixTNowXSoyhIML8fWTD/bLeyz4
lxl4GpbrGGC5TmKeG43Q2sueyiO5EAJIxxITR3PME8RggqZ3BLqBBTZoa5xRXSOYgyANnkzUxAxa
ZGrfCBvyQjH0GPiUX8mqFYiVD8lbvf8pO8lpDxh9864F+TJDaAfk1meHAhTO02fpyFBsrchFZCFX
IwJdXASYg8T/HHdMWBOECTYkboLGk6sdjbJFTz29pjWwTVx2GSnUPkWrmKx6tsm892PjI/tP+FYy
PzSDGQ/sN77KqznQ6l5rYWoAmVMay0tkWsCJQ44kO4bEzGG6N3WTdoSvHJJlpXwe7DlNbPRHh7N6
/WQzTs2JTfH0MTmfmXvKt1MwzmKADWRHCjA20HnuhPyCHjbFL94WCeV9PjuOGl3IRDLmjR1JMIhE
cUUtqrxLaJRCALlu2yZMe1AjnmzPyZPVd1RKI2kB1T0mpronur1Ntd9jBvcVapOd8f3xdyz3y9s0
h411QZnyVWrBMIQA4IK8Sj3qdb0YXRlg6XHgsa3FBESg5mh98P2emgJFgw392pqdLPEEuVAyvvP9
2CqgCLWqhg/c8g03EwZm55TrxBPgTPjne//EbnJSmNAGuYhORnncS1PjmdO5uZ7iuHQatwuXO6jA
iiWonjVdv5HN15kg1KOSyrg8nWdz1pzgUqBqJVpyc9paQMPRk6e8maLIZ6oKivM+PIX8SudlrUa+
1v1rmEIJfY0WDF/tNIHJOcvtQ2XlxC1tiqACLwM9U0R7b6vz7UV7c6UTflLgE4DbDQi9tVlQEUHL
HC20ki0U5P3H135nyQvUvLZ6P68dwKw6Xph1TQmWZJmH+el4Cacim5vTDVXcIOm9Ri8X0y4ybW2X
dr/DvdX6u/JRjrvJuhGlTm91fkdhQ4Sewin7GmO7cN2KEnsvoezvF0n4pEx/YNlqSmjOcZDqeiuj
t7YhEXO9gc9cls1x4osA/vUc94+BW915RO1xk3YrWoxxRC74ajC+Nh3iPGmx/sOcZLZu7igHjikn
0PMTbvjAhnyd8vZCyGGnaUVE+Op0V3qX7jVRpyiDpoYoR6tCGSQ3G/M64zk023TG0BLNv6a5TCah
qgpSHT06OAFKVGvX52Tagid6IYZ79G0w4lpqGA/vX9X0vjBqqxWWF4fjI1cMyvuI1OpTMsetRwpA
3J1gGOBDbYpBGNT9dD4bTh/tVf7O4c2xJPpOTTsdxOWYuse6+xB1n0oRU3ooXv8gDT49uF8GxPN7
wB5u8FBOTLHQDnjbAQFHoQnoR8Kf6VXeBlywBrrx/jHXnyU0Jpi/0j/rnG18iZ9CdlYO9qWAnMzD
Clxtru0XLVgc83XPItBqQGRUsH0kQv7ZqD6UbLWT2YbrNZYb6Y/f6XqVl3e/qokJkuVOq5BrBQYh
iUsBD8GvmaeAaSBGLCgmm+BdYWqzj3pfeJN7RSM9bA2Y3+ygnFFD5YaLvcft2aBot74e9cZ8eftv
M7RXzNd858IuJvdy1UMDDf/ifMAqutSBmlNeKbUa5DRQD2RKc4QMCVXpQ9YD88VjeAX2qm6B3i+x
qCElcAPqY/yxGO5Z4m7VIC/6AfNptl/I1OnoLiBa9bsEVUg9rs+CsQEaGOSVrz6hzKOny26ps4yt
m7VlGQlICawjmXp3/YjPznHzmYhCu4/Ib89nWFTWr3ORLlh/BMJ5xX3y2C0QHq7GbKgpK00b63cL
maK5Co25v+0ieEcig0MiWjMNPJG0g57D1a6ZVAw00NmU+EWq0lh//I/9YOISqGYkggBk6uM4E4S1
cgSr9qHDWdfYYhBDw58xABIJkrMs3y/tFSyGXgXjnr1Z1pAPegkpjESFRzhXaeKGYQQSlMc+1Bc+
vJ8jDigu0E1qBL5oydYuXVWWmdD3kMcHj2cw8DBl7fO/SGLURP/KrMJHhN5Drjgl6SldAsui51v7
Lkt9beW1pEHQOuVXQC/9q7VdhwJvS2lFD11tIiOedN9s5M6UVPNQq+e25CANrxWW0N2mWiZgsPPw
yI5qtQAi+D2G/EsCvYIxVGMmA7ubzjnCRUIBoQDoXZVGZ4PIlbR4dfjTLh8QEyqYibyRtYSomJpo
4L6a3Tt4TuRPC7ZFQSsEx7UwB6CVQpeG8etgZ26HbkYXHAaRRImBqj72+OYvQqIlk1sMqjhIK435
sA/rodo+xSvMYUfeapscJLesomANgG0q4OFT9UmuZp2SPVEhte8IT4xn1i6DzOlJ+MreeQBYI3ON
baVvl5IOJfsYr13BEiCzwlY868nyVmOyzaZwrwUQHK6OSsxEMyEnrcvlVqEiYDrAjerI8JsFRjal
jCDbVkLS1CvIgzrGTuOaJMZSu3zN3IFThXvMFJ2tefgzuJhBOJ9VxPJ1gnyTvGqkH+fMzlvDdU9b
wWTY3U+U0sjsUk1F1xpvUaHXRxnmmtt7+OvrbJ+cHYCVdn5lbcQeTDK+vt8rEGvrhcdEsR9zmHtk
vRlk/ERrEyIX7VNdemdRtTvAyx6v133gUxcTeumWR3r5JfhOgLwk2ooFTnrLO5Ib/0Eig+RIO5F8
uuFM3lF+STKw9rVKIV0bDKuQfxpSzmPRukHKDBMwNW9V9DLkVAOWdqrZCGBIYYgvnwqiukprDhl3
T5hQNw2ZvsohOKL+zzDXwzGoTSO+JBzTE17DyvfQRgTzu8MSmgJim+bKnlu6h8JSzQKdso/GfCZA
w3kTPhm+FUJaEIl3qlTCTnnqOIjuykqHDN2opC7DplBeXLeqgIj2UM0kNUYP65VeeJlj3pJoJUEc
F+2cRb1W+abQd0irBMoYmKLWl4r/RaNpIw873WFPi5FSn+UwJMEmbQg1uhm9DA9k36UoFoH+5bUe
SkZAE/DCAW1bGRHGQHIN/kAHSGdE+m+XX6Xnv0dW8WZMYe+LvhAxlzZs3ZO3JwEQssMv+Eb/89GX
5EtVLCrZFDlJk+X2tSTIP9tCRLX2liqIJsni4JB+27LVgxc+1qaiVq+HI84ncr9yGTjjz5gTsQZF
SsNtVGcPyuPhP+7HdfN6OnQFcFDh2ow/lomlCNSLyY1KB65Df9/UB7TOoRKztU/UZvc0h/R/rp33
SXynh6rnlKcnJT9YJJL97lc/bMDRC70waQKUDVypt7wvzGXPctJx1uskpJP80dJLQcTYFYnShjV7
DeLsSUH9+8dV9PCKtnRr5wTSweRi8yegEaV8M83HAeOAx7txsUL0SskY/tMG3Su08KCziB+a4Vqx
yejNEyAMlu3aoMUSPYViUtO/P3+g3VPaSvvdk4E2GkyWj6S6YGAg+7dplCwSxRQ/gcib1OOmF/2y
sVP0LREEmvXljLK8mRFvj6p5To3F9wn7OnJKhwnnM7rE0soLcbTSkd3vzjtrwI+JsaZR6zuQo7hB
fANfT+4EtKQJ9bCU7TpMi/f/e0i6bQvtfz0+2mMJRefndIoz5w8M5nvEL+1yeop5IKLbduoicbSt
p20FXAngmxObnK6esaRx1MlxrLeqWIz0HGbv0H3Wcag18AtCCIjV8BXmjtt2E9jlq0uk6UgNeSu1
BKljg1PxMnd45TzH6oVPRPsqtHusQM55Nxtt4DtvB8zcqtIxiFhK77i0ylSzIAHki4CujuO5nw0i
7aEFvdSRH8dUUXEGCQPQQMFRf3bXD/rKIWg1fGIOZs7j6QBmcIv5uHOCHAJFpoZ8WZaabR3tG7JE
jDWWjeHApRiXP6VC1uPqUE0fwYOFz9GLMleYo1HPItnm8vjzSa2UMY1K9AaxPeCtBPlcvEAONXAH
eRJefbgQeafA1lZI4Cg3P45iCZB6NJ/KXLwjpCYY4Mvi/6U2MjYUkyM/EC7/7BGqOSO8deeAFXwY
QgDHUjbWKSYwo3Y8SMoBcZL49EUPmZ+EG0iPkb1an416meU9oGpbSoH20d/AIN82phc4VSeB2niQ
k0UBE78Xg/fHJfwfTt41SbmcYTirhIImTmTVirtUwOuiH/9s0Imzd3g/DNl0ax7mnK9D6GSeUQmi
ZcSBQMfOwLx4yyWQ+ZHFANkHYhJzsZsqKC5vXqnunf+by9XXPyYPpfsWG2Odquw5h7nePTP081LB
F8VCIc5uicuN2OGGqmBClvPJ0Sm4CpnYTqSQlZ8JKrpUZn1B67y6q6cMeZtTQ0q4tcMAMznYyGdW
SswRN2wqb/oN12KTYqR7T8ZgTCevTsH6tg8pfi2w2NWRnh/HKP9p3XkVhWorYaxTYi40BxDa5KNU
8Jlwdpa9XqmwaVqM8x0JwB+5sUqjl4K6EExoL8U/m70XmZamvJyfZGzScszKmfp8TbN5vWEFwVyl
6pTqvhPwa3qE8F5n3M8KzmkACNyfPdLo9yrerC6VFI2dswMoMLXZaHjZJUHZiYE4su+7ENU6/ugq
IWGKTBmyPcyE3iNrooos2k0AyPZipWOXiVrQkk9d657aT7yHgWJRophhxLVHGCXGdPplUfAQMsys
P9TEc+S5iGkTgv/eUBDovXw1meqzcGv+6VAKUwQzLTsYRUPO3pH+bqhdbw3OWYp5ppqqQ33LyJN8
3gLVJYlFk6XF7udmOpZ/dsWJZhINXBf6fqlVrwHqI1tcVup7NUyY8BE9ruigqm6pmj+dNYZoyHQo
N5obAeaFBaFnToaMV/ABPpvfwW9Z4DeSFN+bSzBS1K14exytjAE7Eg/cZWEOd/oHqvgq3tf+udJK
SA4XESsCfNo0x9I24IKbjwGv6QVsj0ot4W9Bsf1NjNWCv0HKv7iwEw8QitdiQcRaeWoWcwpRHyLm
CCEG6wI9KouEfo0K+WT+XspF+13eRsXeX0+Oy2+ED2wCdG5VvDkt2q1tV+OduN+CMNkA0JtBrSEU
xHqsdXsty3kGxmE6DVnlE4e9geyyvZWPpeF72Uy6BjfyYqSXpw/0A9f6u2fRVaMc3SHqD1uNI45K
RfgMwjI0a8sG8efJpwHYWti5PrvycRLPNRBuyr4ms6VmuNvZ75PiMqvuoCqDtFWGVh6zUxkBMBCg
CPcBIERywHDv/pwmszcbpe07NFBefbrsKvF9t8VxuviPrNKIc/Uyh5Dh1brt+Ea+9Gz1UuJqfUDE
ohFTIALcXpca2805WWixgrYSJ1x3gw6cT5b+z/5ZHr+4gemPYcBotQYqcPsTs5v6oreKpbbj5EBT
abeqWKkekg6fa4xBGIBkwSWCpr24cbrIneIndLJ9W8I3KEBu5s/tOAWK5J2qPc8jfIjLIKHpShz6
XJcigTaYr7GP+Nik5kq+Dtv3EsTqK1dtlAm52v9UGaCruXgYeY0M4ZnDhLF3M9orcXlc7ts3sApa
onASEcp8EDzJjpDzPZPUfw7gEPaEuRxKVB2Imve9KUzuAOgtkWIoAHRfegcYQkLdgOIS0upcNynz
vEG8uM/6Q6oPVyGbW+JEKjF3gWndgUuSgiOf+euDjVTJ2tS/f1Ik4hrFljMKKySao+g2vldnKjAf
3JCqHMo62ALg5XRcAngeh/sJkdq7/j+DC8auWPV3WSbNMlQMeBSTRXn5S6neMYtjc4n4QaMcum/n
SdfefINpyYrYIZB+8ZUqfblWsxYo9hwFNflLvWZLbbS8+q7eIfgvP5n7B3fhaFMDRJnIe+9qgks4
kysLAhbF+18WOqAzE+repCHhPxX15UBaTuyq0zGdxV6x+iRUp/dqdAAhnpN7YDWKwp+9ZWfoYrp6
DKHbKTwgm8yeSYP/IOvwJCrGKP31xsqfJkR7n7p1NBn9RnWOcBTJ1uYJNIMPVYYivOi8uPjxQ7Rz
U1nZc7xp6oH5cGGE1MzhvdOs0pko/wbfcQiO7Ws7GHUR17Tp3aWu9FGS7EovIBqA+qQhFNAKuM+2
SWjoo/6MmwLDn51ERbdqo8+wsiIrISScpO0jo8cHFcOTK1kvzLMMdVQeuigV6s3YpOXN/vnm0sP1
1qHF+DHXUdtXb1xyVCxZ3IXOTDHg5GdENSTOcaaBjF7JrdHwz1KKDI11K1e4/tgk6s3Xds71CJ8I
WvhD/IfGCfGGrqoE6v2Jjust++zHkr/ewS+fjiUenCVe/IRaqhmbKqEpFbrT0/0xaCQaJjVaL7kI
tc+vUd7BB50xBJXPUXRF1d1hUnTmRpIpvgg0K40MeuO/dfwl+EtcLh1oTe1HvwoxSJfGN4f3RRBx
OsO4WZ7HDkYcBm/BPZnIjdxlXNbKIp5XG3wwPgXJ4zMgXWnqNFVtxLA2TG/4cg5SYOLRcmi3B0/7
GcaYr7fD7kethICQbFTPNI+tB7SUKcl5LZoGeaafKa4CfLcw4leuqsA4ofzw8ff/rxWwYAZ9yjTm
FiX/Y+MX2MNAUvBTWTqFNVny/nqpqWgJ7ZFaXX2f9m8wByz3pgAIXx69vADLFDnSIBlbi4n6RAwU
a3YaRM0FoSaRfp4/MahZ635bUJX9nLbcE6+kbqNe4Nb9WoYNNAOtyM1fpaFl9Q9Gq51O5qmquOM4
c5ulc1VFhLMLL1M8G8PCitP55310+qbXsbdhzQDw7Zagw12GhPDLdfNWb58PHM6tbFoMYj1GRg81
JreMZsO/r9o8xnK03Ok7jwRKj4nJEZaZM6rI9N6ka9wkrjExLm8yGWc+lCzph7++r+dKi5kzboX1
zioFvYdny7RZ3GksUL1g8ArVoZaXR6h+eQ+iki6f8Y7bp2K6gbvvSUzuYiOd4SUaWQ2uMN+fKOzf
lFO2tlkYLq/Sgg/axboVp6fxJEOyd7c8XnzcDY3ztlb1+pVuaCVAzAnCrg7cimUQWBKw8LgXvHMq
Y4/FYz1Np8FWZi5Ny+J0A4+58XGTjCHD2tLxOxD0c8qbkOk+QBp8EraNgjUBC6yEWCGAEp5TMwGA
HfmMPM/A0dIdvyKjkOBDAU/0DT1DJHLFIA22HLqk5BMSOAMizbY97yHRcVx78Bzg7zd1N1okM+qW
FZfEJ2RhUDN3GXPHmDYE3Wf8vwgZxKT/rRlXIjAcw4d35c+uJRQ88aMw10UB0EMOU7ddC3ydqYih
zX/HcCmHTKcPZMfj7fIoBNVpo/RXyZGHeXMSlaZ04sb7mWZgezSdHR9oASp8km47qAzj4rom3Q6v
N3m/2NLwdL3VOTWbrx4sbW2/Lx1neW6abOd0cZOpUtsM4H5ILzaF2eb9amGWqNX3yqSuPCMe8s8+
nt5GkGzQYcCjEYB5z6nDfjRL2YUWx35D+WEUinu1wgmGaiiHsiW5XSK9t5Vhf3AiVx8KzXZWNYWU
gWfmJfdPHfhlB2wtFF1kWiOG6zGET0G58n/wzOrPTsnwKFtmbIQlZ+TDIGA95m+vO1Q4OwW50NnE
rNPdl6Jr2kbW1+0o0HA4H3RtsFlgiKwsokGiua1nlj4lDkPMySpr8YHOSEi5Gl88Bvt8Hkr3h7T2
Hg4gNMzwmBPlHhQBUgWDINZ3FwAAiTa6N9bkqJYewNtSXSDFoFA8jHNCW2G+hMqe900I0UiFd6fu
NPgUyzfP6wV+TqeR2DYrBuN+B9q3v1/wLasZjkd0AWR3TgYdYHeh8uKkkQ/WJ9iAzwEcaJAPPj2j
ITCclyBiQCtBNnUXTu1WwdADS/VHWljFxb19uYgGjhkB5B+YmdnU8pwzRZJMobUuTH3slSmmfl56
7YP3pIHbz0L3bRsSdp2OG6XKCt0lT0zNgNdDpG5/5N4e3iWGQJDY5+HCj8HtaNcpG3dE5LtSKI+f
s1ehiiGUDIRxkPFLDJRHBNfmpGnv66F4vKWSvOU/OvncsxKJrrutw2rbvS5Czap/odL69zpLfztG
+7KYh7jD0JGCSfJZp3Ellq7R7TCk4BoSAZdoX5clZTMiLNHogyRlaepl+tpFiLyc4nT4NbHN7S4U
prdt2hJySoz4UB8M3yyFmCfJuzxmxN4L0srFRB1kptfRx1PbchaAiDwaNlbcrWwm6rVBnjf9P0/1
G5N+t988lY+emRlv/i3WUjhef81VqjBZbxjk+uUtqpO9UZG2WlbhM+u9EJe8U9SYa5xU+WRhBEqX
JY4YhRoV6DOKiHUtczrxGIbBL7g4iBj33Lnf744Ipzt93VmgLVAcazDoJ15ETvXI8So/X908nZ3w
zLsqLEa2Xu1lTmprLMuv0kzN716nkJQkeDVA/UfGJetm7pVpH3kdpkAxLHHXnr1cBKaytzMWMMts
PaeDp/TtPBwjT4/JWzdYXfI3vIVQEJzk/+mnkkiDEmMCO/ARYb5keirw+NRZj8fiWtkjzR3uc+tP
6yc8pCePwwvBQwDxemez98mhS86R21qda6xBKsDwaGlQjewvNf4Gl8Y4ttpI05NhumL8j6qw/us4
18jPOteKOhJKfHk2z+XlByeHCQ/Qyr+xY3AyNmtr0iraqSzwb83oK9WLvyE6ziX3x7QJ4/J8dEJI
f5vnibRwDpUr5KdG/oZS0VEoKGh+VqsCbjams0QeUKqMkjTePyKMmkEyfnZwdr5MY298T3EPXulr
Otn/rQV6VMDAbBhiU+gKu52srfSOzl3hf2NoU5E8yNOPOoIgdjiF2EppaequkqOm6IVGboziEXuD
1uffahaeFkcvM/Go1nSjDH8Pi5QXmjOogR+/FE+SwWh0Rn6eFdmwUEElkaYCQ4EORV9UzHH2ozpm
fa1LpJUvcp68NSstKPOAaebFO1hulbOePMF4NAZYQcsaNDt4JuzUNgbsV+62lytur6Bhn7BGEQAT
CwJX75cdtPxHl2DzbkcQixUDyRZw0sVeHhaVmE1kuoAXxLw+ISnhq24fpGkFf2bRmXMMcleCZxKW
XBmBYjIZd2ap9IHEFmfk8YyVJN5d/3SuCVkkMloVCJdqN2NOHsV+UfNzMqAFfIJdH1oadAbSNV75
Ii2Bmvf6XRgiSH+LzEHerbc6pjPQsgjWcU7SHAluxnDGI8pUoHHX9SyOoxrfFC/jhuzYq1IVBA04
ZAMjlifApEESu7Cd6f11OtcMEfuVJ785JfHRwfmJS545YPNX38MIn1XcfpeyinpF/+p4HTXw/vzR
/25tHDUIc34ZHZAuFO2AWmoERN77e20UEse789IfPonV8lfRQLMmMZON6IyXAxBE2JhYb5CMGA2M
ndnZcGaV4LuxLFoZ8V20qN+UU6XZb493BZMRvTN/KNaijXtabYWYcNpzmJaNiq42jq8Z8XfcMVGu
9xLiHqXWmtqT5NaKZgzxsBrA5K/WPYZzjoM7kzm9aYsiBS/S0Jvg7MUX0CDNPdTU1yj4/Op9pT1o
T3FuoKJzd8nsY+43FUH9u/9Md7y5/BsCnqO97IaR4tkEQJ7LoqF20gv/MuiEYXFU5A3DlW11ZjfL
4eq6bt0wjosKQtuNzQC8ryTGnEYKSg76s13wAP1RAbPX2Av7o2t7qMo/drxtSe26+Db8NnVWPwAk
q71S6M7+D/4TUBbEogGWeT7q5NaYPTOj25/bo9nOs/+r2UTY+5k2plTUi1wJBENY9Ooey4MVPxx+
bDS/+aZ04xGJUqYKTsoeXplaDz9l4R483HuxfzTnGZiejbWLY5OKQBQCj2WpSSfyyNMs2kiMAxQh
L1WgFA+hbGmcZYFuVgOc5m4cE6QEq0612WPaTHaOR75M1JEL6zGCrQn3eGXsL4HphxmPXaA02727
LbCCXnjpBPXscZLFFDyB1/DqXKbgeiqW+KcUiGhf+jaAJbQfkR3Hi2M5F57vccAviPDCD7lx5IX3
1Rhj9QW5KoH8tVL6dhkCe/lLLyNfqp/gGYrKlZDsI5FbFpuOYGB75zn7OybeCNyDxtujrY5mOAZS
OtlEaGhU+2pVLQDMrwfjCkya8GR8OXaWbW4TAkVED+6y+tPDsU5DGBKy6WwgV9POK6utev2qrM3q
mBdh84rAl7FtPbacriBncVNuPR7v7BXMJbsanWEVBqqm1OtlJ1seR/3+WnkoCu4HRaaIxs63T3Lp
VPTMlB/4f3OBS4qB+ffPH4QtWjmfNwvMK7MoB06oCoIHOsECUKHeGqsUKLkiX8V8/CfzgSgxkNaJ
22HWbGtHTOYlm8xyojRelKkZYh8e758gQZkZSlhw5w/xYQ1tbSVnAvd4x6AJ85vg+plle1QpwXzA
aGFaphHDkZpkyPOB8JSadXADU2HuuHuf+/UjkcIfg9ouQPajdC9qP0K82oizlGvIKT1eVkCWXA7h
rrkd13tD5qOmF8q0TWBBoh+LSed/gJs/V4pOkcNBjZ19OkfcbYbw9XSQocJkpnQ5kb42wlSsrGQu
Yb4TkK4hFl7nSfvWk3OQh85NRX1RJ1SSG977S9u2UYgeLA4G6Cpu14Q5J2FJYd83aRjjcKqvUzQ8
vA3p1ZPCxH0TxnjavFgk0fe4jLjchk5iAWUp17+aU0h9TfnzoELvPHDf+tVYhEqj7CLU4DVh+jEr
iODyJkU14jPuJ0uuQAOfQFD9kKsdnGVjpoi3Jaoyvz8IpRZyGDW/m3uGxfkY6x09UlVYt7PkWwQK
PFsY7SIvTGzfBNtOOlNr2zEWFluIHrNvrP5rRZ7y6CVuMQWtTfR5zfjm1lRcbN06sMXYAgNWx/Ul
qKM5cX8+Y3pu6hxDuK1czZGtYU2u4obUD179zmO1MB5rNK0dlscvdToA3VAZsawxLyPIIwvumRO0
d8o64juyhaTlyz33TDebrDln4+bu4wfwRZ4X9YU3WXY8msTl07qmQ3Gld20h8JlZ7fmlvsumLLdy
TmmX5o/RvPXoRhHK5MVq70yC6eXVG8HfsikoWniZi3EbSxDA0EkmqgHaWdR8ID8PLonItaz3H1af
PbcZO2yaHPYEJNtAWgnVpsk4oRkff9Wh+vKMtotRZWtheWBR8XTtdupdkVyq5us2HJZq4gx0CN5v
2AVxZt0CfNwXkbSW6HQwVgM6CRsuKIobIj12joeASz1YgI4xIeCiuKWZokB7DWdkn2JZniJVTbxB
aJI6Vfx85Yc/w5DuKRiNiC+UT0WBt4XWMZlGY3Kd6y8ri+Rv7M4S2mkfgbjQd3diTr5NZAoxGz6t
z1sA78ohmpJ+WTif/ZFnV6U3gQZRkhwzszPCpTA6Kfzi7p2OtExUYsoh5mdOCPfRxkygRfEMEbsd
Mh0vvilBhHW5dfaVc4NH6HSvhoU9I6PAL5snu89512SYQe3YMsFRqkh0R+vjHm2yNx9mN1CTuDab
2Y41DXilRoiWjbIAOL+sVETpKSgOdFxI6/LuYjE3KfWn1S4REDdiIbOYX3er2bAXmlyRS3k0Xu4z
HSepb2mC0H/hpgMhApo+uiC7JQv8Pin5fUUH/HYv35z0+dlmQLTHFQ5nr3QPckdVtSLhtcl5NJOt
C7ChM1t6tKZX6vSxZQt4VG3UoDfaFqz+M2nYa9UX6cPeUgbhjFNUYRkr1ORlSO9yRilVb8soHwLy
C+sGyPyLIbKGgjCdTdAWfhk10ev2sQx2PCX6gXHLE7ieEN2MM5d5iBMG5wsXFpwVpsw0+YczPkSH
1Nsc3kUuaWCqhtIp2VLRGEMKBtRhOGHUIgvI7aUEEFBp7EdnuAG8EsK/TTOb/BmcP0ZgQDbPvoZw
IS3k8watiwC7IZs/guJSqiTwy2wzVFbO0m7OsL2ODdrPf+uowGM9HHzLb7xL/dX4SaXTV2fbs2Ca
vcTG7wF/JGYCsnV/0LWSyxYMEkDGHqIG+drWtLYFlw36eqm9YVhn/y4YVzqp+YUkBStnj3jrU3sR
OwsyiLtFeD+3rvik66sml8AeyhSSNDM0ZxHuwfDviJIt4oduKKQi6Jg+1FQP00j45PGa0aMjJar8
Vka3uJQNSqPSnIszqbtR3titGEYVUPzRnIOWn8/8CaaQgffx0THPyKpjP1dGJFFavLQqUCJgBIo7
xsqOqPwQkq5096PcXBnKkfJ1fhjS3bnxaXmVYgCBwNFb249ckNrbXkr/e2GiZ5HmxjaFNcu2HK8f
cwW9mwG8pmes9jMytlzGAtvG+kdsUMswdiV3b7PZyCsYnSOFejMFyFI942zPMYumj2vw9X8V3yEu
YitLQj91siyjkl2l3DsGv341bN901bg9tqu0aXclawu8orxVcQMO+m2hXf777dbu2nyXfuRx3wWp
ar9scTZNvyu3shhHj7jNkfCMHbiKrBnY695HQ5+IqJqnFO63+oOAW2G90tFAeNvCZnyecEb2suzS
pDTDOjVG+P8fk03Fv3VqCk1HtxAGlZK64y52PIHsbFiXGYsQHYYUVEoTYEdlKEOVcrVKZ7b8GOJ/
rdQ4gKJVtm4giAiCkphipm/yNq6kHXa9WB5ccQ5JObDY6d0+N8DWrKSJXDSbuT7d9XgkpSujtFk8
kL2fiJXo0chRZe0niFilf8A7uJeooi8wgmNuGCuwlCNk2Vk+DKR156WkCs5tGAChTp72dTDlab1k
oNN4wPY8uadMKrMlLENofTNNq7Xb9IFwGZ72yqviT/T7Shb2dNmNSMRUksCSisxr/7THRUQ+mL2v
ZXmg7ebBMYhS6G/TtpUOJByiwQUgf3KqPWdZj0qyFnQ9r2mw6S7sgo8IPUYlUJU9OVBkGq3SeI/N
SpOXLlkZODufPNVHTxvKtECJOy9gJsXwHM/NkuslkfMx4nZC7K0gPREApdiA8hHxgUlbDNqGz9sE
D2fSWhjbEWk+DeOOE24UC9UmPs/o6SmEz09+NpbEtZnEo/rAqDIO1iupMEs4kq7BxUM9PmVaSSEE
Yu9UYa6ux3dk508tSjOwFIXX9/yATEQfI8T9xIH0vneXt60JkNopmGixwt2qPKPPc78Zxfgo9aPU
MtURixxOjwJid8imcVrovKui7ls2mAhX92AHepFdt+aVi24EZJnfFH8uMsQ8+JqckB4UvrKytmsv
EW++do7GNQ4xwHEa/n7LIHgEXwMCGQWAPNNr5tHl06XwbkGpAJVD9fs7EYq3TyiNsFdiPle8i0Kt
vIsi11YTylGlaURAIAW1DYNzJmQqZPSu1LDEiCcVtwpGMHQmnyDr5Z33Bz/ptsJ32wK948Z9yBiR
at8TkwRCsvN03g+A+hkEUZOwHpOMyfZQnyXUtSL+TgKZrR7Rjy2XgyRpubD+i5/YWMMjBwpwM+Pc
BLcnclIf2PPFvSRKA8O3d7N0rMK9G6O4ckF7pV5DqygJ+jsqxVt8PK/2DCY2hnZqoFFPkAnNcbrL
Vo7lGygm6VKEh4LHFozWMwmdo8D1UcYKeQx50Vpf1KN3QYIv6ukkCUsjLHCcHh3YT7ji3Whir8R5
9072ELrD7GvBNHfKvAAqKJeT+2JOKNyvgPDCddxlcB1uURh9vhrGOCGIgcBgliMgAN+B/7RV9JmC
R6+9oIeFoPak+E7kgMtCxon/B3EQyKeEU+83zF3AB5PW2iNgG0ExdIgu416MBU8JR9TIbqLMjPJE
Q0NH2eZcw6m137hsFDnDRp0e2QmCBJm6A0rMieQ6PV7fO2GjcjNsJDYVDXe2UiLUqLZv4ZUnBsTg
smy4fRCmFjyBR7fmO++hIvXvfHFgh8uKxQaH3wLl9nuo0ipM3G964wTweXSejWTKtRjOvmV+2Vr5
HviwiKotm2lxITyknnHYmOy2mINdwfmAqO//6h+zma/C4Tn/6y3ZJYD3Xt9EvFxYJilVoPcqbGlX
jTh4bGLLu7tIAVIOZ/yNBNHN7mN+O5JQ7u3NY4HpS2WgK2hJHF9gFfqeIBleRCwBSRbP5sO2comy
OIeSF8J2bKApUnIF/0h9f80AbmDKtWP20MDTSXdwgnBPcjIMZPqIrmsJg5OcgdMHAi2r7TgANOCw
SEoYv+zG6T3H4FZBfzhW1OMUsL1uuOlwOiXn2EUZj1+/bb2CefkZDOVLwfrsTeyMg14NQ7WnQYLT
91uBEmcKI6F92ItS+1xrRMKb4wx3311HBYX+spZGIsM2MX6uIqW4coCDBRUoqnNgi9U0l2JjEdbI
HbeoHtVQLpZA3u2Tvpt0O/KwiQf0rGDv+3mxYdvJ9cPjPgMe3bdBSc8LSJNwOpE200OFl5rbGFsH
NW/LuFnOGT6C5fuzxHE1ZxaPeN9Fm8OX+4B0YBpAJ6ux9X7WT2U2wWtpx6YLGbHwb3ZpeMrcLU3Y
hdubsFp6Bob5tmxRLMWh3nIsEBbyWvcGxvksF2jYXu85k4k3mas+425rUXYrjGx5ov5EHGRNKop7
XniypMMfVpYHSsuKGdC3sZwZ7jw+alddTqTy05kcTVphpWSDcao7LIVyoUdkPZVtBaaDlrqvJUh3
gAGPOW2g1E0s4oQNWjBbeMz1FTQ6iVFOD+MQId2g9mgxgfLXjgYgYz0QXM2wAnyvOlBEUM5lp7rE
wGKMnVAofyN/ng+o3EN7qXaeQRpT4wnhog1OB60oF9okGMM0v1ZWcZBvVauuuKjChSY6ulmLPPIJ
t/4SOZFk5w0fFSw3LZSi+rMO55POg6Yvn6CYXTTBgvvOLXkMhLA4CHP8+TxwsV9dx1J/YFjwBUyt
x1ISalhCdKKMiA0QRZN6zbWWeYOtp/iLOfhduGtTmyGGR667LdSUngXj5mVeOkOSuUe92VltLJOZ
kP82btU3aa1e6IdwreKlUCrKMhBfwEB7ELkdrprXeYuMY+86qIyEP2hA4yrCD6yIy8yc41QmxnPL
5YoFV38JPNaleE7tklp5+z0KfqwLTCXONXPMglNNdAvp0a3I5jr/mSyGMeNJwCtkapFcNdE+hrfq
44uK74GwZlSA9pGPLmrkrd9+oM33xgDdnVLhlrZClwpV1S8dzIoi7LMgsFy8OsLa1LLtf3/H0A/b
RMt+BgkJ+MtdRT0xZic5QwV1qN/lUDdidjtQNpIEJbmi5Xq3TlNzgF1WhVPUKgsnzOxistDnU9xr
XZDutuBv9rHk5B4TJHQIJ6n/citZoR4m5ZYO6T9ILGVa2QtiNVaRgaV/OYWRK89wuqkGE+NQ8qi+
zOFnK3BBHPz1VP7CI/gUzTbGLS7fcZB1ldMllzdPfZfeOvaYX049MJ/fDy/Jt3aq/K/edqRUKAGk
5UmGn43UIDBYCKkMPoJwEuMUwpEAS+l4DUM2q+XccdDvv9D4IFBI+mymnUo98kdiuq48WeJzJVWe
wOncNRTL4E9ZvCqB1m0dB4kHl1vwubsUmPhpffcHCL1liQAXVi/OX3XdBBLZJ/DAvlhtpfSEpANz
AIKELo7FWq0CZFczhgwyWIjvHlaHOH1rZzJlpgJ74rZzW2kJoTSmB83sY/4jgMuGoFi0NSXjl1hL
SIiptqufk5SYx4gNweAUVILt0bbkohTgYrxfXyxb2WOW4hBUAOJYI+HY2bUgrOryod4/P31h8R2Y
+yPgHYcNkvcx/cYFJV8tQmmNDPgEbYa/1EUp88RfTGU3Mhg/u3ejGSEcX6PV6yQMNNfpC0+xUSQs
VFnLFipQh5VUU8MqhEiW8nsLdLXH7TmFjRLP0T3oSD2NxtPGAsvDFoO8QFKjGGyKBam//7BuaRhw
aMX00jlVZuu+2Brn6zx62o0szDJGwyjJose+Pko8Kped0lYUqBrDuB5kjySPKRnLenwY6YYUuWnU
Z1ZP6ZzNMqEbJ/dSmR1HJ/NyCquasvofWeauXnvgM6zgnJjlM+kUOWBOFv3RhypDPabXI9zwaHcb
YlAtiN4l9PobMa2YACTiAkIdm2XbP3esjS2l8voRa7VbmndsMGW3EgD1HJt9sRmENRZbx+Kfzg92
nK87oDIEzxNbrqOGgduLCNf3BRROhAT+Btjugbf4pyV6rTJLaoEPjPn1PxIkCc8IhRp77RKdFsIG
eeotA3/bIl8rt5VTZY0d2209ajQbsiztzpwBLHc+s5lPoow+rJSaa9hTX1UsjMLj0iymmjSDKwwo
JTw2WYRf/EtZhg4Ohhr425sL95AyNJjj++wvvMGKtpadUQLI35IdGB6JlKBFCQWi2MfG4b7oG1Tm
W8hjJAiGuObdIx5F+UBEl4L+kWyKa48+W+Q6Z/mKypzIlFTaq3xlAxoxCYAiHPr4cBVjqJ8I1BkX
yxre9EZdPRIuKvm8VzzwnAaavtQSMD9mQNEJzAGGk7zrvPaieaI0d1KM88Z9k3jktFAsfsl/Ounl
92UOZh193jqN4Vf5pqE+Vex6dYrkVEb7KMpfvzlJ2/0zDyWhfJ0vl5vYkbXr9rMzVPo5cQ6pvcvT
lvb3dOLwzZGxTou+1dNKBot/GdVKOYChJY17no7Jt5Yr+L49aUl5BIbTm5vwsHxtIlIM6m/817/j
xYrnFxryYO6F33n1xKpKcnpskkPJfQXHfUpwfpbYczN/qLkvdIV2CfGGD69+uzY+olfkHfhinAvD
Wqs3eKKftZPZyovtJigLHV5XlrkUCQ4MNmAXM8cUafTzfYmWi/aoyt27zcTAoxWpV9A7ZCmVYrSH
kTT5lRLA7PitHPLyxcaIMT3gZkV2QlNm0wmLleTsvwAdBlxth1kaeXapP4zhVyMoDKrudLcvwhnn
xnel2vkORbuXeKLcD82athCf8PaugGTqsrem1/P60lI+fRWQVgSSR1yEnIcrxWDhB1ZKRREA9Zot
DoRmvAShvD9c5eTtm0lzdzL7E3PDnUtrv3wOwoowW2Ppglg4tKUM1NYDv9GGXouIH18hxiK/2EMg
78RaJnwmQiY2VGifSmyfowmA0iuKO/Qz5PPpDm58kUeqcXpnDou/7m9wCEpgC6Aqm2+d3AX0wJai
+9r4tSNbTpWL7oCXfzvFizDi6uUryBMFyK2h9XVrtv6uFenrP4Ix6EdKzG+dr9oESPxm1gKkYHF5
R4wc3+Ekl4CJ7RAxG9iDNbxw46ihzTT5wgpsAQGofJLjnornBwYEnYYMCTHZ/kawZibhOi0tTYMP
+SGpYfrga+QLJNU6Fp+iD4td/gHfOMS3fdi5/RcEu6SBW1gNrLhfhIG8k3pfQwVs2jPTYuDgWawl
aRvC7Q7J6Pist9ofnx/NgoiqmqibWUJkxXi95Y8V5QtpDUQ9suSwyxjgOjMHjHMRlXVxJ7e4Fu95
s4tbE3YsEv19JdIuWkdSbKgBqZmee/LWNvplrm/G6lqBum/E6SC7YUSvO383y2nHXZBrqoOmzQmX
mx3dJm3dP5imGwCXNlH7YiM0YRODSegyzzmUI5Pj8diWkIgj55yv0pKm386Q+TwbyCixXTZ0iqzN
pabBGT7M9xsnJ5jTOIb81hlikOpBO1TQkGOSs2isBV/Ye+QxWTB6xTSye5S/BqTZsGAL/mrasw25
amW03YjK94VkSltegMNV75ypL6O0Sem0JyCS+hLeG0+V7aLL0Q604cp2QzSbE9uRDV3o4CsOO0QP
Tpvoru7MQcK3cH8cN5ZqlKCCydzG50FzvdJnPfGsdL4mJ/CPdCSWgkjywfBKW2S9n3E+KkTnKvvJ
n64jAJUrrHqTQskQeZhWh2xyKLL+Nmfh5Oiyf7vmrEdpZL9jxPkhHZnwF/122oydAe86OiGR1YwJ
c7WpQQe/ZKf2hfJ8RYLNqc7Fes193XxHk3ijp+4QdCBcSEkCbkxBFNo5Th+3JUjI8yeKWqCbC6iS
agUNfJ492omA8QO+1sMJE5WpEWii8u/46DUkURKaHwcCtB/V+yPc8EJXGEQK1/mZKmejkgGMOOGx
5eOvKWJV1TgdoKI0O/wNNbNl3zu2T2Xa/29lRouvVwnEy2xWE78m3Er2lumIEidO3I2fjOXbwxvB
G1sIBaRacsd558CQqVZX/0KRSDZ2lzVloEuaLjr12mpwi/SKoJPWdc35AHgnUkDrrqWnXwm8L1JP
fx592kG6d0+tl90947Y0W6qqCFFyf/KzHNP76IPewq15NrUTriYT1MQ86oqo99uGsp9G+NLeWONp
mlFfAL+yCZsHlGgfIgkRB7lAPkDzcNGJoMmK36esf6xSjLA4VslfcMy4Unw+xv2sX1aLBPg9KPr8
t5g1axNqqTuQCrHzJvkFaS1wJs9gucLYypUOkv/yrsxKbeG2hD4xGTreWITFXQLSWK1JBREeo4Y/
VQECjJAuBtxAP1xbCCUAXQLRgipK/PcUpf4KH7eeYrL2RkTrUihx+SpPgX2dGUcApjnF2K0QwKbh
QUAuUdqDFuYUohvwkXeFL4605Fz+1hZ0N8Q0WHqSjZS5kH3geeCGj5APRIYtH0zkPAp5w05Z6Tjf
2W4UZjKnzsqwFmTng0bginrKlPkOpm7VKZQvssusgnmW+mSVXkVCYgb6Ueesdxt/8wFnK6aeox+o
VZFrK7MoGQQ+Ro8J6+sgXApajY6OcVf4sASwjhN45r8cdRuIT3WAT5fbDx3IJ6NZTnaw4wRIrs7t
39ZV5KHEXuhfBQd8A5R/A6yzBcmC0id/P/kDIvhdDYphio/8TXAiJ/3Ic2n7IcPy+HwgXAc9KuSj
na/jjVNs8nqFEYP16N+enc7QPXMoOpw0K+8jUXex+vxseZOi4Gj2gQ0PXJRNhdN72ZmTkVzBTYl4
CubJ18liDxjrsOUCsijhTKPNNxM4H4bDCX5GLYe3mHva9u1d19xW34xm3GgQQNXgdRVT6qrVM7NF
d8cJYVmJQnR67IbRxdMxOlIdW/slhJjR3OS0cFK4oGcG0CKG7NtaWpIqnAXqGdpKiFL8xW8NeHmF
E1v8yUwIaOaLmsiHFuXPSn6YWL/v5Bise/6ss2aTpc1ExE8CsFpvGuPT+7OGNVZKyNLazFfbBKLh
S1ApJZ33/R+8DJ3RU4Pr1HtL6rlv0RDKrLYoJ7vcPlsky1RquoD8Mok06D85teNoDtkXJ51Pbc63
iFz7DwZkdTghJR099zYXHNdzc1l2qoofPivdVVk/0b5LXbMJ8U/mAWTAwkkbgiDXHQ9wuCUd+wKS
8e8UDHjKaakWzbQCJ7Je6Jetditk1tvLAeZLJ4lI326D9IkDX3jru/dCki6E4p6IDoXZoi3Q3ZOh
PyZxG4CjoU8no+dqdimosJa/ban4GRJf/3u9s2p4Ym3AQ7kAAGEK/6pCmkyIcmeHwILKD2FmmNTT
Cf/eJGrd4zi9ZojLmXbeyXISJOsm0H43T/DqTG6KH5C13gZNumysN9C/Xd0swyqsLwyrjGvom3Lx
QwznN4D6A2MwfIsoF5Qon7THaleYarB4+HOUMGhDrQerz01L32fOUUSBxdal7haSiI7iQCYnHh+N
mL2oRs/ZK8682KVGSIpaUruQbXJvRRZ02HF6Y1jHNNc3nGddkDLfD7hcilDhkSWNlDrDKFtlnm32
3ajqqTKGb4izBswYX/CFqAj6WeKslEp+AL8DnOHFoYtdTczTWxBi9gUPIp0WAG+bqg8hQWFzH9el
V+9aMo2hwqn50HS1xhmPep83hL85HR4pUixPi2ITOk9YIfGyWg+MSJO/Xfq3f8jUUAiTixLfUtRp
rZKkNt7a206jy9Reg2dCbi1BxFDs0duaWBWsBSIftlbIGL2wUwyX03v1N0HxD6XR+NrOWAY3m0Hu
wM1l8rvDBCI8cvAWzla4x/GAb1wJ4qR/IOmALYzp02h0aSBAXZXV6/WWtXV8Dr9k87NPyVhBIZMh
yoKLFQa0AAZl+jpjA5VQlJLXtFtpXc2xA4d9PEWeNQbiWqbPkqeSUMPL042r0mKmLz6QoPKjrXCs
6hmN1NWu2/MDczzozIHo1tMV9Uo4hHDuqaGYQd8v50MBfNm6cPysYLNt/NKyI0aJExd+4LkivGjw
DZUWgp3PEOciwDqnepmbofw+LGUjguHiVY5K7yBrAZpJsEmtN9VZWQE3djhZsWHn7hIlARzBtJo2
e14bmQP8kmp/fqKn/+1MBMfNQb0oolbauikKdn2fGhBGViUBKdcZcP2lgx1fu2ACrc2s8SIHRxNP
M0a5SnLcWUZMJ9jbhImX/WlAlsZ5ai1bM998TTN3dbUzchuMq7+GECWZI8giXEdEcAY/srSvFSzA
MxmbOQSoc2UZkatGbmXLTIbnPDqORABozj7Z5Qs2aq6aXAwwNwlACQnnA+rmUW3RPA3waMqbhbDz
EJr3Oe/gmyPqUPL67btxB5aa+YITYGKkDg2a6MO6joe8qRwCfGg4+K+MC5sU3Ps8F/ITtL5bxQZO
DJKN4+Ql/bXsche5c6Wdvzdp0dmcTq3BUOzk45JLfD1HVb8XNj74gaxZZBZOKdfeD7kCKf2wrq+h
IBIyBxBx4yEM6GHGWGbkLPmMjFLUXmne85VS3KhBrRSc+uRneIvvSKIkqjRf/lkFldyL2kO12nl5
K0SsLnux9LqEp5Z+YmaaLUmza4anTS9+ATxMS7odxoW7mLMtVuzHUq9W9FboJsO9qNyQcuKzek6n
TdPlvwEBM/F61xsilYCYcLY0toDC18aHWjkJ6HOwZsAzJ+ou8rUbNrkT8OjsuKCTr+QX37u7Yz8T
yvIuNn7E580hGtNS+Joro1yPZBWfUQPVEVZrbINryEVnJSBjiljT8xHwhsbBe7VCSVRjge53XEBt
mV/D15dydOgFzq8Nu2MxAvvMxFEYGWd3Zh2TbcIA2+gzuYHNPYU3zpAjOSm525Shtha7M+jKMeAJ
cT2M6hTIww9IUD5+kgitzX75oBuy7uurl3T78OlxuhcnJG8bP92d07aRFl1fdjcKPi2osj5KgH3u
Fi2YM5ggI2+lTrwUao0im56/GsGdBCNy0+aiCMPuYv4d6B6mPkczIrO/YUe46nvNYMN3K8JzNLV3
k57FkjnVB4aKEE/7ONVI4LhKR2RzzVWivex0FLUNY7t0RoxyTWLRr0ousriBxXpVo/ZRQg8WZ+Zc
NlvF96x0wF+ytuibAx5cxjiklvrhpSfN41iVOR47xZ+ku7rXcmTzzLS6gwIqYrZVIjarh9+mLALm
dfGhT8S2EbN7rklIdKDYLJJQc9c1lQhrt4HJN4Ctoi5yvynHR4AtoHYcMS6ANlh3WcCxTMro37iF
2V7oxS4ww6N4slZDis0/zcKn921VTcdj4GNay9/FSYDeeVkkpNjEfTcYCPIqL9CA5DkBsq/L37JH
AKX/vmC6zy6qZ4165gP00yMy4sKcP5zv/wb6RUJkW0hNYbTRhr/JtvVpqFX4e9IBCo7GXcNcvrn5
7qnlyuIC7ikhldABeBRZDT5GW0ccWTHDxMAwuBUt7b4BTl6DhS94/8FZB0Tk7fpiqqc1F3LK46ju
dcWiJ3vn5i/B8LblhyNIdQ8nS1BZdC+cAR6ouWhUz21GTthgK0UMZ0E1j57BqqyyhI1+eLWwPpRC
Qt6FXPAj6+iFBWJl0Hh8b2/DtYvfM5i7fkOIFqsw7yw1LQj+aadAr/uxH3F0Rq2pjP9XST3Els0+
aEzlnr8c2xQdO8MPW8DuEmSxZQy/jIGe7cGH13XmU4geq43GhtNXrxqKnxcYPa6duAdpuuacfhvX
09IDIJ6iWzMVov+rWqsp1267NdX8lmSE7FyrJ5Z6WuJ6hMM77zrlGfd2GMev5DhxU+xa4TyPkkq2
uM7eBjo0ab0B5dViPSWNfMlsvDgPYskBC0N5wV162lzTiEZayOTEaS/Vs1iRMabzZL1sJVeA8OOW
Z/kKRXPrNHrNWPFbsZloYEWj0C1hICGE+mtQ/N3iukt4HqQL+QBVCLFE/9H9FBgr2Hf0BL7foBff
GoVL4gPJoOiw2zM/KDHCHOz/BkbWCmhyouQHkNfRXhMslE7/GKKcIohPTkJUDUHSCUp+Rbw3zhtm
yLjFNGJ6h+yK1MziKXgPcNMvHzP8JT9j34+i2eOM/KlORBxbqTwyl4Ly+pbUxycZMM7frlfjLctR
xaseWV1NkN4OBifbhWsZUzStpKRa6SijQA7Wz+jMB2mtAy+rlSXNTE4pA78yUpPOeQ24+s2mHyuJ
r/JLzDx9sxB2IWHcz9PKk2q91olM+SGzhFsmhULu7i3Uuqcmtfv++2+NX1PGznLLFApAdzvPkiXT
rgvWIY1pA869QZAQsHyl932kYqr1XnflhbC4ZpIA9qjYFT5C+qv6mY1BvZTQzBJFww1YoPVlK+XS
Dns5FO9AwSHkLe8gRp9QbhJSf76VTncNHWDiKMvqdhzRYK1RW6AVmREaWPqBzMRyGG+UnLfIAItK
MC20VB3BFIq7NsKKdEhfWdj14+E0WQG9OHVpLhmfWUSC/9QyEs22hDsTwqKVyGBTPuB2hNy5PrvD
hRhGISq9vslK09LeAzXnUP2sYp0OyLo21i75o35KKKvhF4CDIq3P/+xfrZ8/4Uner2x0Ljq/A3yf
HITo3S5Zn9s9jcJ42TfMyw30CSs4yRFNO/V2d6sd2xAlDGRf+r7rLyWSr4XLq7mspGy5WQgCLJwz
RinNzsYwd8WqWgwjKmaOJxsMqhfclb2zUb+UBuNFNESBX5ASHDbxXPto82dxJWWCD7+9qmePy2EW
cyGLoxflvyS6gYl307gMHzss3UAOL+ZX1RcWpT/JRFi0tZi/yCiYGebK5TlwiYz7wTsw9IL/DA/S
Jin6M9bsLkKAm9tZKXdjFLG0/rcwSTcFXcSD4g4HPrTMForhkwua8S3vxclxv9tjp7HDT7rBRdXw
MHbSzfRT64xtvormXeb22I59USjp94pjNuri6U/iveJcJl61ajr/JbDISqZ2WVo1COcc+5zMHIQW
Wo8euGu0l5ojyLnQWZ08wcoSKaBQdgVE+pQSNnYTnDPr4T3j3QjxtnaQt2lYY9B/8MJ8SyvJKoQg
UeZtGzZCVOqIBPDQYZJtUmxLt45IHrc6/U/fTKZYzLNNfwHnj4ifKrx2VhJDst2Fuc+Xjx25WiPe
9OGIZFOOyFyHdnEemRXAa0JsBv1BbdSPv4hosBpe6xjpUAs8PxXkXOtHQATEJ43GifF+ynCrC+jF
JztUMm/ZawrXVbsdjRUKe3CI7wJnInm7QJZ27Ec4oxYjW9RDxN4xHavqy246I4Bq1q7upQjrhn1N
kjqW/GWl7gOQNpAJvu5wuveKTEJKuR9hYnr/JIQSQ2Zwh+uC1BFGXB7DQQIAhjzKF0tqgJOTeotH
gT2if195HmElvRwR7oUxla3rRvUL2WsKBrH+nidGhHzrAjiavvv4zF6BorWGdDtZOD4a14cyW5df
BLmYiaw8L7Jev53ymUMQHu+lkXiN/bGeeQaA1qAuKkkJtmvxEymLASIt45Ht9TgVfANzzA3ufcpe
VYAL0NxPzhaRgnRVWb9Xrp+PL41vJowl6FxZWvSp4rJVgnzxUzCLiSvqxxXNvy3uq3qKjLuDdy2f
bv+QypG87XV1hosE0xml/1Zov2GCsBhNn0WYP1iIX7K4a62e/x3ifG28N0wRWLHRJ/G98bcGWrJZ
jVfw+gqpFTXnCnAJV3sbzYRoyecVzZZDwQtLTMx0vLZ8HlqoNtttoG5Po08ytsc7NN/dERTwKkVi
JchQ5Q9bEkxO9bQ1KYSJ41rwKsnEi/oAIjow3iRCe4NlPhJ0rT5MAf+AmCERr2EvEQVPtPuFO2Ca
Dl883AXYvQ3zXHvEU203NE0C5Y5KowQ3bqpHC+FPOwavlBGgcBnTwJd5zCevWsO4TtCgw2NpIzYl
sEZxpafAajBH/Vwb0kXFJxPz4QACntb0AQdzngZ8J7hoM1siAVoAU6Yu0+CztlQL0X9Yyhug4rd2
lEc1Dc45yVR65BABCT5x+N3MIbY8pJ84Ll7Mt0d9WX9El+FKd/YJFaAokIzKm172IG7cWPMS16hA
XGXpJUnx0xIcCceHccjby8J5JGElJ1C4ThrojHVZ/KPyf3BNiHFRo0XmrdhUODTWV8J6uJpLsRy9
1GRTsIXOfGHVDuijqpu8WTiX2zWLQt/dacQSLxvbpcrMRe2h3TYgEbvt5sRlsCjuZX15Qzi1kl6u
PiIq+gWj3JMC4jLpo0FobUhhF8cBJRhVPUdsQlIHubcqn3uWVbxzSsece/q3sG86veQueNH1ip8L
capjCO5fCDbzZ7AkM3ZnGZoEGF5h5pwwLVm2igzqPedp7yGnENX4XBFVby7hFlUjPN6dRmNYqFSy
AagVPZJZ/+ljMGdjr3WDdYGslzjuLRqRJuS7mW01cfMHFyfNUyOvtLvIWYDrpyYTGrrrRstO8vTM
AAzGmxodD0SuzW1ZckmDxWp5XSacbz2ePRkur0PGnhC5aM7uki0XBF1qGkJh8MqYeNBVw1VMiGNO
irfj4oDgwAZO5CWgrAnmVT6UiiNro7D73fkf2kA9H9umyfBdOseL1ZGj5Ha72VvEZ9VWEtyhxJMH
0HOM+16PDks7mW2rKlZtHzSfz0f92wKmoklMV8NAl3R0x5/qWgmE26yBQ7LQD+DO2GXbagKv4y7G
MObuiMy4+yn6ZVAtlUlmxIOZp+SMSvgvUqMrSvBQkkQpQLDqVMzqarfSsLsNNMYK1JDL8T24YINB
zwutX9dCpdAFoc4oC9os7JI2QJ7I9mzhP/ngnh69LFXNBkTwTccGZprb3WAr6bfn+jKSrcchg5qs
kGZ474tJu6KFMrGA72cC6JbRjAyzSABsxaKFg3brw+UIIWzccXI+NVShtXJHC++0dgs6FzO6bPq6
PIsjThnhKE52+ufpYwW7zrAKrMMdYyjBk9ydjFvoOkbzPV5aFFkJ7Xuj7B/SoYZF5O/dII9udBHi
VfKA5rWMEaGVYlqU1R1Wmdj+0KCXlKLEpuWChbp/Ed2w7I+4S4L+ViDoRbLajJ/7+VweFaasdM8O
STJBaUZhkt1Mo/BViqT3lRVke9upzoa7hNPvhDZIgcsPQ4Vh5FUeL1Gp5bhM8e8GX3RlZrSBuZQr
0onrTBBPdpIuUhXPm0wHXbZAgkBw46ELjHWYA2vRvNMTC5Ot7eAJPtzmLOmGL+aTw80ZjxBwx70B
C47+ssv7owjpB8XqjfGKMeMIyANsR2+DYLaT8jNveai4AC8u3e4GEHvnrq1uTlQ7CSCO/6I3s3fj
aO254MI6jTXJLmkUJiwu9tTOFKM79eKEecWNfyD+kr2k7HYKTq/yCUzcxjPEMbJLTa2ew7jAsHkZ
pLJne64OjW+jJvjPzk3P/naa9b2s2Gv1k5wyKD680oXesyjoS6oHRuYxLDCAGbHG9DlK5pvlFJVA
wmf54b9vxNG+AgHKTYqdV3oQ1lQWCNw7nyscYiUTTZsnSZGEGaNb2GiODP9dCpvdxjuJdPG6yawL
xgHSAhq5Wjunyk6YPFWBpsclomeubq3ll2gdtQwAjTnccqBT8z/7W5xnaU/2gc4fd8tn9lPgbv1j
l7U0vT7LF5eUw+Fir0prjNVkskyK8oAyXaDTBzmiIc8gOMOPFOMX132twItA3EBhTlhs2HZbIp5a
GzVT74sFtsahvFRL4xeUP0uDBFwvELo24CYQpCxMRNNuP+Lfonb0mB2o0V4byM9mQVvuDPrmnwVd
JuweTCjcVXphrvKOtC+XyFULT2+fh0Cng8nCgNAh/SItjsnbIzpQwZAM791cCvs6lixPhp+LdIfW
3DHYQFPnPXrRDMARe9pEl8SMMLgGLwO8tKMR9O8eo79eL4oDcXKmDtX+JthoKU3aQQz6qGAtB8DD
6rOwbwKiTtarnpiA2AE2x7A7p0w/SrkO+hEGnZqV019ryEIxfILmEhWsq8eJ0TB6s7rhbdCCKm0L
jyNTtxiZYulXsSVlT7iM3WHL0lvwGXT1HK4sGe6gVNfFttqhgmeCmfSediEIMLlXWKe54arBTtxZ
kUFzw14U17bJP7lQofd3feNryb0XXUzyuVwXJttAzMrWD/UgQ518pFZYWVmqvsRobjf7n6XqQXzT
bA+ZuoRTOkvU1HTfFoXlqxUCeSvux27EnpoKdNxb8XbtPJkOulMZEjLhkUxQSf6eJUQODFQrKeaQ
/q2WHhNP+ddvjDdIsB0GZs3R2J8x2GwpLSeQ16ahFgaYiCGwjZdFqPnpCXKDEskiw6JXWPxGIy8X
+558BOCiTdQzzluPXNkkm1BNd6Vt7YOpbKXtpr8akKmtXzn0lJqCxI5u63BHq17GJBlVsLO5TFRW
bh+TigQfrSUl9Cl4Sq9WftB42W7mz0IAR7pV85J4KeuERuGhy/Gi8Yuicfjz6u4M4ZfTeG5P5xKv
Ag7xy1qSrCbaMjAP2ZHTfrrrdiSOswnO+HHQwj7LicMLZ24wlYZpcRf4EX0VHyj6O0tsm4TQVGxO
05FrzTp2GG74r24gfdMdSA2EIgEXwT8y6G5oiJ0+2j4yYzVmu+rL8Wf3kooxqvtfCucbSBc0wyzK
DKBh65v2JkaXfa40J+m5/plQq3dHWzu16aODYz+M56U87rrJnhA9/zn/Bee+RPOQ/O2wqoJvv6ro
u1PvgrQTOrwdSa1Dqnr44xxRQQXU6gkG5KU8ztPS46LLyOD9vEDyNBa4IekkhyhkUVHtkOax2qIS
J5I/51JTd6n+KyOobqdxbsstn9dldguhzs8qJfl3fRS+6hzYFGyWAUcXNC4CNazoTmnc+LFTH3/z
7mC8pn+39Cu2Ot1meCRcL3OyuxNKGLKN+eFGkGaISU5FghSpMSd5f2CjP2jzOns9Jqf8Vqi7xmXL
w7Lonvo499DJYey4wSfvplrAfuO0Bu7nIBg2LD5QXuGqzaqque1veRRREnLFN5vfvxmeHGLdHGxL
AOF0tkLrP84rQU/h/i4hAX8wHGWt+kZB4bE7NLav/Msjn60vm3Irz8TWwjuSUDTUNJGGhBBrJ5gL
2F9gmSqxEO5uwN7b5fkl2+XfHVGaUrSeibgBmoyFlaEj6oBKIODNpsCZkp11KCvlgVA7FMCdZGSw
ptqTJIgzoJiz91slCLSPt6o+ZoEt+gLmuMurm4wtvcpzMCz067AuPKYZ4tK5ekH4W6aZq4Bf5zts
+8CjgmJb8Ehu9WUhqD2ZwHksc92aq0jMIfAw/lvTN+fZ0lRCSfEknfcOyJE8r+E4rwHZI0/Z1RDz
SrY5TUFdjPK1emvAXlKxkvx94aUT8iwG4pG/OxBU4OBN+UTy866E/qAx08hwqzHWSGtXgi6OewkU
9ECWfVDqFlqM5osE3CTEzlt0lyzvT902TgY+H1l45FxeZ6XiaIXoxlQiDJYFPgoEcAuw6V6zZVSG
cWkAvONmLo6witARydGiwOgNRifl0FjK240HvrawlFTzc0htKbqhmuBjwem232RKqk1CwkESoD/K
P8LqoKyw94A1Cw1RFrQkH6RLPERcOThTqRXb1+T7nk8QCiRgrAoUvWT4w5Do5Mdn3ufNaL+zdirm
6mHNN/O+B/k2JDx0KcRB4FikEaZHNQJ+GTWOQLrcIAtzwXDDz0oC/zTyiQozywBgd+6CtsuzPjdP
KgXsD5lMS6ZqeEg40OwUAeOKje8+sZvUXBs39QQxDbg6nkJWImfNODPZTb7svNXmFuAHM9yKBQaW
3+1GSGtRKqwIeDam5g/vZKJWl5fmClVxXIg6vvOPxl2odhyeIpp65KE996rPQ88CNKoKz6I0dDWG
YP8NW3fNfjpkxeQgKHSCITAtQZMeVLkwI5DBdlEkk5YmYnmswjQ/hsNWVBliZ5CeuJHArACN00jz
8oPmq4EJUNYxTFlHID0CIQaiQi6uSoYC95d4Q1XZrsh9plkRK9AUURMFRDnlZ882ed/9raet8ARe
2L7iiCMNCgq4rxhKdX22WdAm+r8DWd+qtoaoO3ub8lfZpYV1Tk/DR3feY6mIXbfAj+CSUcamwpXY
7GBzx46dSowUPiw6DiOmV8ifEv7asyi8nI0SXxLLOPnwfkEGVluM0ER+nbQNNzEUL9Tm6GW04dKT
0qK413wlJAcZ+LKZsE9GmrccKJkVL4Thvg6gf7AbIOPYBNejsVPtUJWYlxVseuaI9DvgprotELNV
G2mSQbm/v7rIYX0n08ZHvqFA5ecPHC5ZbZAmDLI/tAjHGvzRg9HN1lZVu4jOqLkmcBIRLqzCaaE3
bnl+IiULVrZLEYWoZqwCpeCTJaMFcAqIOFJK0XdWP6ydrtiP2fR+ohSBZMEzFki/0YsoL/IS+Fu7
GgoDxnGI0QaPKvs9uhPqdpgEO0FE2VwjL/he/D55Sp6KZWg5vbvoCOKv7crgJlhG1WPVwZI8TukB
aR3IcOIJOjRAnFE4sN+mLkH710GzBzKQP8Q5QN5NG0Rwi6S8n6jsO4Iiv/oBlTV70li8OCVDXTf4
yHGdVCYX0HpggaALLYHCJLPAL+Cvuks41C9rugJcSm8teFQqpso954a20NgHH3JHbyRMkogIZA5K
zM//ZplQ9pf2pippUcyM1TOqXGdrvb3kgJa2sCaGVeczNcmUEEKc7koGbNyfsPHuBLJ29vacIghC
IOyrUpqj8hJUkrwubqrqh5I+x7WW2mLynfHeL+DnT5Ms3R+DO0BgCe4fxJNLu1hqlO/+6Rutb2Bi
FxnfvFLs7mCHqf/N/lKxdLsga89Numdsh+2N/Cyd2TqxN2+IkyQQfGcBsVC79KMQyGHHXqKBY/Cg
msP9evL6p3k0iY0RkuZcWyg2pGsCHqO8svBPJi8zfRzPAOOpTnBgwtl15S/nRCzn9ttZGHQc5rkF
7e2otQkNLrP+gfZ2WRqTSKcLSIbO7qwFRZvhAYmc3rkNJXslicCMtnkv6sqwD3J+iQTx04Jh23dg
yRUMS/r9TTq6+j1A/kGDofNuDoIoyFFaRnRLaR+DNeVoCJ218WzGi/K2lNXOkikHodDvCXkkM6PR
CHKSFsAEqu/yeytVtIGAVggFCBNKn5HW0IaqaH2GIhscPHVqFaFimaw1/AA0XKkDG0ANZG4sLrD3
0TpZgw1bI5QE4wHzE1iReTQ1XQbMpGL0aUvpX9oHkleypWVDHMNDe6LDnd2PYuJymvtCQUu+8iSk
YSuYOta7zIJogmvuOJvoUAdalDgeN9bwA6t2C6PcvVQNY0LQM5NSqTio2+WpwvxlM47qCTRI2/2L
3flNFbkW8ybncm+iCFuCUeiPzPKpe9KFM4TJXLZUvvYZsVL4eoguTt3ZvHBKAaPPGuNGhXgOlFnA
vdb4xH7q7JNNIEVaqW+WkO9R+SR5WYL2s65+z+4EB/Z00Q+OYFzX9pR+Y8WtZ+QzYLo2eOGEvOBF
sXkUw7Y9cVdWm57+WJEhQ5SXkh7GFmY1ChsCVqpxHDZ3cpnHo+AHYogKvwS5InkldFsen/2fzoT6
Viq8kbIucvL0LJOosr7u2x7S7H1gfmeXyQa8DqrpvDc9lUVk+wsFJUR3ksmhxMSOu4rHlgR9bQ8/
XiMsFGoKu+Y2NEgU+Cy9JGCtz+rPVVPKWSOEBeia9Nh1zFbgzljJYfdz5ERiXY/lVOgMdhUO3bBQ
hye2LncPOfLOGKMW11ajfEOhWcEDuhE+in7/zvSEy6JnFKk08ykX8AjtTpDaO+4Nmr8imi4JcIbo
b5Z5LpF8VDatbZaLmzvwSg2t315lLY9VgjB55JaHdmowKxginq2HuWxGfcBu253Aqg4iqnIDXdOs
N1SFt+1qjSuzY3ZyvQINC47T/41vJtq6tOirIS3yuJWLx3oPGIrhAS1PaH4Qss9Xid4ALdTo73nt
lekIXPRTjEWtFvlgpPXp5xvSGygkm7gVpk8fyhXk02QHWy31R53Yv1kZ+fX9nf1ZxkKpA4tnVRcG
WUawFLPGVM0pMePE27DhQGYIVXdb9lunGxY9acRGGIRqefeQ2JgkNyjb1GksAaJxhK6OHuGOTqgU
2KjkNpEmd2PRy5Xg87sA2sAY9vAZfVtJ9ZkxnhqE5gORnKaycbQrUH4+Mu1/1ZSxfITZ1J+Uw949
09Qd9Hph2YCfwPc/rR/31nnVWy0ssG/LR4FXI/FlbJs3sNgOz/g9OqBfgb4ZECIzKl9FOnb74C5x
Vi9eSsnoDobNNU7w+6LtGJIxxjpHAj71MAEXAo80vaM112zqGIuo9tGn4XUTt9kkvXh5ZV4bUUar
4CmyU1ndEljL9jW34Aj5FScS70d+VXM0AXclKvbNt/ajwIZ3eTuyQ5qQ+3ij3gaHw4w2qMsXAr/f
CZh4eHAX5kmzKIxOvafkGJCqmB1AzokBW0Vhxs5uX7LdHj1oQWXKTwlMtABptuMv4f59UbrdnqzC
wn502F39jjTQ4J0Jt21HTZsH3xh53MSzKscwH3m6zlWkhCH+X+jC2iaqjM0OSRFUVmVAKSoivvu5
yQSrguFY2jVxF5Bbnx396+IAZwwzNr3TBT6XcsHgWvwdYUnv9K/tq0dJYatrhY2UuszKS3YFC1WY
D2H74eyjGd6OBgBKicgMgsp1I0aw6OrYaHkus0VLHLFP0frVH37Ly/N9l8UpJtPLEwG0bNk0Yxx+
b0iCTdK4OQ9k2HkCvf/5WGPGqrcFhQPthj0CiCEiGcp/jjOGUUSHO2BlUvSrL9HDwWzRVCx4fx4u
mtuXgudi5dV5OwMPBUFHedSh4nhSyN3lyKqaGUiJFu0S43rGz42/YGqWdfdhQTjgQdTONRixuXFN
dqZ8jeQjPVYbxdIt+KHcewNswymT02yfQMEL26KTzsYPM7OxMMqnEiOvaur/ABiM4Z0YX1aVfAxe
DOGOMeRJvvbuQI7cdgHkQDQ22/lLEwNdMa9+EbBALgQ/RWsqrRmCrrM9/GF4NCml2ANB/1xriJlv
HrgNddWjYM4ODtAH1fWymkWVbqX2XmnqkoemNYc2GAOWkph0Ve/e6LyDLhtnBAkU51ZaaTR2Rfar
UvFdMVKnMsLfZdR4hPImxH7C5pElp0tarXckrjiD+T4iQt7hY1n20XBTmkylQoX7MyhfzzYSFyLl
3DgfQhuptl6UFpi2IihsOpP1l+TGzrlXilWCTdduDFOqVGesEwySCosd5gv9/0MIvEXXEwr4irjJ
4/gPpr8OMDZo/z32V92AXAYXt+KPHklyuIde+8G0jt+kr4+/Ke9MPlhT/I2VW5UFK44GRKH3BvKU
5OZJMjOk/5hVnaHvCCkEZYjtXLXYBb/K9bAj9JUal6aeqAyThvwK7HTPkcIUKShG6dCFxTLn4i8l
MxRYFhIc4SG8Y6oEKK01eCoRkRx07a1GU0kUXm2MASTjcrlPZNOAzCBF5kOanYAPe1uYwxMjfHx/
baN44bNLkEMbX6nFRkUy8BJ0s+dpgj/q/XL3BpGHt9n5sE52ezGbmnt+m12OusbCicgH5HeXjoqR
4/u5TRqgTYaUwXpk58W87I1LUvy+PW8Xk2BWtSckNzNqqQB5sUoOTZ99ih9HtxhqO1mPgbJ4MPcL
X1+0xCZyc3H9ji9JgOWE4F+eSpjwSWfjlRuJo+Dlv3AKT3iv4N8x7bnsp1c342sU3nvU5JngR8BW
LB+dsTYoSuYm0EG2KraumnwqcaPUhH4pPzTcGKtWzHEDWNbfJG65ZmeL+25skhV//QThyBzcvAea
MPqLsqUgzpy7E5FqbkxN1HVQU9zdhYwiPowLYq4dn3wRv8IZ5UnK7dGPsxiyazS2JUM27cFW/LgC
X9QvGI+DJw6qVgk6gi+RE6RyL78VQD6jBgT2s1c23Ju5G946n4hMZNHyQJd9NyyR9wlpkRaYIx/a
gJ7fIaimLbA8QYyYD8V4tAprKuLkIW+zjXtRN9V4GF7FfzOQ1cvBpPQzuadFu64Ly5cP4EE4tBd3
KDuU9cW0aig1hHcKHs745u4Z4DQs7NHBc+h2bGqJlvUr/gavp6wntALDH2VcDVNkJQbiAWBg5Nih
j6cQhNa7bplJnkjjQiULjgOe7MyNAuNxnVvaQEYpSIqWZ3pU+pZdNajXt3jyfVztB5oz6GFqPupR
pAGkVAW1ZRI+3u8LYUTgUxz82LTTaNtp5umL3S4epWV0lj2TvcjW9MdiK9S9Qs+w55qSAsJWEtLa
xzC5iF7b++7N72XLgmqo67dI310OtkyddmXYkAHn6+k+Yx/rl1VmflzavaQURslbZU2gXUpCpMo6
uV0mOOY6+ZFkxJRSPfHAGI1KNgN8QydddXuaSoHQw4hixxHpmE76SeRiFmmEiU7uhU31UT0+yBCt
TzSRJekdQM4UKgCmcgYDfDZVLfMJIcd0XVg6hMC0yei/GZKl5jaKPbtsO+9U+LzD0CLv1v4zvuoq
CYJrKJb0gwInJxdgldLl+RwY3TttUJYt4BAXIBQVE8/uNvcROrc6BjUFGobpT2S7Ad6XStJwhQet
UHZ65MA6tp6f4TOKnIkmHgGEtqMPK+zQrw/ca9996ZHu4/oWyE6Jbb/xVrMjecuCIW1uI++mWmlM
D/AIMQr05EQ5LSH4lwMB2rPC0iL6l9VesXua/+Dx4KoGe7wM4UXwiwGL3avkyqZEBy4Y4kmEuFn+
6r//w5jEWlbEiZtp6vqDk/Kd9tNORn5vWGMUSb2N3cDZ84YZXWFf32MAOfWNylJuOun+kjq1/uKx
snvVHnDuNC6UI2FrqLfB5xyAIcGC3KRgKg2LWL98TUPwnGEdFjMzc1frxYBhyPIcZfMs0OP/yfNP
p02B6CfSBSnOnRmxcv3vZCSbhW8qeB14jBIq8T1AJ1iSLDDfZkDv4QGIUllDCL9SPC9RmkhzsLa+
1QKTXHZ1sEkCePKxW7I63ae1Az6hYj/IkMVzB7ER5sm4OhQA4wxKvmPhKFb6yZJF2yoxjhJgkYGX
vJIpbXubVh1wWVwgSL7Pd9EuO6o/6otNlr4O8k3BMPRtQmtBxt9ofQWQyHXtXlboKo+T7hTba1nO
DtiM5Dbhb2rXJAgnqGzHaVFVTOf88yNGBGH9EaFKXYB5Q9a9dNSnVaa2ycKFUlobiUJb11tGWFC8
lIGiahnb0ljZVSiNwI8+uEl8yFc9DfnuRHbBov5iCEihC5ueCgf4qM0guy6qJNILs6fPh4OvUyY+
zGxus3PvsVMXkqtYyhUeb/1RuCe2R6N8aIkJS+fnbMh86aezFEy6+bidUKYwc8JZNpaH9kBC+ztw
bgjgsNAmlsgPgfbEWCv+6Jjh+gR7v1D2RAe5ygJzVpV+SnEKWcrkbRyzxkvMWJlYRZYDE4btO5Ez
kaFLZxz5A02lE+trRjzy2AxtVOjKgIBiEgtITcISUgb/N75pxaMBefPB1zAtXZbcFAcDIX9Z9h/Z
hPRYEOobKOIZe8OotnmhJD6NLLKqecBlnW0Pnl6iJAqU+jz6oKy5kPEGSCXJ/98RdKBrbq1EJbhi
cnWcE6rZXlub6hzFTC1dNshwlPo4odPiMbadfBkn5oOM+A9mpOyeI1tBoKVLl1lLlKuHu2hL2S4k
ZY3IM+O5+55gCdleu0BQOs2Hs1xFQCkFU9V5zcWS3hRicnNn6zqxqyThkr/Zd9+VEm1JtS/qP7N/
fMcE99hGm6oQO+7MqLIbwC+iBhBtl6rBLgEo9QsqM9X++9+NNGUOa5rQ3r6QPv82AOZVer/qgMDI
GGNNNFMET5pUtbEFKykUhXDUxS9cm3OQ06ih3hCUZodsGM29x2S/6KUnJL9SjFM+pbNLUW/HR+Bv
btUl2FNMh9uGOiSaL4DKHfwaF1z03iX1ftQElOrpdaXb0g7Ixj1UVNOkyBYMMVgUeRUHAuD/Mxdh
8uhE9sJD2vcWXPqMTB49UkcIYOl0Krx9SSaes7hdusj9ICuZCCzVZn6YJlvZeCV45CVF6TmzFoen
hgLYA8hsqmUrlbJ4wK1+95O1QYxNsl1zTV046e8+zpoPyFhB2PhvPZ86bxjUaSJlbQOTzcszB5Vq
gSWgYYfOLTO5hJLL0swjET7sLyhSSJct29+rnTr4ZefG0YvQzSWMmEWFbXQ/3ssr6Fuzvv6lHYIW
QNt4uFXfMDYDuUHtQYIWuOyOHWY4TwK8LscvucihlEwFff3MVUUi6cGxg1d9Uhl8CQLT7G6EoC2F
P3sMhvKxJt3HFy59lyaDc4odW0vaMhcl6X9ONo4iOzERxxVvgBe5jwlsggFWLJvY8N4XwnH1CQAh
zUVf7qvTgqxWKmjqqbW+kjZe6W0JQSBDnGGYoCtxioMseK7NxSqmWv7D6pAcQSt9/KPd7s6Xhlm0
7sYdToxgvnoDOsn8kWZXlIqF2PMGLM8z9ltFndO6/gbMyLp/vR+eKM3Naz8x8nfXj5H1wwLTGpgI
n/9H8eG4e+Sb8w7QtgmwLRdbD9EjHFJG7eQ1amdgQvdCCG8ytLN+DH5/9rGrdhZTCwUAUaNhqCVe
kX+q9NVK6Ku9s5mebU6GEkq+GBVRu4kb3TmTjsQO5r9469pmSnMvmUVt1++QwFk/NdEbEDi/gCK3
J7zJXVxTGrYimJ5wHijdqiH93A5slacWdDA9D/NSe5RhwFIKoehN5dPDJCi+6ByaxdIX2LpsE/tR
X1/E3D1l6kMFPUunkNPcvMfrj9W+osbkujGgddXxCL4hl+8I1nW0I8/opGGL1zA9/0ZXirJHJdTY
Tvv3hfBy4tW9dlZ1uOYGlzsEEnuMM+HAzFXHeTtK7Z4eQAMiCtuqj5yqzs/sKk2HQ/alKBwPMqJI
uchtgAfHUsZ3VMubb9lo/Tw6mJqrxK70WCMwOilnKKxyIldvNh3HQG8JPWRRLIfEExV7Qb5kjjIx
nqHq/VCF7NxCDCKDwPwKaLtRRtIrTgecu0isrUFNVfC0+2XCNssrkQscXbyYQoWkMH9P/OX8zIEj
CSSkeXpWh5UmcddD+yWdRXbYDI4+/F7HQ255ajMEYnNAPboKSHKmMxCuuxH5pDqtQAcJmI6eUaJs
O17uOpHRQ76bybdqplOjzUB0Yd4amhj3N5z6UH6kZeInscRUF8lQpNgUnaWXPw+94K0f2K7CUR27
I2vBihzOHCaKSFafxbJjYdfe6EFHEBc27bnGSnuD7o93xlhyuixzvO+vf9Kn3fgqRdmRl2DVCNvQ
kdn+S5ZlKorBLp3FdHFvJrjN+5x6Jsv7bSJH/xWns64O68T/cHcp6+RskJipmb2Wd9s7qBo26RpF
KcNZyUzQsvg7EacU0V99bgO8EIw8TlT43O5i5DAxnIdfOaLoNC9tP/4xGfKho5Owjeob7Rq3ktTv
Jdm466a3XbpHoAPPU7cTo/Eb0vcTesVySf29KZnftVGloWAw/AqNlTQPK8k+1Qj/8vbOopmkrenI
qNnkWC6kkPWg6QKSPCqpkWEtTH+zLavdgjG4ijud0hs02mbmgyKOZRuOS20+koeHY0rHk4g3gZpm
YDXXTHkMIPzGCbOkDzmTG+hTv0/MZwKIeMSxPN61zZDu83H+s16e2wTjQ06ipYdm8TwPoDcdOvv/
S8FeqSMKN+GiaC4ol5cIvw/Gcu2pL0bITbumdDyrT/1dvPxhpq5pVw84JaGQn2LQYVoIQIQ8JKfC
3pKfnEWm6VbOWH3Lp2vt60sQbWP1LN81rmn7A7Gvs+maB2nx9ttsJ4hq/sxFoOQfpFQEyLGDe4Az
WFVUhjh3YNel7XD1s/mmRmXhdJTXSuLsZT1AmuvMr8tDWBEZ583YLs7WYM7oxSDI3RqBXfCHlNBO
qRawJyHmmT6WclIWZV9qi0feig7aQ98OVPhdWfgEheLrnoBIfNDKi6hovZ/SRBJ+gw01Ui/GR11c
VhGJ6GN5Xbk5nKUMajWtL3GgVupNHwWWabnHDKosYEI+PvcbudkRA76CgYJscXZD1MYwaHmm+bD8
3PGTxpybw1gzWVcd9O5/T+apqd/UtqijovnT3jkhMJNbgn4mJYDieea75cf5UTvWFkqHK9hW4nFt
Hk4JMEjEAcXrLJ5diIIDX2TH1p/9B5IFaViIZnME/ariLd+HjfGzaC6XRcBV0nDhHaGy1E2sbthT
TTaqXdeFDFQ0Fm3KBYmXOqFdzj6L/GxDgqanM9toUbUJMbFm1vXEoe6kHne7q9Pwf0nDOz6wiYpi
3qZ/nzCNB8v0E0wIphrbeGEvmKNoJtDTIL6GH9dAnHZOZ/pbyxdu1Xm1mu1r+cH7IHq5WnDBeZ6f
TgUKAIEhJH8W6oi9doOveL86hOc14k1hcHzZZtsmF5L7Ryjio8aKlFiMjZm12ZebBZPxmjjugjO3
lsBlHDc+9+Cwbw0KS91RksxkY/RK8rxCp7NZN7YxrddPW5EbaQLISqg6OeSqzSIt6FNaCjjL1Et2
OAriY7UcbL7jyhZlfNvDheMv8Rl72mDhKVO1lVch23XPLNaXwFDMQpTgC0T8JWzaXlD1liGy0Fe/
0olU7TaWMMmT7TsKUlm20L9xcD4Je95C0aI9ihjfm+PsQVLctyEN6nhVxxA2Rw3o6SxAwMzU33uQ
ZbrujbbHvWl3u9TVCC61yrSawya6NkyP0jPxsPAjG/rW/bFp1+tfNYy4UzMICE8yo/vtlj1eS1j5
ZftOQFnhjypMjFAuzP/vIQl33STbUK3iBw3Qpig6408ur2cL5FT1WVhSPn8lbP+pgR8hJmUC+cPZ
BVfxME45GpDLrlg00DLgT7MWysog8auEZmRaSnqpG+4EpdLuzPsB0v0JHT4x4qSeSak96gPtXxx7
b7KazJlhs2kkEsqNiVYj1zpp2BlVreg8P5OUGEtAkAmZlOaH0KepkOoP8DVXwnskZsvb0d7yL9CO
S27aQx0Uq/9e5k7xTW/Z4LSxZ7qHnfvlz4flFS9J7aVCBzQq+eCV+oXRQTYLlUI4Z4FlgBeCLpyp
ltzE+ESfJLIZ5hLu6WlwBTGMHuWSG4NE0C+XTKPVneO5+NaR2GTGpYFtYDByZ0Y3WK+e3znTc5l2
/7Zr5F62zrkv08lIIN+ZSOtR5VixDV+vDP91ma+hrs0p1e2IDEHk/nC5WvoEmxw/mPSdLmW0LvfD
mJZKXKbiEDH11j3021yd5Y5EMA/gnYgMRZ1ZnhqHD6mEuJRVxb9Gbxs0ZYq1e4wOFcsr1lOHoVAJ
krG7I3xGm1Mi/A7LF+EEr5cGQsvxWEATUCoH5RXdkKvWHcZWvDohfHo9Wkken3YSMS2ijFyolj5/
gINM1xYD/9sUcKI9xXWEv6aoizwzKL0JoVDjhYfG5Wc029cIgDlZdsngQrEzxMThhVBAmF/9O/t5
Yjcr2E9ReUe8o5rB8rigMUsF8Mk+iY6emgDnwUWZRbQedPaMGMFMBM1C0pTJ+cQbZcmLSatIR0rO
2yxnr6vNrCkA7yodoMSk7CdW7Go0Qb5hgtXsouRVwNygQ4wJqceB7H1t5GcToUK+ETmryX+Skeba
PRcPgX8CXTFskkK2bFvKa1GgrPTBABzV9JDss6kZyWAookEKPw8x+8aPuT1bpsQ8hxpzT+Vmbv1b
SvSsBLtSTpgikPJOeLbMWnVwtIHi0xcUG8c3u5doPDkbOoZ/sK123itnJDjvKnPJJ0i7KKLlr5/Y
SFVBoFMr9LWQ0GgYptNwRFD4cFxbiXh4DaxSnxtHZqWVDKlT/mAz1HlH16WuC5dBYn080Wy1itS3
jvQlk6tC8h4nO7tcQIDNY6CEH6VbIgjUdEyV947/Rfv4r5/AaHMyayYKtp45k2VraFsfSY/q8vuG
NMiY8WyhJQo+qaXrYgGcQIJCJG+5DRO+Ysf+frcnY5Y7QH/6Ks1VWzdOl9tjfJ2Bf7cMfhnssryf
s0uTQPvFADGPhbADX6VwYaCpTzidk6IQAMWMwD4Q22M+2xqIqnEtYmMjjEqfFfBYifwmx9hrYqsi
Y4cKNKfJJsEOHcaZed+F7pGtp1Z0Q96Q94RpZRDfVfrIcQUy0FemTC/hERf5LqQRZeuAM/9cuuIg
a+cLGP7pLeaYx5QuKy0rJtXWIuBqllNs8CwDw/myQTq7GtWLkruWgT0a8FdJ1IFQQhsbUqQgTLNZ
DVjuNwS1b7pUheoby3uhpzuzYLu+Pj+5kpSQ0GQJREvYEN4rkExcXQD+Q2iRNLJOFLgLcHY0cLxY
oAuMfeWfP3iHQMNffqt1LXkQIeviB3iWEFcRAV4sRsM1bhKH7jRkABEbwsdje+1e35K3R/xIn86z
g/iCRT67jAFabR0yo45vDISfX+fFdYcyyR+7qvsTRM0SH9OT7r+sYQIhUonVTw6RFs4Sm8Ha5Sm9
tRYW5cGP229J70ZlNxEQlAROmS4VVWWChwVGLpVNgn8ersepPT/RNSxOlSUpi4kmUiaSQIhCSFq6
rNb2jrZezHuCd1dL3H9WHBjrjmiZcl5UPQSKlaHjCx2I5k1QxRxCMLhgZo4YwWA3EHq9CbJK0xGt
BhwUMXY6EweUTiIKdGZM7nnVRABE71q0M8la1WmKOEKn5F//CKczuB8qbGYj2xRRBx94OF2b8sJX
s1y4/OW5mtbmxNXTdMxH866L46eQ5w3cidJymgrhbo/J5XIkLO49ztsE5l9ux9juAkvW0meSZdeW
b7P/0L+7PNU/F4aYVqlfz3RoZOMsbW+L0U7Qs/fxVo4OttIn25vQNnx7J6swPHy+ZEwJjuKghwgP
0MKNDmi37X9TyAYG5I83jh3XNSh82DIOm2AL8mTKsUzjrGO+I/ylv5t3M2Ofv7K7Dzack581N51H
Hsv960O5lWGqAt/rvNTZTcupeJnP3KMPFQT+PesJwE0s5Ey5sjA4TLvMhXrsL0wOvtRgJCX6QrvF
4xrgfs/HqvHKEzS+V0s/sQj9Sbn2sEC1IM5bkdVD+yIgSjMR/OiL7qxWX98UYLqALWMgoLH7rfUx
qrx+qzQ7ZPPE/w++Hgi+KwmsNAdgaTq2YB9xstJg1lNvQFQQ28UTMg16HrFTqISFoelkd+5eLHX2
mC+t4VJsVEM8+JOu/O3SZPBX6413iW7vDTeHhAp+8TMEcgnn0YoWAwRd0gtk86S5lwHgWfPakStB
rKiRIe9pZ8D5YQkSUreyVIQG+Kb4C2ATdx1ZrUEZbfdIw/xX3WPIPn6w7lGqdSz8rdjVVIE9XmWC
QIYWtcLnB5Xvp4QwDGYKbA6Xe2QvVP9RrNfDJSra5bOdMF4fkqLwW3/ngEvI7UmnJxvxXA7194Ih
0kgEATNZ1f+1Ne+bZyO2SxIPbs6OFKAZbW1g2ssFEuto3ADoSdac1/Hhk58eBNcGYRP6pfkQ/Sub
66UVum9k0+GTjX6/9VBtat+NRJwgrZkB8QGqiiy5uz3PGszVgCC9BBVIm3pcweIAYQ52/g0ffYrk
bDHYE4Fwrww/cZOa5oKMl9FHb/QVvA5vjvDVOt7zHcOWquUVg1H9+rOUOYjEl+O9oZxvNqV96pYF
1TkzWXLVltusbQF4HfH+MCaiEtt4Zi9lm3f5GmaPI8qOx/Pvs2Yk4oAJfk2DjA2uF2oo1RmwQ9Y3
Pedg5hV3ieAKTuOfwcnHprrRnHbqbeDE+w0V/ISqiNbLxwmUa+cAUpAIkTLfr/Sv/gIeULL8/GkI
pL6IzhmhbVHrYlRkDUGedMoB0OeC3XmgZUFCYJl6/B2JTGpSwq3a7GcjxZcSC6p0FFI9SicgLBOs
+3Oq7W+0f6XIjcaha3Y8J5Ju30YpY2BXLLrCkeA/j3taFDLr5Hh3BLnQy6PL+lbrdS4mu7kdDYZB
4fFFJTlMSK5znzmA2GCZ94moCWi+hCWbf7gjmWACrKeBDzfBfvjNBPSVCp2IBzbwc29mM3LhsR4v
cPi43hWaZZ1ZkbTWMdO8QIHO5ewDwZWmBrbF1keuNHfssjnTGOdF+sr0qJ+hrgPaYx0HFArQSTKc
1ogEmqDFCfI6L9VtRJdkd0TOTbL1ps0VJUwsnMzHD1s+H1XFXGysGjTdqQXHmutcgv/U8/K2djl1
gJRHau6NSGMSay+nfl7BER25Kl/Mvj5RE89leNz2503jHj+LpPAg4s+ESRILbXdg5pSMc+RD0bTG
Nd/UKxBfnN10EKIsvfKhurPNpeNuQKo/PfhBu3T0OCJxy4BCmvcmQFqw7TCueJ6VofqepLpMB4aT
ieHV6jT0mvT00lGGEg9RNfIsao6AfDjUrmJwaIdQMdcOQLvE5s4iMMG2zlEaoXkAPS96ccZqz85a
/bXWwdrpehmG6P8rbFXcwA2wNenOBqvA0bPRoVJi1qXK06rGYdQN0Us6aqewDL2AzKwS/rGh9Wdc
g69f7bOS5bo8frt55+V/unY0BBKxaDk0Nn2dhZCPQmOSXZF/+k2oQeu7GY38DlFrhISN/wrRvixa
vvwj8z5IFvkIKfiWroL7U+3uKV6Ul4OpQ2eeCb75BgfCXAfsg2QfgPiJmwgxisYpsCXEqidU9xkI
Lq3K5ianQVSPKXJGDklsboL0wJwSgUJ1pX1cBIdGgGF/jAYxXyLKPDaQuOPzvuzEWsHum40PMe4a
zKlnB5XHkQZE6+HnBAi2WwS2WzZh5g1ID8NNfQHLOQMalulErl+pcBq89+u/8VbpJ/Oe+0UbgDjy
Yq0JkAO1ieKQzAjWl+Bac/TwMmZw4JbfyxcUN2gC/hvc+L0fT5GD2NT1PmnHQa5RBnpMFb0rgWFT
EWWn74q3CGBb7lYv8X5Oa3t3krzkq322sz7MruRg3Mbz5/s6TiATDOTMS+HqToiHsV437mSKpLC4
kMKVMQMziK8fwAyP87PpGkhNbT3HP3Bzw9t/xk1E9sj94Ixag4exs1kVTSngYgjES9nUvDG3ANnS
FkJRbIe59D670lLdBWYDLYYt51pdEQrzfA+KyURkknestnppinyS8dQ3rSFaonJ//rdQjaMRFznF
UHXFbAZZkpFu4qzrRo4TU9OUXDCQtvDTM2jWmJrTg1DGWA4iUGtoC8Z+84YeFOszE0M1YvSuv9r5
A6lsBkjnlWId/km42NGn45DAg+05OIpq7e6C9/NzoquDNdPy81g6vc0hBBcPgXyL53+PCRaRf82V
vGNk6jBOVlTdA/qSdXIDg38UUpsbEAdivHMOAR1K+aw4u41bMWJsWdtoaTwVUCFtjfKl57RE9/6O
8K+IdFBMXytV+d9zG2XzLghcwETJCTcJQguU9oMfFHZsYiDuo/ABQRNiSn3V5U10GP/LRSrsvRHa
kbPFzVDXLoEXPzV+CrS67fBps0xt4mdDGQO0vDzUS36WBBdAh2mShNg9xc8+ByBB2f6sDvFRScwV
J4j4omMFXX1kNOEVKoCLlWXYbS4+wYI88Dv8exDSbXzhF/5X8RBaXUClG89z/+nvG4OCa8a7F6xx
RJMQo9a/CwyT1mB4K8fQGHxJZZvbJg9KHJC/qrP7g26YoRZKQ2CuRZvrOhCXoghoI5rW5GTH00A1
IaC6O21/uCdSo6HgGzFgJCaIO4TL493XTDMTCH7z1gFlB5VK1VZch8mwBOBE6INM1vqf+Gp4s1iY
ce2wP9xqGyTel/a6/Fgsoh3kOaKtTwhldN6u5M6AgrtelhXvpoyBOgkLre0R4BW8jlfTB86lJgVN
SIhGwHDrBOAu4tLVr8Am9LNBU+jxp99qewTO5Y1MtRlCKwkLArZeWPwFl0f9DzEi5ImG38QOnSsR
IQnZYy2fA3rcobC0KByI7iqg/v1eEIiPh5k+S/yCz5et/gw9Q/OVfswSL7ofA4gTaZ14NSOhJLma
Fo4aDbev4KbAkIFvywqYdP3fgKEAF727CJMyyVaTDYRqnVobL4hCssbE59uuKAlV2lgjWri8wdlr
kD3JXWiWD+o9ugV4S5I2nCv8hseJzRRxGntFCTwLYy1bglmtMETBP0uXaCveOMSBaOqRmlPCXiu8
vi6XGwK3PZz8pCnTY3PIr3/CQ3Z5hZHdgJarpzil95DpQJ51HussjnnSZbpk4Bn53laq4QLbq9Wu
OroQGqyhIoVOFswaibDmP1P+ftOBNRrEOE4WD2Rb8Cei/sbtbiE6dQ8ECbR4Tb4Um9h+ZnTFNtML
Be50vVSNnXmI1rGypEq+MeTAFQ9vAeOH6Zjy6ntzX5WP+jq3qnqugwTO8wy+K/WHaPWXrn3OAw3d
ojKPEVz5vgNW00amVT1rb1bf7cuEl2J7G1pO9DCqAYAbKrDvpIHoagNrvVx/Uk9Cx2vDvRuHG03/
gzD4BqOAwSMe8YaTjhCFKmMPachEjRJ5pu/4zqNt4ohZcfdTKVrIBQXExf4qjFaNqBVnLyt8xcQd
bnMSjzgtf/01fH2leam594sr2N4DQp/BKqgkhwdfhM6cVCBvxI/BTNy6p9YFeNDO6lLUL0SfCc+i
tJxVSh8bDG60Ad0yxd/FNErB7LhKRxN4MLwU9LQQYRCKvDOcMKb/qavLD/AhtB5G7Wcbjz9Fhhtf
02VFrwV1u56Em38tCW8JHpxUia/kEigiw29Zgi+ldaNQuGrTBwVXEJl6p88gbDLea98TZaDlzy9j
utSDmvFNQijJma+h4WdDs8OZviGH4ziKVQYJ0+34TF85ipbtapHdnVC342JgXeHtGHvCosApyHAN
Y7KP7P/gDg1MiAP4WUYEsuEHXAWs4gWbY+IdMLY+v5VnHSTEPXrgR1g1QTFY+sMUsoF8HlNwzFpo
bDkP0v9tlMpK7NlrT8eqNvHI9FJ3f6dF6ePMdsCOh9jA6OPheTeDbM/t+z2YlVbz4LKayrJLbsi4
PDySFIesiEz52H1EHg2xQpGT7qZ46YLzyDBGNgZNo/BbvpSgq1Evg1bXxDsksfO98rIrrEnqs2Nl
kLsXZY3E9x45Zz4hlZ3knXpFpsSDee8s50vCsvgK8p5oO997tNAiJhmR6BNfW9iBAfvLBWHhz5b9
RZWh/bzxixMV9NShAGc7pVwot8VgU8XWxIpbYlDbrOlmM9OR6uji0473dpDdjbm8nHB9sF+rVjUg
6eHN4qAN0A/0/EFmancLdwRa5ei22EHW8PkP4fSXiiNBw82XLf/sRxYLRe870LOKTfG7HLyJTnPl
IBo5Q0uS1FzlW/X4T6KUtpjVQPqIj8Kepz1U5nov5ZP8kTBMGS428U4/nfMW6aqiV2W0ie8U3hzV
bcnQbns0YaA/Ii+hfB/iFlbcXMjwPPdNyaGx6d9xYCzK0emYb0GpFJLmnUivrsJuRr/EhP06mjc+
+p+tY7/XlmmDCLXRvrF7FcrnYNDJrSjyHBxw7gPnZkKGQDJEK+x2katVHh/Y578VD2AnwigmZp5d
DV/mmE9I0eURsCVQwvKRU1JUTd0Bjm/E4C8elP8+e4WyD5Tt5GVA3QrqU4mX0YuiVaYAyQFyHOCj
v/zYJ7kWcrNbdt8K8rXCS9pCrx/j/KMeaN+0NGM3Gs6hg8TLTtkCYOwXhbyF6Dmho8BM7KoHKl8A
ILSfU3vRe+KyNHdRfEtdQo2fLZgSSPLG4mpvzalzz3T6jyEshjjJGUgoB7pavzZF8MKz3XCfInav
WGBl5f5iFDB5seGrIw+xhrg2EnZXHWWxvI2nKvxnKRVtat/TL6MySyB124YeDlXVkaVC/1OzpbMh
NVijY9mIoiq/Y3iK23nJ7gz66m0VPKdw3t/Ue8V1P1tQqdd0gPhgkUh7mihVzdEnqfuubdzuOhCU
HmiVteppHs+I5HnQZzNkdKMLF3vXMRXbXqlcuYlcmFJ2Vfzd0OlMs8+oIKpNpb2OnRB8tfvA6i4B
VNACWYGYzTX3Mu71eua5Xy7YoxSjmGcjZe4f2S0dBECpomOs9ra+kt1xTXpZI8gbueAmFTWkg7Oz
cx6dLfB59W/k3V0afRd+zYKDlMdntSRZBqYh3r4ffybO0CIp6uoCY0uw0q2HhfGeFQtnSQmt7n6n
6QoHPLnheB7/D8dfYxVKpRA7xdkPnxBzL/Ul40aNc1tkJQuESLkcJvaz6d1yqhyqIDH+MUoIZp6V
EoPKJzdH31R3LD/WgypsSXEMWv7Xs5Pz/z1HzzUuX+La8HDXF/OeAYUCvZcidR2WSvBVYo7aje3m
ByiEvgSoSei54mFm+/SyvuCVGReRoZnGld603EA2vZpuhLUAJUwKvjHsskpVZksvEkVj05hWVBbN
Km8RT3cjO6iolj8jnzR08p8hC8I3UgB05hziQwvT93FQAs4wT2CkUBnN3CY8Rz9ppSspAXsTN4iP
1/IzkAx9z9G/GS0u77Hgusb7ouBmIr2ZAFZe5wSCblIDJEscWvpcMzevUlEi8gjpG8bp1RM3bnaf
ZUOVg6qbDhpPLMVF+lnOO66biFlKPRW1aFKawo0gQyls1OJIT8gcqE6rlVkEKr7HSAt3apUWqsp7
1ly48KrQPZqSiZF8SaiYcDTVqziraJJTRAHDeNVeIs1AmxBzLRaxUR8DU5mJjlwa4nSME0QhS9yy
ov2opsR2ZCnVFXEglbis1KON39EUp9WCviOcHspH+lw3IAH8XqRPT0gx9mK2DaHDu0AYttcMdZVa
hLxNPVhPPuGmIvX0jgFSzskVVB8C/thN3puRRxRY3+fHymPgXFsPp2QUgCA9U6sYeJzGopV6ph9h
RgGcbADuqd8NA6xglRlGcnOX+WDj+cEx2lBmj5IiPg1r18zZ1kgXY6j1PYzSbD0nXlgjgqdmadeZ
D81J4IA+yR8gqewuPCUluafWc+sI8k+9bPl56z7aYNYMbKLGu0iMohmk3U21sHeWBdp04XFSgOMC
3pQeVYxqh+6MgD520fvogs95s1zbdmcBIco0TREGSLmj5TPUuz/QxSO4aQus+pA9WVnil0/BF2Ba
uHU7sKGQjlgynfDt1MF6Iv7i+pQt2rpYZXN6l+tEJM9PpAc+08Kn2/uEMDQOk022lQNW/r3mkEmI
oj5eBR7dq0lBTXRnsLF0K2E5mukcP6VRYhMQF1/+nk6K3bQmtnUhNjgL1yI9CowB51RbyxjztSfU
JQI8KXuMoH/dgX9ifbfcONyjRo24aQDfL57ec5JZjHWxEcdb4iZsJCDQSRJMmXHbc7f99WJe/oR1
jYMedqANismuzn6vNVXA8kZa8vUE3z3Y+JNUxjVp/lQxUt/rgDSzm+xpTl2hQ8izyF8gf2oWAb9c
tFdgdKtteKQ8Gk9ox32Qdg/o9ili6DQuawG3ukbWes+f/ZlwI4a+3jHVBETW1LD1LvqdgtIP8fdP
HWpe5a9MapKMa88xXn/d070ooNg70lwNm3FyTcR7CTk3C4hVG65HI28K0hbBdbIyuVrLXxkAERRx
qpNvtHGzJK63ZEmnyojiskSYiIlclQbnQjs9d8Ht6E9mcPq8/gXFmY04on4trYlLN7Azg7ees1dS
BbWWmxSR1z6FHBb8hI9HWcEIbXL5Cp42BQKQpmtnoT01D2nz6AKdu0GfePFcmFwwfKKc+Rm3QgoU
R5zBQfTFh/SHXnXSOVHogUhYLugZOdepr/7wBQ8LbCMmbveyNcEf/yjZFyKKAcXgd+K/4IttLK5s
WPBA8i2dxYgsJW8IVPG+xRdO95C+JgjaZiQOfhCaOgtk3ZXoIwheftNgp/l/UVNxcICWzhvIT331
6AxkZf1LDlypoDQhk0R0C71/dLwWE+tdm5nOOHyZC/7E5KwFdSIcHPiq/vXbEG8MbInT8DwAMzGk
Gfd79vyRqGFChaS9o9FU3QctlrP0vzDNUKGXZMQ1rfewkTsnQ+lM7CiFJ3yaaP43LhA6FzvegKDB
5buqIP/In/MeMYXle4OuFqUm/8SNC+mAVGjdIurbSzrGHDBqjWx22cU88tqqk5cbAI1U/SJWdza4
X69tbUv99S356b+DvwXD+rqhCcAwl6MZ8AI3v9VvR4Ao4mReGmm+2kRVkjOD+DO0PyL0B1bMlmE7
C8GyxaQHr6IsYGBCv3QSQ22TrTYxOgcf9RBx1zBAsThmG24e0vWwP1VficClN+9c35074zU7Y6JH
xT5vm7iPzN1YPOclTPPNblpReCW8ItTKvC5YxG/1gjVgD2b2r9uouI09ixLhVOj1rjpjzTQXqyfA
qb9xd6EmfsxilCLziRAom+1NoBhOZ0u7PRdcU7Ud1EefpVjVHlNJ9kvfl4SOQgydBWc1ZJ4to++Z
E7T1tGO7ESIAtjzSpRVdXYeRri9qZzAEYvKPjIih7NF1kBVnEIkEmfEQaaYTl4GU4XdRqRVd8y/0
fCyF6k8X8rLH/RFIc2YWZy7S0kHNQspwQh+2hgE2CA7RwPE7x5oIj4fqwvbnrpK1BaXsvqkdfGO2
0tcoUcD3LpZde9RdOZrzGPB+O/W4O3izhO8i5qrHbu5Pw8yar1NJbAJidDT4VyzuzJbI2XzRymW4
xdRkafxJLwdLJpwwahPHn8bp68Q01K40qy/4g3+RSPJBTDZPNCQ/ga64C8fqvsG6UIKS9uBXizQj
fbT0eJV9ettVFai7Gc5dPKXaowu/Cr2dytWtm6TEhUJ1XQUB4TX+zY52laxgVn6y+oS+kjbJQ+Qk
Z4IVCA9DekMFEILKHuVDZe1ccHiQo33nB9Ca6JDOH83dc40Y89y/muxwP/IrSbYGMEU7OE7DkCrg
/NwQLxOzIFl6zszqxeVByt179w9nc8jdGjrgP1SFGkqYKYb5ivYw20npE9edI1klMQL8RJMeKxgH
NTzfaprx7EsRGeVJbHuHy6UdG0WYLUWdx+KAa9+jFvl1H+p6CprSlrAnL64SlcRXHtdyKMdANwMa
CbuKHC+bReOnxQVLWcK7iZdQhVjKt6QXwZC6OmTxQLbH42tJJ2YvImjUvohqxOU96rLFsF14Z888
eGvatLGG6yZUG0Inm64aOnNfSoWtNDCubcnHx4JPnj//0tNvWxrWLaBUfmiwh4djW33JR1B1fs12
SD9CNqj9Wo9qjQcxGgV9+VmmGDx+MURL6hfNTJRT8EZoQ0PvpBYau2K71hvzk0FoQGMnKuBQCxSd
hkBE7DYjrbaY7ET7r+3KMRM4hTQ1+vzOMyNw1y5k1p90mihz3ZbKL2zJPqPP/iGA3pnoThcOBe5O
q+sHKJsqsH/G7m4W8rtFGKPNOg3d04JJFjpvMihJsQSmrOpvSvU96lTDuwPfRX4VWhnb+6iWD2WZ
vTLCR7o0ryX8A8lMYPG0Tr8KvEdmx5hGVVQ6dzyr3OfL2TsWg/HL+uIMf/9VGOaVHER7TvT4HJzI
ThGSr+HYYnRThk9G/U4NlPBsUHl4dEeDbWc5FRTBb8+uG0lym9ND31tNf2kzzOkto+YsEGmyObST
L8Ot9c862fgUwfJqFJ6sSIUpngdERmh62A0mgxC6A3g3FUyf90jMmcPPC1VMf188Wu6TJufODKN0
saHpJk1r6QdsDAAptBoeEoSD6KhDCEHwKSFLKEuyc1YZNO68eJmOWrPyrgd5ZQ3ZnqQ71AMEbDBG
o3GWf4YEuxtfnr5wBRNXGbWwctDUrYBvqAnRX6wGdF3d7KuFhX9kvjbRCZJbSSq6pv/LVq2U+pp9
Cg/ZBGmm8Gppsj8R+zBLBmSI6CjXh8u6a7zdfrcWSrilm0hS/6rfe4dmLH1lfI5sfoXXC2x6sWaj
Qx7flMm/fEiy+8OCmw7mCAZavN/U3Ik/15KI19e7qgx2flaI5MiHHHPV2n21j99kDEgkFp1k3KP7
uC3B6eo0+OFzAnGKRK6kpIgjULvhVgVufy+PcT0AJ5xUJLPQT/9lC9H4UAjnFffLD0Ms+tljAxwT
b9CbG3MFU62ypMIabJ6v36nsvDthidbN4iG+lhWs+j1JAEkFrCwjSSMJCTNhlgq/Kgn/WWWM4b0o
r+r/Yczy2uEJyz+i2MC/qX/EDB473IYmMqtrY7ZNoYIuCdNVEtLNyTXsyOyVnGCHFLQCtlZUgCRE
hbyyB4OygqG2x1JHkr2d/80EsASjvaOWqTFKaVqCgU39VE8DaOOXVVx4yiq+AA0exPeHCF9qJw9l
nKnzDj+08OWuI8wNlEiXCT+BwrwAtekD5+Wzfi1sdzaXc4ir5Ibw6Rj2S32EQSBJBIkVFWt6jWX4
t2roi5zNBqCjhdrzL0QsrYthkb5qo7Ln89xPvsbfieX3C8Juwoaxmw90TjPR9IsHx7EPAj3s60Bc
k8kdtc58HPe+kRr/eontisuydFF1ADwxnwcnVw2GvXcfzVPdDLQKR1cei5av0zEdvDW+rcykgsj9
U6R4PtRa2I791D3JDaio6J9X5iycX2mMDZmE3XCLzQaXpTUidoIiI2WmOWh7P3aDB2PxVHvpC6/R
XhbkakwrEf3mIE99tBhg3P1sc/59s1rcvVDoDkKhJA0IKM50bgx1ocRp7tMYVd8p1sVixs7vAoyk
qWvdRKk7kutqY+1vNfziCYi6v0OekZ8vzzmNARAVgIl8eCiIZQF6BZwLsiuAbP7w6HsQdUpRyM8p
oDnpt26F08dMMtC3V/JuZWRxn9Exebia9c6OwhCUxl2fjenDygFPRmKSOxRdCLwmVortjmdjCEr1
bKJeqM2G/QLWlMjz6zR6sSdgHubFWVuhys6VtWtB3EjHXHQt1Q2BLC71g6Hnxsz6zb/KpFTCh5fL
f1nROQS8z+0uNrSOupkPqyc2pXUz23hIqrb0pMTd1jdItfwr2/f/YJSqtSZX8fGJd8MIGvoahTMp
Qzokx62i+67MJmITVvPqd50PTUjRV57dY0BNjh9V/WxKJi+G8UAIRUghtc8ML60BH5cfeVXOkYo8
zM16TcTnocGfP5cjU800IGAJAgZGbNlBYENS66LTeDPRb6KRiXj1z/jQWrrtkQmk9FqM3CmEEuci
v1JnblgYH0XPDdDaWDdf2Y6PDfKSgZKPNnN7a9kE2L3ZHZ3I6Vn3U7k1tQaTqJbDvrQYcyitkPkk
BKMW079/2uEYMqOgvYMQSB+dlqYLCWZT8eQqnGPayX0N2/+XVRdLpbmogxSh9fAxlpajH8xhq7o4
ZOlfgyuYcGFCz3iqqU8KoKYllP9pzcYVXs+DeuWoAfEvUTl4Ypydqp8EErvVB/HljTtnaAFGHJfI
2CXDJAn7U/bGVUKSvA3ew7G/Rsn+ylA0J+GKkC0a2NtB+cdFXR/VgOOPAiMkdP7wRFeDWx4we6QD
j8A6VZNQbUfV/teSXQGWy2x/fOvSrhw9VqWY/arbYLAB5PRSzQR/NInE94YVpON2PorNx4Ax5zjy
/vjyRbMniucBE3mgI4hrcvc7jEyHMlIX0sSQlcZhhOlOPVb94SCtK0ZOtOPNRh6FH25r8QPVm304
a+ElMH7iS1HwzMbwBtN0ZbRrq9d8wZgNgtrXvDgLjaqyhHObXmdyD8BIJjoFmFY8R6Hk3iNhDgf5
2nKgi4BWvX3U4QwEYhYSNeAwFnL/5BiLpVZMPcQKnbS+Pih95JO5fTklUwb4g7QJRmc0pQDjY89W
IrxIiQD8O8SkOnnwLEcYBNe6JfrVTesOl7IogePCEZcfJtAmaHl4gyoP6zPUrMippZqAk4lbb5Xc
f97QSqqqSRSiTsVmHdtQfSTzvQY2okM5XByPqLhVHQalpoVLDZfMb9oJJdBQO+nbeyhFfU4ER9C2
YlToW+fQCtMrv7MH7EWsRfH8mekw+JcQ5KX8Un5CxIrY5SHd3fGMk9huUEF3b5SqENWrcSi3Pn6v
FXms1RHbEGGnAR1cQoPlyTHaP34DxCaekLO35xlRvE5Na9t/jkFZI72d8nRgO2VqZI+8DmHSmdu+
EU6OdJ+qz1gYTtl4EkHznLSMm4sXZUe/A9dE75wWNrPGqzx2pfhk2Nhgdffujv/L0VkzsHY83rzP
q4I94OJSyn7XQC1ACDXyqnFo2j/1Ug/PzgZ1INYXzzf86zWFwf6/Skxt8XySvSXiW0bLfC4eQDlS
0//BvsEy8oVeq4dRKuFjBo4RklW7iaMLIzpmPGXfqyfYsvRGkpjokzjyDM6FpSA+7XJG0EtF+eJO
EzgR7K24Xc+cQtSZygFRqa9NF6FiQfbwiZGNGz6c6r/aW+MNXILOGkiuo5qMaj6kfHShrVkNnBci
wpgAyWl4cAYwHbEjzWrt7Ev5ps3cnABaAd8c9eRhoHffUetXys8A/UFlIxg606JUz50ueTBAC16m
h04RUurqGMUWV7QbLu9HwEZnEcSutqmHdPdBZ2KrjNnBWqlNdHWaXes+lbdb5R2YmF5kghB6ECqq
8oXPruQ/3VBudCnOnF2fJUMCCTjEQr9FqTC4Fx/WyfrX9+zhQJIiE8La7mD6Muqqlid7lm8aizO5
D034WzkiuHXL4guIikjcFgfbSrGj/IDwrjAWcwe/6g9TdG4QVHLqxtCRw6SPNQ+KIrTsA5cya0Mh
VVdlXywU0OOaEbmUd3DTHAcrZXUsx/Qql03HiDfH7lm1BptXQPvJ0b80MZlItpGMVfdMvzQ7dF3C
sclzhVUporMKkjsrYVcdv6iDpVoouTqgas45maFOFobZzoe1vnmls76PBUDv0NENQSU8dNDhsabp
KfJoYdQc8KNi1C9dtFnh2ZATRaLZEB/LmGRzJJN3AJccf60c2A2ZmU6Bh3BV6xH2ZLjT02QH3SLU
02HMqZjSH71SRfvm+R1oPuhIoPBlr3dqMW9G6AYfB4fHuvxaa5LkU79USDKpIDJZO6YzgeuoIiGX
7WuyZFd6C9Wh169P+F1w6v+mQS5GMk+n4x3+6lgNkK//RPZELCnRDXw+Q+eQOhe5n1RuWqqOTQez
umsLupk545R9ubRTp3gdvczt/VNQLtx5hnjEcQfJ+8PhQeSlwvqHF2Lu41VgF5j1GwRoo8RB6xlQ
RRy9yDqz3/t+tUPJgN92Kpq+giJWrDqduT8ILJImfP2H8ReAsuzjPcBB82k5bJJFYjUP039nfFSz
XVZS1iiZK1sIIydE0skTS2PnF26ugU8X2GdJNvq9df2iE5kEfHZd9cnuuZb7Cazjg3751JR9oQlD
RaGehN2XmaaAMcPwjzI4n38o0l4WNYo7HuTIwkYLym+Wypp/Lo81AGYflX2B6kwvM0JRfSuLGyk7
Vf4wmpWmN6SUuqiMgK+pGo1gWepdzdtNOPDv5+mfA2KRupgQbvCQygRlLwLkMoAjP+qauj0eFrZJ
oopaEwPzFxDqGoRK2KZMvRtdNPZzukoIY2tpEwwTNxf7EPDobI1h6+iASpVP656KhGpRY+KKdls3
KAuCNwU2B4yxZG1wohA/gRWrd5VsvAO2iiAjc0/hLGutu+uhW43Tj1dKcAut9m9MG8G/E62o6lNV
k9C73dM3QyVf1+uuwMYVqZgiIU48jqMXw8EMKtkAkI18TmyVUZza9NopX4EDuZ/uzirYno4+gk5B
E5e8VOQIskxjJM0xEGMxZsV+urPQO1aRwJu4cPkGlLm04U9y5KOeQONUmB75SEX+YDubLv1xKUhT
kj9msDforLdh9wPyM3xMlrFzAuRlBy3dUiLgHpKFopIqL+gSeV3bfytIo9pP1Tz6O1y7LBz7hejo
4vsyMqT4hWYwUs10muH1Z70NA8jk33J9egyHYS0Yef3EkdJjkwcVQS5pZDyjug6U2AsBfR+LALyJ
y+t9oWUsZiznIW7ZkWF3rBM8xnco4cFEpVBEBQIhvaBZ0ZqN5JMeqNgF1HRSoPwU7K4G1V2hojyS
L+yR8LS7hGUVE2dxNcdfhGcLhyM4UuDXeDoyRKTk4j+IS+Kfmwgh35DBDmhCR2t/EHO0HggwiPKm
0cTwb54XapjMp5+VtY8afTEWuseu6oAFoegSxnsqDEz5m/ZEM+eLsp1kGK9JXRV5IPfELXZfA7IL
it3VYaSBFmXMHXFIBCDm8TYhlAM0aAHfknGHzrs8g+AuCtS/pgrqY2PA3bruTRc63a8m5pJ7osbh
464mY3IyJ1DLHH99JzBx1Z8bg8FjQdkUNGrV0e0zkMSytqaNM3Sn4holAe1UhJ0bQmDCXGWPhjYj
bmHL5ri2IFGFkfKztpjQBZ2745uc7rw6x/zlZgJPyazt+8asIlZiMqLR49zNJVCE+BWprJc6Ni1f
0ygShIjiNiRnQ3p9EbnClxQq2S8dHqUpNt17VHDA49dpKdbS3wD3CT5Pd55u/6cx9Uihe8lBPVvd
CAgF+69Qm5l31lmBh63w0D9R4Md2fKsBqnex1NLYAwM+QMJT6sfvG2J+VfdmqGpChe6a3ll29eWC
y3I2v2ZQBlOvcdiRqCltgUuE9ge2KeMhF8Nx+/sKGAHNBx1vgONQitdllxdpHQAcQYGQaPNRG/Jx
g2zeFdLpuygPhpR+5IF09B41KSZwPGg5FuiCiAWpfMPJGEfuLAvLvcM2omd9nUEeOfagPzhukzkO
TZk652iUrosb8UzRVq3NJP01LHKz+xtyu0AagQIfs0+e7E9aHlVki6cMLyMV6LFatP1Lw1v7nYOd
30pEHxN3Y0b0uRK9GXR1XDx2BvupBLg3TjyT6F1CQnj+1pDuU2Izkov2881bCl0fOqHRiSuY24x6
P2J7E8XHlg87sQ4hLS6wxOUuqX9/YC5inXwAwOVQCJyIDQYSv2gK4V8gPzavOoIAalJpO1lbls7V
jnNzPNFpMtkEhWJkc9JY6DoY2oyoZLBGTFVgjpF2kuA7gWRWTdfXRqN7rTIPfnIM8CmAj38qd5vw
WXGCjTIe3cA3vDAuPky+EMV1pvnPJ/tN4IAL2nrcE/r7f5y81Gthvq5bTb9LSj4hU4iaP0828iQQ
5IFqT5C4+mIGX1YmZN1AW5qs5M6q9PGfBAsesVZF4RM2nH/jZVGm5mSJWyhFhvw3VI5fkfZgGzgU
8XaoJp5BpGySxV13TuUsqpFDAyad30WZpXxeEgwilfViptNjldlLfkZIpUqHOcpt5mR3oXJyFSNN
qMNlKflx+YsCY47v8L+O7uvRTwtvXlb5GvK4ICW/lwQ/yTUcJE2KYiZQeIGW5Db5MD0Ar0+VIAD7
MV0nuO2b9P1opWXloFgDXz8G1aqA/IdhbrvCUXn0IvoP7TzAxBMtL2czZsNnjGdbiAtWP+3kVo08
KTnS1tWfm8z1EQK6dGt0iPgEubCP/20QbV9+aeIhp3r9rKLZTLXqYzYN1Lhbcrag8W/6yj/glQWX
TP9R94mVl6xST7QNWwPWEcPfkCBM8Bs6uZX1ps5MvPYkOAO9G7BU8FK+vwTpYgkAk7tHiAevF9pu
o/1EWlTSnO+0uF8T8y032+pRZuezW0dhwqg4BuZjhNiXMrURDpERR+v8KyGmq7AJZNeZBmABBFN+
2USCRB9b6Q26TuKy2Bkz+99HQr+K3V8zlyPLnoBWSIxaGxFcTCVIfBprwOVbRJm/P42/2b3K5GFK
7bpu/0XnTOk7zZhQ+29nNA/NJnQYUauEKPUEmDj31RDq58ts4rYayM46W3EChFq2qQEZNzoA3cNT
KkLLPNUbQ876tLqpYhJ9qWFRQ62wf0r9a7LqPhHyOtEaUYTYkCtju9omq294yZvnH5t8Wplp+hXz
C/LN3/M7Lam6icytWRAO/mPgFQAOYM1Pt8uws6p7t4iWTWpuC7gz7oybqcXeFrZItytjUaOP/iZm
0MnWEm2ZL50dmA75lu2cL4in5nEpJ+V8tUtiY17zI3eqQeLJC7yBOI9vB6VypS4ry4BGo/GSJFXz
/PUzOb0d6XE89YmQYexBIYN7UCz4lgqBMvLV8kvyKu+3FtfWVXj9/s3GvO7FSLa0YmytFQ1bhEOO
9nJsaKhVhZ8U2aJUBhILwzjTLqI/sy+nN853iQMu1OhyY/LMiISMSoZvyipX57YOqIoyuiY31nKW
aP4YCtse3fSLFkrar99uKn9guzbi1LHQ39BgkxRxagmL7BQ4LkwSFChfXc7U70yHpCapEO2afHeY
977x+xpkb7+ZP+X7Uq4puIbZU/gZ3NwwUMYe/1JDEGBBe5gAQuuk0H6yLz7FlKMM7e4A9SrczKQC
PZhEF6em8glTN5xalHO/OXfv4e2ZjJMFdWiKf6U5Z0H7+4Rj2Qe5WoxFw55xJykaGjjiGA2ONKo5
hublgeleqGPBE0xJ47e3zZ810k3dwEceb13GrStxeLqGrtFSlKxhShb2zX+VS+HXD6Bk36CtdjNU
tmZz0iLczxBxNOhhpdjrTcZ591BZxpWDjRH5wr7sd+Qw3z0y52mq7m2myBqD8M0/E4evvUnHkeHw
RiVHd0/IDjcvuCD2Q6V4Gk7syp6jUHguQyETeIjb5U3iMpdngBsNO3egCi1PlbuRU7N7REL+9TeR
7jl/5NkV0G/MG9lsEBhApNXmz3bGL8D1ffIcUkXhKbp5jgV8SvA0NvCIRuhr7YGqZWvBSDX0wZZa
eseqpXaFlUqMQed8/0cuShzifyQ25NF5jYn8YNq3x2EHzFXM61O4kJ6lDBsuf8k9eRd8GaiLNufa
sHRN1HP82feKbz4o7e6N6C+ZQtHG6LEYw4SXDKRahtCdob6SyG+LnK1KIn59YdOSKsNS4aaJe85i
IrvPNdY/ROdZ2N4XUPRQ+QwTGswGGhU6XrJYRcSh7ypazupjch0tWwk7PkqFBm7L/atdCr01hhJV
Ch3LAD5FFHQ3vrOrw/ruNw3bblBThz7dqVF6Dap/o/OSXpJvVx9v1lzWcfGhgiYcxpbEV5PsY73t
eZFCKnTQEZx1epxtZkNk2S/5Szv9FydfR9ovitb81WKWgWMtLrHn/2OisEoQSwa5Sloc8+4As5/h
VE+0KWjKyyJMUIwoIddnhYRdnVbDqDrrcm4fqK5XAOHaN54DplmYgbV8qoInKFZvcxtrSRBIpTmh
/0GoHSwP5w2uZLKszo1flRcF4UK9ZZBvXjf1C5yVlUqcRT1lN5bvRrpuqdjG/Yj97rAU5a88J+Ex
E4Xvl7X9KsHla/PyClFzMGxyONqfgUFcJREflXWKVzG1W4OLeJ24bRanrE/kpJX4OOeoh368h7Fl
+sbEdPhJw/I6odCdVjnYPkSFo4VXHCXnVcrIcKyBRtTVY4AYiSS/k9Il165/R0zvGaJEths8ZTvm
0WWT36kmPEPc27kj4BA395D9SHbr+hLdWiXJSrYDvo/MgBqIvXQAiTgLuAo1kCHDLpE0bRxa6vCl
Bv02xf+FgHGHL3AxUYlV8D/WyCP5e1lpXoPPiKduX1eECCa65UOnNo9DJUCcqjw0KJVLCdHz9vJl
Ngrc5YkfMFq+lxsJvmK0DaeIFzx7Di4t73r6D9XCTk17DtyDdpUD6bVZ/vA1xpJs5MehSEFHqjL0
iMwYfLvRn9+ycUA3G8yf43dyjJiDwaAPg8q2aF0u2u4vlBamB3OwR3QdJ8086SCFPbLG1CefDBvx
0QHEXAFnscJNTM2SFhMxe9WM0tgbkQtRnQMdAM5jHLt9e8wfuIQYIplkxNzTdBHyjU0LlTS5i5dt
3gFp9/6DAncokbsdZToGIHj8sC+YQ2H5wucptIn3ZM+xnVp0EyY5mBc1XsVpLoOekhGQBvvWfpxo
k7N73Ic4is5H2SvGYKJRVb86zAUJBoXmxFOFedfum2GklFmrEJT6gvgHfwU2diqzcwzCRpjgpm0Y
5cfjTjqPHKzOOJiFwa+GYQC11Zft6MVv0UXVy/chJIGYQ+YGoAssU8njuaPTlktyNw+U/v2bcmqR
zi9Fv/iIBC4TgTIY5LxK5xU9vKYQEQZQuFerIVwvF9kpaeqwXh23w9x0CYRB26netObv8xxKJF46
J9i3ad/2QpMuld9xHRb7OG2DuxXvu05LRFthqwqqWMiRQdmR/tmCUnUWffuHJv9h0w2RcQIInCKn
Pr8p6uhGp19aLexuZVp4DlZTKIDCzzm4525Tv54XjJD1qodselE7AzqkLi8ORLIETgS5BjHEyYIb
1yaAXvG2XXIRcaSlM1Hrj2ejcPBp8Ncg8mUkpB1+Z/6aAk7UACPKpJ2zX13JKoqwoeZ7J4ajh6Dm
JssqdiGVZh9ObdQ12rlXEYnD5Oez7BPn7LZjpwlgFNRaKmsyC+2gc/OQhGrnaoswoSobVAnhy07E
FzgXaR56mNZs7X3XaAFFdTl6HGN8g6b1oRLDjPfn+NiyIkFbKhOnhc8iliU92467EpqKzkGhBSti
oDr426D4KeDQjZy55UrAea1yUlb6ZnoMdSOJImEjv2EnyxTt1ebzwbuHb8y4tyiY/SPs/PLdgfoF
dmpUsU8TJjScK1jujaB6pyHNxpjNJ8HIGopj4v5HSXyJoRy/K/kQQVEWwqRKX6SZKes2SoerPgfs
F8uvwqvGARdA6rMV6iI1hQFyVP+sMttMjJ/BYkmqV8NtrDUWbNSb9TihBCUoYTRqCrYjy5mglPAY
5P0ULjtDxrJuJT5ITiooP96UPKzSDKVnjUavr0QlaLVCqOHdRtxL5/FQeRWR6c8Iw0rUmZCaEWPR
tar2+MoEoxzSpk7x0zafaOda1CA6a+MLHlUvfPdAvO3zRZ0rjn2bPhg2wdmI7G0kC/AnhXp6AzeZ
GrU6tkHovjizbncTfmSELN/wIVKnWABA0Ddvfh3TEez42x6TmeA+21iO9dlGn/WZJOYUqVUZ+TZD
3vGIS37uG/NERmU1OK0NWG+NlCegnENbCrSghzK5evI91HiF0+q2cdzoBF5IrkgUc9X4Z0sF/zbh
vGEIm/RY6jJMC2/NP+2/RXdA4MZ78VQlLSLFfUXoMYbx88+9QAiCRkZ6JrioVZyuHdh0kP/M1NMe
sO7ys+vnuZ3VJMiIJIpiR/os9OFUuHe3UmH08mqw1aAqKGO6eTf1DPeBtyZggJaQFQdQm4jAn7mw
EhHOYSh/PzyLAdYRmSfUvdInHZTHCnZHei3n8VYNtD8ycUlNwQ2+y1evPDfLvUCnx+7meVujnkqP
gLQnNi+4ozz11gZ8FiKKubcLpXI2Rv+wKs2qUVq+yFLp1rF8t2fHMF6jf31DNuj3Ont1uioxPPS/
bWquSJ/4WznumMgOlEbY/mje9bGaZHKGlckvb0kdJVYy05hrlVVSQ3vcbzndwY2A48Dr9MEx3iNV
nZdVVllbFFsc/vOV6isVnvNm5Jlg29nsZ9O9mWUqYrmRlHwKSeCAXZ2MP9uL4j0risfD6EIKE1b0
nGKOHHgmv/ZYJyaTYrksRrkPo4Z1u653KGs2tgAkQJErAi2JH8M2D/YbxrSuX15MyA1J8xXd49ih
3CokfIIXJ00q72jHLP/KZsLGPNx9Cydc/5rXPSQnhsLVflnkP8aSlMe7Jf4NrmDz0Yjz8HaR4/4o
vo5vmNCx+fiI+QoxIGfW9p1oD1TtjoM5KukcUjr+ocX0s71gPxb6dsfDFpGnuCA6mnILm0NRtMt0
AFplv9YJaK+zr7gEen1OfzwGNzqM2skRITlWkimGMiDUouDwmIgoWat+AKiyDsvT6Er2OhUWfMg1
ZmcdmlKChzzLbqNDRvdTFDdbXcnAMz+pDaqdfMxULVjU5juTPpwQgkSErWccWrDRhPf9seg4zAcl
znOyFzdYffw/fXCvM3VVrrfw5IjVNErg/pDL3ER+BvCvchEORxiAiJwa6afoAIZ8QyPn+r4LGN/1
lbTWEJPZxw3qJIk4NeBCVWZGXfdJjGQF0t8Fi79N1TwrpXB5Kyvpql0/9yvF4Q09j0UBmBRvaAGd
8xLwqu6w7J76hmdU0DRcIU8S/zNjj5FUmaqFoIB+m3Xqpy+tbtwLrtfXyBhIxwr3yGKhhm7trb9+
ocz44EYqCZiY5Y7XtJNvd6VvKNxzUUyj8uWg/DNKIzYuy4fX2UVVyMMaIoMtHK8/4fkvn2cmNQhM
FF/RP2hvcR6zOaeJUN4nHiNzSS3ITLGacNSpUNBeYZZ8Wtvs09afsHHHVq/wJUIbg6WFnKx5xP+m
su1clFzOw6ekUT/TNMNdp9/bQApB6DX1l3Xb8JpEv6oBeL9iukb4Uct+byZ7QxRDSaOIdPRv7lyx
jFxKztheWCVYvK7CnZ8omBjCh+neoOCzzNYyLOQrarFS2CkfiOYj4YEinlZbUnPQPZxgVbDwHoR0
F7gCosiG7tcJECKsdOObstyBhPXysXNrA1rL27GwqNirPDKJnRhRyVkWqtn9fTLWj72V0v3Kua9R
A6BcqkvTjCWLgoSLf8KewOIN3hPGWsnSLYsBoNaBFG2yfbfAPZEoGeyAVEiH5g2BF5CS8juQbWPt
XTBe4ceggZioi/yKYU2tNlYCY+WpKZg376RyWJUUKDHu9wx64J8/hHvuvlagLwnU1v49Dy9gydXu
//fj9VetFETX+Hnv89slFWdEnHhc6nsPQANnMu/cahX5Nr9tpLauBwYJ8joOt7vS2oW0s05cyPBG
WIl5nkpdVZoXFWXCbHpoQmc3iI2Zu4rsmA/ER8OPlsy6jOQnrRHZ3Z4Ybum1wFZC/q5QMCrcbGtK
TjEk0FR2YcWXt52h/RbiHutFkqzg/aL5/ZE1IqOK9cgw9WN6BZxK3XDkaQO3V39nqsQmxudto6Vh
zStkURDf+OQVJpd01QIDFN7ySEIS2hru9QUxNEYAjbMGZxX0wsvTMbtlJIb2VOfaVg6y8MbrEdAb
kFK4k+P0EnseV1NB32FXezziKwhqPsBZNPWPMSnM1Q17V2jgSXe3xgi1sVGFd5i5uP+9EbZr3Y+y
Xfdy3EHEjm9hP/eOmnSCRdJBGGJsPMnQZanfS55zC9F5qfA3gxMA60FzTKuOYqsrTj1knoKK6tmZ
5RP2Ey7PernxIDK79gQulQ4BsD6gojXd1LZBVDey6UsxTTPZxMMZ/w8z61e57HVYr28PoOQGBb/I
Yqq7rq/UsXgJB8YM2evikbnDbA3MqZFNaRSa69qrM+py2IWT6etoyxxf+WkUnYBGf4XzzFTEeY5F
7/vZNIkjx/soyzzkjv6MjzjYPhmDibpMPQbhH654cxVeURVzdkPP7T1q3T9vlKYv5aWui46NShl8
yTS97iDrrOIN1MOukH4U7CRMdL8ekR7TudWZtFjxr3hTh/KER7lY1JMppB3UO+kHwaLNm9r1ayux
o1LUHdh/R6MqGRkDc50ZpOBUVkhGolK6uRzuYoOhy7KUl0WAV18eaT7D9HP+RHRq1yPpzaZ6WI6+
qtM5yuzg1fD94PSnLfjTDu1BLFQVfWxT8HcXHHqs5QWdXqQTrBzu//TdnnvyDTpfGfjckrh9c+2P
Z5pG22FHkZE9qovy8yV6HixE7bYiEQAjYPoo8qXmvx/4dfPcw4bTaXdvv3EBmI1L8s3Vf8RsdN9f
7WivbfBhiECRWmGFYe164dVhhVygOMSNrk5h13e5m7BY4phnOfjjZ7vTb9KbOST9ojRuLdQtfZiI
LZgMg3BOBhf/PGwSI3sE0E3iZ42KIecRfyKgVwEgRmr84TyIeQRPG22xG4QmywnDvFFEJfTI8GuG
LGZfCCQG2hqxsQj/ZbL+zC9PWIX2oYCuc0Z2Fzi2DijwnPSRRg00BAzFB69tDPMv2EL0h8Hh6pB1
d/Zf/7pC32Z20HT2sSRU/neGv0CTuDXgMwDJweax5cJNa4yi/THBvRVgI/RI0YS5ACn54D06Engu
22dm1P6hUcJ8Zz6w6vdUA+Wj//nXh81S5Zi3djdEfi+hOFqEWeSSxyhz3sL9lxq7BhcFL2oFAjgo
Wi6H3gtOmHLYyGTgRDkZPZD7VeB7Zfn9QUtpNiL6fpmxVY670ySGK8G6UGiBbok7OANWmL1Cbl1R
2c6SS582yqguEN25tftNrvPnFvRQ+YSyqegFqWhtHc/f5dyBAnh2Mqy8jfyqR8cHVjmxAO4c13ik
EFGwQx0uV2t39TLCoGEXL2s+njQXfDhJiqjlbJeVw8lSQkViVSe2aJA5W3+UP2FEjrKra1qeR6W2
IuA1FFhDuUdMZi8RQ+OTqMTyA9kkzlqKqxYc2GMcBdlmfRxHoQOctyWNStM7FQehyVclo4nz22l4
b/Gk+UDLsXEhtEqwnJu9PC54flIflvsujFYgh85hvUjH7i7oYvIYV6NIhHuUeKqYiZq5c2igHDA+
ENseMCMbz91GwX0YjmNpaBHHFlSnrQRQz2dpXev+BD0Gt1rGqcbUoU1Ox9TvjrT7E9VUwp+xEREX
AnsqvB/QHs6B5sKr/kaSgcNtC7Ieov93Trg5ZuRPP6dgJohhELbHw5bIqWEFQR1f74RkUslzGw6K
TeAI7ZyfjwFyaeZX0wG9Ooz3twbxkYb3vL6PD3nylOO4gX5eTjrZGAN/FFIxeUi+qaeb6GHQzCQ9
ReH2WI3a55kGQzg0n0T3HoKKnrZuQs22FYrkPHJ41DoWuzJQyh6wXZ7bTi1wuenXXM8zhnsr1VJ4
0ZnciSwH5YBAhF0kh7fE0FOlDJ1i7StlPAP2JfLYxEhIicu2lv4Esz9wDWq6LnR9ZYTE3EBifbeI
r2jg5uJ3CHfXp4DX3nM5h4rX2cb1GmhkIdN2lgTgXCn+smoo5sp2ywzYtcIf96ecE3+DhGrOzXJF
IcHMrVEOdq6KsDkwofKONM3sEfVfjbu1CCeg2/n1KGBuihfTjMZ9EVnU4IqRlxBGk3KQUeqtMdw6
tRk29ItJBO2EsyB0/OHC3dF25zA2nq+jcwAz9uOc7xwF0O8baZfT6xME5MbB80U1D9FgZQzFfzCV
X0mqVgpwxJ0siesX+J6q5Uijb2/bELgxsYBJ/3k7OxZPGveUULqzjz+6Y0ADvGKFROUo9AHv7X3o
ZykRkDZsonYHtgnjw/5VOAjRMQrIe9GpLn5Jggdsqrdf4Stw2bLdIREFd1sKyt7m7FWNXK8PzOqn
5I4bzDOE8CNckjvmuDRwajSUuSTeFK5WXVGc4XYW2ePb3ZFjBL7ZmrLjLOrBgcHXcR+fZNBmV/15
ATzKUYSFLjCzBFClS0ZVhAKcl0Oz5P8k0CbZR7xCbQtTGThB3olISW/nybCp8tXWPhjKqnCCtBf+
OYVdo4NyYGwPEAVQ49BZyldDBFSrETs/+7fBxXeBd+FTBoUKQwfXUyrLYbyCWi55vbjrYzmX8Rc9
NvkWuSGl37cuV4XX/hnqk27vARPU/vrs5VUVhVu1pLMAIgmJPnLPrXHaZCDmB2uLUjay69IH9TCU
C8x82sVB73YYxz78gjwrqTVl6q5kYteI/Y0o8ym1FrYIpTUM6V3IOpxq4pDwPPAY0l/k1LE8npaV
QKsPDnHJ6wsmacb5p3FY/Tf4mH3rmnPCjo6IjFJYi3Sg50Dz6e3eWacfDqLObEBo6A52YFt+D3Fz
TY/cI/CR4Jnaud2pqUWkyslvirGnQSb/krpXNsN5N/mhWIXoteFS1t5/nZLIZLlZJgc3VQlZQh6P
k1ACGRPWyxMHn8lA/V7iJE+8RV04ozxZBHo7rMxGEVeAij6cBQVDMQyUFIeEPYdv+SWtjALEy7WJ
UWmQPBWzdvMDcQ+KAxs8FQtEebgpYoxkayATuPg/kySrbv6P03qEiVfOTADtZ/cPE8f++26wgjZZ
0IuMnYG/xk0kCbODtKWQbrdBLRWx/4ZBXc7yFthzv0Nffg4sqeuKgOqw1ZKxEJskVBkFfM+VbzUI
NZqvUD+CqcH6+xFGj+AOJ9zko8Z45gcs9DkCkOcmYV5voqsdsAoSZcAm+lIrSod4i6wUev0CMr5F
kjm6LlebknyJ1aQHLA//+qRDk5RTn94bo2MtkPH7BqNxYxmyLlOujmbJ+zDOtNfPPZQTQ9AoSisM
kHhIVMjVhmfpHMkoHveogM8aXlFM8qE8UhZv/71p+eXpE0BhvNeZVbYbnNIHPF0RVQK6gut4zR1n
eB+RvXfR+frCnJElDaQWzG+oZwVTDWqDKZp9d0i4lvwGZgKGl104oVk9tBIkREiSf0KPSHztaXg5
u/qQrBnb5i/Z6DTYGVuQgs0B5JiaMgLJFBCgSflmfWcD/V8o+sUcJajGtdInKnX05N+MqqveoTIL
Dww6yWdhP6IGUBWhdmXGWamQ6nTGYJxNcDC9vYGtu48XcbsupsTxBYInAmzdHkAYDmRR2IyTBXDm
FhUExmBLSSId43MLHCaCWoXYZbQ07SVv6GAfpwMdVDCEoNHpX+b8gNhENrcmUknC21Ku+plOatQh
KZF/4EQKAD7rUSMDnSEneinr7SRX3px8t5aR3v76PPqZo0/Qd5N0kbRvpMY5MJ3vFKdz+/VaBwf4
PqBZEDLkyHc7n6iaolkbU4zlUSXmGRR8AaezpO8xmbbLgUzBZ2AiFI22Vn6q9J8UgGe70uWOhYoa
edShhhoAUsLlZyoTnNJUT2dLTEk91PxNRDt1CIsxiPkfkARecbCarRF2mZDabQonxldBYgyU0xXj
T4JGMPerEIqMxuKsd0f5Wp9mvyrxekD2dDcYgrnRUbBWyV4WnMLHWXuEKI/GfI+6FGs7zEU9YmmC
ysMR5leyPiicqFFXoWmx+r2DG6Y/MVcw+27Ok2TGwPqTOia9bX25sJcdLyxA3ffbOJov2gB4CePn
RsKN8OC7xVrv1JV7S0h41xu0XoiBTXGwEfGrDxIiok/kZm1B0q6VPhuTCULzTwAuNGqmLj7ATZ/H
C7U2pO5X//ZHBFtEP/AcjsFQqDrWQROLXAmf1hgUYgG6RPupX6fxU/SBTdWIjW4qMz7fB5jTioe+
7pPaoQnaNghRocCt9qQ5URMqblrsRFVLqf1kWU8EAhUoTaOPeKQWMKHbbKbPr2TRZTmrq9EwCXnl
Y4AlKmfJTGjhEB0bxfCZCXBm6iXPafHqX3Y5y/zS7FX56B4DGLDInr1mR4sKjU/4laYpYvPNFY99
GR2IU2pEz1Uvbyj5GMAXZ1oP87UDXL2vyEv/Wa5qjtIo5XWmDSsfJy7tst1EnFRgK8prDH/0vx14
kxLusQ0L0aoRwn8/MTupjT/CtSV+wlOEPkYQZ6C+iel6S2CPIPUUtUO4OuJcyWwh8I/PwwMA9uLX
nOxNxlCZt/JxGxgtUmfVvTQxP9vISsJhSCpA7fL+v9hxQahbpARyJrqoxt7gte5LgFz+bMoLwfO8
Mwg7YxwNsBepIuFTcZP4T7gW06V5E9jSI5AMDjUkpxst/mT7Un+T8M8J54zz98KkOQJqyd/2/B+a
+ZPV4UpBPWJIm+D7vIxZqPbUouHcBixpJ0j69sUJHkZM18Tvs+PwYk5Q9kRgmpKHPUDt6t6kPL2A
O8P+hOKM02eOqj6nwqHBCSYFbM4Q8tyET4XqqnHNE0r6v2OnyDvjSl+ZvcIYp/IVRSkEHwpBP0ul
V4lwmd/MWesClqg2ZBE3wtnaMcUwmH9I7cB5NgH1jU9qdcoRZWt9o9bGvCa79bcBLxMazmvE8fC6
04HU4LZOI2/9k8I0SQnCEqlN58gxeRCXUzU8EiR/no8EZVyL8ZLJwhrk4QU6ZyAimdAyANlIYmzj
UQLzabWNzQ/5Wo7hvHElm/z2zi3vy+/2Ddru8N9mfFvfVJ7DWdGM6FsOdHIvLKYasx2KrPxAyVVi
WEEgktfCNrBXK6chjATDTrMsRmdhL9fqM03mbFioQQ+BnkzzEYN8lu+ipmVQjKDyKfclkqFsxIPG
AFkiGWMjvFeBUBr6mqWxhJJjJ5OCj+bxS8/hW7MGhDTU99HxI9OuwmsyKRrK0cqEBla7A4haWyIE
mEex/nvwQatgU95kCqNJhovFjZX2wx0NPRdl50w910KzETEHKV+VqIcb6REWmnPb9yw34Ing+jSM
ZQ0F9C9TKwBuaoUPl9GrNfC6JpCFB74hNwFZuLdUb9JT4HJNdB61ZiLKNa3s/gxTIDa0csWPk0ri
TppH11QevuP57B5iq+xZbaNC0dKR7RUTT8rtFZVtH/Ae2Ay/zP/zKrHCrcEpNLVwJp3ZCXiaVY4n
453V6qcOhAErnO3oAiGCZ5KISaB4SoTERWmQd2x3a3QZdCm3HOy1Upz2uu3q9NezTR71IuVLVU6M
7mGPXvsr9xlYFhhV3lqUU/a6u0e3R2RdD/Im5YGetsTxOL2vm8oUpURSU1gRVfcWQUUrL6yuq8jr
Ky2tTvaNA35HvUrxi3fwvw01GVQ/L55elakc1TMPhMG/4WWyQX5vzvm0HD/8Kt8BvFlQBKfdiF8T
B4zhBgnMW6osjG9gUFZD5raAJfH3On7cY2OXxMyknStmLrsIWblAIHtqH4FpUzToLQFpCQ3ZSMFi
5aUfOHTfDZ+RXTn0UbiRzHqydh0bTBcsStNrXznq7E1afm/4WjIinz53I6kGWT9aBgRG75kJ86bO
r8QxH9wAEU3qxO1VSRHtoGlE/N413PWkmMBhFGyX9DBkQDPQ+7bFEe8hVihb8Km3tgMPSiLNcGU1
0Dt9s+878nCeMX8/RJWUkB9MW5F56rlMZ5xicvCLi/Xz0ulPpjt5k52oV8Ks76djy+ri0mO45vE9
qv6e+pi+2/kcKVZHKRap8hEU441aZKhyxC0C12HZqBPldZ7sPikzHnjJ2IpbDI1ZwjcLXEAwEI2X
BM25SNU7SsuRJPpnyModM31jP5jyP60hmNWakSk6ZkjibiMR3MhaMI4/lvj2kAzY5VYuV6SM4COQ
l1q0Mnik8lrWpjz3NqFx1FuihOG2cn6YXJW6SxORPLV9LlJg2Gy9gJZDeWn0u1kcngZI33wTG7jp
4Njlb/2rCjHSU4FeZVdXlq9+xFjPUdIrJmrycQ1BlIojBTB6QQIbUrQD4x0w4/lHty5Bxnn/6tk1
HcUfYdAqPYy6jjujtA4FMuSgHH3n7+Rbhvk7qeG2Zb/0VrMf/cKR5V8s0EQ2aORbJ3ler29FRMeQ
qVceF/eHO5wvEppRxRmIGOGaGx57yvqJizAzzRNu7Kaj3KpebjZ2ijNdPO7prYoc9uF7SB4CSfKu
1tqNj7ZhtQBDvhGtJb2jgOpJ8Z7ZlFsgG0CMvYb440QZNlvuWNFJ9hupEZy+Uu76vOiyqPydNDJo
R0A/HkVPFnSwkJH6kfgXb4KZ7FHZ4rUDHMPBcpJn9JFZc2FSvb9V+brN/5bJQWvFTZdpiWHaNyEN
1V1HLYeks6CoUewh3QI+ZEbSNzdPJtOKfiEFG2UAtBaF561sG0ifL4xtPQq1p1mpP+rN7p3anoiw
QUIcNHrPzW6kH53KqpnZN82nx6X+LgpCbFWpYIugxhyCIutspJoioDwdWTsK7vYvM0eme9qMiC8+
OteXsrmMop8JsjhvnYMb3hwCMc8SUMN1kd0Oj1d2krIpsacrtFvOJGvYfj4qn8oiHhI9U06Hmwad
sKziiXTzYE+VBkBE1zAM0lIURh6OqTT9LkANJ6qwRMX925TtUYNQ3iuHLgpPyS9dOGOb0X/xb7Jx
LN3QNgao/uRDvfV8fGuxJkCMUpMTngGZFzIG626zxhpTB+zRYg89N1PgW26dWteTZmK9FhHPzdFI
cExHg30RU7q2WrwoZXsQJhsJCJU4VanX3SINbb4bRQtt7e/ngUL+j1zyFEL/A5Ga1j3rpzLJQUdy
87cpcXMciGYgsVXmnyyqIbW3IreaZpczR8ik3w1ZNgiygzYd064FXXiUIyEwkUg7z/BmKYWWI/9o
gc0v8fS78stgCLGMowe8PmaqLkq4Iyy/YuYwdWQ+ac25WnJFeMprnkzZ24W9ua46ZX9D31KJd63d
SdrOS9PY8xqGdmCKG64VH5Eld2ErUUd7ejDB+uEhCZF5anEThO7OAXfrf5ktBuqx3RRpDqtX+zW2
d9DUV5Un+2BYiLtyuYg+OoI4dw0okFXvWn9WR7w6SyheFloq2LWlAw2jcnfzcwPtqPMYdCu/RNXU
LIjA0hGEqtxBTFbq9SOcmxR1s+xhRRN06o3wDCEmD3sEkGSwtUBY/sq8u236xTCGT4LU65O6PH7x
3xr1R/NflvNB4MptPAryODLVlTA/iq20YLAf3B2gEfwCF0xF7aofqORJihS8X3MTmqWJ8bgqi9kB
zViGI43zT0uuIFnuBZ5XAIXrlcWxO0T8De3r/QGDbh8CDKfUnVOq3TJydBhGPzfC8t08NCr0t1nh
8jOxHV7w3gqzZM7F91/oq64XEOhcgizAZ8SHzxJYbuH1cBEEyk7esw9cxYnX7Bo5+p1+kKUZaDtl
jZMWNCJsxIGpaRAqY9a7dmOWz7FufxgXkGC0j2f0YRpSERQluULlBsZvkC+iQ05HBrssqLR+Hmjp
bdZe/66pJ5NDVmwtx9JGJRDWc1Wb1K8BQdzL0evSQ2PT32W29jDlwrRIlXqTUu+rkU2FANT7z+xa
aCw8JWgeQxoemI9n4IW8+jjO5gckwDcKQcmG7i7v50e58rwlVKWS93iVSitwg4B9SmFrRz3KFUdW
T+u7R0QGQDGTp9c3K3niDAfY9C+ltVt04YpT2Uqe+3nkJpGgtL8d6gvGbnS0TlSp1wVHNMfEOzAQ
J91katzKDJpAguLFIkNgnZSzpIMonXA+4sCvXgBwAY+2KzOKd0ZzeS54sq5pZQ3xiVPAB4UGjgBK
iukaI+og3N8XPonAfb2u2qJ5WM71mLMy2xnsagiVFUrYv9OHxhqewCTnnTq+yLyFtbB7QwIARGP1
d2/EFCv1T0uYxcXwgLKXXdU5/XJEy/0E40fOuwDlm79zNkeRUJfq3NYjrOxl5RH0e4rUL99lwul1
sdGqp1OMC0d3B5SIiXXul2DOAB7B6I/eUfoPiyo8lNOIn55fpc84kB+rAQ5u+CRObPQFkn9rriP8
ExEKwim5kRAUPQRCxzcY+uCSkv4CICTkBFJFsvLY02NJSu7Zop4MOq3d6Q+K/iU+yde0XxdkifQr
zrxPG/jLeh7NXSE9oZRUyz1i5+4Gbh1ilH2i9hNVZ3bcYANQqpnctMlj8wHgdhNuVwTEHx+Nlc/N
5+fmTixsPSOdV2bfVJFOd4R0TjPaNXBoUxnbjX2/+Tsy5HHEG1f2lJWmAfG4fj3srcv9CTDWrcxD
m1Bz5kLfLUgAKfpr9GtDArRuPgvNr0GU6+47Z9E89DFp905l+IMr/eYi+m5rLwn1jCBFI9LsupWV
aJAe2qBcCzm8pSUiIff9lNgZisVDGivlrKNCEJiGuAlq/4fLaGEkmzX7wdQYBy+D0s+JFoK+9wiN
fSJPMnb6cHTOuWWuJFrlIPDmq7u7zmbc31ZlVJCUkDup3Qm0QETiBHYn6hvpZ/zanoaA2+OXbxbA
0Cl6IGb4NsRD5KGMM2JY12eMQ97JM/cC42/ydCUkhJvs2KmGRMotUcsvrpR4lx2Gj3AO5+BeEeCI
oE0WfucxTChojCDWsGBahMNf7giJZ+eUrtKI5XZ+csO1AMtqEZdFZlx6gpbYGYLYmxJmYKLj2Q7d
EHmlvGFW4XffLusK8KWRYZ6eLXTcz+gupek74VdoZMRPCYSDqmS2AXmUo7HiboqHfjMMG1lQiYNr
y+LwSQAc5GItOlNt1hq8/cmgnGnTlvmT0PvHFbxtTA6VuXej0QVLib/SNDD26VhfKoI3pNDyt4y2
ahbmWkocH1qTik2I9nr5uArLwrXHEdDrgw0cOrqY64+9vCmWLixqLTleAQvLT5AiqluqzDJ/ta38
hoUdat3kx2kVDhhRJVzxrj5n0XN0zY+02gvujvBJI7j1U+KjfActGa7tFUx+oToh0nJSC7O4LMzo
nazvacNsvpPe5EbcXVY/jo0zD31Q/RwEeuKi+jUyabJ+fH8twvoYkAhCpLSJzj50F9VPTai030J7
g5zB/Q0Uh2F6We00RyxFsMcB1wz366cVz16GJN1jgZc/3bNCVZQw04lirmOokKPoBWyO8U1gCvdN
UlDnemuEdOarsHc2cFA3wnCNInVMFDwmPYfMYooZNmy7BO1xRmvpZQRcFcL2anCRWiyOyLRTIrfC
lOKghh6pjH0y7kSLa15QRhnii3WUjec/YGhqQv4h7f/3YLFdvnyIu7LmkcNXePDUIGAvZ/ZxbVtC
IKO1AVUqC4V6niVjQv5PkRYjW7pq0GiGHcEYX8veQP7vFMNOZhIOUQ8XCprA8UEjemaCt8CWxA0+
Y3zm5Agc3sEmZxw4cwgowZrxSuwoOFxKXPCBEUj4eZkZjsk36u49nD0pYLLiIDbk6EYT1KFT3//n
pat8w5V76SDMkf6XmP8LFlK6Zuq1sKRWQatiFIyjGNysxGFAPgO0Cfx1Xqi9g2F8NuODNccYK4sn
tIEY5jZYucIijWOzX2jhZ1q5Vln8rvWoXci54htNz9hwXMegMYzka2RjqEkK+5CCv/vbZ09w+GVz
QjO6lQyPlQZenjcR2TImH2yYvIWVs1zMBv6vP7eZa0UrQAxusw1JQhFTG1Fe0MeOp4SWNbrNUKoW
AwZIcPrRGlHKq1xcVr+rb2eb506LyZjfFuoCA6UaIMS5FfF9bFCMvxE86IutJ0qm1HnVIomQKsTv
dt/mEOVpUw3OKXKdgGdnJgiS6UPzZFR+8hOc92WvZ5i3VhWFka50XDPXZ5k37qxFrMknE0JnNJZF
1S+2P1fYQpSPecRiHKA//eJTLo9AhVFpLD543/YizAFwMyDkkYfk1E77xOk8eCRcKoocm1aPKVaz
HzdL5lwMrEvA968OI+lszzX+rEUC+RfacQ8jG+b94IdowgutSMlzh8/wFHmBULoAYGz2eAu4yPh8
SUkvAx0/LSqaaPoWl7APomfFYTzB74U8+/zpjdAqG0YcJBECvGJNprSQ6KWF0QoUphDhHZuBEZnx
kEqTvSk2yLoBTW8XeWX7drtmlMhmlU2x7Ueqt36D65+sJOv+K24u436nvVGKv/GooYumgiR2cn6E
CagEJD1rIp3XxeDASbogbA+zAc7BXBkLV3hKl7J3OFb6HfaVNAHFt38ppZF2ek+QRrq6lNtfoSjM
EUFNz7O6DrdhwlHKtdYdcVof1l1ew9hACHS1kgIwbHooHKrnp2S6x/J8R5S1t7IMz9OKwc3U2FGX
WIuNGUr0v/XfrpxuhY1k5w+FWR2vnleUXNmSQwkY8XfIVOtHLm2T+RNNw3Mh+I2SmowOYTXigKYm
2JmCMLtQMUbPRX4M8NHvSgkKNMX2MOnEGrL8GobP/mof6LC2Ug6wQRHyJQVJC2cSbqNafGldiOr3
cS2M0lhTUROQtNBitfpg+pK7jluIM+I5NLmhUSe1N6MdZZQkwM8lOWjATVywjWbmaPdLmgL58RQx
kWT5VBAa44bTLbPq/o764QugSNJfk/zXZOPfZuQvct1nHk5hxUdrhf5nYUl5e4WbzSOYjv5jZNDN
B/wHWMyZEf1TWRsO4k/foS23s5WKBuYedixGFPNRdXknVMnJv9kcmXFkWiH8GqpTim/TgRX2+tns
eSfrMF/0qlsWVLJ1dwPYR6FaXD4ls+nh5eeL/j6VTVmYvWnU3sV4cuRHUakLV28Dig5CG2/CgS+G
Ju8qxPuHFl4/kkUlmD7eTEuQcAEQV3+lBTSuhR2Dbkhjzg2LnaBUyCm4n8dBvtQNIku0YXoiwtKS
zQ0xjXOuz7GGOBZ4zyjBTk9YTkSYWj5vLfG5BsZ+ise9qSlougIFoeVyd7HDqVZlTWoyP/jchLSk
eiTgRjprCfq8H3oC2OujOe+DDAUEOFRNQdrafNgyw/xSvk6ANGy/FW30W9TnF3OS2fxyaTLZjWnH
HsbALDrq+cpzOQq/rSUh9TL53CgNbC8EBxPShLssDk/9FbXm/iXRcspsI7OtjJYrboLlHQ/JVuNZ
91gWZTHsdRSQtUMwQb/UoHiyFNe5TpKLdWbnCdkilYVYpH+P6ELDNkvSA86QG9r3rU0+7skgQ34y
AQVGA8QPUaKP91dSvKG0DC+L4zI+q5V85TwF8lxBtiZz5Ty/93kjbaUGAJbl72Cwab1xwCg/7unp
k541omi5r/CxaHdLzOlyp94qEJ9IO8vT1asMwyNDtXACRZr0bkLsptTlwVCqf0WK3GXkZuvKO6y7
ZutSp0pyi2iEhwdYrz93Wqrrfsuptw20mMrGBeepfCVjQoEZOETd7/xs8utMxyEWWEK138VqAbBo
JPWJ7gF8jaLbT42kFcqvqBXjl8j04plU9Cuv76zSMUCYVUsi7sJw6/wMBV9SAXCOk2oY6sjcvW8S
K8d5GAIqvkA2ta9p4ruRtjxDzluKM3LwNYocmAXmalfRco1sfWlLqz3m+Cn5YqmbDMOBXEvXHWxj
cWpI5dU6wclAE0WFX5/qp7anovZjUZmyZh9a7tvI8PnBXmQcri9Z0hSns5QKhDlXV5uwDYLwRSvX
ygnzTC4+u5zkkVJKc5PW4WkwbpPU4KRfu2AcpmpWT1Rz6///t4JgaOV0z5B3EMzwpTv4uyL8QhFe
ThbIbtISBvjEQGpvr496pcr6Oe5H+uv8cqXZ2dSG7wBTq9SKB8d+rWrboKp9l8Asjm0nd1RA8/Kq
fn3WMb9NxtjB2775BOtdcAx+LTOB3QjYSYoexx5RcrnuOkarT2eabgPsqSFAhOwBlJtzpQD5seQ3
OQHl3gpAWilIJPIRxw/BdfuNtipbWffmauxFiHVGYetPpKv+TEVsiWTN2zLvo1BuFiMTaj61954q
3toE5IF88zIvRRpHBphzeCl6X4GTABo1Jg2ihW0DBUBlLUGwjc86jz8/+1m+9lLt0/VSz17MVLaZ
rvVaRZN066rnB1FsE2EP2YKnyEbK8WmFHXImEdwIP8nDdK9MkK8hTs2ExHIdb4HDLru9XzgTp9Br
DNpQUP9dPCqd7TA0Pu0FCHKUy4ecmAiydLdvn0g5RNtPaMCpFbvHY+8J34WCr5hbFkfSxFMYVKVz
/7zErfFGOMv0zhCXhqhxEsMusAPHXId/KQfKbDFJfJmrnAEtE9K00ksiwfNnJLUSmKWVx07iNaLo
KmuTVuA0Yyp0HdrhVBtkgyv/bCLGS2D6S3vc8uXP01gXpGnqRxW5B0YpCIdqjvnCLK5U5IT8RnG+
B2CjL28vnFbAIKCKyh/uStrrrLp//8lC0K505vb5xeuczK3zs72GvgyFkSjt2dwfUVPJfpdfji1Y
1eca+pLnPQ3oHbjxJ/xoIuWLMDDz8kwLGOWhqpx3kumhIH3vYk8B3wxZlF9Crbm6phOw0RENV4Ky
3ldXyataqPLMT1wkErOzTpWKvkEFGy1wjinn6ZzOW8Gj8iIPlfB1VmD/60JfaGj8M0wTbOzwDnBB
aBJRHDg55wFrJnUEbGswHnPFoejDYuZMT//xZRVtxWSH8ygUuFKM786ERgDLNjX5wIrrAwzP5vkh
h7BIgah6Ev6LCo7tfA4SAhbrwxjUeIaVqNFi/dAe8G/aViUP7Tp5IVtC/Wp5MoyateICxqhzcYwg
qYYt5536qr4+w8JGldT4y1wu2Cgh2cwN07kRp6GNYYifpGA72Q7ndb+Na/+C6Xrh3Tpgf+XQuzr5
6ee50SXPk6qPTnG7sWjVG3CDBA5Lx+vZXjQLTZsYc8ELJPSvuL4QGy67kZao5wSxhsekBrklPmWI
Vu70NPg7pZsTyHwR5HfBP2FMQn0wj1xiv8iNIx/oNGxEoGRLe0QA30Kzmwh/+YoCfia+uPCqS86B
jEwPXxlzxqid4xYa1it1Ezv8P4woCgWdsnc61nFprViPBxys5525nnfjjDYCYCJsPz2QpFuDHYDR
5PTxdcll97auRimh64E+6oQwBMFt1HgtPcLN/v+g0veF+JptdQQObpCKMqHTQHF8PdVSVZhb5BCd
UOVfLnh3Mp0guvA+DNJhsWMwwBULkNGcVl9DnTrGtiGECIsb3BlfQM2q/QWSUPf2xTLIfn9EuXi6
aHr0cuFWyKJIGMOzhc3nqTsOHg0gOMdK6lAVh3KKBsVup3JtaKE17dBS8a2sN2nIgxB7G9/ukT4j
mF7BogPOwhBG5kT8TOIJBKWf8lhOUgLh2bOU6KJ5EF62ZhGpUfVMkaWfszjeOlQkwJWhWVztaSnt
8pcyaHMRjoMFR+vxwal+uLo9ZgEMeIRIG1n8OBvxWDNAmsxdkzQczTei/iqtB95tWXH/kkOdMcnM
FeSQnfPIIFadkNOEZq2Ssa4pOJqwwkDPxD1N4FzGO4i/CI2gEvvDYSpdux7t/R2+7129QF+plV0v
cfr9FjxcupAcVEiKMIc4riZjwLDB9xg8dlhoIchMrVzdGSyCRuw5r7SEuOhttmkqQ8R+xMzBXmhy
rxXciQr2VE1I6my4Lxhe3NfdGa7HljqDYEhpZmiyBMxF5zj9n7zTKYVov+Il+311ylkWBj9F6LUi
SSIjhjXIB2njn+HARR45SsfD6BOtI/4bs9kwVypWWW4sDpLf7Q7EYQO89jtEPe1/n0hGOAg9ocrS
E1RarUaiwiHaFWGe1xgWAeq6Vg2ZDj2VJGg0xvkrFzjbb4LbVsZdlkPUz60PXJ6fR75Xv8SM87Qr
m19H9XrCB5FQnnzvS0o4xAcPs2XYohxFec1v8WLxBsNM9NsBpzSFyDo+An7agcIYu9quTScdSUvw
3QJaTIIBfkkrjj1+CFXPW8Zi1L7kICj7+k13zRYAQyJdJorrlmyAHSzoB6mF8faO+VD+hwVjuSFN
9+avt+WkHOWaUZDNPhf26LZiZ5KRDVHFh/kPxyOr+otsQ51kKYQjV6hRJCxLndLC+CuH71Y2q6Ll
Z9KfrMP5TSezYKE45NumAzAqznlbbLFOK6mWRdDjZQEB9JSd7ujjRkMdMRBVUWPYoAR/EPV236sZ
EUqZpAP62/uAf46QkU8Xisf9IXL4WgLNhVXve6gNW8OscpJGGB+1bOv7wZ8WD1eX5sTzaTvBSM6l
eeiA+JZa0t3RvevBfXE0vXxJf/hx0zwCCjZTkhsO9GgLC4rxJGFkFkcup8/731rjW5qiKlRnupHa
0KUshmC9p7PA5bOU+uacG5WON5pyi8XKAp3ZQRtqFLmcfMXtAfbs/NKywu3p4vAk9m9U7Vj5fnEQ
aAmEV0hdFfFc8gKeE9GexAtuGaB0fEH+rV4mM3SHOo/jaYWp/ExaBcXnRRlEshdQHFRY2n6aHtrm
b15Fiw7tvfTVjqOuPhO0tDgR1ntG7/iP3JJGz+WhBxXD02tkJ4eIbzgqYB4FILr3j5rWCsenHBcP
5oPw4yxvOdSyuy0u5Y1bN0bC6wXjgyQNglhFro2WxPIOQfLB3mwrSzT0mpe/wIQDZTTLNPDq5PZA
S7f5SKNG5T3+oOAklXLPwd1xWnDyCknVecrBUmigmt2KQ+fEt/D89anMT2FqeyJz7IxvC2qmLLSn
Xkw39P9yfkGfPRJZafCym1FZIn6yJVaehdibj2QrJIAn6tUgRPawKztpXV06jU9QZgC9fMcLugAC
c05ZAzXa8LQytVHvqA0yMmfrQ8ytdlb/chOJSNN6dpsZRCam2vGl754+8XWZbq3XlPQm3f1gd/CA
pKRkpB//kAruvlFG6DnuCoqUdKYcKypkgHc2w9dXUqH+p706SDdyHIYSJyakagh9KyhuZ2thplk4
N1gcNuZWSnlemdVDJ4MiUhiqW4Nk3fd2hkTN/9NwNtA7lwRMeFJ72UTm2CFa3GE9HPTmH5w6MxQk
pYImO3uRqz2KsKyRc7M+VuVJy8WEQplqsXTQ2vbmDVSZkLCxVkK2f5f0776uAHQra2pO2LTvFg5j
K0Jc64MP0tMyg+h1CnvO5Ns2rjDNb1QW5Rw+LH0O20w17epUzbVwQjbGG2NdzEJKnTGqGPB/rxqJ
FYu5LxZeH2dLr2FTVG8x3fEbj8C4nUIhr/Q6zjZ7azNGKCUFtwlTVQPCn49iwuevEdrxEeoQ38WR
IClcI/Ri/cyCTSJuOYTFOd0HiGyceVw6PqKnuYjjfGMHUE2juE8YJlU/PCDjKdKcvZhWCHRLAdA8
tSKqkEzzsmzj0inFMMyz3B7lzvdUoVHylEKos5ZL6LIDxY0+qNvU9IsRVRjDEdyruEyG7GqQmR+Z
YMeG6DIIF9aGGHG7akXGkSzK1+Of3rTiWq2Yp/6qdxVF2zqCIy3oAzvK59wyXlE/EF03GEwO0879
+Yuwn5mu+ldVsYsGF3YifR9SFpXpd7ePCm/vdRpLMAsnTf7x4EYrqDSOK3wlBc0np9Ji4AIzrYrz
1ZeUBdCQTWgSXJD8vNWi2yV9QHomThIkyvGM149gkuMPqtciq51Jj6mXnxAKJElocyZpNCq6DtU4
lw8WoiBoid0HbxGjGi40i3qbD/ZNJT5e0cMl0cfcyBKnriFIenMgDMT0LoKWp1iw3ONEccOV8fHt
BoD7KoS+bVhjDZIappdO/S2uRt1PhgenYW4lYX1254HS3oyKLNFOi4QDxeyCsMCDU6n0YEgj7Yxo
KSO1crc1zGCG+9JZ42JRovdA5jUGlqQG4TdgvZH03VfqpHkSDVk+Mp65Xq+O/24W5tG0aidD7n36
QUglx87Be5s+c5UIrpbE4sACwujGGdQXummpogGdvdlEYAOeQ5R8eriy6gETR5j/fAgL62J1aISI
gDlLRyS2zlgEwaC+2KKWd8MFO5Yv+UBjqB85pQ7AibUgOHBX4Knc/oQoOLymqBBjLIK4hBUAyHHi
gPAEiWHzfN0gqhOaZZTeGbtPwZ2yJcGuSF2A4dy8GKU1HOy/C0MYLTau2PfbGEbRX3qAcldJJyij
VOSXWlMqV3KpQFiJZfr0s10Z95zrTpdQRgGkKnGaXa01YhdetLpwQyIA7s5h9Q4gfBAleVkrYPtN
mo8ji7iocQCrFUaybTOjOsUjbiK/HlfaQAtlQrVzl6bupjhLKsAENhjHXXAS8jvbG7xd/ci2/D3r
O/DdLmAQja2RPUGtoR7oNWP9c8aWdAad65a3fezUb33vx0V9OeoNpN15pC8oU6MP9tqkyZLQwYem
AkGJ6tgwZ3JBGYvUR52WBPqgFE+HRx/FHhbg1h/7jf3LgvhQOmn5z2S9D/baR/54z2nXbgLSy3Q5
W29NdXh0TNPc4nMGnmJvF1M+LurzEyo7A4hti1EmGZh9ossiorkjra6Q3uKSkeTBJZUo2cIgXr56
r2XmH0d2WZxs6f760sQX6O2kR0GfjByOpENcPOEEjIPUJ0M4TFU2SA/TdpQDz3WoTkWxPT5MxScb
Cn41xDEd7CvqdxNECDMaLJhLSeByUQtcFcxEiKqEedHlolrs/POOX8HDy93xzzYJGx4ZhlVEpD7B
4KWjCHs/YbNIXyVTfPz92khRVsNvgRmTZldMOWadxyDhO6Oxrug41FtD3XdU7QuaKH1wlCaRFx1U
KHYblEF+dgt+wSKtcS8dSCuAZ/UG3DjOFXgwze9v5B8N5/bKGK4ZGffqk35Aqov3+7cDlB588Obg
D1VjfbsXiaFQeLvV60ePiEFH3NUQTfX6L1Uolv8+TfCw159/8zxurcn9ssMR4Zr8nPzLR4xjzvT0
HM7FZ7f4yQUYJzoavRihhbZ2g3bTTAJKQ4L5G9Kc92/Vifl3oQJnWnq/p7qtC1uTBcTqnze06wer
iesjOeq8P8XJCrstNpBDsi9l6jnJsT/ZNeWmBKHHHjCEGEvNlncDuZZBgWPRxuiG9nOY6HS5dxxC
woMIzAqXWW0SyPJ73XMwGpPQLBmcjHtZQi8ggiQ4M5sZ6j2a+LRWIIAt47J1Cuq8U2WUTa70L7rn
G/SiAJ3UD0pr5B8zhuLnRPvh5/f3oscbPzXGAuXZ+9zEPNhkLYHtso7PvC3z/RemuA1FHzewn3Oa
njCTyQhU6XqCeAVlUUh0AHP/LPQRZfB19u5GxQyRgbqxhGN8MJHMqw1pTvHuBCBMui6oEa7OxDu7
+Nhyf6xM60FbFvckBux9XJviIS7+uyhhajERW2vKVx7K0I50qS3JI2Q0Es9WS87+tYwYbeSGMEow
7fMXk/rt6rKx4sSLzIUOqRkrG/+wZgHJWBYM6Mg68PJruDI8XMiOVU72aJyRjV+0Xt6R6NhapmY0
V7vxXCuGssxbmXkTlA5sJGqJoKkYWtMm16JpcGHxxw52G4q3hNSnLeESpYhcFnjVFqzvpXN2x5s0
ffZPYwI6MYOIeqsd4Bc+F0nQ9M4ykYHRdMcGbhZ1/CrO3Zg+in5gjUUknnbNYjYxsnvqbMSaluhK
gob5W1hQB093JemD9wX1ei0XSN9mMKQZmzkZxSZ9SNFgFT6I5Id6fi5tLN5QwI4BcEvpQnKCvvWX
am0SYtr39ssn0N2FKb5s6QKYqaR6M6AWQMKnKdTdQBYwVUR8Q69TetMJ3MA0lK0sCwgSk5eWqlk/
4hQ9g6YQN/Uk2Nv7mPFpfUW0m6ccVowrapEEKGjyCiQ4/SHkQNWutTnZ/dxABFt9QZ6OV2s7Jb+s
X8NHn4aQLz8N1VJaOVkfsvoFs2rvNHzxjKhJ0k5SIwoKcCIUqWZkbRQZtC4iiSG3YLC46bZ/jXxz
X6pLILJJFuJRIWPn7hHeqXeYq4Om4DDiujN7EatOnF8tFtNkNzgawq0v9RYbXlnMguTJSXB8roSf
jXYAvnl1igavf3tIwMyV72Sqer9Qp97Re7l7DeSiYhWWvVLZl52J04vCL/tjeCXLstmrh9IK3jpx
C72eunQYu9PjgwMTZQnnrHjOfDFpLwBnoefGRq0GWj0WYBxzEW+b190ncFrzNIufirue+U73yvVv
2s5aRuZpkx1JK8ehAHCouVPeKMqzA6ZIPMArzpNDkWcIX61lQzwJHdTYJkrk5f/Y4SBpwqqozkXM
1/aINFEJ6dKM86nkuOFAiDoC5nYoZI2csjRykRk+MEO/wR7Da19yRFCQ/rgzF1WTKHd/bXVowLzZ
B6cOs4LyUHZFhu31gkmq9Ca5R8wjUrvJ/KbWWTNjc52cAlZ7wBcZ6NMmHvCtqyCLqbxeuWZ+YbAT
OwOWZFFN9EVooiquO3BvVpa3SAtK2LwLsao1zs45+4zg9Rmay8qQsQHlaXvkrcXcQSq8yhvWY+w1
vZC23+xXXx67DdcxCn+dHGnyZF7b9Mi5LDVw2fxKSpc1iKZbUK4/WFqx+LI3o8g8VHeJGkDhzuEQ
0D74RwjIGNfXrumIYkzSAOEtDBycd/vxHpuojIP/XLQZ1gxKLFpPT4Ue2A2nf4cs5jb3JQWQTkS5
mnSijwJrxwavN79o8vf9XpgiXMl1m/ViyeFj7UYLzV6fEFGhCFDOcUFuEVqEQwTc1Vr/efDUgE0Z
6nshaF9iBr3ZaUY4O5LYzV8w6nnG6YT85/cscWdgJrGD7GfWeuSo6tcf8FIx/zgt6SOowEmttIK7
ohv6JViVq6z1OAIUAxggz0CFe1gWN1Dn+u4dimioL2UzMz4b8TYks4+Wvq4Ym047L+/d7lc4jC1N
HbJcVRzvazcp9USdip8SuMwXXKxBOVNU+lpXuGIsAR0WBglVInE1qJCjU1H+jJgFwv0sBOm5k28B
YzCJo7uouoMDTnuC/FwDZCgYs4oS7897CdzqBHyTxgCFdooqIZRO1fj9+5Hiu6nA4godXhz3U58g
ySOThijpGjIEREcjBRnGiDTUxTkzYF/bR0bG+re7GdoqXa/wYtwyWO0N2d0aRxvDLEXL/XRKFCb2
c7TKf1iieHwc/sjGUmMW7mhEotdWmnkPB1Abbhu1JpWXq5r4W4ldo7XXXEEJWKbXCL24zTTsiugf
88pIKdWsOVY8n+tFze4RqbG6hpZi8PtZ/z6p1pFZDPdk57M6A8UVC97mXuOeZd0dMcFQJg045qQd
nbpgFFf1Rp99EPn4F0Ij1BnBZBaefWBRS9DQYfDCDQi97r6L/UO8kRQuDCwIMh9xJKTOM206lJH0
T7xZw/Vq72dbDlmZBoriyD7IQrg8Ck2+V7I9bu57VL3Cb7nUw31bC5UO1E0HoSgiNKUIpGkGzdTA
jqC4cTWcKWU4nXiVa18VcoModxENQN6UnF31oxi9R6ZTaoLW10xjMsqWB1lP53klQ47eWb+vHq7U
eLJPcKZq6iAf2vi0kW/a7jsPPUIZEanPXebDlIUv+GmtggGTozoAq7oVVlBCyShJeDPK+C31Jp2l
oCsgCt/+rh1w6gPgBVVP8Kx4pH4g43zmbG7Q+SscXeteS1yxCbd35bQYT0QvGJiDbglON1NUX55x
7tso7soI08ro828JLC9JOpDombn1jm7qDT4VdIy6Zpw6r4HQP8ISMhWdt5/sp8aIU+WVvGe4B5RZ
/05HaIirj3PEDlSDl7UJ2cxQEhRct2GYLprRWXzD72Zp2k1RLphqp5i6LLpi2stCiulNtfV/se5T
GEJpeB+WKTonZItit1yoaj1UOAQ/6Qt9F10AB6JUSFtHw6t0GgjFu5kErljAsbswTso6OPkK6Trz
JS+H1Y4W6GxgoF2SrhH6i+4t72YAB3VnnaPsthS1uXen83gHFjebCSDPGYlndQ38VA1usPTCnzMj
NiOStc24BOq4r1qlqjHRbfjRAylOb9Psw8xoZ+ZqwTsExNv2bXxaaxOTyHzavk/qteVw5wFYqOtJ
NnnPa7uaqYZeklL6qXoLrp/xj/0kaNrq6E1nuRECw5yvrCMBoVysmySD+SI8dJn6qOkxjX6w12c8
ehrzY+eF0ARMN7fcnzTR9L/NvSsGjOtKo1kIl/A1QZf5RtAdobdWRWOgL6wcl6zC5ItLLt4KuP1l
oQtVwLIG7PPS3PlNnZHlT1HllzfmsZK3s6uTgGBC0Or8qrxuSwwQJPZ4pQcjrQhkswxTzvBuzIPQ
j1bTCIUp4C1nNPJX7gBRVvawQiv3ThVR+7cHBxcDYGBkUzF747F5Ia1lHIpMwO6Xon2j83tu7Q4+
gOl70DmTre7jIpvTWhb9Dd3T+APL58ovmc+kg2Q2Q53mKqtcRcXSZYba26Z2vZDMIDnbzUeIK5No
OiLJ/UJ/+WooIvHrlzHyCoJX6CIYlrnlg1K9EyXxSJb1BQQZWqFf9sw9cI7bvRLmfpGa8c1hYIIg
tDKsGYUXAR97I9noSBoQBZsnP509OvKaisaBmgFjP5Vg2ogX1GADEibLhYoK2JVjum4iMprIXf54
X+eaQMJ8MgQMYlUgKV9HMB0e+VbXz58JWBh0Wd5p8KjjLpVXf9EEi/YjeZAW6p3aCOCzchbuObMP
MSv53vBqktJRXCz0tbJ7IDIQITfFoaMlwakTkliG9ZLJBrJxDtEY7sP/CWKpDPdISQhMlauQP8yt
EHw5ScXdfLSg4pw3+qiU73NPpuQF25buttp7u0oIdfyEvjlOy7f4y9kV1GGM+LE1juDbdR19cNK8
vqT0HVMh3kxtYY1/ZSSigCJ1FihCjX/uYQ0v2UR/eDqRXBzy3j5kU/sICql8UrJb5rdVoC0Mm8uX
t89Wr4ZcpxxeLPTmvuhJ0YNRueXa4zIEzZ9uNxCu+ajdos28bIa0aJfcg6usg8qeNqH+hvCd+R8s
qrLYtE0Ht+MAxSGjshyFqvO+fbEcw6RCHPmnjVSJWRdg8NSuYKi5z5OCZ+vs0IlKLNyiRub+VgR3
IbxHD1go7Aijl1/eTyF/egSk03bCRFw6lagaIKRzlTHTsgXiuZtraaxdIAwRks9ATfU6D+3z2I6L
ZhVOG6IF3BLZiKJuDAS8wrqKnpth4navuXcJOu787bgb6kcqNBKVYGhrUq+lRXHhtPSEOCY4Fqxm
Z71TDAToBbnEu6fsdIUuFDsf21y49L1dzp6M4Z+hOirNQzkZUwaqBA8xdgB+7pt2/ttJ88r39zMN
HWR17dE5FSyFYrOkeWCKHGyNLYSKfNgg6j+nseX3ffVH7jMr+WNs96y66OEU1VQMGh6a27uosA9v
W3kAQXkyLj2a3T19XaB1+w5PYp1LQAaMwmKzTNcaPRdEdJmtYMyed0nKoStIvDyfq5rhgwT8JOmv
E9XiIkPl0JcxQObM/0yDr0stUmqBNFj3UzXxGUgXOdoMv8/qQiIJrxS7C9Jx52MbTPHAx+pyHW2d
O5VUMamAP9JbttTEp9FLJzPthTqmsAtHHJoJTcinUxXiVSpTFJxSMOm9b/Z8Ecm/4ADOqr3VzFts
eLgvT8wsQdO8X7+RjdwtrSf1aJRc1ie976fhmOMW7hsThYq7486dbWxKYNqRAl/FhlxuF9OnXGFa
QEdcQz2pQq84y98CWz3DJUbPHEgrgVDcX65XATd1ndBJHhC51DlbPL1pawvWK7/eESF8QgiF8ZyO
RfDi5Bf5svCfDhKo/OSvw3f6qSBnKKDATiulsUg3KWAQVI70cSOjtBNnJImnK1WfM0e13ZlnpMuo
jOM3J3rdIdOyRzsc8Qu5fCMeeM0CUYKeTQJfoJM95r54SwVZJCpZyCEwfDJcPLwrrZcxPBB2Fgze
lJP/dl2TgYIiRFcXTVeHMKSnKL9r7ch3tVCOoOuMPHaPhdSwQf6fKq8/gCkSwjRqOy48QXnF5OYx
ET1jzXMkVq8DLHk3+cOdbH3c9qGZQG/U0YH2cE3W38UX+Nx+AzNb2plcX5SRv7k4hzcm4m3+FQg6
6E8vlI26G4iAdo0W8H8fOeB0pDhXOoM3Pne4tJ0hJuka/1Ws1ArhptIBqtiQVCkRnGGguxWpAAMT
fqES4IOAljAteBNOJqlckOFX8DSBR2uJAYTCNl9UC78ZdAr8cY6egaSOWDg26hEaBmyzeGcLb2Fr
cRG4ChK20RCx4M83gV1iBHlUmaxjSGvId/bBJitgpyB9gNPDWrEDYkBZpFG/iNGRUjim9WuhCLyN
jeJ2ZHcpYrhllWAkno8tQxWcsO9CueOLHwrGJBUvOYSwEElwprJ7Y+EX2c/4ShJ894yT+W4n0yPR
JbqFwUjqm47VRzZbCKFaz+sbCkLAu+bB3EJkyE1RduqqT7ZBCYcMJ7Gpy5VReSkVE5BX2Q2HoAQq
Lgj2Jv2Cf54t0YJYGynvlIfhQYbsaZBpkhtmImQeQxfjMUTYWrU7RHZdTkMimsNR9fpE56VGU5fw
L69OZ4o0u4fiAQmF1vngQrZRAlcGmygssO35kVBk2C6QBj9n3K9d5/frCim/vhPVGiknZpw4I6eh
0U6NfnL6KA4bYTGFuC9xJkixSs4L9vA5FyMBUqmSlYyYsthfz+5qax3DVkx1xVSTvG+fkx5WkLzP
HFYFHSIVh2qh/28dAt/muhZ1ovlGEbIdCbspvv/uY1RuHgsfs2mmrbR5g9u97HFIJfT/1xG6HgT8
mzk/lWGDLdQXXg2oJgIKTFg3lp2Ye9g+BpTuxAjB07tiWsdeSUh+/czw9VnZlTXOmJ+TCIKhlbrM
ofXFlCVVSLiGEkoXTQSqzbRsmYAm7zRohPaOca+zQQZR8gKJ2gk9fP26oRMOIaDVBMJzkK4sFoNa
7jKg33DHgH0R2zZnXbLll7AvgzMRN5RDj/Xf8K4LsxqO2qAQa2Jaul6Z9U2uGD8ZzIDZh9sJ+7Wp
havmkkgdknrcDg+xHtzUPgNctvaoWw0unAGpTGl7HBf/lOZNmj7XIGKEJIUxgUr9pkca6Zi9MNtS
Eme2nE5cZcGo6K2DY3Y/eQYv4csOrkiT4iVvMJiKZ1ndSPyXKJRgf0vL8f9SNIfUbpnLPzisMDWi
HZthn/sLlUfmbYuWo7O7QfVaV4epNQVQyYZkNHs9B5bB4kvACgklAvktwsI3MyNCWFEsghdM92nN
Lc83d5AHfrNhHZe6exbV89mQJx0DTcVBltAUpUbSAydv74fC7sM6djWzV2zYNjYLDuVWjGKLengN
TLNE7W0Pn6uGfYV+k2uAdiM5F9jw6saSak+fKcp2FrDEYPzI52kPSjVSQkejk7XyCrBeqCeScQ0n
Dh8rCehjCN9CdPqSN0bAJPvYFyd9i8oGA/TThDFS2ehsctLxAMEweH2mYyiDsjQRwXWVv8yDbTx9
EtUfWAUkauHnn6l4zAm5iCEedoo5SWxXRwuy4uIZnXvb02odXEmiKRX1TVgB8wGa7R42kGRSY6q7
8QnnTueCWS6HxchjukiyCVKNEeZM2NYIb8DV/byIk17dyrFkHxlpMurWBS/y8kwtWm5CvnJKLFYm
LIlwmlOdv1pmAMJO72q4Z+BKdCANRXsZugweusmRtu1PnHcPKsJxALJaYYKoV6sdc9b+VcplL/MN
4/dJK59KSHjKpUuKegec07ce2Qtx0JKmrrj5wEdXIglomnyquCtJ3pbuYk/4ok2YeVPBGJ7wzWW7
cZUHfkRJTKayDKuofmPlKRxfAgTv2V4NGApLhwvPb1abjpR+/l5p6rCtH84REiS5B8LIeN4ELarY
1Nx6qdNS1Vjm9RM1w/b4TBzSn+GXP8vHMG4kkRICa0fKe+4HSUYoW54IesfrcsgE4wZ7nKjWt3J/
H2vDzxotL9CQN/Wr5RtzvtHtOE4YppCJKidT+RO4F6vJRWYOXJmpE+NlvT5Pe9uFFhqNPotHnZp7
EeG/jS1Lp5sxmzagGyBbZGjyhDyNSlCLU6iKHKlZAU13nYIRrxVO6dE4kOPT3F3SirfWP0wvSNB1
nGtoNTbdOtwsC+eoye1Ns9dn+i7PiR+YXWCQGJdqv9vsRJQlmdEJ9o43CYnXCt/KKq70DA0lG8oP
lS8zFAjKznclfGcQR+ch2yEZtXwohdHqIu7769TFBwEq3DSOCuoWMEREsUwlB9HHaiJwiCMFVqOA
RtDm3V7bDh8gZgYk2FDYVaMyc48qEh20At8GUZF+AUmemaEhZuItCJoGDRnMLcmv1HC7Y/iuUw+k
ldY0sI/ISodOcCYlZg49h+AIdh67e67AzzqXUSS9+Mt9qV+pABk1FTNz27B7GaSG+wDIGtryeYcn
mV0VRPoAv3pK2PuepZl8EwL9IatkcHyv/v3WLZEGGsnl5BfDXfUMo+bZkaN02ZmgZW+QxLJm5MJy
DLYJIeioYccuZtcBgFox6iQARIY9V274mla13IkUjZf3/hN+c8yJcbAgOK0G9krb8WvGsB0cI3et
+dQRzucu2Iq72FfP6PTIse6do1IPwg8eD4a2XjtVQI66SDH3nIykqttbbTukaZ6chWpubN3Lznmx
+i3cc2Aqpzxno3skjb6uzAx/gNsS6QIxYZhk5SUoDv7aUc3RKOVm8GKpEXDsI65XG6bRtNRxCgfD
vsc6fphOh95+8hDjTQKU1P2E5zKFBfqqm1LcmGnkq/Nnsc54EUoeBYt2Dk+0lG+EjkezdfcTPjKk
yF1bbKLrKpakziNpkFKVNqOG5bYcbm05tr4fa1qUogNUKeaV4lW5Q8vJUlv7ZwSpDUILzxL3AVsu
be3doGVVUQDZKHooVhvp48m0if5QnAlri1iDQJ1H0r5IjENHU7EmVVr9FqPH4V6LLIgJeYCp8Bfx
7E058d3j7GIKRMEXAkZ9dXHoCvcHtcESeAOc5Vv9OEgsfVTB2J+qE5UgHf1XlPLOmdKr9BBf2cmJ
AbAis631iJtrWnavBT1F493r/kw9KhWvR6IAYO656ERD5yRWOp3Qu3ffN3ok/7uytXVXbIWmuMKB
ZCZTGRagNuIdLvsoOxmtD1bdXehqicujZn1wVLJCMUn9RPrmNGPXRziXpAYuMQA062pKCvWL2dwj
PmqXMgcHtCQJgyj5C31kYzrCnQLRJ4XqwUsg72RZmP2Qn6r6KSi7zQDF+DKMWIQ6h6NCuzSypqZJ
pRXcs6W2BIIqIIfSRjWErhPNgIYGP0Kd78ytHWTWYBkwbnAr0jB22tN7ttc7NEpcsQSqm4OafngS
geJ88cAJsqKMJFDv7VtFHecDffPI+1f7vu5ux51ChdTqmJYd1iB9SUIWVLNgmnaemHj45zq2KEif
OJgKgz0klRwAmPlJlEb2Tqea/vBBYpMywKYZwTPc2O1YrUlJwgn7fo55jWYeUW0ZialTE47S7kfc
Qt6mj+9fb5r7c/U7ToXWtjyi7WtC+gI8QV5mGj0mx+CxVVgQk6ShBidZVdWAOICD7jHS/AA8A/Pv
uVBOvQXrBUWxDC+5NpM1Aigc1oyOh6riBQogbzhuRetl5SonCfokU2YLDVoEWverpKRnSPPbyxKo
kZk+6RrtovOBkEASc0HQ2GHT78RM06m9Tm/uuvhomh9j4Zm0MlKsKphrY22OWx3I3+qqqtoywDFN
z8sf6u7w1PYK3kjOCKET99lGI+IU5+1op4vjfhD/1VRA5y3GlUvTx6QShA0Mk7XZX9vykK7P1KYF
/LGp1cXWN308xhbX8cLaLRhp494C2xB0h50uXmP3fJqnopmtEeLcU2PFhqbM7ZDpAF6eN3hh3v2/
mPcMnkVVCIfhRAVmWAjQwyD9Dhsk3N0EAJcSCfss+ODZaaIjBKJ9bH4zQCEH96UWGsUF9bY1Vu6O
NtcgIx1EsNxR+/xmUuziOv2U15+LGCp850hpZtfj+RCvMk27pfSCtom02dPRU7lF/rNDhwX4bN/x
2uq94N6sYEoh6ZFL58H5XYpM8rsej/VEk+8BhefAY3OOstnMXb3poOalIK/enGBFV3HYGue8zADP
e08ZhqQuIZMeD9/FJzfaxdksdD8b5PH3BKADRVI8x/Rafk2VhAph5+1U8hLdBtUy/51euBa5jNrl
gy7bj+e9OW1J9rSTfSRqwOhuiTqcxVoDq3D8li4GBGHB/jdGMmSlgZ9VJgu8l3/hPk5VrUEU3hwa
RLqAQCyIKflB/9U4Q9L+qchLfEFupeuSKa+1YgVztgarVaqMJ2O+HBEBFCvT9cjLu2wZCh0NaMyn
mbYHZQhXGKl2rWHXlqhSUS0r6YqEKryLfusDJ05e/NV6XhHxAiz1SSnKIqeyEXdXk35tJSl+Ntha
Mt32V/GuApzpHcUdpAFYbg1g1ZhCGWZ7Hkx4tpnF+WVD0osCqaxoQvDQ08KjfexEd+ABMY2KMRcB
OH4aYCb9ytoXaUsR1R+RiTjx7AGY3+IuXv5Q45KAOVKxDnM0jYfv7YxcbTIu1w37ThvtN22FB1VA
rD4Fj1jtpv06riaGV2EBQ0OAeyzDmsvYbREghhX+pWDCR67knl91aoOOWRzciYpMfoJh9QnS6e3K
uR3GSYUf6zuEh9zKL+gol///oI+Su43aC0UMtNqSRPoilHfZ6hYQt2XS9KR36f17HVy2x4Xl8yXb
HMcIZZWKCvBgjkVRjUPHqW//ZqpI6eQaKYV+yykumJD1ofu91Tv93DXQWcxBgdffIYnuMzrZtMhY
yMzuXMOMvcIurLhgZar2etGWI6L5FRrt8IWgenlXHNWoxnGHVQ59VbCqI1hS7MNta/XNBIgwGz7Y
FpujcUMHSLfc4lR+pYZQ3QdH+d+sBPjsPhryEflXSW6hL2Ye18ydS8YNM45qvFKEt4uxky/ChEh3
ZIZvKDPJtUXDWLN+PMQETo9PoCyYIL620YqHGnAZtCrSNmGbhjxbIHVUVhxgcrZlhJ+Rmrv20JS3
K4WbfITv+l8EpU5qrZipV+Z8KLYJdUM+XFzOuBB+U3q2SBEsdjuREsMuMNSnnpEajNJV0jqrB5VT
nWk4vpFqsdAihpBZduUPif+Gn7RauJ54u+EU5L2GiCw7sQH81dQz9V8Z3+QHio7n0raGP97ZQGjU
JIHzqqn+ppW+so29tLdq/RyiLnsv46ui9q0wqqj4nGC2YJiOpPzn5y8dMRrYDQqoO5vobiCdPOui
mZXEH48Eyzgd2Lmb1MwES9QzFbccFfnxL4ZVoSRIzvr2bWJwexCHAUBt8Pl4DEINpnVUGz7ww+I5
mqVdbsTVZX+NTx9oY3oY2DLe1yuf7kvTQ57ueMUS9UP/uD/XqjSr16YnPFTY5Uuw32LcZM1aMCjb
s5MlAwt06yadaLwQUzg9JPswJ1YxctB8Sep6gf2F9ltbZht4IBIe5lj9TcfmTHS7MbI8H0f6CQXB
gzvC/3+CgGMOCyXZYfCY8KViG5qKltVXDFa5wIg2MjaOlaBuBzIyua8cQuJfj/ZvLVujarADFq9G
lVf9qZ9g2o4gb0RQwY7AA/lI7vpoHisTyBHLvQ4xkRwlXUTDXPdD+qkfCiTOZ5pMsvTKv0DWaxBX
xlv0LtHGXdOROYlUoeQ/BG0UGwFhh71YovRr17uizIeIAmomLQi+7seepkPS+I5wEbo1VwZO+aU9
v4x5Jb+moTvL9+ZRi9nCtPqKtpIbu1HP/Ax0nmPFndsbZdt8Z5Vf67U/4OFpW/DNT6ZfMGZoIf6/
EptfYcPyn9BxdKdFdGZPj7QxEOWwvAvp/+FPgbegwTOAtGTwPeCeywLnrqIM5wdWqw1MAuFe2Stm
1kz42o9Lp0Ja7kTSGRMrkYteCcLEk4m7lkTIgPq1PUbJXEuQDDtOaCDtFTB3EvT6Ui9hTp0ULlKm
hPvVFLLpwXOixfO3ZrK1t4L7dW1N+JLOr30sNA82PcS8NAaFe1AJG8Ix5Ht8u6ScsdclLvvmK7w2
UA8J93sAPZ+YlznyIZ9f88R/YoAzIuEnmkWrBP6iybTvvBE75kHn4iuaoToIBjhNkwMezNxvc+FT
pxTS09l//N+w94lXmWVNYhEvSPChyojpISZgGp16RNTIJVwFhJ/IzfCOfIEQRB6OTFqlDKWhFBgE
W7OYyaumSScYpq5kgrpmJuKW5l3/mV0tylTDAywm5WS7pv+t43Yq7etziHjmPGb9/14CHnCC7mJg
WU7UZsAb4V93QSAfbBoEchc/shYar6FigcxBhyVWijgCoRO4h6pGa8Zjy1lhmVUCt3BFPTYmZIGR
WRDRPHBNChJy/TbfSYMrmW5piT3cXyoduE4N10ijZX9PJEHiHPIo9hkTRPLGziSmvLl8Nw59+Ekp
ayiPh1n7cgO7dLBTzJ700SdBVk3Z3jKTtWd9Fge0VINmqtqTsKKQrA4p41GE2GvLxW0hNCRMXqqq
lpQJaKXgn/ix5zn/eq8KC8/4NPZ8SA/L4Tk9huRtmN2eebDbbWsU4mvH41ruvLInRtqUtHF5TE0l
CSvE2pa6Hu+skrcy7bCRCAHIik8fflcOSWC+peF3U9VvtPVkfCj9JTMxXXBW2VK9SLWymkGf/xnk
RcirTF0Dtc2k+YoLLxatY3CP42+gUu5D79kYOXRN910jXkoUH+oQcbf3elHrl6/Pc60RhRIgUwNR
kDkyQ5Qydh/pc4dxA/HXtiMcDpnB5rM+TiO21zQXVS+YX6HDyPN4bt+3/cYzoR3NU07COXnXqurq
yt6n0Afkwfcj0seqHmHUipl19TRjW4qbjf/3Ca9J3O/GoKUIYUHZSmMvjmrCr+iV32xdbFwOCBPf
JSvLzSa726m4a7atZawI9UiFbTuBEuschqq65Y9RSwGxm4MVthuagc6k+n3j8OyvrooEbmQO/p7E
j4G64FQ04PYOzCJSF7DXEL1ulnU5S4E/MYhuV5RTMclB8cYHCao/B1GV98d4w3BiumAgwA8QGUeN
uoLixbkUU33LhnAKlbUFyWNbbVqaQJxU4hKfB2QFcKFUdRrcha5CvMN+q9kDFIIPaSaltfmVglBs
Cn1ddTA/jwmG/NvEzsHr1nxqpME0N+5eS/cSAjKua32aSlC3CuQVlz3CyBDWWE9RodgzK1IF/53o
wsnBI1ItHhEeodyeoEfupnbUX+j1bvwxHbwWflx2QDS8UyvEtEbgY75NjWn3Fo7dhMpvNZwPS6P/
9O36agFAQqs9qclTjsiiLfflPSRzKoxbUO+c4n1p2ESYydHv/23TorxATU8QtaDCY/bGQgoPTBij
ID2xZ5bZUCEt9YjIU3oJAxuvovb6IR8LfPAflUNJRUkGZ0fhXpC80ppM4Ut7f/0Ch8ld7WSgTBOs
MSUAZ4MWa78ccpIkfhOTQHDWWtK+7q3ruSRtiVqQavR+bJBSuwOE84w4T0LPl831wpRxEf40J4aQ
ow0sc2IOajCaTE21qaeH1t41AvodbuHr+uLnNxM8jOBPJoRKJk0ScvVxiwUS341Pz3quyBwQe/1Q
N6Pf+EZz0g+cMa0YR+hnDI4F9Tpn/WUiMZ1dpP3Azc2GDz/NBTjKCvC+Xtl/Z63ENnf1G188E3up
Wgsve7yq2JQqjss51qWgUrqPjKbzbzHf6RVBTE7Gz0+vd89w/Dgr9FmJ+jswpyj/qvSmamfXAM6Z
aWyJGSNZCYeTT+G4Wzi/VcToGNnq7kt6hRF/Cl/aS6xxzTnB0HI1tu+B/QS+dYhVAx2IxRo0wvfC
/9qiGp/7GystBGiFA4+oooldh2xjHiw6MkUj7wAJWEffDxF2c4udzLXcwHtKA++yzG2bCdxxfKxz
RUQQjH4asmn3AjZNRt4k9KR2UbY/misTWWh948v0igTcZ1NH5api/3F2O758oZzJo7KcXFOXR3xl
QzOLL2Xu57F1WicEipHC6ki/oKhe+V2Re4sToxi/ENQCzLwLGgMGPDTZ3yqIcI7XhJ9obt6xqP+I
kHhO9UDUP/VsJTximAiNpisUhusrwqmHYYPXsaDsZQZpWAdMwuoz3+LNdzfU1xKmC5iZhaxQ7IHz
8BBEY58C1TxsjW5Gxqa/PdK0cpkAvEJbXIXSiIpAprkO1BT6wWOInplOM9H0lvNtNSH6KalDLXT1
yXQDrH2rLOWb8TARuHtWi2zzJ5R78ou3CPTswrjSsEOsHn9N6qbmU9+SfKjCa6E4pT43yZ4Lw8Ux
HTxTBbHEtZnl20vUzVG0qo99nceJjakdF3GuQni7MgTsMcDmnx+Y9B9Ombt9V40sPPOddzJJhxEl
4z77OGEIoIYohRzcqLPcLBq6Io4QKTm5ThSA1h2FagdzN1X4Dxpfn+lVejwoSzaxfWsIG2X8mF2Z
XcHGbU5vmgH94dMt9Y2CIhpknyD0b1rARQ6NngnvuP0L/OyNbTevvzRMnWOtqo0A/ASD5IlNCDj7
qUXuJH6s7FVWEaq80qnAjhgekX/Vb7N/7Kdpc0BTZoxsZkzQv7vuiD5Cav83LiIXDYMxyqauJs0m
2K9xYGiipJ6Djrj0AwJ6K7aorviX1aPUpWER0wV2+rzhB0KZEAxcEWMGo8iTVcjgHE5h80LWjeOF
uZuI5MMU87J/jmJ5VaSnz/7WK2VZRYT8CcnHnYtPp6MbG/U/dE5k88acmBvhz08ZVvIbcfdMbS7r
QSNjyAH2Wbag693/0F8vEcLN84K61K2X/J7D+b7ysf5fd6+McN/M0/q1oMieRoOgkYRLoeIpB7MN
+SwAHvyEW8yaR5DlwXkS9BpTFEIeaiC6Cu8asEOVxlDsEKt3TrdruG8UyKXCFd8xshBkx+rla13j
0JnmUfEufO2EKHfnAoSUcyVDtNQOEcr8njuyAxXZ7cG3U4zjORKXcMKFWUdUJjhLGQBaYmCD+FES
GHw3jKnDWB+nUFJvyFTnKzakPz68TqFNcJSQTG7qOGzEVr3G2K4INZRj+AXyRolwoVS2K0Sfp7V8
XKTnuwqYgK0W1DuUYPq13LJuDiZHILgXQw1ZqdCZsDJY+KLU9PxbAcEgM9iZjnTNpwkKBt2vPyjf
VoCcNLsKDh32Wmh6mysPvlcXqYd5ZnkpTlDy4ciqrnKQz93BYmf94bfItjCN+vGBwu6Sa/0qtlmA
21XIgWCJ+AAmGCYIH/1LNDBAtM8Pdk1tyw6qTVxqEZfMsIBvYX9FdExRiXgCv8hndHQRXf4FZ2jr
UQIJBuyHnPDMKdji4+LKL4wj3Uu5pikfVJx343xkKTjWJB6KKau2k6/w3ARTaW2XIe2kjX1trohc
abKYV6dg1GrdkBWGOJkq1neIZM7whEJXnimkqV5tOm6+Tlaym801zBSs7UAvkEEF8dwjD4TYj8hQ
IW5Bx8lRHLsP1uiQ3TSGSr5CeQ2N3g5Q+chqF6ZCLVVwyS2X5n05h+BOe3DcUrwIzdVMmY6laOL+
tzyvhO4EErf2o80xXkFcDD9zEipnDPZ/jeuSB9EXHOWC/7ucwh8lJBulS+ayqIXvklaOWrlgB+9n
FPgh/ZErd5vKKHimI6JaFrlv54+/HET34694Ajhc8o1S64fZv6T0vtGGsi62b0GhDLfPsFTanyM2
Vr7eIQEVjRRZ8Xxwzs+DiHKypvlTNfdvYieEzJm46w0jZNYcwo9xH0prD7AMIEiKaKbGVDYqxb8c
CPM9hJGHlokmSYakInyQxcwnQTAcZ/EDaLJdhX4VtusTloJ2cE+JdQYEsJ2vGAVQ+ws6eiows248
g+KR+hi5cGc8nKQ0HfSwsg/uBOkeQJRSzYaQB7ye9eGrIOtRlKXiMzJ3/3p4IWQk8PsKEfOenxqw
uytvBnBz7e9CSRz+UVsBa1qDfa89cC/7LsU6euw/S/uirtH04kKvBULNkyRhzaCZNk+DLd3EfG0b
IPAmwOl1YtfckIJTX+qLo9ypjEsY2bJwS/Rp/WxrTBt8ki7uEKlXOMHW4en+xTZXsxbQpqIPYvLm
EkVwbWMZG4OGlCeqU6CLU67MkQqa4LuEbnty6WTrsBZxQW3omB5OBsMQ/vAksEdtk70L2nCmlo36
c1kLdoe72SbaDksOYs9RNM+7ZpuqqcK6VS/YBXY8rN6sdBwa7UHXGuzcyOdWVbita0mM/2ZktSR5
6kJwBTu1S0Nxa57VgNWTJuj/h7PPlUdb0ieebMYB9a/noHSujw2kBKCbgoLNBSq5c+QlwCPlFk8E
NkE4IBNoFc7+oCLLd7bZCxNKR90Q27BoUaRpmAmlWDl6Eea/pzURx/pQNICTE4mwbOSqg2lyKs/Q
KFbViLe/h3bfBdxvMQGzpIE+/na+TtvaivGGFLWDUy/6WYGnSUBsufx/32vtiDv7tLLqB1hhz0jY
02Cvrmk0Uhhp2jEQnb5wMy1WPIicS33Au8WcwqiAMw3rl1r/9wmjQSmcnrZpO+hEeQtL/Vor+cBK
f7zEeNckPkHe5YLgGDuJWCo+ROUv9iVb7khOhACsu/HHGp1NVUp7lHqYAqcBNgQ2dP3+H7nt8W4j
SmlWGuhMgVUM/w/Cv23BlVJEI7b2aoTDG1LwQOwt/Ft7ih0fXHLsvdnglzpCywetIrCzfblVcD1Y
YucbUhuSbtc+a6/Wq0CbW74rzdgeZ5btFig6k4WkwJDOLV9KUjsa+7LyERsj/5dEmMLwJTLo3nH+
NQyJKo2VEGsOPppOceO5AUTJZL94C+ulvUFW6nhTA6vlNk0ULYohFCMTAjanbHXuHe7/6OsVXgD1
T+x+stSL/q+Zo2hUG3VWJJR1VHVNtkCsFXkdzym5xPZMKxsidnmNONilX3+7Z95K72xIfg5C8trF
b3s8JFGPL58MCvJbdlHzQKV3Mfi3a9Ou6SKbL5N7Ng/0WGujmIwvaJ+7kHDelTxzjtu2oSLLD4Dv
LQwcz/gdYeMCorHdmWS5K8uFIrhOJFnnAhAEv1KY6L3h21YvJPRfwdJQpEmvnwUYmW5EsNprIMqm
GcAMqc/fKXB1tVzh9MBEVjAcjqbx7XONJlWJIAGv+YX/6qW+UzsWALA20Fw6FYAuAjeMdALz3pkM
r4c+aMBFu/csa3qZsxMt+vpcNd87DE1BHKsJMW4qyIGLTJkyPYd1gpgNd0g5fIgWTiNLHUZB8PuK
lA/xE4IVUkmIieC2tef5KsIAuWbPygKz1BITgeFdqae2nNAjg35a18+Oh1jEa99P1sZ6DxK8iDFJ
SYeyHAbmPK59TrOC4wGzeNk2mQmHN4oMxkELsZ9ahGSfCMA2MMPWcyG4hc4wmzxQPQCFPSi1IAwb
HOdozQhJoedjRkZLhhOzGXB1V3kTx1QGOhVcN0yzd6I2QAgd0uDYPIpAZfqip3cHxKZqneeiZU+Z
PZPc86kewZOj38Ty0KWViNf4qxH4HSQZxnFtbaPuabckA6m5qDz+kQLIfPR9+8lhnBBWCNygkFW1
Jub/jWF84/MR6D0kgiqAqX8MlAIgl8yvpQC0DjlFE450Ba/QJCPkDRB5Bw5+aWtW4JnXHXJTdtQf
gLOdIUO2g6KzRYFJfIcqTkDBCOy4zZcNBSBY504vyVccD9rr41jSKkbMyCCA/yvZLzl8Wso6s0Jm
vPk0Q/+LZGW6+CxLWILAwZ84TYHZWPHtoYmkzlEYn8lqZhIpf0646l6CVdALMR0eTEnPtN6OOznD
L31970O31CGtbqFJfdcPHoyqXb0nKvntOMBKJl2rCUBnvB6M+bOU8H4wnm5SANeyYfYT4aB6FQT2
FWSJBIDA+bC2WN39lypnwVXFvdKT3i8OT/jZ6684I79XDGkRhSiVyfj6K2BgtU4WmlKGdDs7EjaN
aiFd3D4EhVvoPUZfMNCbuE1GrfRH+HMsKWm2ocFMJB5ZO8XkKc4qIN2KMP2hSec2RWMJjP8RiVGn
RtAwR6l9dOwobtARJHGO0J6iITcFB48i8HGYywtfpFnhjyxZGcSM5X6xXc7CZtdyguU3zTjgPOAE
qdAF1fvB5gmALfGkA7aFvqWSo14F/6NicJodC0119PuwfvOxh3xqLC+8NOAbF9tgYZ9SCbAJDruU
wD205Xtft8nuYs7krJYAQOEszLIg0lb8p2RhphBsvanpLSQ+TW5ZWLJtZlTIu1i7+YIjzMG65VoJ
EnSUEHPIUo9EbUAxofIAl6n33e7Q3TRx0ZYoCApHC0TpdJJzjFY9SInGCKB9S+ab/OH8G/fbHN3d
9hcRtm2m5Doo7EPGiQLCAgpETZczryGJp1P9P9B4TE1XbOwwlMJ6CA2aNj3SS3TKJDzicjs6wPjd
D3gAqN8dVHTe21neFc5l6Q6/nI60JLAa1KlP1vdVO+T7KvuGx9ic32qIoGI/JWTh2fnoSH5sYBN9
qWeRuZmaZiQwQNwVckOyZts3NaMv15VOsDe6FdxwhpKvHECWzGROZkJiW2uPgrMjU5N1txdWTlqx
ZwN6D/yrUBkNGhJFHZXjAOqKnA9KLkO0a967t6l0TU1kTY0XD8374o4w3dagZD2/Ut7/ASm0rqGr
FNPbwUiycsAjuAfRwfBNQFoQpWYALgXt/EXWfmZ3Vos1OErj5jjuUAPt26AJTovOEvJzrjNdeCH8
MzWhiC0bTXlpxo7uA+sm1aq4vKJnhAAI7tYM4/gFAqh4r9VKMOm9rz6eaF4bman8IdmUINS0e54E
Rq74GQqwSlJREmbPHYTX1Qdm1VJsn4RNVQDvutTk3Vf3nqSZmhZxpo5lKAoqaKMrDiN6K4rPjA0y
48VaSNM1mF0cUiRFoj1Eayl2rsFRPFq4kk8thmleoqnNoQCQFnJh6c77kojIzGJPJRCOth/Abonn
/hQB9No/AqGzKnD9ZXDjSUAScV3fVOo8VpYzRSjWHoN5qbUx8Us5XehVX1k8FXHxS20elEuXrgTW
bN9Nvt0pVP7RjlP4vFFYcglh7xx5CL1HyBV3pzaFR0pSm6epbzlgUd4QPlT2nY3Pr/bm7psnIWeB
pMD0gJGiXCNQ8/VXu0dw5MgJUR8Ru7CCFcUZiGg1i9BkxU5KLqAmQ7bw5QsrCFH8j99CtIWe7hhL
vG1cXQYBHeL7Cff0rDf11pPCNwmt1g3mxh5fpwh6G0M0D9UGXlaIF5wwWzKGljKm/NeSNi25sxPY
e01OEtyxdgvaRS5j50c2b+Fo/y0TZa59lnPNUvzXXZeX6Bm7IU6jQyJ1kHYXyIBW2XZidXUw6+nY
Pd8uhJl2En0SMuQ32pLCXvvNy5Y6UBl9JNboY4XvnJOtL2FIgAZhS1Yfp5yvm1QJbMbpNFkoCoVM
8QUXomsGMxvDFjxkfBGhaVxcYI+EWYzPoNN5q1KDAs/tzYXrz6a60f/psRY2aB1jePJ0JfPeUFKT
1Bg06V3yfo8Ub7ded+F3z2GDUFeDiZFPLDCyV1neo7PRh+1ao517WMJ2ZAmzV1VXUxnXKafi2MGX
J8waogvpbDFx8jg9WyIeTIPHeJSbi1H0aEaHccWrMbJAaHpKVEKoekwlrlAmDLXR9swgGsIz73A+
2ff0FnJIltH0O3i24w70RxUIB015cdp355C3OfBtu0Ktgc2vCx0JZRCkzOeDOOXxX5UAr3g5NZf5
aNmcPfH4iGtgvaCWk35zEOOlztWt+WLdB7OYtf2q8YZy2T5Se+NMp/tlZASg2WQS3SYMcD3fQOjP
7vYaGE4Tfc9LXMIBn1bFIfqAEkhiXO/cH6s871pSaiPM2o9G+dtCMi05uXjtSWcaPMMbyDABBUUT
GP+Aj4pl2k1VYiaLKGg75IsDYONpiwBgj0J55f7P3GIJrqq+sgqL5FzJTIHufM+oXcshm95imF+T
+3YYGvdYqt2khbEzhAl5cLscY3i+Hyx6PXslmuSR+8AcNLzNUBQm3BrmYuskuXIOvOPKHGwnPIy8
X2jpVqfEoee4NIKrwpOlGhIpI2r/jd5/io/pMil5zIXhPmF7uajoSJyR/c1LcIVXdVFjTppjk4Ff
Y1dWzlYLTyJSGcMAU2KObEbvJrz0Oto9aA3LUjDbnXDq0V1DF/05bWkq9uFvmZ9xYP/ao82KKUBf
oBQj38c9/rD+x7zWNdiKwRR4Kj4NtMRc6EuutVjkcNPJ+lO2i7lt5kYBpT8kqOdVjBEzPSTtKrNl
heM2Agx8+YqxwJUGykDRXB+KVyQs4tJN/9SCQl1RNZqCb0O7rUKvcjwbyCyUoMhRjiejD0Hu+l3u
LnyDHeUU6KpeuphYsICxVGtpDMxND11RYd07Z1l+IdqLvkYNIOnODBA99DrHQyY97LwJnfXCU0b1
YDUw5KpR5sVlKL0UU6G0aJk41N2QJA270m7kTK0qQdvomL3r3riklx3tzoXq6xQOI6ku0GVE4quF
ij1534BG+Q9ag27bLREK+CI6J9F8Mx90lyTK0+PlWTvKIdyPGIwyebtwGjxB2drxyE8pCO7zGcf8
rhVePeDeG8d2paBdZW6ifT9xmeKkKc0zfOqup9vH/LkrfKrGqnNLo3EXCWblId5acTIqC6DpjCii
GNtp31rWRj3cN7jd1LH9MCf6b+Auj7uo0gDXR5UoKisSO4mjWervneh++0X8Teq8LzE9W1bsIbxi
XLVmV8qDR53ZNuZ9mXx89rUVe85DeUar7m3nze7/Adkfrm2HsAeoDj35AXq7pliIOIkugURPS8ze
fxx4GgmUR/d2V3CoUWjh2RZpZEiSvA/I1VaDNCdHIfVxqsvGFEpd/Ncbd0R45um+CYWlHwfgU5Jj
gYrt88dHskrYjqjoccUuZtNnFPUW1ba92R6wTfi/D33U9uoDr+tviICbIZF36gC9hPrJ5nXi2iOQ
hgXTSPiyIlfm36mvQI0SMdnLX5ljGorHJ6LTrzz2T8XjYyEstiY472QL4M4V6ehdIZ1kxG7CUeVs
Wnh+uNbJtaD3mKdvZDas5PDVeB9o+q5l0SYH0rBrvSQJC5ojWKo8xXbpAU4vpnpmGs3hOY9NBQxt
ExR36SnBGMQbgASir3gCKqRtWlQYIEKQF3MGiw4NG1snDi3dgX1Yw2CYzCBUMTKwScIbtam7inne
JK9jOL63Jd2k9qlLFHUoEaDGsHqIvWU82RhI06ouV3RnMkiAmaZyp7yttooPkwCL5gg7tzYLwAWn
sFjcYSSZ5jcsI/Jf5oCrxWFdpkCABym+Ny2kHfDBLqrS7RDpO2GnyELwoP/7Ol9BmPr8xXO/+wOO
7knh4Rb380ctQN+1UUYcxFHvvT08kjdLRRkbtYgYD8SBT8n1am1c7gYY7AS6ibK6P44FKRU8NL53
6WzHiPOBNtr6LeIFCBLPU0sd69vuKHURX6RSYCMl+wLRs8pLYis2CeKd9anH3CYSvwsdQ9Vz858d
EQdcd3kKWnOfICvtqGcCJGsN+1koibEofL+6mG92PnnLMx1018srOmGc2AkI4Y0DV0qP4BXPgx5J
Nmq4zvvXDwEfkx40s1LNrT+sVLsA7/tWpfTJ4MY6id1KpFrszOgaJqjTxDiuxbOXre46wuGmISMp
fjAZ9jIXx6uNUGOi8XNuXFYhDLuDL/jwAkEmFiivyd6Rp69bfppRHrLwody//OF/bz9s7y5Pf9VU
baDo3zEtLJPbArZAfyMaTyUn8zTS5cQoZE/UoFdxq6JiOLgPXOOFk5mS56LPviA+Ly751jU6IuzP
u4NS/kOdoGbmTWULqN3nXPbwykfYXMUdiCtqhkhpmYQqCHt3Sqstv067PTFCYY3XYZ8GCZ6v6op5
3ENRPueSnzVj4ANJ5VVzbnK2dEjvuNwb5zVAG6pM6rh3W11W+XemnpIZ+6XMgMFxQpzbVH+CVnQM
W7dKyTs7rXZidtEKtSjNfNftykCWdfSEUydo7uAMvKaOj18ttYMZAsk42KEmnSDUidMWTlbIDdX3
cs3Rn2LDvpF0S6gUUX+qv7rgOBziE9LzDpRG/fBg7Ib294aTkjJ9JC9V1cLI1jEE7zBIvpm1nMPM
sUdQNpxTi5JB5EIRlh7f9SVVX0LcBUybA4C2ytNXP+Nx7t+iV6HgCAD22fAolN/u3mpTf1OLnmCa
6zK1L4JrlMJY7t/HjGVJtqfkD5TwnIueMumoIayfBQTlCvJGw1aE+39ouddiY6DeBie86mpSgQjG
aU5Kh8qsRVg7tphJyoHNBAE7HUGk5memO7WTjAQWWDTFMN7PF9aCx4d3T41TWRlCvCzhj5MPst3o
TgsUpVL1Hnru7GUQX3VaztJW/lthO7lGL9kTelLVk7LjwDxOQ05hQfX7+sY2mz/ba0i1OTxQljJY
1SoJzMSf8VQBqjqwqOAOZI5/X0iG/vws6BL3XS3CXGriY1C9t2SsYpYim1BmRTkPrT2TyC9Z1eji
gfpoNo9q8rny+/2ZO70D4297/NaU8r+4McSV+qnvgiurZwo54jU8C4G5i/4g0A/AGPVEkrQSfmdy
Kri5Th6W52Su4gZMeMzXr8Mj5v7309/bz3vHTwUnf4DCkXIHOeC/ki5Mf15XDhwcv/eqSVUKw94V
aj/9wTbmnG3Sw83Fv/uYfOzH1KwPefKEPt2hNKPlAMBnWhQhV9+XXYvtarnrCb/MJ1Blnh35Inf7
topSeD5gyng+DfgNihgaaonNIuPgmzR9LZdu0haZTtTpS7IfJfxrBTtFXvK9oWa8uOSKt7JTkZZe
q9FJWxsWt1ocER5huUOVIkiONvD0WCtCfQcuZh5ZaIXpSsacaXwIKb91MdhWnn9AEYaUDgbOnp8M
LRU1f2xk6w3c46TXCGdZkz13cGmTuUANZExXcIWJ22Lm0JnYZEYfU8CF8qmmxgUU0ZagITILA7vB
3xWV8wlb3yIV0aWLMwqw05ocu0/EJ2o8i0GFwGfo16SXmAoC3eiw46acJVn8u71Huz4CemYNcbFq
13Cy4eJNAF1W9NDHdeoK6ulwl182zuYXWi27Fpt8dgQys1rKRFzLlbLCR7mzQPsCCgVrWOudSsoW
5CNP/bPNpyHMVMqkXPnnjhKzoQMCa/AQD97/AcDpczdFiI6rtOH4Ff6YsM1zBuCzKfF3xNLNPNi6
2f9WOett1OOtfTntTq8e0gGgQ9PihH4wxMpZq9Iurh3btoRGfa5X49z+WxSLQGJLLk2LvIjCM6v5
tmCnC8QWadaagFpXBILDZaN85HvrQGbNdu+L2kUWVbAyUHkqZsphFtEHqUSYfQf5vhH2QEA47RmA
1FTo7LRRwhzSyS7kme8QwPgf6uKAhrUCE0XK5TCtmsNpnr4TC2llL5yw5qXjmZKLSHq2va0Q9zwk
XHstbWSxTs4IrNTiY2kJi1duhXm8PpuZ5xlMa+NEuYfJTjQFHXNk/wAZ0++so9BsbAWLr68rKKvK
ETz/Seo+oV/jCJUQrkbYUEo3vA34uNIlvoyA3SAFjmHZq2HmQFHBdGivgxMh8vDHUYFDXEprT+Eh
HX+xixzGjbds+69h+aX7gRAroHuX5v+KTP+ZmlWutv0Cit0Zkwbmux9ViXONpJhnf1l237InabNg
2ZB0tfi9extqsb6ecZBIQdB6cfEw1z2HhNGpG+FvKmBLcY4Kd/2FfP1RZOxw4tVmYyz6n587t26L
Rrm2Vjk8Fvd2JKy3nIIB6ecT74HCLTHaC3SwZRkhwtwRyxW/SY6Ls0ki0un9GuvST/m5PHxkftsd
ZS6RpoRzn9Sa2v2wxuMiYbc7fJpjrPLxAcnJ8bPiPcym+UoVADW8d/2W7Z3sxkt/SXAKFjEcV4Dq
Q8n/C5u6sUMQ82ToiQw01n9aPE3Lt50m1DF57cJCQ2txIJfFin1xT7GGq3gxbf4brm44ku3ypeWK
jztFobphKJM6oc0wU81h4f2veSzUaSLFpDqJj9KFyluqZiRViN2KzqeyMwoeEmekB/gg7wRTJ/+T
RE+8QEcatgzHRTmOV8Xeyc6w7ZBkL7GxX67gNV4igFC6YxByJTSAR38DUGRvKHC/eUQ8rBn2iR3m
XHMjs9IfPJ5vIcBzN8U0B6kLUl6OpxYXSE/FuCUvAjzKY/dgy8I0o7k+doMXNnKrYZ9vYvt0UsiV
wItfecbfRTHz7t7zYWzfck/QGALaoY7BIz+MyPJyTj2mVY7OANFknOmfN5vEOma+By0f1xsaSrv0
J6gvlxcS4H7fSCBh43WCLX60bs1j93Xc8GPVrsApOhw7trBxzhCUztXF6DL/9zchiorhcrpEt+uc
OfKlY/HiIrK5kNYGPtekPQ/AB6lHg3U9KXeti1SRb3pmw+zaMCX8UXLYVxyElt98LL7UTkFIDBxL
0fbCphZfla6MN7FiIt7Y8idy3gQ6zt9CwaQeWkLBbCBBWf6GyPIO8IsNGii7XfiqaIfMfgIEnZk+
wfKztLIkQ8gACcXR0fGX09z1mCFORpw/4LGH1jTYsTlGStpG/TwpZbpT5qMkKASbGNVTIjeT2CgZ
U+Ut7yl6tHBpv5KiUeoIPryxlf/nS8wRm5Fez/n6okMhDHBkNFPi0iZVawlbAV0eRATfTzlM0Bdq
pozHl7LLzez5BYSfI0Um9ypUvBpZr9Ddo8rqBmw/KcruNbJ05h9rEEaWhzkIqo0j6uboGY2VOrnW
vkikaGBdFLHu9ePHE3/8ng/OfavZCDUwxfsKzTjLwfGUQQnFX0q3jUYQdXFaS17Mk+RoepNStsUP
1QavEUtAj3Di7W0YeWQ/Nti/j0rV/39LToLh53zKFYX+EOx0RfRHF3UTypua/wAkeJpUlk9/+L59
a3sNxfmb5bBacF+Rku7fxxAJCgXfQdE4V5wNFY2vQArxQ0PScJQJEvpQXjoWISem+Qldjlc1hGom
kWuBaki0l/f/LtCYOqrfujYKIKGic/CqV/eKmp6Cbw6Q2boUnG1mNJBIhh1DtXzaOVbdgYn0lFr9
O64BzTv3sQPVrDKlWYCFgOvFDyDEqLzmea5XHoloxTqgaw1twkTMfs6P/86ObIczOXN8fGCo5kYF
lcw9no9Cbh2XyniMy7/Pbc7EcMkEFMnVR2KE9AL9CON6aNEcEFRcKcckjLT22GxDPs5TampDn9Y9
bcRkPplop9zM0tDsxcBZyknwj6wPqVcg2W+Q8rS460qWrQupeqY6kDaKuCgGxYyWl+aah1YCzBCV
MDxTxErXf1qKSnvm5dzupx+5ZDIYVlyqnKmcpy9VhRbZ01gjBF3wLbiK6KB5H9a6MYNPveEXjJd7
itFEnT4CycjpsOM2kbpNaKbAMJb9IK0NNBeo40nLjI32UMBrfB+bgwA4zdyr5GhzeEOEPbIsQqy5
lE6tUsJ+gfWn8TPEtD61mUIu44+fKFL1CXRP/pC4GNCob78aR8SxkWnoVB8CUym/XWUjOfRJTLkq
+mzDB0xFVal7Ey4LQpM4DXQD+4G1D2gGsyaI+ahKCjfVWHr7gWDkH6vizi8pSMvuDgBLb65o4uZf
oTHdbD+HJQnfbO1R9YhknDy58oVuSsXJhcK7GXEuL94fz+jhbeDWZlfSPI3FtlvZeYHQx4bs4nz/
xcGruSxrLStkyO2/W4R9OG9YyH9TsGxVl4ev8Zl0WaChEbwwXzLSgh0uzas7WeqiQNWKwE6LorcF
0O6KgDGJ09CNvbVn+hsqMVsKVLulZIhHjJUIxoFSHmisfQmvmqYeYrXzVOR5qhDbK/mwOOs+xgB6
AXMRukpJcPnlaKqs57HbVazBrkkyAt0F4Qu8fW9gFsadKk/eoo5ntUrlrHfbmEnJ7jzpbuHvJSXh
O2XRi6Ys0+y4FKkKkh4LGEYm6z+qwSx3pqTOG2ar6hCLBYPEbzLx75Bkuzg2IkyLPq2OybgY8h/+
eCvWHwYMpwQAajIgyND8ngo2ZSQVa65VsPWUQmzvT0QeGlPr6ClPVGSzUaGbSGehDFclQvS/vBVQ
erWwsbI/c0C5OeFpagUDhZePsUGeJMb+cLlHBlVkYPd0hOtJBqGmwIEQ1nWiFrhiuJz82ogN+hYe
JOB8rktoxNlSAKgDZdLFN3MlhmD9Q4b56J/5z9Z5oy80/mb7dxTrVJOgfzAghcsTbWfU1LBtfWof
c3Ra6licTjBczSoK/eYbnm+uewxEV2Zj8ngb/UpA8IGqaXLIeEH0TRa7UCcGVgrEnQ1qbJif+vDa
wAvdA9bWv1TL53CtLCIugkseIcqok3/ZsTqwWKem6CQP7XuDGFFoMLNnJriV7RRodkXQ+N19goOR
VTHFtBEoXitWEO4q703nls+71ELXUalVNaPpWq7xh+QxiwzYd5/9kWW2+11dIyheRE8YVHESk/HP
NXXzR8UUO4vq0/ZCRUTt8YUbm20dC/JJxzrPkGAfgSuG1ChnEdTU3Mzvwpt2nEUOqSGd+TPWvw2x
xXL6KJAuvbi6O//j1Abr1Dy7qv9tv5u/jrmbq9YMkvGLEOkkiXm7JtHWK97fHS7CgSzeLhsJOSJ5
mRhx2H23/2MDVaE41Dc8RX4TV0sIq7chTF0zAXbaJQenuNzN5+IkPdiG9lE52ip3czFwmmTaG8H0
02CqcYDDTU3vjOQivGo07JliuGoxiXgaq3HJmC/Ap7KcfPWy8HGKKgmnU3oSEeA+CdzS4x3gpHHu
g5dWuD37k+sBgIUP0s2bv6EjJxrUXiOwe5VqGWLrSpCegZE9OhkfbWHoTXTeUCrJpDOKWloETMOZ
PED/6rhTqyzsHxqMCz3ThylhTvyGZ9HiTFyGPDIrOA8+uqfAjXSLrMpUSNqALNY30Qmb2hnMwvsv
VPcf2gNwnJkQlpmNGBlfwwW3CpTJRPE/AOCbg2UKbHMnZkvLEkuZg2RMfacO5/5nYxBClJnXJPrd
nP8GCIp8aPH6vrLqKMqegZAdfRYmhukUItS9Umw9JaKr+UA0lT6gzNHJNOfIQhtaSW7lHFoWvz24
ErLE/hbfdqZF9EcMQQmdrKOTmdDL72N59f1DaF36cOSyS5WPqhSKgxT3NWtfI1zRriGVpXuG1C3A
BAL9SRuzf8y5zv1te39wAfu6MiENJQSI+q/ll/yPkiw/HNOY7H50fKaKHp5tcj3xHuuIhjq1hz2P
7XgPVRcNpQRMdSc5wZklQAQMOkpYwD0AbR5Ar3HFkz3phEl4GCd6XJDYxBKe5ShdyAMx9ZLFqLpw
/jEc25up5lSd/m/AwHJ4DQ6VTgmspvse5uJP3iHtmsDvmB4137mpFTgyvGtwuBBDAMomNB2XgIR4
7vFHTAexroQIQxLO9Oi7lgPlvhqpj0X+J70PGqiB7k/drv771J5YcKuCU2HEAfkWPNjyLvoxZnsJ
grAiSc78wSnLK57NV19toPHgeTZmw0pRGjzbPq/P1LcSX0OpETmAZrpJKaY4OryYHbMqMMxKI7EM
QTPk6NrWFvq3wRyY+wAJpXGTcVCqMRWF6cfB/yhmHxusDeDiWSiafR/f21A5EJuURUt3xn8I0rBe
PMrvr4IeEJKnf2ChCeHfVQuhZoei08W8zFcS1U2KqowR+ekzP6nIyzgs7pY6nlaMacw+7DC3DHdf
gh1F5B+nYXpMQpS6+XwHILFvJOMu92FBpclS3zIMJlpFlvvRPnGt4Yub0cgqps7ma+64uu5wT0mr
oxAbqDqnZK25q0Wf9WSRMOZuef++JDoz1WGLpsvL5Y4gaN+hu1oAkMtcLt2g8mqQe/vwFiOv6zaK
IAAAc8qb/Rq6pLl4OMZZSYLz2J1tZnZnN6Tk5t7GQTB5gYnU3IhBVfAUBs29rIYc3+vNQS/2N8GD
QCEdJnN3wvjRRnBcR3XdPCi7tQEnYcDSThBS7DVuYCkJkNF/r9I3SNrxWc151tUTx12SrZaa1PtK
Bohy943GBwhg8Lf3/IOtCJCacE34KU5yr6LAScte2gFZ/TTudyFLw706IhvJVGLX7aMvFTt0La/Q
zmusRCfth1y2LKRYM2QhxgXmRC4zA5lR9MQKWbGlYAZtbn7+vSfX54vQgmqD51iRX6sQeNVMfAx5
JR0Uj5rs/egNUegjXmoyDBsSPkwvbgP6HpXf47WqAudZo40GMCy5C8t4DGFxK/Jg+RDL1A40ofIJ
M0nOHN07SwUJRjkfjMh6CPHaPZKB0HBocD2PtVtxgh/1c+m+GYa3ztzXdkAug1VSGl0iqBbbr7Bh
odrDRmDINhKatLSnJonWpgLaFtbFNC3gTY9wBy/oAMKnQuWYZTzeycwjo7F0Kiz82wURebyh0Uj2
0QDJF4sb3qCYSjqv8gACEYRCeze3P1P6F6u2ZWahECbEMfiy/iLToHGe1bZOSNIQgD7RmtsHWJHP
wyz768XaFRi3GPlvxYDNghmqhmSWNTe8bx/Dvsez8yYu12NNbxdDER/VD49/WyRp/RGfsUy2A54l
RaawgYLSReeQdeH3d8UN8TvCBZaTFtPDeWcZrq2c09Y0pdvv2eClpNLan7DIuRdc7OWohfXHatEf
GsD/mI4AAdHBflJVCPn95IMv8RN6wg37R7WL6MQ534cZ72TkH98Soip9U3HwvCdPYCcDuQkwnY8I
TLXh9Y2/chwpAG9DpvFLsJMFSpU1sfRVE858pHHoBlZt/EVnun1mN++t2cKgBxLITmhx3aCKMdmM
SDJtU/GK6j0rX74X+0sQUFKzEzxeDUls8YI/lJNdrtfo0TWt5ks8ZZTOQgvI4SxdHuHMGC/iWUx4
2Zo/Xk8CiOKqwl09jHEiNQS7zg3vXU7dd/ZToOeKNiUmlvcakw2cIVEwhCpT3+Psck4bThyOJVeD
/r14dAju8O6nyfkujTShjGWgLHJefG0S3R16pK1o7frQgEtt9hR04O8EFtgbnQp0MNc6V3LDUh6o
SrxBOva2PGR6G7pygDDEs2xHGBHFVCOFYJJ3B/0YpUoUo7OA0uGQB5A0lOIpezlR28khaVpmM13I
bYr48rmPr17aK8Gc4wTRrXfjBPymyTZc1wPJCLxhPtzyhRwGkWypxMxyEYxAC0Un8IEu1Nb2uyyO
/fKdMOHeEb6KsPhDvxWxhu44qgmLv8nzy4o4ysTcXOu8ZyTC3e5u8ay+OEJDgqPtEgn6Qyyq0/TK
pNPPVfMsa2vq5YNDYJocTeu9Oi7492Eo1aQEtibm/wMMc1ELC4SXhk5wAb0SZfNiLZeHagtwRs4z
W484kQmiFVeabAh2r47Q0p7IHWjYCcUqw+H5O57+llIJoRGax2H8PfjbzcOK614MC9NPV9RlDQf4
YlIb/WkqwtIZVE5llT2BjKBVpVPRU80l6txSkLq0Mv8Z9Z2m93drvKtCe2MDoAzTlZyzFOtJ2usP
NNFndA/FEFyQmNridpzhoxWOa4mb28XYOm3pR9uwIpbstp6VPgv44r6RIORF1OdYqnbGXYh1GjWR
GVvZfdLcTehOjgDVzzgW4tZke23+C7rjLjDECqpng8lV97ecJeO/1I5D1LnJ5wUS4ODlGQiVTNhS
2FMo4pZvN+IGPKf0ayp+gRNF20EC6547J1kqr4J3CmApIDHMU1u70S7Q0HNs+TnGK55wO1czrXNt
Oy7KZZXA5NBm71F4+GznfFN4Fz/RM0vfM/Ln46yfWatVK7XTHgxVfb6i+oPruWi3pbH0Sfh1kLqD
wGPq0MCEvoVm8hDrei2jTYiV118TI/lZNHgVWAgZcMWZk5/lZsv4CHnZjkFXHTVFg6vf/zIPU+9B
JYFy+wxmScHrP2zdTforO3hsGOvSI80XrjTo3/TbSk6uz0pXHPGRb91rSUQaQMw6uybR2fLZUm2T
DWajeFZ347uOAWmirLEMaKKGgfXhUp/zFmx/ho0uFOoIp17o3sxreYe7U9YIOqGOiVz6S8/qrnNH
T6iH/Ib3P8O1X6uYmgpF3SpJaftXZOe2Id4sAockBAKkn6hEgdBp23hbt7lmapqsPU0Z28L97b7q
j2mD3Svi7Ukj/wP4DoCfd7KMFAGG6hy3lVl4sDCemtO+C6qkkIVBpnXIHYeCxAZJNUz8AbrIK2xd
if3f36kHzhkwMvTbC5mKOgkG3xvzlbltyxDFIR6Bu9PdeHzQlerkKpNI6Dtldyfcpq8a5jJ5EAly
35cvtTt/0SOvDKIdkiWaX02DYR9z5OzhCHuDXngTubT+tA0uASHURMrqXvB/IkI1/lq5QYrdUoRt
/JhbAKtfSOh6kxoqcxWXoEbqdWG9HSu3wD1yrFehl6pfH/ajsmIVRVG6sG/s9Xc6qkWG0/LjZ3hq
eCfSlixJSAfr3hNTQeMYc3qCcB+iRwFkWQIMvyaJAOsHVEq12fnAwvj+ce80+UKEUqn+/WoSES8p
ud52IIGrn9K0JAWrJvC0+QU1zZ5pcafmq7COEUw2hwzDMpBP4e7GSFrYbscELHtLt81KQiqMRXHC
fChFpJJdngbcmOWarn7ZFhlEuIHGnQFfTFpp444Bjsp5oskWv3pfjFbdSXIS+37aaWz8qHxlmRXK
ugrf4z5PeLzwT6hBk8YbdmxQM8s0Ki4m3l0ujyRFR2DcttRwK/vD6vW7i0mooUAG9yL/T7kpcWSG
+tBNBfCA8rFXpYnMciUoG/gjLFuJ+uYejJINUuZ4A4Hpuk8KXcxCdizl6XH+rHx2mlzIOX3Bd4OZ
qXevPrEeEmkfTCuL2XfzVxN8VK1JHaw/bCa+kRj4vBv6Ta2XHNKUztNp5A9sKgTgV4zGZQq6jKuN
wq5sHJLF5TS483Qmur7X8Ys01adnld2YDESPwTEHmqnqueEY+lPei+Z602YjjZqBpAxfQ+JVSH46
cCErABP7C0I8KZmBka25JU+s3sRwbfvPQgCelSfIlOr72wv6iml7f5G85VgvLpUDmF3UORFTwKax
CJaFGT1QqY/7E/XX4Wmq2Yd5yCAqd2gjpPCHlcflMPxJQRe6J2iMxRwvlsTSL7b87e8ona8tvy6p
FbPq9Ou6Y6r1qfJ0EKe8C+h5F/7qEW2r30hY7rri4x45i4Xm7JP498hCkbgd8DtKmaCvnxrBQR0f
nSdKhXUNJWzrqSsJAhVT64v3OjUjWWjjBep2UcsNNQgi0HrUtJdF8x4t4EwE7MEspR0b4x/4DsEz
/fyzMXYOFs3pmORLTkBsoX7xdDyeMM0fhoJtbMG1xL58lycu89IjVcy4ClVyg860OPwjsTwp443a
VjlLEEZywUN5Qi1I4rEini5n1PMqO8DsjqUmt78l1XDfDiaCh91zazj4B9B7undKNK+jjQ1/3cTv
aG0zeUrP6zAIOGpAvetk8AQU2AJIlpCCpz0tLn57ya8geKXsV6HGm88pAbx6+8ryNQ2/ZXRitVA/
60DHdToizJaPYGtMoFXLwR5hbBGdLKQ5xbb3GMTawoDaycYTjEIM+hcuiw7QZRxkr8lZ8T11s9Cs
PgmowSIrVuoQdhu9eORz6WpvCq/V6XBJnHgSj52eYqY2XVzqeKQkwzx+ni1uSAfr6Lq33VTXmJ0n
ztDL3ZCsCjZJPaZuEjjLUjLcfms1oITx2/C+WAm2K6AhJXMRTGQFVE9i5iQ/C/oonO3zO4kMh2DI
4yQYkBnBJm3z3CNxzOGYXFE12qXinwZCIGQjpNPKAqF0tO3T2cmgSKLlVfBV+eHQDscm9gqNgJ6f
MqiqXGV7xoVNPqdNHPgeCJDNp+m6ysx+XxlwlSKoFap4Jx0VDWH4F8jV4uEIAb1Hz3q3UM0FzYgK
NXUlQAv+I9MDUxPxfjEyOXD02J30uSZYQdr/0fMlR4NZIktTILhBbvq21VsYZKt9x2eNwJoVEzpC
hd8mTbsJ5pEArvko9DF2oscZLxCXzAgh7wF+WlKSIqCi9OHZ+mVUFILOXWryw+6FhwPlcwB+C/Sv
gTRNp2H99IhP0DS7+nTDP8Noc6fFZRyDNB9+Ut2SABW2qJw7HdjLDUI5fwFR7thlN01/9RNdPrMN
ArtfOgBiETOwZNWaBk42Y/MTKIDU3K2xuIvc9sotYx2Z2Wp0jaTwPKDbA/STI5W/ohFe6/ybx/D/
buwdYALeuEf8k44AJHprDe/mVPnzsagBdasJZ36x1qguE2/s63Bizp48L2kx4vDHPNO7gob1O7og
58Cw5YXzDjWd0O1JbYR688z61SpQv6vpLMKPjkw+TMuibsQgRGFIn3dFORNu8FRV6F7YEDjDJYKS
Agpfoi/N0qpLdE6MaxrwjP0eg8/GzmkwSSpWMOgCQpzpZHrlcusuq7U8wFZUkhYr1bh/aQrgWBmS
nnUoKCHP6xPA59I7MgE3nVh7N5HozxATNwvjbAoQKe9l9G4AP/4jng57XnfTDECyUenGP1pg2KGa
2RDfuCe/m5enrfxebMFXRRMrzKCBXQXKSf+ytJxUy0T4yvCrHEONn841E36nyviQN5MH+FKCF7K3
gsrfoUiqK0kKMQe6kCnssZV6F694+T+FwdaDf9C91F1dvjhF1RkJ6lizoM0HEjhPgsmf5H89rZgz
ffwdJKOrxRun6HJ8Rfn6Oa8jJwaFVHezyYHVeQGigOEobVbTqFHx8h/uIdYkEeuhJVw9g5jLe03a
zGOx0YtDyg5+DPmh7nJ+7JuiSug3V+X1GJozhauRbfrlgqi/7q+1byclhXZHxkamWrlIfrIIXQ0g
Dajifr3/STPY0Fp1eAF6yeIcxGhw/LqO155ur636pJZMm/wPjaJFlQ2MA3qwgZfv2Ms2doGP0zdA
8yNrWi4JcJelN2R/O6KIrQujvA1pKMQwrar+IOFeBPa6JPuOa7Te2O1kV+UPb7lHP150dXBAmUXS
jU+DJWTTn7D70C4KAbzBaj6p34EaxSaMZcFvxfJFKEGldWoEv+K+uVK8q7v11BXr5SLpGgPjKSXN
6TsQmIBylAH50gazjbza9Uu44aAOKiA6EsZryAKkBxbt3sR15wNPr1T6NPeRBaPfSKMsv8wnnMRv
yjVxWIa9ljqWthp7xiyCJJLjJCMXejp/xoPAzggnkxoqweJT7gwE+LD6Qgg/gzazNsANKQylXhCI
fQItiyshDXBIQCyaiM6ezyFeJSfgvJ/zdVx5g8uayLRICrlaE22pqpE6KWxRcN7IdsJt1wNVwunf
Nejxwx0dkY5WF7qWDuAQi9kUiu46wVSh6nji8ger+c4tOBPe6fHIS7eNtbqvqntBdH98BiStsH2V
NaAnyv6FlaytnDTbc7xqwce6Nw81HsfDWzxEgohVdjJQff91UcUtMXfLcERXu+fnT7PdR4he/n9s
vfbwYRt55A7UjVhVGrFpf8AeT5y7HJ9tmToWFLzvkSqgzTl9x5TBToxcSkZGNkbxE2Z5qgOFyRbH
fJ9UnoZTgsZylpqj6BCqKCPzJrcJB8Xe6OO0XMGzUNmY5PzwtvW8Yvg2AgfGhttd6BP7lK3KZEwV
0W2Ysa2QhuraspfbGhp7oKGbGC84ayCZw6eXhW9J+5eGs9xbDVM29ypLTpdD2uhao23l6D95/Edq
p+jnYlL0jeahX4Nbbonylgxhfnh1KyXmOtJzBMh1N+PcXwVf1GqzkIWsqjCZrcGhKl25H4mXvSb7
ZJMWezvhBn5+ZtgVuA7eWy112XIDDqWwShbcAMry0pCl+OWFyyDlc61wnoxkFASRwda0DWQhhjls
uD1hsxqmlItPnPEyBMQUkmtxlPtVPinlmo6GPGxmb9tIZ3AMGNNfS0mZA5etHYk58GsIUav4eB/j
y0QI1M9WcHeG3KZlxNXojZdiwsSIwz4N3uGW6ql+QJ/YKJb32Sb2eP65ltSSyHYrgSz5+Nca3xBh
uY571vYWLv614vH4Fw4HXCHpuCtnTepOVYPfvo4rbpLRAaX/Z7GjO59edJGm38fXmkVQ6/OhdMEM
ndju0hHFJxuv7G9VrGyMQyzUlf9asoQ6zqLZ195Lv1oPzr1Bysl4RckTGhfF/fbwDgg1/uP0okLH
CTaCwb6VjnaI1Zr+AnVKvgd+c/oa2pnKBXFYeFWhXs2EYsaRRZBtwJc2NXtktAxHNosJPl3QHXAy
ASCT260gkXCNPxBVmotFRNNaAXsZEnfPImlUjzA+uxM/kdJTHAmq4il3x4c4g51JA6H4jtUFK67O
Y0xQZVX2eYLZz3qSAquj3XJwJMIUd3AH2wVslZ0pQyojIYG6lZW6CejAOG63bjtHLfkYAAERLxNK
l25a8u8lAsL3cOvrhGwZ0OE2wbrxjmrH3DURT1wuFNK5XC6kc4AYo71uV/S+kKnd/TuprZsOAbJi
+FQv15KnsyURcaP/3uSMEj5CKciQano4HLhyI2m3KqooINnXEYg27fWx1CzAdvcmNWwahWX0iaJZ
pO7s5DbhPgU5rV35omKjyBZXJ4qvRkcA/Eap8ClFpm7QhMfeixmzxDCWZO91mhblipmwLOcj8JKa
F0z/DxypG5fm1fYRfU2boDJaaxQefsWvBvA+1+XylitSfnh3LcBNq6IG/wVFrLqz+RePqLMYpBQM
yVUPkUi+IAIc4TwpH3BEFnSsH3JjU9ujtNJRilSD3EIjOZ+W2NYbYEFJgODWi66H5zPCj07ON0o/
jV0+L/M9J2h37CUUlEozTqDyeA1OmfFSGq1bay4u112QoOnjc4usp24soQA513oLl+ICqXHCi/a+
p0zeVLKhozpptBHkT+E8wHHggphX3LirgJ++Rk/ewJN6jn2x2mQxK9JJdodg60cHKjRTVByx4LUa
Y7v5/1PuG/GvjZLl9KWFESrtn6ibzCcHRgkXMpoIpNI9GLC8oIywnnucvyHRxWkiv/Gvi/1euWqb
9Y6s2Zxg7PC/Ofl7Wpf3fNJn2XNStEGaklH5R/w+kMclCxZdLGEkZZhfXiBeWVjqBcKHCYTFOB7B
+iOrGGKJqGpb+nia2dQzpLuiE0yBcQnUvelTnvXPHfAHtg5KiwUpWvbaMeGwgpq9WykYbCHyaqmi
2UqNBsbr2DavP1LQ0n6iU+jkT0CoBgEh2YWQ+4mC4WdNpcyPwUqqIeKUyuRqnzKCdBsOMITqHObR
BuD2GsBCNjcDsTOS+KoHCF4wNwEdUQxEcsrLCSbMyZjzy3m/HpI7Ezln2SEG1dp/b43cQbBhTshE
s8+5PRZ/KS98OAoYOpZQCakxCULrHMEABakMsCacr0BjeKvBNuYrrak7tcrhBf/mHqu3O1hl0iSb
u4iDHvkRdgy7/MFgaRb0Vm2i9ehv+kLbMTFgRrocwDwBCMylKkkumBEa01/Bz4MI4YGw8XoxqwMH
hki5Kb0pUgPzAOqU1q2FAMfWrJzs4ylFPrXij8wOeknV4baoHgJ91s4eW/YIwf7PPIIIjhAGM29/
V2WDR40TM5qXTrePjvbKUZhFUm4VdEQ9SFS4g6s+jbBF2ZeE4CdxLqeXTv7DVqBCz4NHE3nkDR1O
1iJI0Urz0KeJxd9MoaxSfImlHXZ+1M1gSXycLeBzENGBwklM6Yi6BR8V0wXKJxmeuI5Ckw0xJqCU
R8+/HfjAcm/3i2vsLvYIP6Lx+cbrcHZ4EZH3QuQwqkYFKtyhI+gQHujMwhQxfgkgSCN0HFUNkndw
PEKQWMhto3+vmjcL7ZdKbXotGiwODFCGbLEIgOcFd7X/FrIcBrqzK3bBRXvTYNyfNxRB3C5C/c2E
zZawLZ3XjTPmhA3pcPuqqLF7My0Wtmrcskts0k4jOKDXCBEcokBQxzNuKBiVqZpwIoj78L1XTjWV
fX23+QjYmEaajkUgsGoyGTVT4lFH/SV2/YAPlHAtlAkzBLRoVeu0n3zqVWJtn0JAHsijVm71Yqql
5tqIJejBlJX9MymZuuCxslR0YhsQj3LphmTVebN9gWboJdQLMN/K23/1bbCVpYcEVaZfEU0gdL0e
8xQUNwkBO3LNEXoGTmMhA211kkT8Wo/5oAtKuTIV/xaDWTZSPmKSSkKtaKhW/4gY5cyfgablzV/i
AS1dPaq/bcr3SnXWc5o6XDnO2vW0PZovVbyrSB5tVmhXLE62umrUeqs2AGVT04+R660ec//rsOk8
TWfIM9yko5qzz8DFn13ozKfJRXDfnGiEBoHfqCZerHLGpHDPsWGqRBO05pM6fqOKzf2ZABT6lvSu
7biKyFizC+EZ5Ib+Wpjt9Go6+Sp3BpehewKhXM6v9cgrcFCzhaeLC8rgQ4AvAPUcQLFLjx/tfEju
qRwbUmKyyQN2aWtFGkcVXdEKFpSZdeCrSZW6ME64LyakK85BV2j0QjMKnJXbLsp8jpuOC4XaselQ
uQ5BkJuq5QwA4ED0IycNcYIf00dVfedSX6Ynm4Rr8I132O6BvROId04QZazgu0m2QRJGk5ZeDj/U
QPBLzp6yXuHufl9kcXkB2fwUMqyOCdc1WaEZ1NzcyzNvt9nDLUfj/jJlEA5UBDqwRE9/H0o7zOcD
CfgliZn1bF+3ZLEkqK9xSnLR+N9VuM68aBKPKTiAhMwjHmXq6qK1g8ci9heDNbUw5Lc1s4qjEtjd
Nc8taeJQ3UXBJIHDd7QJoCjZlXrowE4UtJ038ZTD0cIlrz67HIqNzpraSqko3fz+t4+IHJAAyxcB
L9FlR1jvXKu6ShPGtucr0WrnOMmHYS4NTsLf53QTgB3njG1lC0LdiRM5MGqvZRxgEVrwjCn3eJ3/
mqoJWm1PtMB0oKsvUFSTuaLd2Dbmh4hCjDY5UdmEyR7mILESNWhUNjXM3wFhkLzBftYFJBtmcFgC
e8kkBcGDkv1QFc316/UuC1MPfiF3M9WDfU9pZonWIvR3ZiWxYbnb60Ft+IBGjBKy4eKbN3I6zRxn
hfX6w2+LUBXKnhNc46fBBXEaKpC23tKuy4tfxdMImz3/3J9B1Lefya8R29PehSNGmN8JhzBI7Dj1
RB6MhppHPkRSEOeeRFhIXIf+4ZAhk2uzWu3Rkb2ajjBbQOvUY032iqiP0JxYXtuO4cjeUlZA9ohl
X2Jz7XtrkXYx7zUcnWaWtzDSDrksushEuchYhhAVdzcZwV2P6rdI/jPA0WZ54GPS+CxymdDeF1+F
vE/rGTOnfVQeFiVdY1Pe/8IPNbz+PsC137vuK0urJ7fjpwIDvsUVyOKoy6VE7xii6wKtr5T64Vb3
U4N9tEIqkGZLHsMwROdo40e/ctVP0jzlIUCWldzRFvBMnyRRdURY/NlD6jW0OjX7BhnKIuI9rLuq
cINL1LnKP/qQmNYMSnyjXtRDTeAotQpeIRZv/FfxQNrg/g8TpOMT4zcauaxBuMFrd6XNniquGh2W
DQ+NzNXgLlQ6XX3IimvFALLzYgqxO6ty+RCaFz+OHds8xbzX8pqyJG+SYDhdGSF9Hcclml+c/2g0
pmL1+PY9tyz5cQYyKkwJAyeEY8SQxfMGzhbG6SzXRqDFz1swDcny8z3oKMhlG6HT4b4TxthJyGc/
wEEtpoE7z5y49TgWMJJnAIC7yzhifaqMux3qcPWGhBwE0xfo+YHCWX0tQCnXgMvciZ3l4mkCe99a
AsTk8vgVz8pqHiWSSzL3CD3heIr8yb6cbPCgYakooWg4XBnNbWG9huCpFBBSzui4W8pf+vCYyesk
23x6gPUqbJjz9N7lUgCm5miOe/182brjbMy9qhAlciacwoWZtMrHmIc7Wkz8WF08zNCmGlqpDvIA
xlMWGIEf9g4tOMbvizqb780TzpO4M+jKuVrtLrDtTT/upo1EKq6o8rMF+uEeeHR83kZ4zXcZ/heJ
dVf72y4fnKBOy3EuRNdjs704k0DsGe0c1VMIeTYTmn19IcNAQl2HHPlw2d6R7QCSrLoGInN/6n0X
k4k4r0paL6fhyneJW01dU1prBt12u7jiRkynA/LwQ0uTmFS6tR6za17NVIBF4iFa5UDcU/Dkz8ko
/9Us8lW7TLfFXV5ZDYV4H4MYcQrZ8kE3e9lRS4AtgjwD30O5kTHQ562QIbKI+25SzZ3WsZ7abA7a
2hIZNHwhPYNCdF8bg44fhgCz62aXbm8MtKR+owX+DIDpy8k10hiW77qviOMeb/uJd2+W1XQWgOEM
CCzKh5g4V+0hEO9/fYWnfyait/z1Jm5bzvKnHBAyRDJGvxmVl6KJ14Uw6fGwT/vx6bGesOAjKrYz
ox8H7weNjsHO72f1Jpfsy+PVAGJpoU4QUA9S/J7ba72MCRjlRYrKPY1gFQoULCgtvUC4lqkmyJ6X
PNJpvPsrFAuQQA0hH3uj1s4aL5FEcpOcajZURlWm3Jtm/ppATlpgx1OuKxcvOASYVDWJ/pFGTxw/
EIfIP39+GqO3bzDMdfCxSDw9lQoPAGa5ZUteooBAKUP1pLokxk19lrclRF7y/6Jbr5Pz2wS3XeE/
qGgGxOEbej92JzskT48Qr7Swiiz/o4ZYvtvgxgPyN9dRtZadM9lNva46SqEFHpcWmJWI+zfgC713
4M3JBV/7tKTPRmDMtdsdujW9SZj3wG8NKDMkB9Hms9XKoflW1yZ4a8MonnRO1oMHXtNqmcKjTG6u
BJalt1aOWJPbbiSls8aMEONEuKI0CFUfp+M/u+LwCMcgfwWMCT0Kq1eshjY2KUXARTHGQo8Dbkd8
SxE505xsRV27ucaDSWaGR4E4Vx7lPpA+MtDAB2HTaimddAsVb2OEK2qQyR/26gL6BHBmLGDYObC8
U1wVYCtP3pwDLFw4k+M/+TL/VAboneN9XtI5P/Hha4FS4euU1lFqylwV1FLQeKSp/2ykCGyRV+/5
YOSnXQU+UsBxZGc3tzKoLzyF+EBER5OAKwhZaS1Vn3leM89FZ6Za4yuRmtj/LYMYLCMvAt4oXrBd
e8QAzING8CxBTQm5YHPUr3EKkyzncOPUlBx0cpvSToYDG+o31tfQprnj0A++OUoMuKUoY+HHSnVB
1VVUjAi3ofSMD1Xg6xnOr+tcgMSw5xb/q9/V/oAU/Au66eYWz9jDNrPUnn0SDksTfrQKjgwNWPzp
CadAI9Gl4TtiNAWSju8a5sdLJEPfCN75MyyuFDUt/4EslHHCVaQ5SsExC8i/SGCA3l8b/2msPdaC
Vl0I7J4MTYGRvpjSA1qiunf2w/12rgX60ouPet4G7eBsfZyX+cAHHmPbDX3z2xpaR9bqndWdcfFA
posTbN2Id4l90HfYKwABkDKRvnYfCdQPHjnUFjt+LwPgtv8bpLYz/zo3bdk6AfS/i9uVc6I+kvoY
DY+bt4NKNLjUYKsNFDA7iFBidoZzK4p/OG0/fiLwRzPYDb1p+ETO3AeRNgEIg5B1uy6dbQ+JocSm
ZBHf7MhtGCJwYhc5oGw5XvU+v3l9PskRPoRZMB65Mlfd8OcZCaJxXDNRFBNXzoQ8+kTQGHKFGkJ1
WhZDtrOngLjad7PKmcCeAUAubc6iCQXIGPIxKniYSeb8MT/XQmq8hAWff1bDzHu/uDbhhzDge4gm
eltljwKb8OnNXyBz/0qxw4bL+7MW6m30ISyZQ31EpeHrmEYS+DC4aU+FEvy+5flSdhDTVZr/Tv8e
/dNRLLwSGmS1GNsFQHjIHBZICdEV8schqpF8Uaf/g6t2fV+MhvOsKjuPa0Tk2BbW8fqrRoyhPom8
+g95G2tM/0JuW9J9xWH66Xg/kQGVadplijkfBZDjQP9gnoxqJkkB2+Wa47R91vipfL9ZaSFiwrPx
xXsVmaZrr1P8leIvp2PpfhFXWdskmUo8UeSqgpi0SfT5jGoiP6jtSgzdJFGbfwCGlW/I4kaVwmAO
wUXi3FY4a70puDg9t9ANsGMtqvG7ByxFx1drOB7gglERjwGQ+5axM3sHQytWG0bsTXxroLoukesr
a6j2XfcLtDkI18wUSfpWlp2sqd98Pc53UjXr/gt7P9j4+IY+Q79vzGYYblo1xWdhxno9jitqq32R
0YmdhpUi4rcfw5TqglyLcCEuyzGgMEWGNfU67Q06kJUqSGR2Q8V5AbpLS5y6jEb5To7GUIV/fpqn
L3LiFxZ0Who7E2tOmcBMr7zmohZvOdJsrvBLghkc61WHLPxQvmcCfye9t9bJgRAhBjBhXRpbFztV
CL2KBeQRcxlqaGzdasM60kJEapuY63n7XZGa+CqVUXA+l7NC5RVfGXU165XwshiHGHdNUax86JOt
S38PmPKiMt6gvUImlqg+SGZ41VVFHwZ2Yl03PP/meP7715lXLCorBOMlLOU02rliw/Ub8QkSJB/H
C70sUeiDZ3JfbmIm0+aj2Q2qc+OH4z3dUQ1LMF4pyH+qPLJ73aKswBDHdklKTYT6471vq+ZWp8xc
CBvBlsKomZNSMTFEOAqgb5fc1wBgk3BN1RTXQrog1wuphfVVLqKuv98M5+dIS155Azk0X386OsZA
HKqi3/vQ89JDIq/P2beZte/eiz5MkupdqgWKIYBE3G8YhZ8OdA/bAUilTemGika684r9gZ9h3ugs
3AauYRiz9B/kOHZzYUW3skYs2kujYoL4ogYah5+NUSR5r1bIZ+CC1ux95Vgi8Nr307acexAYJBvv
Y8Xc6zSIb2fOzGObiROoR0radg0smLwmm+nuqoQaymjuDjp766oXQpEJv4Ah9mlNKSbybj8psNyk
09i8qlke0z2ZEmBlxL2UVAckPTgcugJ1yH4PB0dCAW+jGvX2rLU8mglwXog45V8SXMZE5OU7qvpb
F6PIDDTqgHdkXMCBsTxuAQnE8zNpteXWWyKgDAjSX9w7r3BZo5WSChDzt7PpyX763p7V0rSphebf
4o38n/vdqOyfqZRFC2vcrZOS9TKEPtDli8cJoCdMiEh5//kyNkxlpjNH6Rg/G+PEi5akRcybf5Wg
2CUOqY7zCUsNJK3XXW//kWto5jGsu5H6g64gbZPMom28hJ+i0AMHOxM/e44dHXslQGdj+RIf8nYv
mRoCoozQ5Wa1hxBRq0shdpcmLRnNGFPS0CrwQVtRlOiaUk6Px4XP81WIFBWi/4ehQyH7maVRZTi3
2ZE7I4B/sBFxzB7wcp6xkTc+wqDEElM7qIEfdsP9FMxoq5105VhsxbuTXz/5c1C2CBkc5tH8UYOG
ltGpNGV9rCs2I/m5ALr6qCOdPvaPmHD9ABwAfPVOJn65oACL/wR78V7Ktl/RkJvdX1Bc0+J0dOKW
HrP7vmxsjnWhVQQuy+2l73RaaaYWWhu1MLeYNFbXw1kORvv1sk4n05e3RtkfDWGMTFfQKtuqRxAk
7uxzIF/HKIpRbPQJDqu04BY3rThE7SaP4MW1qF2qjqbpXVYZ0lIKIFiro9wtbv5kDbOCqFDCFDy1
+kqynBF1Pf3xtEeMkIAN/roFismycJuNZHwlv8Cn3fsckTMtadwpukSLvTu6RLcppiVnAty8scst
DI9w9LqxkSPlu9O8jA36Df6idn2j9ek9bSEYVorbsvg1Yn+Og06xoM+9AbGUuNMgRliHdq+34/Qb
bj6zLykwnHrK2MPvp+wEuJ2aENahxuV5qFWNRGQkGIKGkQd62GDBGdQ9ttvO6zBrngK0ZIOC02Qo
df78EQ+Q6Ymutr85LTO8Jbi4+8wZWOGgcdOL0+vYbjBzau79Z/BFobf9lbw9ffKC1fJI7YJHOLcV
Vtrk+6SI8PWAm9hIpwuc7wlVhGJer9T7ysuUCZBq51fM0h4tJkU3OtnukPhwQgRBv2rULroWAvio
kKKqKMZCUzZnR0n7pC625p/BmV0fjTTQzfTOXza/lBgx3mYYamag0G/O8n8Su1l9xjvN21eNM7Vm
WFqz9L2nUOavqZstNgT3WWD05g6Phgw6K7+6FsR1lb23phfMxHy3AubZ1podxxYFAuzPytnfV8KU
+uMMfbSVIh4+kN/fVL7u76sJAQU2KrvXyfaRihIyYxmj7AAzUQgogC4+0ZZwWrFAYE3tRFCF1aou
rpLmyb0Ss+KpGIQWbKfMJMggwPH+SFUzMWPFf/TJ37QzMF5kludX7Y7GT8WgDo8kDnVjf1lIDD1q
5hQJCe+Mr3jNCqMphq10mQyQuRbadlO6WHJHzyLGKii4aGi/JLFDfC2yEuj8zx0n7rjA4SNm0qh4
Zg5C0VWmPLvV7TvZ8p5tJgm3o1SwKRb5nmo6ATF0rQKNuOU16GPu5futuFMCV3mk2fcG7//JJPmX
BAB+RY9EHI5qgVRmV051T86CNIsm4iTmIUKY0JopkpRrMrUvQdw5wCvZDX/fxh5PVbx+ueQrm+4z
GX037pIfv1wJsDa0ZS6vJuk5avzuc5xC7kRrZSqdLO4DX1kN4t0K34cJDgrbDyRhIrIj+oMIN0kM
yyB6HIvAEjiarj5q5+joZ+VQJbOnS1vyFGjP32Z36Up90rCs7M+zrTodjOJyvNqdLuyKtPghSwk3
luSTO3iC0ePgE7eTk4RGAmH1+C7xUc6RVymv106bjMLn3q1WurSE6Bx9SeI8jQrRl0ITYIBB1h28
PE5lrhEuIZ/5ZrC/cEzcoXQeKshyvHoDEtSxaHIigXYOQNaGxSfY7QReujjV4vLvxU8s8JxfipQk
8g2nq9/rOFG96+RTftihly6JRtdHahc70ERyCyiAVyggAklvZdbOpD0QoidKtVqUbYhKN2R1TKNU
VJUpIH+6AjQdAv7XfzSfUHxNOPcekQ3XgYHWCAoRTzg+MSqtIp9dwiwCvAsTcDe96ZnSCKjqh6cN
6I1F4dpkB46RZ3h8RmcyUSLhlYXJUb+cLS2TZC0dCdHEAOPEceasMJv3mUhLDtwhEDdcXXAkTLMJ
BH0pVFReZ7I3rSiq2HWRk3ESWoL3JlA6AOSyVXfp9GLvxwGFpsO9/XphwK/nQsKHME7UaQnIhxG/
NGb2SynYjrYrJIm47WSBE7FIGfb+WjFt6RJJIPpCe0cTeRZQdbzu3+vRrMJhPhgBDfaQB7FLF8qr
99BXlnb/1P+OLef+r2Sj6t5g5JUVq8hMpOaw5n9jdZgR665aN1EX6g806E0A6N7iGe/OVgIS7COX
Mgtnv4xw7szj+ZwmMM3mjk0xxtlhyjvcJxyudxjSEkaX2kh5D/coBJQJWOnoXD5Tp9sObZOs3MIo
OZNzZDtNJHaUvSvqCqA6/DrnZp1+v+D+snXIfzU0VKq6WAZMaftJUe5bzrDsEpOooPoJZ7u5/UN0
mwTQS1Qm5mF2U7j/fZUzinPnNCZeoFM/p7gx2LClachWMVYtFJ6DjQcwzHFhPMuC2ojrYasAin8E
YZQg0TFk701y1kAKQ9JkF0+5Muw2wh8lb7DAWaYiEX63HpVe/QTLqObnnkPUhpDxGCO1VlYs0oyd
8Gxcnz7RMcOTzKVcygLYTmm0RSMHYgnTjDBREc6NbuqAu9QnsthtDjfyq1LAY4EmoyG2u0U1Z2w+
8eTa/spXSuoJQCCZlCxCSUuc54+xJjek6oqrpLc00NFebp4DWimWyCuYdVaeyNfJdVFlfQeoo9fr
8cjgjQqhxk+3vRGKqAySoqXsIsEOk0FIGJG7EyHJX2sdTkAL0QMiuMCZtp22MSPvvdVVwbEHlYF3
iUGhPhQoub7A62c0R0vwHwBrjcJa73Z20Li9ZTaZlvi3oMfA9qQ2RWKfqjKOSuIIJFDNgCYkh+dB
D0npOOkpQrSu7YTKKV4fv+S7pz5yyiqXNH5dXJdr5xdknwFkC6VubREWpyzjqJiOr/al53Xg9IPD
cR2B8DFY/Q7Cpl399oz3rkKcNx1ljAASd03YzpP3/xXKT5/jqbcHz37sbbbr+z2Kq3UQ+zaTIwo9
lDXCSHnLsObpFXGxpYdDK2QUNhIpLYKisxgBqMzWYBGnZWWUIdMBctuE9sDCEUXbVhrYbapkyj4J
IYFcIkBctr2sgwcJ/WCHlA4YU79MsvqRsAMrT0euwOSEoIoQP3v+xsA2AjpwmaLXEJ1pQ3SpISbf
2YzXm78D5LjYoXpTWsJ5CHRNcAsyvDAyq46is5e7tfEu8Qc60inyJOXXBzNJvnikdjOMjDmCsYiY
4pMgr7VqiDBKAXbJE/Q0h3nmHu03FvlxYUynIgDLh1qFj1P2iTmrShX9Y3ptG+47lUk8CSznXbIB
xWQYmdM2uGhxqV5DlyTHEwuat1F2n9eL2hPwL0TSVN+k00aZ5Fzv4ODf5E23xLERp87M/U4mf7wH
y3pAi8WCkVESnL8iMdgpK8dg9BLVdKqWrwCNQvzkQL8PpewmuWGpf7VTfeD9mHUAFFo65Tf5hYr0
//yQXKX3VLVrR7ZWZKzk2C1l/zr95jEEHydSD+3WfmL0zRxzvbhGzRGUNVr4RJMqcvRLLGC4ghJR
a0ovjgsJnjX/v4OvvlRB5bV+dwJhmHrLUKyk3WEt2z93Q/RLR75xCBj5zwKD++K3bnvSkG0DmSY5
GGTrtzMBCPfjhuKIeKxh7OUbOVTQ7w5UQT5pYsZSbj1/thDwhtmYGK6k+6aV5ZSMOsmwlFI/chJ5
fLpd/Sx3sPoZDLl8GRW+xHSvSl/rar7va7vspgTOpGZCcXzZ+TJgw1nSrgZesF5WX6joBbFn+pso
sRgFWyxOmDWkdM4u3Qqg1M1p+a1MKElI5P6D6P0XLGT4/aPR7Jm0KLaht4wsjmrR/H+HdDuBj/Ia
zgCIH3nH2Hz3j65lQxv7zVWCg2TqC+eqjV7RJ+xKkNI7Hv1mzZcpNdBsCJBOy0xPBeI2dCuwVds6
iOUDDqoym4EU2Rn0jgFTQx4L9HajG75tvrIib4f9wI7XhOLtzsFH5409rgsmuAjmgnPHFy1kiG00
PnV69yuXT8ID72eEDPDg8LwmZIuQS4Ll+aYEqYBOw5fQzWnUwtY5+PZXtUqAE5Xr95HjDpj3E23C
okDO8fRKMxySnKvF27I52Wqa3wj0JWcUWNIKUL95J5q4IkIlC/ka4QRvZQhK4eRqIINtEttl7UTh
Sm2TwF002In4rt2YC4AJsvh21nXAfVEL7T2L7HQFY2eYnajliPpffImcHEqlN3piN21P5XRT3QX+
tcMZ6IJQwxdicbFFi3KU9CtShBXM7XZHHIe1F9hhTMv3EwiKKPog5lC9N+FgUuVqz+bWKXE9ONT6
72doKL+J0zmYh6JZCkHb2ccCPY9E4ctztx/Cpuoz0mM+QkvnSsX+T9teSal5ACDFk42R8MRsf/D4
MTWzTt5OZkiBnXJ8uFd20+8PNC1cAmT8oY3WXWHyWDzIbAzieTUjRMVsqfsyXxUcz9Z8XVR4TGFv
ja/nyAhcVtMjbXXisEIPfeoDz7kinHz+6bfx7HotYpDU8iS+xvPC+YGWB/gQyl2ozn9+NanpDMg8
kjcZoaL/1ORNAetjS8xPJ+XeoBgdVtpeMWDF34Y37XdlHQhJQukbAWs8+TuRI4C0Lw/Ru/06fs+9
1pK3JwLyl9kppnyEVnA7nvcxNMTI4c8bni98erLFSXR9EaRL+Spf1qvaYpxkoLJhV9cgGbV9MIHc
izvYlYULtjhcnpe2FoXHXSDPpj/dQthicIpc7UI2wz4mFuYdbthFbHnyFlh+ywtkLo7TKOcaZE+9
GZI7ALZ7ojWPKTKcF+keMRsvQhAjGn8NFcRcGb/gZ903MDDWO922aROoE0zUzu0yAcRvLHdNWsRn
EFXe8jJ16Gjt4xOHsYqtCUR70KIKW3Sihr143HRzm3itJp2m0qTvrkigNrQzjhN85L5EZWi4PqQ5
bYJ/dQ9kemA5VBif+AEf96lm4rwTls/sWXrfUCxTPMtlDBn0Pk0OdtPfboRs3dCZ0pgpHLWj+g9A
8vHRQPOOZwhIAzM1FqOMLOjxSCzpspRwfleP49sIQFf6GbatM9aTWIAifPO3G3YcCcumj+28ZdYn
pC3VxR5WLOMqq1IS0276Xi2UPZZlRT8x+PvJ7WgIeQRWViCYtP5JMZjgJyXhJhjwNuXjgbV3L2ox
x6/iFjpk/7LNatcjrzmvN0Y/Q+rXh8ldrLuKnrZfyqtXM+D9mSEJueLzlARj3qXjmAWxGgfBancC
fL4NwM6AdutIeDFug7jZgqqm8+5nIHfesuxnTCZETLTUB+pMU2zgIOUa4/5bGBjJgz5fQ1AjapLl
Gyr4x6NO3q6/PhTkp42ZUDsHkbIUrSr1zB++R3KpVhqtzmNJ/mskRF+fzBLsUHGpQEmn60k/0d+y
dbykqTptQQ7srbmziseeIhBt3No1ROVRq3JrA9+NSLt5FG2qOlnru23bFhHXLBaV+Udh+AK5DqBr
pKCUloHZFgIjquBtFqnEISu1HF4S8tyPtbvvdAd9/OZr9uryC/91jLDc0rbwIrnpiwJoMVCUdfN6
DvaS27RO3Jz7leyYUPW2IinXr11mVAhHXd7o2zUAjASv1Sq5ILNLdTc+2uCmlRYkNwMLrqn0wIT8
5nC3LhKbM0ECSE2cmnC0eoUwsMd+VmKVh/EoyEv+FSYB5eaHeDsvlthncI4iqfS5B2goI7jdBgFR
9SAD5XOtPRGOdND46S3PeSCefeTd5zvvvuLnPWydh8j+8DCVIBlIUp+5lS5G9n6PAnZIj5ymeDUX
CzwpoEydIELSaHNg70W6jqd0vY0P5bU3+46w/ohexz3eI9JoisdaGPWg35XyUwEuxZa+8LzZ1yOW
IKbYz5ZJqJZBXRuE18Z40fJR67GC+crBlMPH56I7ajcxX4KUO42dSuaf5NVl12GaSdVI/h00KXLp
W5lkoQVisCR9QLGrpekyzy+ccGHDMSXYegt4Xr9tsg4JSg5NkOW5n/xrXW8Pv+JfaIEb0Ouso1Nl
KB4g3NJwW1RF75LNldFEnKUoTeo2mdJn7qVc1IU8Oo0jf6e4VnppDKfV1dk+te8lijLdkBtL628k
xn7K7hHm/D75+sX7dK5nHpRlqA2aJEdAc4PKbHd09F3b5ZMmE8WcqOvgAcEwLF0cXmYaUIGmf3/o
n/VsnHosjMmYJoOYuYkwu2z6/jBd9anb2PBMXt6K+zSAd+aqlYU8ML15QuSch/x96LY9JTqaACOW
imDz1gvstRl40oW5VlWpT6JIVs74ZxhemspgODKxCSUaDWc7CRgSjPkO6Z671Y3k4+bszTux2h4G
4Dx+w1TANwhwA8a54+NUMTyYMUU2qf/PblhsvmmPVY8P5MJbx2VAx7mDsMuA/wGvSqxqdkegVSf1
6KX2BFFNuQa2zupjJotzmMP7XydFVBPtVa4iCuabTinAK9ekKT2LiAlpfq2teKMGfGL8GPMMFSyl
voExg5KqO2s5vEG1Dg/tshc6Jda92B69JZSv1IY0rlWeh8vMeyP5clk6NzKRRsQVnQX11tgbMsvX
kq0uPSwOONiSDj3ot3YQ0VDGo/bDUOlKF0Q8ttv+qNLZ5KCu6OfgnODIKxzZk30nwtP4lKJjFA9I
Hro+UiHWv9wtu02QV+zL3EShXj0F3/jAsHghsu92IepAWcjxO5deanSwIgqTCU+nsIbLzmrLcI+F
UOtCYtnOkCMLvVHOBOTyvCoG32+8ZNfUKAaZLILT5FMhYr3P9c6U5OUKr4kMOER/1M/O/FGJ7mRl
/le73NahirSCiXwG8MgERBi2zRsEZvbmviT9vm9m1MQbCooOvro/kj8IURAWRtzc9qwcxXfmhetg
nXwVH5jJQFMFWBbhI5YYAW01HxrG1p4c1Y7gmEfRwrr6+C89PNN5ykqtuB8mMPpMvb+2S987UbLy
dbi5MBpwTVXMDyuOruTDomj3wFduWVzD6R2aFPE6mecsMKaiC/lHiGzPY0XItRGtTDeVW7pGXDk6
RyvEhm1H6RSVsTBDnqlgwf1oQkeZxgQ7fzIOgAjioANcEsNpGwZvGis64fITYy8pMee+50kMPoFr
ojc+tQzz0D1VgNNYtFLS+IfRdojSBINTQwsQDOlTPU0atbvdJMOLIoKqt8hhEFnBoY2FBS5sTo+r
GjaoP1wCB0iq+zqT1MIKmdhHaHBnO/LZ2xaqcQ2y6i4jbelbpqRLxkIHkRyYbvGG9cjCJ+bEoZpM
QyeqEEv93z/ynT5LBC61A3Lm6IrIV8tV5XiQHjqDZq9WFXjZbQyO3O3KXL7ukoSyZFWsrJA8gbyR
RVL1gDOgLde2gPGF3X9XZ+2prU7wlgmuItFdK6WAyrRHP+lgQmF7JC2x2BuTolQLsT68yYnNIjjx
eNfdAvc7WhQEPjjV0txc9RTQYniaTZXjmIvCVRSy+KcCpQHxLhcOE9qG+UampwwxtDlDDx3y3mvC
c88sJ6pPZhaE2uU90NxvoZx3XnUtpe4DB+8lb68tDC+2mpEHXiRjJybOnwudBI/i3D6CqZ12kGOD
ZbpRLJByvzpJyojK9p3GEHw5+SLzBSOsjO1BP271PVQ6mdapM82kLsAisLJO/stZQSNr40uR4KMO
xdSAtC/RtpbBeQbeUK+NH3JCkm7dS4vFht4ML79hj48XgulyFqg56PN2F1kqjWGOmh2z++qSpnCR
kPX/rzJW9O0v+WQFw9dWRdShc645M13YlC+Nyy3ozGkJz6WMJcQ3VyDNoJMegYj7IBUe60v6kwtS
osHAZcZjzOH7Zu1L/F1tzELLoYjGdf03S9efHY3tph3A7MLpe7+kc67WR/RmyYKsBGO78M+uh+VL
xAHYYpb+O/N0aMZyoLSz66zRnGdx5q2kxbIl7mZSGSPrfij0vLZB9Fj6wtS3g2XlEsuXmGGzUg0O
9DWyby6w0WC5mKkfzrJVcMVkhkXyv9vhaIIK0HfJQA3VfPjap2oQYzF692tTISKCZG6HjKhWJjD/
75qXFqzLkUQ9l3m77dI0P2FWns8t57dEKSA9Q/m08HdXnh3i7S/sv7yMhhlfmllJF6MHt8vCR4nj
rY5esz28L5WW/4FO/JbzfhCrDH2xahn5D1FPq0Z+zTLhan7PFakE1QZofGMU07tnDQt+Q6Q/smki
X4CDmhuyudr3vnyeyZe3scbE3W3Mb6ktX0TuhPCiXiw8oPNoOSGjawEkErNoI6An242fxm9TLkow
/J5A4wYaRBcLgj1qBvk2wQMt2agfZk5/BmO69fYcBKq8wZzAB55ggE03NPJkwyE0FtiI5JE2nOZj
eqiSpjTbRv3fboGkIL7gUXqKKJq455xmSzL5kwEI39EHitLHUaCBzDpLy0u1Gjxb+FGNpFrU0gV0
9LLVv8SVcgLZb4IcU9JNRH4dXksNGPIs0H1UBGOJJKcjymc9HQze/HtsDwDMxH/67x2WIXMnpiIh
5fjS3FOfFCBqR+cfixUZQOBxdZjSFC0uOvQ5xXbGc3dOrlkOb8+KiweLhS4HoA1u7QGNq1D1qJiQ
knny86GDWyTuvhwRELhkcHgrr7kB+RE2aau9sHUIzs/cfVs7H8VI0b0PSN6OqOMrwQw7NwRzUify
hUi/BvxkxfWeTwYsBAjeZQNTyxVkVA7Vh9GiAUoFyR9Zu8pRztIufuL2XHunnqJyoapMNi3GnfeJ
Bm0XmNQKxPiIfht7nPZbiEdOGj78C7IiiXETYXPoZbM4Mub8wC01Cp4+pbYc4Rx6gEW3vYLWNfz0
rfKkPDDWnmfW7CaLwb0Tau5EFTzyP4ifM6813PXWwY99hnoQ79k90ssSuLgI7DjmV9qxv8DuTyza
ClGoZRbQQAJACWZqB/A+PSTw9x+4mC72lY+8UqIrfthBrA1UjOdmv/Xruj1sMKQiHYyrma7ngg7k
1RvpM3EkJ/KyF4PQp28rQfphRTBf9u2FTC5oB0nsPTZY8Xe1UCoVn6wWkQu1aq9qEPAe7VNN6ZIH
0hTu23XYw4pN1SALp+wo3w31ZlUIgu5jmaLL0i7Y99MG+mlD8blP8JhvO/wxDe+iwX1plnZR2gtx
I1NA9f1jvCae1YbvN42GGtzzQTc/o6mlimj4qGvQdrTn4K++1IHKSSDI/ley9qHXTE5uBhGhgCGO
k74D6bpfo/EX+gSwiCGRe1W+DYcqr7s5COMymlsJ527LOz/EPPKJMoF4aNM/KSkBxgWN86Dff19+
ESyYDpMnTbVyV9g2IjOLkD/JYb0ETLuU8iJSLO7lmY8aCovw3naf1NnSZMs2yirhRUDWh9S0WjgC
TEhHI7WsLzpB9/rZJJSj+D6sb1oVoL66+24R3P11LDrZzFdfRI9cVGleyEfQF1acilcXPzizmaZc
EUB1OKAFX1bnGLRKJTO03mSyJNV47ZaT6hQ10OUyUOe7OtiUg7g6yDWwY4kxY2981XmgZm2CdxG7
+gdPXK4q5IgT0wwHk2PBvfYeXL9dl3kgPM+IxWHnl5/peEPzIUffMHY65W4MjXVxJxxAzY6Blzxv
XrmApMxXc6rMp7E08DVeTBQ4n0HOx5rKISrrFQ0alxA4bx3w1QHOggJYJAPLXfMj8iwktdZWoVPu
inCMcVTUzWvTYSjuc0XU3fbYMFC1GvZ6yzLT7I+aB2L2Y/lxaWy5Mww8ZPgNlwEWJ/EwOrvaeU0s
MwF8WntYVyXDMSh9HhXE0GY0Q1teelKbSgPbH90qoXxPXN2WxHQbuC5aiQJmVG2T1UOQLV7fjSwS
wi7BEZLhb43lqXMyFizmC6wGcBEl+pZngB+xnb8n0NTutLg7MmGYHaabdn9nQ2aEjYFbVW6D4V3/
1MNfNc7hoaannCmVMU9DRtTNl75ZgdebynkVDq6xMzX37C/1hDh5CwhgCfOcoSO2J6calbd+9zFK
GtlZb6tY74oWXrefbFgpIZ7hL9+oaNl6fijEuyF0ytD7hMgWwws144iJct4crz3gY17Oj3e+NyQm
qodlJ1ErOIxj0SyszxMKSUerPnCovikOOQN1upXmBAenYXGEniWwy4S1ksCjRiqzJWEucDtcgua0
XFGsp/vnW9/2teKF4P7KZwluFcMCgaJyQrQ8JvGQVIk81jXOJa1vD9+j/bxhcOFYEAUgg1OoDRfg
vgOF1mMU3bFJdV+hoIRww0HUf2GSrAlIr0ACuEubgz46CopSqaTqewPqJNgTyq2JXGNmrSJ3igH2
27yLGOWMlC2uUmNOsmsMPCr2LPTeRPrm/QmVL9qtwbAS+5t2l2Fh6a+xPBRVZ4yHjJWhS5mLtLFP
nf6nBOCID9R4RHDD7jKcPaEHT5T7FeQPQu9d++wXLmDGIdyiwf95lDwAOwU0mmG6KLIosVkBUaeM
IXhU1161mJX8Qqn3KusC+Zsyhp9l6jAXA6ZNvE3Tle1SWlvtC56Q1772Y4SSMR+JaF6NUJHTGOLY
RC1WFDN0TcukFlPjK6JH54tiA3aNpeG3Rs2idYu9MjechUV4zUNnFakS3M2wssT992qDMQGCxQB3
6KEii7RQmdUuQONxvszpaoqX/1x9tsJ0tpHp1giExJGgbZJYySHw3nQ0FgC3C4zmVgc4M6kXpNou
JbMJFIOQ1pNXKXDCCP7/ybe4TvvP9wg246Gk+qopsuPylHtRRxwfc1N52rzhVRqAUPwiPiqWt2S1
Elx7HYTG8R0Fr8r1NFrSpjHs446tsSaxZtIrm1R+VCbjRNHonQQmrtr3M+Fii5sExHaAofJtOuqk
H09GufVyGPSWfmuKTfzG7WdDBnAcEQLXGEZg2vLXxN/1CvId9jcqFNU0rKGRfrxrQIfNwL+jPT9/
HK/ax6sAFCkyIUsV7VwLMEvM7iLKGBbE14F+hl5TCAxOz0lqBAVYrHObIEnQPjal8pO3NnQyo2zY
ne8VhaEEp3pHfl//OqYE1ByOc/6CG5UMCDikISYYxGl3yi9Fxs64Y1JuQAqcDEUU0Tjo8CFePKDh
8PjkmEbd20b9bx1Gn/qs2BP79VTEqNRfS81RhRdwDRtuq1Zss4Dui7aGeOvvfQkMizMSMPG2bb9U
Xlpt7ZiqHmBWU0tm5AvmYvqsyqv0QDiMVPaK9npAb6ADxgING+hVBO4fl81JaFjSJna+IP06VLBF
o/RkUIAFj019EfNak//feWQrWczQbKvif0qawKHkcT/4a45HeFrn0e0oBb2CC5JlodMagRtmE3BQ
x0LA9GeTrkW6UkGVb2H6aGA7XlKTYbuGb7B2wDcUZqzOD5Ku/Jyq8tBXXabnXyDhyU7gH8Tv0KnP
xU7Lutnwz+lLkC1k4ik08HvgdxeVKDexJkUpqealjxoa9euCWxJLhFv9WWLEGMIPurM2LDKSPXKf
A8GqBxKY3NY8pcAq0j51BsgCwlJc7+XhMqF0HROwmc+RgeASXwchclv77/tt8WzPx+Ih7YeToO+u
WYsdrFlAyKw2JivCAHbD/S+7fCWpRdChJUIdQifBIWoREheYXSUu2qoMiPU5ce1UxwaBSIW5sJWn
tJoTt4L1DjPoZpp0jyTAWV0AcpPfSPxtnuMlIU4bSr1izJBfw13hwxsP/tsJrEO6XoipU167rCb5
Hpz6YAAvNT6OsvC9o9ceOy1fuFA6LeO/NBB0YQRNJJEqITz/fxuGkVWIuaPUH6Ba0KlSET2vu4ow
VrIH9dWz2QOpN60Sqm/BSQTqwZRcIDyn6bLYwKsdgc2VHEzaLlNNsoLDdxaQcrx/qGrGnD29wre1
sV9ttAIQgD58loSK+om0rGnpz9GgPm8Pz+EiiyeYJyaK2FwnQtBH3Ud0GACIFbdS/voK7gynq3Z+
377oP2YfGExGiSH5soQW5f3CGtuJ1/Ip4svvprL1bMDA7qvXlp437VylMgiuxYIcRTU49SOxx9YH
WRetuWk08aGmxM8N4Yb0A97JcYS/A8Ywl7KWfxrlwxEBxfmOFRNA0kjWXbD78QN+tZay0MSsY9bu
OsQebja6sK7Edb5IYQRgZOaRoSCPDUGgmB8IGwyYyTf8vaFEJXhNZs8kkfc1DK9M56AAY5IXa2mG
5PgZIlTeR4oDMSy2R3csjoHJcgYiNPQoo4O/un7XlU/9r1upRaeFaH9vpFXprMsr3W1q68wiAyev
iC7jrGMYsXjEAoV6Qi4IC+WWCKKMbk26sGwBrxajRJyJpGU2dX+1VKPKMNNEYpafXRYrWhpFyBum
+8PMuZTgvmhHrzdUvT481NKDOJBztJMQP0LclqaLMe0yLdW/VOJLb+sN/bgQDuGBj84bKYWEkTXF
zrbgz0pFKG1QjajT9aKBcV6Vitl944hV8/NEiGCaXvNlcFBcIH1bu92ThdPJjfnIGtt/cg678vJ7
HbIlnx5icO3x3xFRYqyH552LqC1SEdlIDjxtnuEpYzzVkH2sBqJHIhbbnZHEibTV3nwdtwVTvRUv
40YMxP5Q3gWKtVH4AeYS3qWtLglsFGiWDFFD/i4LgKptAmBqOiVU5tTJrRFe5TcdilDYgz6Fu/Tl
f6iWaSAnjjJQu0dhxcQP5tQ2dcyjUyN0lYLdG/TsVbfU1jFZGT7alpVyVQioif3nh4zNd6XVGGEP
ujrCvwHc9c/h2S7+pQ+lwe7QiI/g3JLuvxfyJpxgx3Ee5ckeC7UG3Q6vzTyU+eYwNllrHJO47V5x
E5/lg8EQQPvMPjqOZXWmv6254ZsjA2lwrRPqRz36rV/oxwHfdNkMxxsoqobsDxRqwe45zUcs6Ndl
exnCplc6LnrR0kMEhHEk18wRQ5EkJ8SwsUJyTQoaJ0MBkKty0FaSeKuIkClCrnG62MvWqDX3kze6
6JoSohsyGTz+ZKX0kKjNG7PQdGWjanC6Kh4htgO31rHoOMa1lAXx/8dZPM8gDNFjUu4HNmhcwwaj
25zQEJD5qkdWyya9/c87+fKTlQZyQSK9PcJO0X6GNgw6SIj+IrXIOYWNftKjsPlMXc0IRVbm34LV
zy0IJmF8YPGG9HJZdZ4g3ria6SOF9sm8M/OU0draSD7f0yFWTjFX6dsrnZE0FnEETZm7rX3D74c1
qNewBsHqowf9sYAWRU9SB6C2XzocdR0uuzmBR8sW9s+T8shubCfDhabzl6t5vieg0sQ6KDHHv43n
nOzmMhXyr3/UGpFYQ5OiT/1bn8UF/pMBnKrHn2tEdYs8pu08WROKSBtAKQNfo9HSq0ygngFY04gk
aQQ93eA/nGFQsoXMUzQvrOGEtPiV8dLNkzSabgzniOXt5xM0uo1XJWXGQjczcQGH9rKzC8KmOCno
IJlV8jaU+d01o1ccBj9dJj0px2mgDpwf8Y6G37u9anS/KQJ/zgaR/hX+GBliiEVX0/xNENlqPhvM
aWd5I/viPoDpGBMJJ/hkJJfac5l+dq0fyrTPaouVhdQ0VldrfW54m2wMhlqkfQ3+j92VN1hrmRuo
UDYQQZiu12Hs1KEt3sL6bcH9FkkXo9lYR7hsaHSWpVmsKSI26OpFSrY0Ag2vFhs3fXsh/bmiLBt9
4CCvbrvvnKELImhWTqRNUXN6sIncke1otrQohm2Pac3WNw9TaLLoVEiD7IpvwnV1sAx4ToSTOD35
bh54ScZBJIulK6omECkMrgdfyLtizehUMK06eO72raI1Cxw6mCIjAm3BvrUUSEktATwAAgVeMxF4
2q5gUXJZ1Bk0yOxLde/XJtAHb+w+x7Y8NOmr5ZfwvGbxxOxsRwi8+Win7jZb1PPYTyEa2kKKS7pV
LrKa6EOfcZaXizyQ7rfb2R7AEmxE3ItvfTy5StKWp0en5quf7hd8gkvzQ7QJZAC8PnmqyNr+ZsRz
gpqvTx8Yl6J6UpXsTX6UHF1YLy9bz7J6sjWmZvtPUNS4Z8r+RpBXYOOoIYTspe7/zwTw+S0x6zXE
LGNorUL9cTftjsaVf8UZwzJZ34l93zh7Hkvi9nGOMasMj7kvbfP1W5GVPyn7WIzSNJq3GvJBTHlm
kTRDvrB2zDOlFHFochL1tyMwFOs8gV21Zcq+6teI2qUVxvvhyPl7cPh3w70GtoFaY/3kC2KEROEb
7huhHiCXLCJsaUAmE5lRhd954EWV5GyCG4wSMyePTe1era4msEzgW5WAQZq4GdElBKhWMnPxSSay
kMuuAqRXorOJpae2dHv9KvOU38iyMKrOQIAYlQcmSFXiE9JCHUucgb9XwJi+cygDRN3k9Iv71wdk
Rxa2C/OT7vNBt8VKI57+zhODFaaLObm/N05Pn5nsue0y5RPjSBG5MqkwLMQVNpbO4igXBpdU/zbF
nNy3UnWZCc6VC62CaVv+bomR+E1XWAWX8uagcskZN6RapljW6qR+pYIgjzIn9qsePs/7NWqWOOqn
Wumi6XLeHXjtHFHjs9O0bFt/GV3ESLtEk9hYzhQRYJ2u9z9DXXLE4WrCPGcncy+PbFJzadRDzsR4
OAaz+gnYohnA5IfQDxorPDD8EFOH1EaFpXehOQFLlBl2gA6mX3Ag7VBvTfJiQeu0MB2d9MQHJyG0
vE5hv1BuYK9S3Dkx9jharl9V0gzCqUiJLYX+hEJM5v7+o9vfdKepTFhZ9agegc9W+cv8HHv8Ftiv
vU2JJOeG/M8dwXaatbrKV/oq/kYdqrIUElZ7eQ2GR2/fzkN7Odpqseh4GPzMu2WuKBAMYFyN0o5L
fF6laZEU9h9Z1Q8DPLipEM8hv1qq70xKX1h5xm0O5a9afkepyVGLlZOvw5nh3/H7dMkB+XuaQPSl
p1606M0aBPY7/9lHuDxgwp5bDviYDqlCAuvG6+Xmp0M4wM6vWTRaKZgtz96TIghvf6vscBHJvig/
AypPb7TMgGXLVspJ3aj8UE1gdqkH9MsLu1YSLTnEW9UbgBONEOkOWvXKug2BMTGCelYslWJX9OPl
rHP1LkhRASDZlvSrpXWmXcMFt+nnkTLpKxKYWWLWUk2PckRK071zX31rgGlktGPqJSjQJliCWDC0
+fQW0Jprx8tROM5yboxREgpk0o113isNp1wPYK8lrJHD3b8wLeJBiZ3YCntDtO+Sp0AGMtaPrnF+
kyub8Bt+1xvJaEaaX5qeu+CAfwq16cVHaIR/vzBny4o2hzMjffe1R3LAyac1oXArQ/lMHPhgfqCH
y+O7TTQtWX4ZzRGHudT53p7DIybTKexRNTNxBMAoxX7qW5Wi1U3vfkwCRtS5WpqnoL0OzKmjpWf5
wEMBb77rgw2OSMRtJIvon/YdN99QSojcJvl4rQFSEWhZyMG++vUUJAPYaxPlCBCmBXYRrDxPEfOt
bzho99HeRrw2qQs7Hp2Ge95W5uMuek7YTMzzMTuIYgRwyKMHg9uXTfypcyRRxYGqFGv7U1H5psb1
dv/Bc7FlydVQezIjbMralJ9oXDfce8jrniphn6B4+MOFXJN7aYj+uWaMFGN6m6CWC0gHPsNoOerm
kiHvfWf3CHmxo6gaW9Jlk56ZutFvGxGB3sK09HaCQd6ZQiJEkHd7QsVa2QdbHW9ojwEhRfA7tMuO
JORDvs8EAXxsq2lzlClpJ2SojSDBNbuFkUPggmvehSE3J4ZRgO3Efq1e5otY29u7nGg7cs5fOFbe
WVp+PHw6iNVMrSB3Wid6K00iTeHYGWbxbbU25m7dHGIJieomZiPqkNb725E4q1ge0lASFpWdtIEU
gAmR007poVOfDUCPdcWSUwaGWhiVxKIW8BjNO+dPmXCoY3R9HfBRKcULFKlA9ixZGb9omqAD763R
jU+qafnIKYjgc3+Oeo1uPOBibJCblWj6tdOEvsaroh4nbVN3+gj25QvTR6o1va31RS/+Y/pYFZc5
izPWLAGx2Mz/xVnDChOtDQd0sFp4w9073W5WF4TJl5W5BG5XXNg9K1rqgs68xLlF5+EF0GHmhGiE
g28i8+zUeQ0xc/0BgtJphtf1ZB6QF801iHynnK1y/Krb6lyY2Y+CWfQC9BhQbiJsgNZWIkGwomaM
cBAG44GN3QR6n0Z6871LwHk3aGNDZ+/NU6tiil/JmqA02V2wFvyXnbaDGRskSp4cK9x4eplR1UB9
30ZpK9mG8NaQGGSVyQFHVhfi++yGOUhZnZiZ/827QKqcRlKeXC59MZwWL39qgWKXkAFsV3Tg+a2Z
KuH3TFlcn9ptOA5eJwFY4LnhejVKukkO90RSeg3VvqGQKiJsNtzZkZVt4t7+HUJTrGriyPm2H4Rk
OtMa6V1A9t8Hm6r6zj4VydIOlu9kpvCv5CUhJUDEHQ17fQazGmhA/xGKRJIbqtXBWXRkxZewIIsJ
wnFnoT1Ag4BO+aY5cuhrVP3V1a2fz+lKSO9r8PiEfCw20yQl0Uj0X9+cRQgsmmf2bq/pMspfOaTL
xF848VrXsHYuvQRczc2R4YNSagKPilM0NFtmskXiLhpzpu7ysZ/35c6VhC3L74hOZ+VJpFNiQRkj
qB1XuFi4YGT3fP3HJGZu9Gffi0XouSvsSdp0IPV/Px6c3NS8tRyprCyC1hE9WjrGlHfrUzgdYoU7
kgNsMRIn1yFA0oYC/BR1gr/n9oc1Vk25778QdNUYvxQyYXLBok2Hoy5F6PEaKacdk7dqO8OcngKd
t3NpxxOZ2eiwK4ObJIrca8sBzInbB6ZRgYOpcq+oc8IqIH4O+qru0TdoIgNRlg9eWwle/wLa38cG
OjnI/4lzAiHxKHZZsZz5Tdgu2r8kMh9beHcQKUAI0JmKs9ftpPYk/iM+EzKmWo1mzaEYMikiXIb9
KcflHj6ujAEnNmFwdGvl/iiNvTE3SIFdJMj8J/vKWkSkuQBGhaTbjhewuhbUvbBbrw7GSWaxSRT/
lOws0e6Ey7d9KbyJL7DoBhLFTM4SVNfpc1HO2CJldHdmdBSkeAawwZHWlLg4VZpF5BGDpmHopuhL
RE6h7B7Oevf2G/E44a3YmWrIMth3/VqrW8fW/HvyBF6huQ7BpXq5+zUKMLEPJq6pxUJPlFnT36T4
gFw7CVOpJ9aCbRT/cdE4zUlB6I76UHO50Kzns37C6s+pig75Adk+dQ/Q4lc/bF68iMbSJv7+dkRM
IBHm8+qWtyZSh+ivt96Ypy1iFMwDsTzDgrdiQ6GRyG147tjYcHBWmGii4Cx2ENnl+x3PF7pUhdc4
KSzwaT94kx43Vg2EVyg4enmDsU3RejU6gVeNK2ljtThJjZHDFqQiPAS6WdGNlY1f/aZ2z87Elh7J
LUoEvKnWgk9oPqUcCFzYZDAm9qygWJbVuXixKrS/jN6Ud6StFRzu2LlF9VBifuYk2dHAI4k0l6rK
k43/Krg/y9Z8XU5m/ujoX26bdcT4NzBcsOOdMxpPpiYqEPFLA5FhG6Y8sgEULUdIC0Ci7LdSx8Xv
qnqMD/g8/Y/mxW9BQjbjsmirQXJ7FT/uRxlDHqtSWQJ2q9sZeUSfp607iD++6pfRN6QmMp6OiuMO
y8ZASFAUyYtZ+7zuyTiTlvIwHq7+bTDG7NY1+i20U8HcNoXNpWRhWdxYL98BXJyvfGBQ7JUx4i+V
oq8Y8oM4f28lJqILk4kOtL/N1e8KwwRvOwxghIoQ4tYFl2x14nZRDwpQhziKiAn09qF1fkZZL3MQ
x3QYF+npFIBHa39GUrisvpsBhlBfNYFsmSV7GLwHR7GDk+d/M1ZXsB6aKc6NkX2bLpYyb8JhgTAD
59CZEE82VSZxNm0m1ia5QAFFAoe1NJD1ryblq1G+YWx0kvgoAqvfRKj1T1lSW0xWW53r8twmd3xi
6hk3ss9jrrgQgnfpmFi7FBJRxsb8GmHpSUvSyq2PqwBBqbWAu33EtRPtZ1IWrfMcBVQILH6p1hYy
hooRCWIpDN8HNpdX884xEjY0HDcO7sDJrTLRkdtQWmNvD6B/t507OMSyuQzNxBcXkFmeZGiwneV3
4g1dORD3RjXuzuNtWNgow3qCTecI6l7eUJzxPzFjL7WS8/IaOCP96QllaGElWvl4ABpgpmX7+FXb
lXlDS2B++/WfcgTimJDC6OmPTmJgmY+1vN48XCQPs8+PW9dsV8cWAYpXoOAGlOikwh5v3x7HR0o4
4Ag1dNRJwNgmmMIFrBi67yZMpqdqQBxg69OruLw/kWDTp+pSZod2CEzeMc8PtEtvTw50nbEdGz+G
HSJvGmMbS1vNRH87FZ60zdAbvewc1WpbBV7BBWY6Hgwj2GJAmjqPYMR5pAwukZ5zzFb8PSZABu85
WWEs+ldnTwsttKozfzwEpIKXqDBRVRecFILIs6+qWrvar/9AqF8nks1kBETbOdNSghOT4bCifidz
tS0EVULAjyVw/bTFYbDtbIwuZzdkRWj7D+YxpQqNz5o5H2LIyotnUThj8hs/UyvsNHW3YL3hEMYB
rN7k/DZu3WOckvJwG30TchNwgOcOhJvo8O2Y+ZmmEoRQi9IDo8Rdog+lhky4FgiWLnS10j5eQUbf
MhlJgL9LaMta5dlyxDqtpF9+8OASod0X0J/Pq4VOjKKBmcYXlEyQ924U0qGHlgjFbpH4ReFSKchD
nfSnZbNqKAsXIliifIf4Yu/CjqSSfKTo3u9dlk8sYwX1jz3FhLcRnvcTF9WpBKYeT9zSqdH9B/OR
HyAT2Cvv83Kwt8YJjbpE27nwazNrB0hKA1HXusiHdsL6Xo3nWcO/WxpdpRRTnx7ZU/3KIcuIRTyO
XNPF9cIL2nZmK8/aJ6CwLVBO16mKlboMEBYE+yeVHjY+xNzMYYyAd6OecSVWSgRUwqsGDR19cdXs
tHF42SNxKL6Blzx7bfJ20i9GFPpXWhEyCgf8msKbDAuDSSXBQW8bLhfgdkHu8CJ/VFG6s8pQWclS
5RagLQcMFxn9qxAdQNWDOvn5q44NqG7jYWueKSpG8CliK4x+1ZtOymoI0rnMowAhIXfDueeW7Sal
Z5hFzKNxX+AQZ/GM6B7+tG4o977DdfH0iyOBoWyWXLre1IQzEVkgJLWDCPjt1oJRHL+57Jt5sYtj
cmC/WcO0F86zNFdCIH/Lgwjfy8qB9D1eMP0FCDYFM3hxPg5eiANP+OgPjv00R2TjzpYBOHAYDG/z
5nBOfRFe8Ydc6P6HGFSg8rW6QgR6SPBMLJRxWvLj8weVMKNYa3y85YI6w/fF/CGtfF1l6KLoecvD
2FeovCnD3xCfHC0g0QYhN/MnsqO+JZoeZDbOVpDSzAXwMDmr+uKho2yz4/OJIcnAt5mRFP610kBp
xMQmDAWdzsrSPjOowddPr7FTmS+tGXK3fE7MAi9ZWJadeoZovCrJmoNIz+WXrqPJLy5A9XDArLLB
omYtZ7ATu3RV6aWJmXw2twy0qjcrw2lTOgHR8e79H43KWaAfEgGbqdp75HX2fjCYmOyQONp+5hgw
0UmHdsZecSDqVgIzIWa6GYLaM7uEvzXpmjXk7VU6t5ynYm00WYIN5HO6AYnifrjC9aZCcTgCQ/4g
B0YxrSEGRuI5fnUH7p+Cn3ZxoFy1zKtcNZhyVHif3+TDyrcbwqo2n4zgpKfvzM0nnFgk/e3vkbRk
eBV6h8FPwsqFreuDt7qZpVoRjkTQEQl6q8LZpGcbF8D0+j5ceKAJiRaZAmA3jczGFts8c4FXY2uO
3VCHbRzDIcARPN91mOfQykftq9nWwLthPHjBnAtqlUlirGlXgNYCz1oMb6p5o0IXtAVvVyD78rHQ
ApsCnKp7jwUpOzbiEEs5b29ceqxAYxPBxniiujwNt70r0+xl+iLTLgj2CJZQG4zDpOxtMIhOxLeH
ka7yNNbnvw/Cqv9qSTPftsa+6W7YWSm6Cb5A2ZILN3BVPI2LMvOJj6yxQO8fkUJLl4QRKwWhDRGG
uEDjd8C3OOzxiOQNdwu35PkKnBk5bAz40J9eQkEaKUvVc+DLwC2o6sTkOnnMjTMyGGELWh9eyERa
x0Uhunwl+CF2T1TQue2xfNulU+khjx0zLjZffCh4orIHEaMmYHtMCjNH6InSRd+cEbNPNKFmmqvu
pu5+EamcsrBqdVtojdgq/vFBcY1tJvwClNuGsUlhJXp9TFMQfyQ3g+uzuRueOuNguaA7EP8F9dVp
YrMvTs5D3ycnjiAxBaMoCwE7vRPGoQ5ERJWz3JUGpt7wBHMjiMZkvcMYMSrL3eTN7nIhRE/sMs/1
y91FVizn3dFNpFeeWJiAR3rqIYdD0eJQaGa8DvAUKGIZ+XnNissM34q1stU9JNHxAp3Qv5B1+65R
OlFWBQMA7HqSkKGZLXPnu7KGnN1hEj0Osw73bjsv8MlHZc/z0G0FVXUOmUPH16BoZKkZSVZRNGnp
9aqiEekChA9YXY1p6MjL3mXFrXDuHDZLC324R6gJymL/HyV2X2S4egYrO4NdfUwFpRpTFqoEVhmc
E32F21F1CtMtlcALdXkyuXVuBWbzhqH44T2Eg+XYsjTZSRXAqQr8TvXS715KlHUaPVvTDHKR12Mv
oPGQ9jgqrzIycN3rHvjE+BNO1MbH/VluaqQ5lTo1DJ35jz0L+QU3KW+PGSMYQSRUGOBwhrDG28zl
eQG6zll1RfyrfRYfzlEE9o+q6tjheFv4WpyRHWPPCwuaXUeQmYrcEHOFqqEozFYeaxutPAngjy2e
hemPFfwOlWh+pEYvGrhSV5TApFa9ZlYo73FQoVKfYcE+Jn/+eVC6RHb+wRJ/N01aUKC+ye6J/0Xo
pfv64KlpvF7ghzzxjQtQ9IjNl1Dr5T5+ubQHdVv4jglt7iDAUYcMIiMvKXy06BBK59f+0LKLm1eq
CRdpTowSAptGOAZqb9u7EHFwRB5eNSrq+Jz+qD5XjUgu2wUQoQFDlqNoy8SpqqoLAMfIG/wzKr7n
GgbYdcWABK61Putsfz/Q0jz1ZKD9k4mXQep3vOK3znNiF2BvJKGohzj7qto1KIryUBnoalsjT0c+
45ciyG5TMRgDHAGPP1uglpgkfkHuoX9Y/XNSHhzZ5KZ/i1z+0A2ViHt2ymf3UcL88/q9a82Kzz7y
d590DlriPvJkKlinQkgNSqGuYVSOjilHRPWjaXvqidslpG0TSXjfWYeyTb3QToN64v9PQkWw87N1
B7RaplD4OuygJdkXhExSXzIlV7hF3AyyrW6PbWG0lt3YZXwDty52y+jy62RNJXFToTnjldCzfadD
vA8og6yJiPkwjgp+PSslVQYwQG1sZjroHJ7iOASrZ1Br4aCs67gAp3FOkjIATyA4GEh7DNr31f4d
i7DH//H9W81n/dNf7mQXDdVLVCU/u2H1QmvnodTMP9mI2wzqRCvew8WSHvaQjdusSc7tmxKyhmkB
G8ALul21onmkmv3MAiB4zDdFh0YcJPKj9qL+J2MQ+08/x78ntOmUnbJbgcuARZfjMIaTuMz5Q5Vp
F1waELHVaEMxFsllw/TBlzTJTyxGstKXLRArYjDL5NFhO8lm5B99IdrpoeG9sEP3pV4l/acBtqUc
p84MV8Xw8alVSyM0IMqAOL6c2gFcMppYgLMAWMB7cI1HxOZUCqBj/o+ZNyAsJsvHiH/mAZdqGWSL
VI+JG7u331B4NFSmEogzgt3E9i5j3ITtkW32UEH1sEIHx/vDPpNmSXNDyowT9cK4btkU30rAoiJ2
7uv5tm+6qjgcak4X6gEhTwrhV3jlCq/oOz5zjP4Zsz6mGQKjyP/zmmcdkep5T0VRS5JHfag+Ydij
Vte7FA2A5zOeQ3ORLPTCqBm3Fmfd7Evt+4BYRb4DoUUJmek6vzo4YqD/PJlVmB2P+NbDMzfKkbVp
/x2ihqzK+vJY7Y0jqtKkaChaBhmV797RfrojWA0/Gx6CNIdkVkWc0LCXW9Rk2PCc7ijdhYF2iFwp
qvP1J7AVWF8+1/Ir4Ksv6B4idvKKDC2Z1EkSi8lCNrfrNe67J32jVnBYUqwEdooYR13tY1sMeyEo
Iq03o08JxR2mcfv5tkZNF3xR8Ab4Uy4PTINjsYE9YcieLb1hctHi2hyAKNAJYdcl+tKEBMcLsdMJ
fzU87AY6OOGRp7st/79szjg6clvInYHMZfTw6hdeCb0zxkgs3KBN6qwNBMhL83ZEe9idX7mRT/BA
VSPPioYzxoU1Vatza8nlo/3bqP9tRI2mt97wOUtiwKi7MuVWQZfVAdBdHQQ4XNpy7zFV6QCphtGU
Fr9K+ekSFQmC7zX+1VFPvaS6GQHN8bV2QjZi4ubQC4mJmkgTLTT+iN+n08IxnnEJVsYq/H+t8Sd7
VBjo4cBl5pvnQImtmcz8OjWQB6whbai/pzO4bQaFf5WGTCV237cplLdo5H88Al+l4X1muzzQwQXP
Scghrrd8mLCoXQjXqeFhkVNTIQ+tmBvRr+wStu1naHal6g+5+/uX/s5ZwgHZ8LvXRzBs9zbFXkl5
8yx0P7SeAdc/fZlyLJSKRE+kOJaRVpSjSFUbxipdhuQ6iktu/Jqdy5mD5yyvg/C/nrMWkeMyuQ7f
5lIozrTLHQOH4/tRX7hlatjT8613+V+oFjd1ObRc9+55nWG9p3OoHN2I1rXRmGsElqC1iJlYq463
Hwdj1IZjAzBkKXTVvWLobf6juEJ2vipWwK1KNXJNjnhVbj8t4xg9m8zLPSExmLsTMlgyQhsTYoXx
BIzYaP/7+QJVtz/Q+xYDH6ZEaI4nqi7oU25oPj3MtPc1RweCE0IqsT4BLIfTolnDUoOUSgGWm/X/
LMWMqv9voWYjd9OuwUQx22UuAVEJqwUKlc4h53wfyXY6MhVoZEZ/ZLNAXkvA6ERwuQSvfxoBbOSz
5KIgVVO/55MEeLTWaMWNva5dXYLvYpfmJF33UUc+i+p5U5LjCjWB3c7Ubzwa9FFjCoyo//aiFAsE
mjUH11vzq1Y34EbXblYRJcJcaOFbqLj9hkeO8YyIm5nFEwfnIbJErcfQIRYBN7l5a58JPCN6gq2Y
W2IGV1khpcxH6xtlOQ31XnUm86KW3KEPu0SDMaE4QL2VxFG8ALHw3VZWvUfnudp63Yznol+C7fRn
p2pHu4mpAQ8dBu5BDUdqHlTqxohP1gm0WcbyQV3kRN+9SBEvOgadiijEUb+bd3fI5sW7Ieat2aKl
WDZ+7bRA0vUAA1efJ9LR15SAiqFW1uIGW1jZhqFf6E+i2FMog/kndmpBh8LZDJKxwn9XfQVgd/d+
dvFKsSBuU97JDvohuhAwY3ZfuAsgkMntGCdfr9wmtvA5Npx4AD/zOKd4ww1MeXaDeAOH8CmzWkFr
WgYskOFA9yKy7TDVS0/QYQw2EzWnV+0WKR8E2D/zrWGORP1l/R8mdLokzupJj3FtW/1l1McrqHB8
HWdUUr6a1GCoSZoMUijhZ+zQfgOXU1PLd3NpxQ0TX7AjMiIc47bZ4kKYnvGNHt8XSKIpknlVasQ/
wOz3kJwRMTHye4Ih/hGwTDVOKK2fUsH+dSb+2hoJ1vAa9erPcBtSZtuQ7SFflRaTiAkpTC7lKJns
DggR7kQVjF2CD+x1SWgp3TFEGQ1NVeRfHcJDClSxW3ZmMWVqwoIIAAdyJfiivhZwu9OLQEn+RMX7
BFKvYQUNb05z4PPeG1e/7pg0J4wSd/6NK20p/8rAd4A9qTBbRIGaXjbN8tjCdjmdRfjpjvj3XegO
BDId4Hfv4NIW7VqC4afnTom2Igze70ZaF+Du5mZC16xGoAU+8AFMHl6Ga5Ni5TbzILcP94qvObG+
fuHwwLguODoRnCHzZRaDuCES+vQxzgVA4lZn0dgehXEeJBJ424kiImnOJA7uqu3rIuMqir2MjI8D
IuvGlVOdKov8O42hit5+v0JllzK0RMRGy3ech8IKd4LPxElnNvEc+dBq34WDWorhOnGzVzk5bETr
6nEjuc/mlt1b9pCVQ4HAfeVBxAMTV3N3s06FFHlTnDDFBbw/c2A0YvI21Txzo/7fRVEO2GMMk8M0
7P8ElxHA33G5eyE/lyRfZzvqRnhGbOk4w5QDBLFs49c/FZkXAtchF+wPPWgljsN5L0EFmOVgH9gx
LQa2BuWzse8UbwtkvAOS6f4oEBEGeJVi394q/GOfwyi2qXF80/EoyEW5V4snZStyVaa9fA3w04bn
ObZsCd1AX1/Ncz/TaHBz8AHsr3V6ebQh1RlFMOFs2ts8edKQ8KNzasAkaoiLjPID55YFL0JlX7jQ
FAd/PtAbhslRX0CHbVfQgAWQqfL61YP9VTWgQFlrWF0yjae7gr0WxDDb4GY5Z2raxNDrdBI7t/+/
G7UufqCCukyx4uRxzpv2G9UaDBfsI/DgLjsD4bbit1tXi+7qZLFhBLkNWR5SJLIDJn1iUVrZpCaX
Y8U0cFBXhJO6ch7UGS584nNuZFrYz5OVJkL8jkezP1N68tgC2d3B/C2F50QJfJ4vzkJZN09WGYtx
j3kwC4jPDXmyIyLUjfvZccm1RrATQUw442JHXIPz01ywG0+SAFS+CAiGpyK78InJ4PMtsNk6F9y6
7ZzjDBVEeRuQxAi8X1lylzCZ82QcjcsoB/HU3NV0mvwndrWtV1wu0rOQGISfUS49F8kRnCrrfseF
wnxhdeC07M4UsNKbU+CpwtZyUUpH3mUWyaqnEdMvXkqFKoKLACS+elmtzzbQAu1OK7L3lUomaxwq
fIV5QlyfRYOZ4cyrwpys7QWo1as/O10XaxC+cf5kw3Uei9lSQPpRVQbcOlvKlhHH+HfbwjIMGlBj
mkedp0RMzr8fNMyx468+NSKcqRYifAtSAIY4BBUdApdRonUuCai3y4/C+PhQo0NDfVApjwB7T4nP
ukraiHlfwCjctv1HZFkud7jEH3Y0ZxaTmk9d+3dDZMU7S8puKOVhqKH05gHkD7NUCn5PWokYXZaV
8VDsEbvESdkp8Zi8nvjoHlWOW5bym5NleQiFhQAIAvZQK5WBx8vFttfibOqq0E1q09wfAku7gJ7R
saBQOkm3rTm6s8weuC+K6k/Rf2qzGgzAMF62jL3n+4nnJ54QqAP+jj4Ak7kGrPZVW2gyJThs8A3r
vYYe5MwqguAL2VzZoT02vdy76M3LVcbxuKDWeUwxTF9GYPyhkH5KXGSISXAfleQDBvHRo/MGLmNb
IH/M+69xQlrwP1WIxzMLn07k67JylDgORNawp5iiXeR+7Hv0Vmo29yUwwmO2yV8oqkz7aBV0wd30
SdEw5NDPYMhksoPUOQbn2pTdD7SWYtBZTuyXL0QAGQdwlfAfnJZKg8IEVR3buFXE88sl/053gpOs
XledxtSwH/OFSwl9SmhLZwxSM2PBYVlFXUfqVz3dQHoq+bliHmPvS+L4Lkvy03KFQUCgVpHpGt++
QE/HoeNdBWRTPCSKbLGqZqtZC+Yr61kJfweNL/yWx8uC0i2tr6ja0inypBkVpOMcXo31zxKHvz+2
e8RgeWRAk3ph+ADPMyFi76YOKvES3PJuhBfWJahgB7StcnuZQhDhWFs9iRADfl9Blt/EcjHjxLdu
f1R/+bxJsZ1TFdm/MNWBTArJPr0cf454ax6WyG2sF3oqEE7rv+3K/lsqk869hQSQwrvC+FpjwopR
1D6QyRPA1RRXEP0aEIhuqgN/JGnQ1txDQA2ylLGrcXxFcV8k3sqY48/iXQCeKaTJfKI6xcaW1UbT
mwzY/CpMMeKA+b7ROBZNTlZcxBlJ0+EbtA7hst5Y2oIEZb6ION8/1C877squ5Tf0essfwWPsXDw1
2nbdgRjtcQZOKvlOI9TfUiwijOnqMuT6Swp6GOuv5UUi2n4GwuGS53yHhkGpLA8EqE0yz52hTOUP
tNKw5Z6xHEYb/e8EGm8aGi+M8wRPrJ3HVGDGtjP2yZBpEYZ1sDusuRYiMj4CaCvq3fZvzdnvTD9C
Tapc7gSQfJuzbFBnN2exjQZ8TbCdN7kUrCwOntQuwQOu+Nj9qjMDt/4m92W4YEgq1Z9YrITFF1Fa
fXic5N7cSvBqDkrhyoB2MM74HBYTt0nvAJ+84Y0MJJvvtJCHGz6olcEEb1NLn5h+kTLytC9FZM5V
TNXFUR8XQLJqfyNAbhQ9456PSd475S/mTTpWch8Uuxi6BnS6CJ+gbqZTzWRcxw5Xe1rB9DMPD89U
IRaZp+pBylyiFc+R2UDXNF48Q+WpOP+JLyjlMY2Vznfm7nkFDGocj+iRCoOD++zZBH+W5Hc+VtEK
05ewhlxnSHcksUjmfDZkZMubEs24s2XCBEYuSxaPD2lXm7uuH9kiHCVO1EXzxOBwS+LN2045o11g
UTyVFCaiyofyUVlF3GkWNR61NVvqhXNPsEAk1U9CgiGn6l71q0t6/ObYa//phNn22U19GzbZ3MXv
mT7qKVN6CvknOWFH5quYB7OP0cQEJqgVZhuqyN6P0RNKSKL5a75spnVI9Lqdg1/E460yK4UUfDSU
8fRcHtyiElMnufEuPq5oml34GHfPxAsTdbc9lei+y2efbVg9UGZZbCeY3rgxXypfwMLrtdrAkMUb
hspALZbU4aGtcwYWE/6Mb7hUNt6OALw3tVHbZwIqBao4ws66SBxSSqp1n495H76zYa3bKJ17gH4B
8j8pHBKxTjVZ+0db3mSny916j4hxGDpS+KJ11z+xcth/QBn//Da/XJrgTBoc+7QcOFoBwjZ7HE+S
bM73o8qU3QotKwRPWiRJUnAgCpeRRayVOrTYywtkqVeglPpXZngsio39MncNg9hBiBWeF/iY3Q8U
jk2YJSvZnV1JlWU7H6Ao0PhOU1LUg9mSenddoPybYidS9/St8f0715nxvoXxPgTIr4x44R64rUdx
Kje83ohRmdUAEAEBiXWqv5TQnLhdUrGwGbYNEQc1ezWn7uikS9y0vFm+El0qavHI49CUwsZ/Ph07
WuIEPQ7GdPcGtgJg7YYDiovmHpv2GaMHJacaCYU/FuwYysOY5VDKKevts1Oq5Bjsm5BTjfSCOXJL
HYV3NDjZUwjwLrmtKAuekPM0+6QRd5UQCf/kdQ6XvF509mNMIYSrXrlH0bUkhQXUBUxKO0mFISl3
WxJzs1KA7stZAe6IXFw8+PjSzGJ0U000PR9IjnbPnotHMlgapWERpr2+CUOzhu/yL3y0vBlzo7NV
1tQSx7YdFO/ZfxUa3C6gAQq9CFGYaTZ8EDe75o2NYg/R1/q2Y1imAWYIubiTqIwqsF9RFNLL2cpK
RGf5Gmku8vmRYMosfmq1iH40C4G5+40Qm0oMgB9usbl4xqV+5Nl5r1r5s/owlJGQZLUMhEgPPbeV
zPR6BLIUmNlCDBxf2z5HZXV5xzgeFjlO0c/KHwNFRl9tuNEVXtn3/4OTD4ZCYGX4gjhw9eCGqleD
xHw8PPdN4qctp8YK2dMFQ2vv1ACMrhaeWMWX09TFd/Rgu4IWIYSxEpp6GFxQyZA0xFE5I4cYY3/S
BlhBsecOaGeXu6ZIV3AszVbwtLf1bwY40GDHKjeCKleiylG1+OtUy+Ze1+Kz3ewVSn27jX+slQRX
vZJpgTHc2wcQNrdSP+pgD/1f9g2G4clNOA7iQJ64Se0MnL1bXNXye1+oolicqP6tY8VSeamF7DNL
oJtOCXRsQWPdkSSKSJ1ZTLdJe/xbZ/W6UDdtQta0etfdhWiHplFuhfgglIV6L9Sw/KEDFArmj7cw
x7eastiQO00i97SJzOJycxlA1tVSXfpB+OI1qZGVn6cYO6oVGrH6EjTjmiK2om9NAOWg1CX6uy0f
vdLMOjftRsOjKu0FFQTKltWkZuGrqMPeuAWdjVv7VgkXF7XnJRoUMRxM2IrNPiyTok/LRzlBQih6
sRDJ/Pi40hCStkg8KN8fAe/w+E6yX9EBNm93b+4zrrMCe2esxYcfBAIjmnF6Gix8f0ndBJD3AgMW
g67Q38chMgAJ8YAC96tMdVd4ASq/zb2mBeLMyvhhZggk6V2/UOoIXVrzyMMSSYewCcTQL5AQNJbV
1BRpDLcIe6EtbwTGs/1TUFovTfxvN2rqEtU4ip1pZaxxLsxhK0a8L/ewF5Z/TVMK8zI42SwpWwR+
S+bfS2PQqYsPzdErUQ/Heva2F0FVRIJa3s13rs1xNN50Gp6p8HjcWNZu1WCDd08vg0kGiNHc+NtO
o71r+e8tgSk+Y+X2kpULnhqEEa7ekATev2nndUg4e5j09tmSSOWyqEBwp+Aw/ez/paTBO8PQ7e4B
+RglDppB7ig86vGv6RHNpV9RPrHbJyQSTRrlBdP1f97IXSdPjngHrYRaBqlCw6STfxqXKpktwo0f
HM1I1XDUrnh6BgNKNgE2CgIHVmDgWHLI36zju+RTOw0VJXivkVJzqqKY1QRTVXVIWxP9ocK6gG+K
ESgWs3t+L/Qh3ClEZKsC4lMrb92aYmiZZZuLwGzF3HH2M51G6l8Xlp+6dNOxkDDfejCmH+uWnjTp
vGYYY67DEqbi/CijHqX+scdSbZMt9830mLE0fSRMw9MT6Oovp3PeeEKtrcx3IlC/VbuJ2HdR14YO
mQqOIjA8GiuG4IW19IsM70EZ5LH8pHNvuk0vBAK+IJWE2qrWqX/f//aCBzAc4NzqXTYNjQCOjzVL
3B+CuSrmmO21TRIX4QJE2dhCvsr+DuRkQx1eueZu1+PTHhQFoQlQzGB6Z7zQ2J8M8LGuAyWDhvVs
FMzrb8mqdbhLh/9KMXVF1kJOLHohXX7QbY5jL6WbbLYwSiw7USle5zu+S5i2X7BPrB9JCF5hJxwu
5tClks/qfyiHDTp5in461UxqjZWUJR22GO5WM3QL3cUWwa1+1HcpnhRXOVFt6XNKn6edfdMvf6c3
HwtYCr6AOWWFaiTy8miXXt3TOqrBYouI2FetA4gjrXIYzrc2BJ/ElVk616vVxpAxeimzaiUjBrS1
bdR96CeEmsjHi10x0HIAhjqYW0Uve9rV2TqurqXzy6FDEKHEQ4CY+8YinZc+BNoqlVFtQR7jW0/C
+2BIo3oBuF4tFP5Onys1PCqJGr1x/mKfKXHZDkCbvR6O4XBlwtK9OpigRPVAkxUI2N77NNe9bz5/
R9V0EA3/iLhcN9Q4Iz6T0XK3yCjhnw9RCHAFR2XKoX/FMa2d3MYxpMQYmh4Tr3s9PzCuDHAnhhcF
TD4dzUnRRk0KbJUdwV1iUdqcNFmtT8Xa1Ad6UOg4uXOF520shsS7TPilIpjKQPy8JHWJxib2gPBQ
FJbnMrD2w5frW+kf6pdU/yXjHvmbQPcFnEm+jEoXHEbjM8hTyqHjbAr+S2WP3qRJObod3n353Hcl
SuYsSWX1ROAdsnurRDaBUqwawunHmo1PaA/qXajDPpMVpe7ar+T6k5HNJeUc+X39PYIClot/i/GL
NxoULVmlmwrts6V+lwjwzJI6U/0IQecGQIfct46BEhyqamJIl355nVyBxDaCdqKjQLQmjlpLUETd
SiwylMlQXsu/92ssykPIl20XUfzXg2bINwsk2b22mrHWKpmTd2pxloB37xEz0abmENGdtjJqDQxm
40EWh2Nejd/TWY9vL6trlYpBc5G65bjEQm5ZahjFiqueWLKlv91BghAUum5VaFVBBs/2E4dGKorG
Rd8FXLAvaWPdNTmwbxpzVFbylRE8L/7Fmpz5XUCWY4ixcy5cWI2A/g4x8e/927K8tdr3WHNylee4
JZ92RFnN1R60Sqo7mRSOBcKQ3wlyOTt9ejNJiPw6+8+cNyfhIxtpNbfFip787rQgAXKgsg/kG0ZN
ZZSsb35FcSZsMkjT7wx4sj4iMETc5lnxNnD8Upyk7mGXSHsug0b5D8eibOyqL1l+saDYScMjnAUv
3Q66ZqKT0xcIWYjlKda/WfMFl7I2hiKbLYW4Ku0Uht9OLKaKBCdiFElBMR1ioTDpd72Smiyjn1l1
vB3fma8lictYN8r4BThspZ2xGNfqELrzva/+hOJwPXeF+jHUl4dDjuU2yBh3pZu5uby7ewc+i3b2
x6HI16BIz2EE8Px6EYSHEVpPh5pn4FfbUYaDVlfPx72nkgXbRNYgiu6Ey5lJ/QZq4zQyxlG7iMMK
IrsILAiGDEV+1s5ea+WC0kbL1fA7s8N/CNLzeQkHs4dr2Zy8QEt/7xpeMo2N9+aSYsAB/lRtd/7Q
nu6WYNWugzTwhAUHLkMBtF1/E9an9Vs28de3SNm9rkxJ/ayXgH+8IYeLQP3BwMXlshXruQknQAEK
C/4Hdh8xdrlhu7+LqlE+OU62TIW0DZVTUZcfCfU25lw+SxhSzmIe9Ie3RjMXcr0R1sS38pZ+h0CZ
K3XRkJQ8haxN9lVNhxO9gVYhTnceO+qKeiIu82UUhfq3ptI8xyWHljs5vNXM8ref7FgO4/7ryIaJ
NHbWP6XdRmV3WMu8GX72MCnUUwZhkIjs+Y3yHtNRqFijA9JMLLeC/vQh6gye9HIHpq7aAwFXY6FQ
RY3awdte1rY3EW+Xy3YTDP6vQQmDyq0XgHVlrkek1E2kxSt+Jyof/gt1Tk9u5UhZ+IiA6QKBYyWc
bw8xgmgkz3nKUFPILm6MDcLaqH/EmW83WdF709R2RlcTOD5BeVF3OoEJZJIkhPplfkdYJDQB5vB+
JKfwOFYDb006j/SJk/fs+GOxUnkxUrQP/aYnHeKjakWRCx3OWprRfqmSSnzM0yJyA4EtbcMeKIlk
ufFDE1U+DIhem6e1EZSCYiO3prBWxdi1zzcuj2DIoFAadz/NLHFHhGolrPe8AZ1TzQCEOjfjUP1s
Y23s9jZxYGbv6H+OYn+wChqYSFpF7EPlBxmPymauOu7PcXKvaPtpHcYLSHclFBzWYErp3OuK4grR
m/PpcyBeV05J9bIwfNPknvriwVl69KEKZjdWCxXNJubOr2aYvP0uCh2/fSCe84NGNMpeig22PCMp
AsXW/gxnRaIr7I4W9BqY0VtrRkVBLAHeXxCQ0SUZY6bxAXpD5FC5TuavBA1BB0ZvjL1ELeXFqiTC
DfsC/oBUEGMbMfinSuLuIcJmeipMN6EgARroyWBJWEDnVt54Y7XFksduirgeWn+IznexXR6sGB0Q
H1jMVoLMWe2jJet1LalyGS577mjgZz4pupcoQ6oZhXFRtjIrATfQ7UOucfNuJyBFi8wdi67OBEG3
MYgllQpicU54efut3pxkxzMqzpO6ame5Lltw5Pge3Rc5ZVhp8rDBfIe2gGSnRBKOZRGcqp+GWp+x
1rRrUNPHSNrt2CZR270P3RWQRMiQKAC8YpEst2qL9tfrKK4pQoX3pYfUJNt9IIn/G3iz5wEN6rvx
ZNV48ja//y2KEWmq/XBp7I0iVlp/D/JbwvIvxJy+oDrcYum8x2IP510qgmu9GL+P79vvLWrq6e1h
JWSkpdy/542vvJiOY8mjnemUByAArg1F9u8xuoC9gmy3Quc3o7MJAr4BJ6mjooTtIhY76/ZhCAZW
pFCnpEf3bhEALoRzU28IyfvuvCK4qJCOm4FROXsli4IlbKDuyhli0yWycCxIVfCs5RbxwAFro3lm
p29mzPIbrJInRf6BJS57aykpYZuWrqHQFcbtkVo3KO0kp0hvK6swvBsI68U8Xg7o/zCm4Y+yd4jA
6UGkZQu6ZfYLetrY3MnEPyBBmfHR5HLRemTO4S211p3mGy/iM9jvYYPhw3927MQRbLHT35abnBF9
+ahkeZ3UNga95ALMNwlEI7WVc699BqJczf4QhoXmdciT4QjKTvnWZ7ME4vCsh22mzzvSPeh9yVLZ
B3vrVGLXkRgnCCuLGZfwrYElA0Z9wPlPDYnz0BreVYYTm9bybJBLCWFXcmYjXFcMG+5pQd2t/u/3
qAp5eSUlhz1Csfx4r/yS6tJciwnFcfPKSFeR41EYCcvvBYB1uN6i4+5xVC3B7hDpWoHC/2UkWphI
qN8cnwX0+Tre6SaM4xf5cQD/ZFPjNg7IfeIqarbRzJou+gMrCA4PVnVCjCMBRc6iEDdrQujHfrcp
L0USQTgxKxqQbLV5zHGQ/BkMv7l1nhksUlZjncFC2m+MC8+b60k3h6JEBLG3OErHg1hpxwO6SawT
ysp3ZjD6c2WPai6ep9h/w00iRErwr5oKSLuPMijopkQWq6MuX7phhoSTaB5oZN7+/x83J93nFbMI
EEaVl6YGdmJ2bNU05ENMWY7Wdei28RMBBIffYIiR0nbZ7Jy1dxvu5gx49JpfMpMCfUjFUwJ71JYn
rmM5/1ecCnmUVa6Dizkq0IYF60ET86adytu7v3Npqw026IcGSX3EqKQV+bxe0OEZrEZX5gUULTbW
Ur3cWyfkek4zN/gyMx6UACCuKRHTGzCz1I5r5OXQQ/2VnyvF5MD1BN7JJiq6bfpDNflr5ig9U+or
qgHU384NYTcEKNRxTgD+/YRRk9hgrR0vIpOgs0Ebyz31AveM1rRKmOHatOPHVwNnjKNG9VaAeXC5
0sIP2NzlfhyZEUK6PhNBcfRmO7qiiloDW/5KrLOKi6wkP0lhyi4rise7DCy032+CpFLH8rH5JNnw
MmYRVCpEVjwgBc3LnCnz2PBSwFZNKyBO2iC+1VMujgu8gngwyb9grw46T0N749BB/b2FBIpQ1qWW
PVv45C3+Sg9ujJSlUs7xxxWnr0OSGxH9ylSv2BbCSBzM1miui0W0mEotG6RbTdPeSwwq9OGsYCF6
hjNIn06i+K2h5xjxQxP6q/KsKSHkDPk9P6emliqYiEPOaaL1x1O8t0RpO4nXcOCwUuzhRYjmxPIc
oeuaLLKNQhRmRYchb6edmff4wcnFS4Px6EWQY9bnurdzK3juHldXlMSdKGqTkACCU7BbImdSldG0
NNoj90Ixkr9XucT0MUlCG+dkI5RaVMcNX313hAuo7YbMOqtGMYg/jtFHIhaSw9BKZTA+Ry/0SQs1
oLmdqHNv78QQEi7JmgAhfeIFewXd9laxM0l37yMlGAGZRn9HHJ/umJTBEAcXxWUPDY0RE2/qpnKN
hrlqMNtC7fiWBW4cAwitbxrXTwjHqd6F6IrLzmQ1+CvtXKQubCdVG/W40SAS0e4yhPG/Yh/pIGI1
TtfEzt2f5/c46n3vw3WjmhZAmJVe7Gdwdlqx+2hYqfjraDfaxUzZ9Kiyr5hpdTt47tK1rWpM2+Od
5YW0jwVFy8S0/san8hSrrko368HcP5nVbgqx7/2ilYmmJ9fgzVkWR+DEjiEeD0KQ4IlhQP845EdG
E9W/IIuBLrrosCXtz3ON3UmDPTflkshI7iNhwlwRVJ28ku8bWCXZGOn+eK6MOTtk3p9hTq2CUfsk
sVTbUuj5ZfoKWv0/DjsNFXFogCchUGY/rvgQpeRf5FFLOXJehIbtYEQiA4NCTFjPi1EFFHWHZ5uD
sz9RzrYs8/0u1IO+dNBtT42PuWrtM/dE7AgwOPR+xQrmR/7o0CObv8aFPvdgeKdOH94Y3JSgDZ0A
NRZ7Vtxt5tU2vmBxe8sTBWj5tiQDJ+UN0DgkczJICQvlfGfoznqYSXrx57aJP8s3ne3qYrhp9Amp
sRH6AMM718G3R4AKoiVaw+HOHWZHzW0k9YM2mGCQcTQeEIjTrj+qihTbofoETQUlCWjFoSWUmRZO
ujSFEFXQnTIQOXvz6sHFlJaeZdBdQF4M4pZwQrlnUmnF1LmCYkpoWQrvFK9kdXJC49OqU6hvJLZV
i6Xy8MasvOO7w64SwwHM/1/GEDPFlaN7Y4yXIAkg1qiT4csTZEGUKhJyPgDlM6U82E6gU1yBE9jH
Ks4TX9TcVWWwzdHxZovdIGi2wn0IBTuGKCUrP75dRe8S5htR5YjbvM7UUVvsix5YuT6ROjmfQ2YE
XAYj5DXSqTy8MkvKdoFaMxssyflv2PurG7vYWPrhnfKE+md/jtiGOR51b9zUryaEtDPJQwd5PPPZ
3NBeHPPCDk9lIYfjf8+1ut26ISHA2RxXOIj3bUYZIQjbrkRwcwyMceTE7rQw+PN1Q4Zzf2MJT4rM
eTy7am//a8zfClz/9TC1JDkjWpJqRcEVt5ucW8yg32VLwTZ/rupcz6u6ljLUtd9suJ930cT58yVy
hmvSeSumQEAzfqvZ/ubtJQ7chGu5Amu+mhJdgNA8DWyIzjO6v+KQ7R9VDqCSYtyq6O4VYfhZ8S3B
leD7ju3pPWfGbOyB7u28XJZb7fT2rsaYd5M360CxEm5rqczCEizdfn0LDBEm7CA31I1y+lX74dRe
I3Hl3mEA4IYu0OYWCI+/YHYkNYe0YvCvnURz85SX7LOHAdfC4HARbRwxlB+q+qgtWsfkwLia3eKh
A0BWBvtrhK+K03i5rGbawkO1kQdA/EpKUOwU5oOiin/fCF1sg6nA0bPukHYHVnwFla9/t1wmfilI
v4CEOrc25QaVuYAuIHszknDXueDxQt6PZTaefLdpdUqIXURerwhcXPgW0KtOBQ5HUE1ifaIYwuaP
GR5aNx6WQOX1PVeUUCoOAQ69KQZrmHKSZ83wVkTkru0UyHPei76wnlkG3wpkNtlmy3bcsVax0ZR1
A/a9wr/STX3MvaAMAe7WT6eTn/ubESvl0usO/jet4cCULjvajkXrjfLKrda0inEGNiMlWqWOwkbe
VqjxPZXcJJ2+ubmh6vcvuMdK3AkJ8ZxoDxDhS5pF8stoolH5HEB6Ze2IqjHNgn5P6lllSKGv7V3q
5m1s5VRds5fgxBJWK/ex6EW/xc1V54rwpE4gBxco7A1hFpW7UdhaeTx7hyBUfae2JNCJLjE7BY1G
ntF6sCMvQ6RRhn/FWXh8Oke+ENBkO98vNrO8qmXDENzmbEgrHs/JJuiqaIcuHGWT+ARQ0I/5yUgR
YvOVigSBOTiOSxDeFibU3UiY+vt6C38DfHFvHSMK2a+2j/Qlct+V4i6kGzG548rPHkq8EK1vzaqo
Z7H5KjNmKruOmbxmaz9bwNN3yqCYZSqox0a7W7VmodxufoA+JrzjPqElyvpz1HNpeovX2/lAlS3X
Uyq5Xs+GiPRMNMWHtn7ThRWMha5QPaKF2AGPUz5tdeo5cfjASOM95ComWsO6PTG5Agod8bv2inV4
Z6s7R8avGf0zyh8ZWIODnXyRUbAmud9gpQiwSaWAS8F9t6gCbFi325KGBS958562FGX7Mvp0yxxo
RTCDdzC3AQ3dDYGvqlrT+A/+3nxX5ZRDUQCjKCcBQk8/749BM3hPqVIclftQLpKrhSQWjwQ+WQ/P
sYPYfmnpcEXo1aCfXBsVXiepwGn6R5GN4TTq3jg+RXgJQE3LmLvnRTwfqnJXraXNZ9EuvBosEO2k
vckWhQrVL9kXOgXA//ngeYZz8Ckmnb4C4AcmmQJm+MYKyjUowyhv5Qqp1hrsu6UIh38pkVL97xtX
RkSn/BdMUqsq+hqjlKtgv3gH8ixkmUJuFXIWDHk34SbQ3hO3IQmGSql2uItI5NQbDmyKpZyrxenu
obYGAV01fzWcVCkN/GBXT04CG2ITl11+bFERhaWEGmgFL+YOFNfOn5f0blmvFyn+s6jd88WoN+I2
l1za15X8oK27cE9e3l6V0uVdmbgx4YRFg//pRONnoJFJPE5N4kN7SG1pfqCL9KZG3c1EmV2c1n3b
ZykZHwCMTImsVPBOOOhLloq2Is8M44XoTXDKnxGvK43C8gzORRLMoRJWLihHG422IcMuf/A9Op59
H8dLMWKaaANI3Dkw3MxJ3UMthBvnZWTs7i5/bLNOnkDlOE+qtQwvroESzHdgWRaLgLqE1hN3o5xX
tQRW4gCa5h4AvZbMt3E1bCUm19hz4R0HpegR9BjgS3H+kOCbJS0o8N6DPFH70IKAsU2sRyfHTiET
Ei5bh8++goRlc8KEbNYHMtIlypfioBvpQdHcCTcrqLGTJeKA4UlFez52RHNxTxlpqgp1+i0tBkeT
W07mm87HRSiLljG1Bd6Dn8EL6qTcBjDDzq2y6C1NheJS86DrsTERUTet4PnV0k4KYMx4/LFQq3LT
nkmpwqXVdWme6fYSydYzZS0kD6twqGtLF7XG28Fr/WQ63dxruGGgHjnXBgOoAomL9MZGKrSeRrPT
c9ZuJe7JjEngsYmMTtz4Vh4w0XzmuCuHVyGsn8xhrB8F19IcH5xqSGYqGvTY2uFiLFHESwEWLUJt
mhLrV1CBzHnQQFXT8RcF4mnaAcRigQg2YSXOUSMTTQfJDSL1d6FLE2D/yWhxoKQG5asKNlIhILt6
Eg8PCwuPia6KpMJbFwaoaLJwt1K+PikqCLKgTAgLAhvAFZJbV/KcTyBVd/PQenOef7j6ybbn8z32
vLZzLx6Eo9jHrcTrEozEl/SY+gDdDptC+SivkCOZvVLrJoh7ZyWe79B+RRDYL77EWbqOM5GWSKSt
httmhccfCXHtJU5dEFqdJGoPGrerjdjRdf4fMjcm5//gBNHtcCKiaYhA338sLgAUgtPS8D9BTwb8
I1XUvTHnUhNsjNH2nNmv9/gF0LAUgQAdGtNgSNxp552W7ykmwzK6n3zWitrauFChHDMUPOJ+T5oH
nj2ysDYImUHAoaUj1cEoYAx8cFyonZn51OYDWtvN5cFlTb5Ksygyqgvyg/hmPOBbE8WsyP5bQJsL
6k4yi7H/61dWutEUtHuC77xm16eu+PwVU0daLGvttYKCKauYcpFUx7KyDQ3vtOA+AZTlImCCL5aR
IrMWFzTcjHPtgaavAQZ58ofOWh1z5DE4Fi0HkfzSDacFCHWUUa00tyt5geDUCa04WhpwCw2nfY8Y
A6k85nRKP289bsGmTAZadJMeWPaL2eAUZwIN2OgwXmQLmhMalM0j4+IyHuapcKIPQAT+FTsk62GW
ORCLE/cFMJbisdXpcIabkovCeqhmcuoTAYhdlluykCznZwJyU9eeglgkeVweYhLlODWsTtnyY4Ib
oT24WVYlxRm7Xs7zR0kY2uBB8uSgxOqhpM064sgJmmmppqkITCDufBUfnpn1+6ZvuH9Hf7HyOIs/
ra5jeHw7vzzHVqA2AYf6+qW9rtXoOo+tEYZjZF5cHOOvhchVpv/+cKYzDqkfp+jV23DJM80X+2aK
pyGQIcm35j0xJSPoJCLAGtrDFO7Ya4fGiGedez7uQQtsajBEPFTBCSCS8T1Rv0Aok3oxFKO+n2my
ywijZbqdxVl3C7C6rUAs008+5HpBgC7ivzu2bXPpCOXbGaQQKeeNIxzZayBEQC97O8gOHxkf0B33
a9H5DGvkhFUCeQ9HP6aNiSg3oKv4hcBVd/D6wCHoTh7SLzOiyN3BwqgqAbg1pz2W+hGTcnT0+Vsc
clbabW/Tp+gpgZSiFKatuu/bkuPhuITb63FEz+4BUEynWiEWgGNBXb8f/eac8o2MbJ2By5W3U/m/
aorKtR/4wiX2wEtubIeJCpKKTA90a+XmdQC0YfOs0voIBTdSlrATdJtiTmvaa6L2tsArRYC2rojw
rUYGuZcy7EMIoT0a9nR1eILTHNRb4VZ96yJNSQ+PIt3nFdTJVAePmu6peNORJo+rxjypLOaWVLy8
oXfr0cIuU3yr772jQpw4Ypzcf0eGyMmjN40rCJ/uAOCeG3cTT+giYd5yt0AJbGw6YNgGUE7t+9Kc
xJvFbF5Myg7e4uDpjxgEI4c34sNMqRTr2zMYUuPRs1Vq0miJkbSkK7T+VoAtBsKchjMDs8T5iIbO
m5Mnz7AWirVjDNFcsEzJSajgY26W6W5oIzM16rcvptDXV6uyR54YzMJnaeLB16bLEtgu58uj/4F4
Em/hvzJkhFebcGifvigJ/UMFN5sxCoGTBYpnPu5rryutUty4jTEMKgzvUZMmc5OBSSTVPRIfdwW1
UGScN4ngXAQJqVzWAprzGubroC732OADIKq7M+JPbts70QdoZR50auIB6+srmxbv13mLnWaT4KQh
zi4y3yjO+jo5RrCfR5+Ol1fYuk+yTGsLMtWyLJKAZju6SCoEFB4FSr20YKD2qKkIDSsu+xznGj9J
QHdYKpFwiMy5FwplPw4jnV5YSY3NB6D+xR3zkVfKS4K+rEEUe7PCh4Z7lWID5PdKzkIluSeSoybB
aMO6+ZE/oRyiEeRQQUayqKqwkl3+ZgfUQ2QS+uE/+ehzkD4YyQ1xvWdPfJo4fQ38OSfWgFuvFmF9
84qgxCqJvf68gnqjden1CDTAtmI3gOi0+6D1mFuseJ1SEmArVUuALCKayMpG990W2PcWeXqsa3Db
1OT5toUxOiWSXtEwfjulTQ1ViYoQVl1RupqIobKkoBvAT78lXVGwBHaemAh6rYUyJU1EFBO/akkT
wwVmp4asJkuv9LzZKFGLO62LHT2bUH/U88CHeDYB35zRc79EnKPIqD1NlFmT7QDyrEgU3so1GOSR
6ruhX4rG9KrN+ZhWxVbdycFSlv11/DEFatzk1DCvyEJwmP9R0H203hHe06yANpixRMPOHtN3vCeU
DvPLU+mF64gfo4iet+VY7Ox2YP1Dfu2nhVspG6lGrXcvwK6dyIAUoIEEnOZT5P6pYm92eG1qHbsN
dKRcrKYeLQedLfyY4d2pmky2cQoHoyDn6mjbKO63OT/e7ihVPD0nw1CezEsiIPoXpC+wlZWx8WDm
Dt3bt9ckZJoFy9k7yy3S0UzQWhGEUQDuRZ7bCrTAm4uHv6je95X2auiQL3WOJWmF0YASL9wxwXga
0uR8Hd4X6BkZduoKe0RN0Ldk3wG72Y6roWPioHBlTcqcKT/YVlQHxpkggIwUu0FOKk1qUpCLagRe
qRQk23O9LrTWPcL0N6Kd5LpJAOg0DVcMQP9MWctCWHq3ijfIYsrp9BjDdqt4V90ws9x/moIJ1w/h
fCRCu2b0RP+1Dyi9KVyb53MxL8qgod2La9MJAiVr30mB/oGsvH2Fu75m00Fvd3x0/MVEtVJppOqn
DddfcpMac20dJ/ZwIJVNQr4zAL8s+bnL1gm9A0CbIETdEA90C9D/r0ZZmGxRI27apRGS61AFNqq3
vtlzkl4JIgYqF3IxbeIDfzORh4XzlNLC1fgPWvF1vppuY96sqeg1beFcg02YPxx5Z4KFd8/JKRPb
IxiMs5qg7RWbvnOkGBQFw4IumRjPey9BvO1Q/wZELuh8VpEy+OxnuXysSCLJ8mLFyvVPAWkodh8Y
R8p4lWkExEYbUq2emKnQWHaWGSLNyN1JoWhf5Ag77xTzXAa7LcKAfa9DsRdrevWd1m6I1q4qKqv/
VvbIDijtVCgVGYsF2Gg8yAxK0vhE+k8swm51WOIOTShRzkrIDjZIh/TaUNKqSuC6ee7alBprmBTj
DC+tH6YvNKitfwTAtcMC4XTpgXNFLnSUG/Rn+5qEhtg2E9/CG6U8N9nw7AA6D4L2bKxAdcW9Fhp2
NiJMaCmR0yROig9Wkc5oCqvTv9pEsbAk1laH+DF1IJOkDMdNlZevRUTLRrbEU3csvALqFhPcadp/
SzXCOx0fe0G1Md1VLFRnC3md3evyexAGE6A0Lf29IZ6QMMfEpXAv/Mnb5al/su6WBu3e0+blXQQ/
OsrOhLHhUJU5iN2ICPGlsBmKeWqMQKjnUoBQLAKa36/FgnGQLUYDHvasY5yb4c/bKY+pdKGWwuzZ
eHWfyCfbR7NWUSfB2wCrEc/aQhjbgk5Qc008HBrIhlQclV2nq3T+9NWYWgaEUB7R56fE5e/A1NBL
FOnGsQfsljXAMz11jzSLzNCjqVzoqs7Z51u/L+AFkIOe1X5IpMgRUhqAFyWeLtiMnkdRPDhwjGBA
3BbFvWMKelB1fj378T0M68w+adf8dTQRg6Pql+VO7pUWCbTaTabm+7o7/pIIRss9nkVKYi3atLrl
JygRP7ikH3pIifnlmPRvsKmIndqzTEdfsqrqfMx1GtRTp0o4QU6epCL3lU1o8Z6wCXGZejVBe8ZA
NZWXjumwjZmEoGFVu/7+MCe8Z2lItTzV4BFsOsiTdeIn5IJ/fj6k1ilhZsk+nYGP4jMbRQrsIah8
L1dzC9FDUThUm/V5VtcGd6Pv1QKd16S8njBkaStAn+R8DYIzKpB321z797B0eNstH74jXlUMkcuX
2wo6iSIoJar3FK3U1y+6erBQVx1G8BA7z25nns4JFfwWWOHtQuUneLz2UbVcNuQhw1mNSbm93+hZ
u01o2pyWrIV8yNuJzCijZsR6YleeKIongsalmrMZO8jkEBXoG6cB3lb8GtSeJg8tI0yJHBYdeeM+
5Pext6/bSWsqUfIqfdnOw2Geoe8RyW5o7lQybjBdUAkAoZWAkBUlkPYX/zsAHbc5z3QptdeZklPg
9t49B7EoAQBzD7us50wIjw6TffXLmi8CjXDO/iCMaUM1y2Fjauknr6fW5MNpCAYwcVY61b0FQHsO
aoLL0ib3sq4Hmm+vyBfiY6xjla5aSPMpHH8JR/35+YJvpIcbYN6CYpc4eT7TCndo7MPYR+vdTx3d
wrKbxb2tmEIFJfMobEgAT3hL3kFzR7VieweGuvXHGDUsjs51oPFvwwPHNqGEsHD8P70g8nlGf06M
WqW5FuNlvUV5LS5ybOnBCJfTc9HzINnZamfHd+f5SHRSgB2U4jUYa//AHYjrpIM7HnkMV5/AWnYc
biwMH4QMi3MhGRobakumtaQkbzyty85MIUFLogxJ3MES9pQC9ogqwaPd1t+QKFyIrn0/aRM7nw/K
HOV3YIBxhE6ZSfACJaFWBmWjWaO3+bk9b+a8wv9vH/s+1NINxveTVpyARU/uwvtmqBlX0mlR8SpS
O+yO0GvPTvdYBif3gVlnQtmFYFCgoUFwBjlL4Wl8f74QjF4PaOuhfYZ5+VXk36ZzzyXM9GhGafjB
sh6wC+Y/EE1bjTb+O2vuLDc5HIUTHAOC6mA7ZW6s0SLeYr8YgXgDUfqQCKhSMk4+YLHNxKAMmkG+
cHORDiAJcncK/ZPUdS+MFDG0tQo9zdu36r/TiddhMDeIwZ7HfvMUs3jkDdAFSyMdXxNPKqnsGRoU
k4dcg01yFp1n6iFI/i3kJ93CBUG3fYDPHP1hfMCilHSBuEyPHd50LZ1vp68Ms1ppIFpoeV5qGKG5
2ItWc4hI0hzk01/BbqDIlqAelbQtlAq9i7i7gxMdlk/5Er1igKTgkVKZoroZiAM2Ke3n3E1V14HE
DbwfmWFSxeo8el5ylTYJAy8dABut7fRHnHixIRmuTpVzo8GaBipBWRTyXnyXMvMVDd2Oz7dYK4dR
l0xt3WMwF+6A9LNN2+OAhugx5vccGvub6wv451rWl9FpisLyAkt96TUO1NMUT+3sBZ2hKXFreWkO
f12YjP3EWlesj7APdDAL8v/c5/JCdQXQg6Tu808vMpdfUh3hbQvfSTuHvi+aujca19vTvt8iBtJf
SGemWfAg+DoZ+1/T9JQPt+2kNvSuWb8x2ng92LUpTfeg2VXJ+N+4qbQL55eHbClg9L0EBLfaAkEG
trd4pC6A6+eCgbqcRWBgZeVDZIFY75AcAana6+tTTI7p1ZD0FeG3ZWic2PApMR8sPOPwDYSQPkcb
nfBZ9Hp2aJeHBwldOwHmN/MMP889z4wuYy5BkXbPiSxauuM2y136G/ykiB72mLL8zvk6H2MEj1Et
TmSNNpKNfgvGegHuJoxc0bceaf+c+Ykotz88oZ6mOAwdKTu/UQ+MOCAnF9z9p83t5pMcJEZm1guC
LyFSEP6+M+X1416czzmEkMYSTOnkLsX+jKjwmkIgC4f8FL4k5BhIoITv/Sh6ThXwo3YJB8f/OAk0
8gUVp6qdMvwQILCs6cA+bHd5Vjec4dKdq5vBfJ5GJz3II1v1Jkxr9SsKkMqsO55EInudDNZQ886J
AOgQxm0UoWsL+whduTDJBrZMXk6zs8iEgrrr/VOPzn4cOdBKA9WFRx/ZMJxRqj4Smx5npT/Alr7U
3D3tEKPDdp5h/Y0T3N2ZfCb1mnvpAPvrUTZnSZDiLwpHVbzJ15YDTHbfxheKXATFDZ/zDyBCJ92L
4KX4XEDShJd7MZtBxfICz443FHWZzHQhMomWCpcFZYbHWqMlx7XLQbNP/QdqcacvhNKYXteP91Ba
tMquTVaWVozSKM1OHYJmanrbQKjEpT7/iNvWnO6bGr8KxRDm0/Y5Y89HfTDtNAfY3R3mbXp+gaFS
+8NDeOM5m5nBc9utcAxqjV3Z3LS/eTELtCI3xZEUzNfDzpgJBv/qnpaOqEyoIavHS5EezmIEtBDr
z41/0C9wxFJKmPtAs00AyAZgiRAfvGYw6E+pZCih0OxfTuQ/npPkiyx9wql95ki1aRJ9o64ycETr
pMrktENTlQmE7jkqKdVTQq1gXCb/OwKy5RslvzJwA1EyZb5iTLLF4JLqTwKjZ7lDMHZUEfeZjTnk
azOxl+4o+K1HXrnJBmYvz4MZJ/gfS7WtarhXamtSBu0cuUmMoKlomLWbZ3D7tau+epZwvFuKqR7K
T72YKlYxq+6vw+dVoc8sgS5PwNEbEuMBRNUesO3RcTt6QeJ4SRrsZcpvsRQQFr1pUOp9idzz2er1
RudeQwWPKhMZ9PMIPI2xMzilAhPY1UAPr8fHnCwKCA6Rcq8Zk8pcSDDQEEPLndwHjG/UPLHB97zg
cvBVqT+Adv0j1hHQyO+ahb5H4cf/+Zjz7ItkQoZzPUW9aqZvp8uNDkTJqhbuPqam4ECBOH0oYbmQ
ymEAFjKrZ0q06l1Dp8B09nqu27UupYg3UA2TgiP58wBnSm2ON1gVBRDN5KTxdXX2y2ICeVPMSj/B
uMecvgmwOIhoSpGrD62WbV7le4WGPzBMs9eKu8TFy63c9aufW9knfFqAupWqgZ7+Wx0Iw/wsmUjh
uHpYFd8Xx7GQpt+RaBS/QLifkHbB/xIwYYAhaYCavmd3ypJiETMNp7fbkyzns/an1tyKzrOPeN00
n2hOmT0kQkYlaQwiYUTj2UKOoLYrmkqL41X3HOnIUu9oNN00w2qR+wUh6IHpYaFcRt+6yrKQSBNA
thZnxH/p9U8MRd7FUJvOhGTOax4JpaF46zzNaQVn11UHLiur12tYq72M7gL0jajCTD8HJRuDIFvo
rTnHdi6oXTQj3I6XdFXsb/XM5OzJPO75KPAkmNjX0MciWfQ5nmWI3S0uFhrBQExyObDbKvIusONN
Hx7pAgKFfn62NCy1B9F8lelsKteLF0mLVvz76Fdq/rO7oAethPArcA3QLPhlxkMqkdaqWHEq2xTH
SC+mcGsKW+cH6AXMc4CLl6mZP2lI+al3H4nbwB+uVzv/2gVVe/NIOj1naJA/qOUZeIQTE7Q2tEmn
pw2oe9S0135vqXdcI6EMVmGo0EGvyBZcQyiKiQmyz2dgPXtdlhgj4dBR902IwdBM8zhkCaMh7oEE
7xAoPFog2CkfCU4AJuWo3U/5uHvtWMsTIvAzhXt7Y5p0Qcy8fyOQCDS2VJSIMT97odU6fObFXOj9
wJ3e3cSjX8bCJBetdbdB1o9cQmDUYuLkgUd5n4JTc6vmvWj23+Og8MlF7k7Oa34upauQNd6tKDsd
uM/BcxA9Isw6AeTAK6xxlY/d6e1DsGq9frLIEmYEbdXN4sk+v/DQbGGCWYclCDc73ELHFCSUtfQp
jR8CTpp3X/FplsOERyNlxdane5u1kteWazQqk0HubwHcibPIY53BMIEKJnqEDC4musnMTy+iJ/8g
OV9fFyJjFmEggbER4Fe5dfD25KjRgqPHR2YhJPleTriq6qoUmPSQW0C3PDnx2sfQdpTCWc79fEH2
5aulUmJPI2fz5VoxvPU17K8T8O3tZlOr2ofCE62lEbv5+lVbLB6ej70ynXGKeN7WWT1sEz3UE1ws
aqC9fKpYVuJIiL8t2bp6pbV8t9acDV8mSd5cq16DTAP5+pzSR8x2V9H5mx3WiMPXfgWERafqlyXY
kS0nC6bNdIMhi0I9kT+9GKb17FxPgvpItF3kjTEt7FR7dhgZ//gG/TGeioDhxu8w/ddavyjYIrH+
31W2BGT0Ljkd1FCulwWdgLLHTBzXKuh1xEHTBT2uaNo4z+2iASIk60RCEum5w42vYhE4QWHUE9YD
WHE+2Gt2MxVGTeyNkKFfhcz+vUBiCDhSLfPEH6dEWQlyRKWVKHLR4QCccopsN2F3NmEoFS973pNG
e5Mh5ojDqiffbEENKeV/d4ID5nSuVCx/DtCJsLqVs9ZxSRxfNPNlNa+1PcgMiweZNVAGWiqHBL3f
WTWdD8aC6u+6eft6ZeEo5zn0RKD40m9oknsNVNNwSIvEogHHrVZ4gBy0rEXFi2vO6cOpEpIwdhmz
pZ7jDC5FOB1Xc4v9ruLxuyQGvpwyGwjWbsB4WcCvPgbOXWcR9hts2qrq2Cxrmawk/+jDRbqHXgWE
SUWMsLVdxLoRXL67BSqG+HvE+kJBBJJMr+BrbKTtlPF7nZKBzQc283tzTZvYnrOCoLsxtkxtcI0T
x4OKgBSRy89B2SzFwiArp/Naib/14VrWyirXBE6Ij+p8rFx7G5EV01iLWPEsGav4zPXg6M9MDoi7
ESvCMVUuPGK19R95QNQgg2aD643W5efRarYsqmO1aAKE+7CsRS8X6n81UH2iM1che6byFiB66q5e
GP/dIQFtblM0h/q+0eHglKv2Yy7B3gub6G/GYxhHB/0HvyqZQOJGukm5OZKhYFncOCSUeJX+PGaj
/svzaYV2QQUpZv5FDYGgJaZZcKwXC+FuoA/Djo7mu/83nsLGCBKLQtbdK5GWpGGemLW+4eleyw+R
zWY9kGHUj0eEsV9N14X/C3Y5R8XhWr25B5yfW6rWK7+3/11RTCeF+/MfjA1Hqi1rSYbZ/7ZfmYqQ
66DwcZdH3t9FcciaNHjkzOdulNp7uapRN9Is/xz4QKWpR/0RmB1AcGMXJiIbQ5Q+eaWP1mRWTdvp
H2cITjPv5Ty8OrpiwbnZZktMp2nY2SA1rnqZdTA6ajE6wwNyZlHhVVeYsApZZ8cv03TaRC3D66X6
W3uh+Iz0/Sav3zBKNNQzU+egBfQYc3jlhMeWndayxbBIn4+Y4yQMmUqFvpi9lmPUIc1P6o68ETnw
CrBSEuhAHyOXeD5Eh4kCbTVAOm03rYO6/DgQBWI3/ngRoPhbi09OrvKB9NXyn70EWVzix5eGb6dH
qUTL/cGhbZy22yjjqwwE6DysBfeJnNw+kIeYgqoUson2otUldD3UcAyIHu0nJSRpf4tyinUJ3DTL
CEF8mIt4VopXHVaakRGH3grv99WOkLIwTngZCoMZbCx0poVibcd5bNguxgP4075y8wn3WMhiODsp
XEI5EB7sMGvkrD9ns3a3+qrWBMWZSBhOAKJNK/p5VHhvXy3dLVaBTGQLeeRMNgPMEhLlcrKmzW0g
oWvsmL/NRdRbBfnEIfLbbx7cTXeGtlqI17cR0HDbAiUQ9R0XCbgOx/YALhyNomv2J2z6Z3dVrRX5
553NL8pt59ae2MEDrHmGvgNhnH8/WDPBHuZHzKbY8aRsGmNR4sU1Ihrplb9Q/uolycxzBQSWExcn
PMadyT/YRJz5zuhtpB/oM+wXcXPIMyji+wAqs6RSNGksQW3kVbcjQFMJUX6lC7a8LdzXehcMyn/c
9f/YLQj9m7ovRKe/4sRwqCOhuLQHF/+fkhN0KsesRCQ71ImVeutJXuwCH7kJ22/0LmVUx3JTWr0G
JUcVk2lBHGMd7ijc0SnbwrZdBaPu1W7BX6Vtd4UAXecktlDCUDvbyjkMfGO+JNyJ1NsCMuPBUEQ+
amPsCql7fJzhxL+RH2iBLauCEOqAZ7ulJKenVmKHpy+KE5VyjYc8LxyMpywVy2msV07aIf87oM35
8UQx3ux26Bl+Ra8hrQDGe0MH7u+WenEUZa/d4aaOfQ10LCY/GHUc9T4/hLrwOOYtRpYGS3LL5jRX
YYeIb1I4wERmngpIre6m2sDPByhi/9jpfRLxK/ZGI12WunPGtxvxNKjbsVRyjL6TmbETcSBQgp9C
gAZNVF4EcNTfRyweYAcS2ctqgY5t/vFNMmaU10G3Y3HNPMAU6LrhA3NocsdJ3d+a8r2iwzoy2b9o
QvqMwbhvcmQT2ey3V32LZX06AVgvP3kiZCl+Ne6Mtt2yObQzG9bOXDZ5Wcd6uUf/DFr8pBVRWHw8
enF+hteYtO79riCIXI1H17Sjw2pMCQqex5wIz4vfozOSNdDB+YdOsXHJJF1kYbyO0hXvftr+duQs
xkOa8UUDlKwyIUvwhv/xMsW96pqYaYHr/Fv1W6eXOdS/4CTrEDCuuWuXzmWepcCMTSc05rN7CmJR
nMquQU8jysYKlzT13S5lYfxL4X9wk14kgAZ7g/H/+bm/+KoHBPELDo88yPt1Be0Qf8aVh7DWXHXQ
mUdlpjaIzkPrx7PtL0AalRaiA6mLx/9ylPn1sLh4iFkGCUhnEQ9v6aKvoWt0Q7HPBzqvrXGt+aS0
bQmk1zCYZFUPOrvKTI+szk/ehkd+I126Z917m55PvfvA/FhIhOlW/tq0aJ9DOsonQUNIWwKEd33d
M3PY/0fDrkgEerSNkcz+l2PjsxqvGRZzTFwYvUhDqerWrzps715fla5dbUsOEalIvSyOujoFHM63
5c2bU51Gsjsh2ugLBEjqmLtO2H0/KLfgvrkQ9PyX0QQ2psoDzgxi6TwAwXUaZkPrrpvQ9JB7Aia6
h+FWpN3wQD3jpOa28GGs1GiQSL5Yn/glMN+vJE1f7Shcn4jfL8zr3RsWw56yrZcnrswvXlGV+5Tx
WAmyWl6TM8OZE0pOSi/c6GaEkue4qX8rtHFH7iXgE9cG4UY/QXEkeynagEJhHr8A86yOAbyZwwnE
g0iso9VLCjgG+QI88IFPUBxymoLjue91ynUZ42K3jxZcZSXR/Gfv1YsFvkJh8jX60nExIPumC2eX
bpy+8gZybrQbPDzfGpwZKPtgS/lNx6vij7TIdocbxXv5RGOi5rDegxPX3OM03F/t6aevw5gk1Foo
uD50hbU+0cjzi9038pLkzloYae4uz6h7c3st5ZfHnqMuaYgf1Zh68rHHuDnSLasWYZXQtBd5Ndwr
Vy/hDjh42Yp+BMORad40C0T49GupL5Fl8oebIWzL2uDRVXgke0aUEw/LtT0btXagv4V0laOUQbLB
260QBFzgwXr6cpp+He2jWOEoIrJYJe1rkvrGd7dJAJzOutLE/DqXVRWpj+vIWXgwgttlhTZV2qQB
rsAfyriEhCEos1kEmCEyVvfsGrdiwtwJItFU6tHbVIv7WOJSABtrefaLFpc/XmspPaLywPPlSd6E
Tt5+Acb8rHnk8sI/81MCAhQLMhVq+IMBKpShppeX+kzAUXecABsCkAERJVx7ruUKvz5PwcY0QazP
c2l5nRn4snPyxHtrIYqrEQnS1cu6ahfi01bUW1UiFoKNhk/BqCNr3iCogmjNfTsJTib8pDJmqTRr
p6NIMKQ/LCv3C6LKravOyOJCZFwXYJussV2m3pyz24WRGi/0GHilY02A8oYO7dkGI8TN6DIynJkI
iY5uv9K4PcOqxGtr/dqyWaeGAjRsh1pfvryAQQX8P+LDVB+/fp8jcv7ywJQ3ohyU4ObFeUSqr0J8
od8FNsIOS6u10Ul0IrVvXhjPazX0X7XGe+qhwv+8I1uJn0fKAmJJDgMaKxlv6c+VIcuwhm+JXkP0
ZgtLPMPfXsv37jue91sabNz1zJnKq43miOODKcb4l1VkODXVFmvWxbA4BBExZ1NX8jJCBvx6qh/y
OY3ubme82DS0vn2JOokhsjmrXTi4WYekMhGXPlvRF36Mvo7r1TswpjKaKC0ym3KXLEgkbp8ketCx
RdYIhGE0rfxyDGVf4CiCnc0+w/mb6r7eopJbxFeznppeA+2k4qP9ecZJBJ5vHEKxk0HQXUFlMICK
rjNJe11py//ZjZGlQPQAYS3kW2QL7Xyc0++uKzB7Aak9TiykEEVFA9dqB9xc1rbsJal7cH9rjFf0
rTMaPO4Xe0bmvkU8Ya2XZOBZAdFinXEgfNVDFzL25jEPquYNZeWP4/4AsS5tL4G/nc7oVwRvh9ic
2znZP2jWRLN5S0RsDvwnG6WNlrs0KufudkKVmYSfvJn/eUJgsA+ZZ7/X3gK/SKxao8ifn1aedBT1
2KS3Jvgg2S9k0JfLN+9GYZPaMhdE3vOe1acanpJcc0fymc2aqjpi3QkjyABNybuLVVw2LPczMGYZ
wF16Csb3CZ3cjbZCotK4OtNpzPhgDb3ZM8mu9TTmcof43O7zo1t2tNWz5dgX7KDLIHHmHIQiQpvn
P/EiIOJb4UxKp435RmnvD8iWTAozNdcsijKXVvqAQSbGmT9EoNkg2VeElOR4U+8RzWBZy+bf0kr+
9XriK3cv4UJS+g2l1zXYx/xz+rQo8P+IIbQFl7yZ39J3cuXyvqKRsGmmvFhpy4P2R46+d+GbmMo8
C+KXGmel99g6RNGStUzaYEgKM7Zhng61RkBb2yI3wOFJE2b9K9nbigV32iDXJ30Rs9ro+lV8IaPS
IURz1EKkXG65LA6pS6MaEj6wkl4vZOWDF4X1s8gWMQS0wN9PKDQlgfeIfJGMQ0BwUZhTjkbpV+Ay
Fxu5dbYbe0q0Z4aadFc9zsC8Wc9NavH+YClq2SJE2eTNLYCdNX5XgEWAekXLBLe0TotKNtCSEdAL
aVnDWAXZVc5oG+MMoJcekHFkRYZk1zEVbpjN8tvVjbmuF311O7x0+vislFDYGuGwYF0bBvfQz8hG
zD5ypvikiaskJhJMm8wuXmoo2OvHIC6YfDU2WUWv84TgqJT4kP+Dlh2Lu+BUiJBdX2CE5V04mts0
BT9GVYuesm+4IhFDSlCGKHEfnBkFVFjoU/WbHgCIe5lYjjt1oqPl9tZyHiDTTqn8hDZjzDOSTAjg
Sg26c6eAvo5Mg8zWKJdHb0TEkfzlpSbI2V/wYdliCWRbPDcVM+QSrbNaDTijO+LLCPsjD/e9F1M+
bre2G80DZBwNX2SYvLzj8b75cM1jbR3aOFL+1z8Ae3HXlYItfFOu7Oh+8/9LH2vKqGn45pJjvC6S
y1esvg1Zv3aJYe/oV+uzelXXmUCRCnTOHDK6fRRPWidMLa/uWkAUL3h3ppYlyNFCqd9r33PMeH3P
y6m/SquvbMjtoP0GZ5JrEerXnbsQBg0+HTlQunVnGtyjY/HZ904pDrSAscruNW1jubNF/HNqsZW1
tFohFgL6mT8iktkZY5CPYv6Ywaci0vDvob+3HrU5X214eSFjz8NkMeNPsJf7+BBspSG+f74E6MP8
CQzp3NEZ9M609+Ktg2YwoulhruBZFYTRdTq8duFP9FaMbN4Qf82pOmtnv0Wd5qRTACw3tuYyQm8c
mT7qROrVBlqB90sEPcwBbqSYdhyQRy0rwLkm3yizIRV7d7VHEykfIT+Er/QG9TfGbJC5D3exMf0g
adgnhGFRQV0X4a5KovgUuBd2YEx1KHboK/vq4UeBKq7zRzr67T5pNSicu9Ku7E85+8za4u2cDL3S
kebmjpYbETgM4I/v4Nd5z7nL3HTrOxf0n9S/rFLonwQz85YpP/lqxrx52onnlRLpU2RrC3lmjY2G
V8ZHfpOb9DIMRYpGUhfibm4NW3ylDKzNZg4h130MDYThl1JmaOqD6bFc5eJZYBI2I/zF64RlBTGR
3x9MvnBgtKwhMYQt/6wMde7Dic+dGX1gMisShzeKCBmRCpN9nSppTqSOcq4apURM9R0ZR543vcRB
s7Ts1iBn5fWz9JGa0pSXRwqMYed4BD+uVU2ZsLfBvwzNymzYegmylwqTFkREsmyD9mF7xcwpm8kW
dYnmgYTQGgaLGw6v/tjixFwHKx/hKTEobmaigo60rsfbA2qt6ajPILjW4GtsJ/+BpHVax94mkpFP
H+Q8fHuhKoSIJMRpgvcoGK/+i/5gwLU8MReKpqLxwBX7Nu6gUjs20vpFFYIGnUtkyGCvenXhWkRg
B15fzHCFESGnn2fdC6Ej4W5pzxJ6PazM3QIW2ofmowGEjyCj1F0t7RAucsw+wXtRD5dJoZyp0MQW
oPOkCU4/+eaqF8K1NX7IXuWpftHo3P7v1UIqd+JgZ+h9l5M9UrembVqa5wQudcsxthJOIAq/4K+d
dBZTN+dRXNUDmO+6w3z2mW13Hx+fgnLfDkJjwAy7JDriHuDFRakIipzecPszOyK5hxtLNKgJS8xO
Y/3WIxMohEb17VX+GRG8FiwcQ0u8jxkPdWOsKwoYzkh5cigQjiHVt9z0xv96d5NZKFIcPAXiQRbf
B812l4Y8f9XYG79jPVef+dVqZerRaT48QxdnW8uFfjFLvb3M8EIGmpPbS4UuA/13Ad/DdhiGkT+s
H6QLvAtjNWiBA/fjLHNzv4L/PB32Huf67dPL19eveibrSGjvnyFusxH7vBgPe8oKvbOey+rspmSY
DVsFXxp5/US/zsByFUygw3b/kC6su0vUmCE/j7DUhAwgoDOrzF/dguVjbomhz37ca0TiwN5F9XJB
pHwatZHzNQNvtm8dCHyuLZ5OnCEgAFnc26RrPY59rUkWmDa+Z4aCFanraMZMu0hIh1b2gFA/ehkl
7YS7umwolDlKkTi09jTBEl2e6t3n7kNtDCcgKIMONDq4LS+WoAPNxTjq9txq+tENn0PNtR0XsA9j
/xxCwIW8hIhCovmo0PrrFunqklTiMR5mJ42+pV0qwlfJps5b2JSteeFRhkKf087sTY63N4i7UjDE
rs9CTf/Ne0zLquhLIc9LbheTxhI13vAqwv+BDgLMeo1xCPvEFpduKQ/K9HeHosWOr72PieVLaVfY
bqjBNGsEJPe9AtTptNoiqi0MF/soGlZLx1X3WTNanjCN+uDdpkUSyv2ROWi6c9QQeEJQPZQc4vp7
x0xjhA+vvdQyZjXb1Muk+svBsJ6ao5dp1kPlI18V8+z1NK1WMzTvdswQFpZKBjrXcPhU9RSQOgiC
Poxa9v8v/S6npDYm8JjVMmT7ofoUEGjg/C9n6YxHsGXOeNyfNxLAILxDYIYX5RCkiwbapoEMyuCd
S/hXUjLohJdWml5S0SPjOuCMfzWDNHpwmPyq9vLt2yIJAXXavgrOiabdDp/Tl5g0/dCMUYTWdw8V
VPPyTUWAqIn4eRAz2mAWZDNL5E8krbOIEr96aPNP/dGCc1vZQjn76ScIBQusIdOsJyX0IWrugVW9
pol1SUbSbGpANMb7CaSIQSQ3s7GmgtQnCDKWHPAE+C0LZ/LrtcBfssTs4UqIWlEEwUH7Obk4rLkX
eEwjIVMyxitFVdFOMEexJErjiECdNrc/VzGyiTWjb+edlFo1RTVNtXgTWatyg1n7WjG6hkw/7Xw4
JG2aF69VivDd15lFyT2Uydp8sL0A+hBDWBgUNLQLzs8334+ksivUpFWH60dylna8hBYYp9exglAs
dcfw7tSZIoo61CkUC4Z/AsrK9DtTowr6+ouR0ebCvewlGlAElp3FVe3aLlkBut3ypEcAcj4oSn1U
7Bs94MnZZZpxjBW/drCFgA+c1/kxHM3gLkFH80rgqRjVvq+RBCjdOyRhCW0mK3N6az34WStX/Hg8
0qSdtXzJC6UxExgxUem0WPJ+Y1WxqgNzlNaR9JixN6zd9hXA224Ge/8DikcyWgRTLACf83eOu3ob
OyYftEbwg0Cjjv5+TSPlqp3InuROXz8IMrC84orOxSL/W+1BU7uOkfKYn3GDmYBIeixcp2zcSpWR
/Zx11hybZFcpPpAzVP9S55B2UDe8ae2Db0PAkMz7FsC+CP40+0MkChrZIL731Z58z7IMNIYsoQms
YvNRuMnynC7qVcfql0h8/3mXM4yTMv7g7Vu98BgovivYVIKR0Yyn4nWtAMYfz/sR5YjK5lg4i29c
lkrKa1qDDsKSQ9u/YbuK1De/0fHPHrH0ABhSRuOHPvF++VlAQW8H8z+ba3UQQckvZ8kCJKXnVSp5
H00zbNxke2XpnstqVRHAyNOKmegIh43mqkHifGLKJo+uf9RI2NxvLlqmFwCaj0hcsVq5HW6M3bzL
DFuRPlAJnxkXlkncKpLXxX5b+gpHzRX/+qtCwe5I6NNhhv9Cl5XKB5hYQIVAoc20CjL9GGUxS09+
P60nERQ4E6hdMl6SKmA1r9v3t8vfw/4LAwAMdrfjXwTCiGHsxsVR0vns4nmWataG8Oq3TBWkPiW6
Usv3e9XvVam+o8jzePTDRDwn26KV8tw1v3rWyLqwgvqIzI1GRXPPJXE7pj5WkpzGesM+cv07C80e
SrsLpAmnJsnq01XA8TfQfCCCWsdfo9xIt6P+SGWf88JZdNchMk1KftU4PnUHh0JAAPds4SZQUYzx
9vfCUy6yU7h/zE/Y5vvdS5UYwSQAt3wd6YmZhBhcexcOpr6Cd2O3JQmOYjgdMep7/bCxNCW7keMC
gzJsclsT4WO4x1j9uI9lnTrqi8BzRdp+dGbThKUmK9C0UMHSKrqLTyx8R3Wr2y8/Hjy/0TkR1JTb
W3MUWddNTX1rHjbma6TaTyBJuiUGOZPXzkjn4zGMlABJgNBpiAB0qBCS1Zy2VGSEvGW3l5XtuLUu
Nlqkcq120MKqdU8L0hoadTzjaHNunnaI4gJ7Sry+ZEz+14HpBbrjEhTRW6fqL6Lxy+FkfKtmXFI0
8b0Jpsf08pdH2wzOrIwzsQsn3dUAq9GyT4uXZ1BQToRtx079vAd7cFTm8/qkVuMBMm9Hz+ochxQa
jMN9Lx7IYqvCbr7y8ZvhMDzVvlomKdvQ+UxtPqpKMiCVHlDgN84Pol5r3WnHZfl49Q3oEHJNZydn
LJanOfdBeUwcIMSaf/tn3Ni0CAJnICGH17nwuwipN8das1cRUOTLA9XOrbv8kVepdKPUulD5aQDe
6j937ojy6ZuUDWfFxLvjateFf2XWgJhW639PPwWYQ6yf3WqnUinixVKsP/pTqYWIZHd5CXolyCmY
Eut9b6jFXzpMdxFdfvz6GuOpQjuZ2mTaH9qAGcSCJPvD4xaRW4Z34m9oPO7xf1m9Rl46PAOEoKYR
zDXU3FAHpTWaQvWoAh+YYTUjKU7OxuUkRwLwOyWgxW16RpUSf+wMBwgWf2AMNi7t8qtTvv6/dXxd
Z+GHmDpxP0d6ZV87ujKb3pvYgcRDpt2MeuX4PyxxmDfwP+tOLETey6PiMthdT1Emr3ueYLFFcv/T
Gzzf4qyXGr4Xa23Zo6zHewusmPkPmAVGw47ncAGFCmLP2CUjf2pnQ3nJPcq8OQ8d+gepIozhBaMo
sN95FrKTa+c+1uqoOvVZQAXwth4H+/WKzq6VOcdey0IPf+H5oclMxQ5BQwVgg7dluTPAcpMtssYG
TT5EBZfm7BGk07MQwReRib5NzNPvWY1mjgDRgQAlSkAvh7JIrC6VIsa6I4v7lC8hjBec838uOMmK
bOJuioTRjMT6IdzYYsyFwWRZI2QPCaBPh85UqjpK6XSL9r2J0kd4g+gZUK8D0tLUwKJt8SOuFPKi
CQuOISOjQocHfTRC/DgvWTyb8q4b3OsDi67cUH3sqyMki03lYvZETbw0s95dsWCzcwgv2deydiCK
Aqda2jN01MhsZwLbyfwxLj9YetanBJe0ua+kk4GKTdiG9yG6t/1jJDyJ7+d5xQD6eq6wC79S9xbr
NZsU4wuIRsRXP97n0deS9JpubAVplDzUvumYnc/pWXToUa1Uvn+PnPlLhuedko83cZT05Zujb2Ls
5Dl+2KYjChZ2JruW7R3XAvJ3g6PRNWDRPGPzTPldg33vTOcZrgbfNx6rErs/t6YLQDEEAeQzZc6J
+f71kcs1ITZUqzZmudY1Q4Sg3jFT7Q+7NH7UMiCHx4acl5B4w92/qiKHiwQdCxUJwC93OFq7mcm9
JyVG98q4r5TxhLxXlUNOiTtDVpwb7t83r3llDXY/gDZS3b2NP/FOGlvkRFVHJK/3axYQbZpbg1+y
hmzuT85I7qSlfb/SuU7LZPt23McQsb21CDRgHTu0Dy+BzmNo2nGHoIqMuJCNXqO+yOb2VjZe4Mf+
XorkEHXnsDMmqv/842OyPJ6ddHXMd7eJvOBIsVzk10jflpNQNlW7dP9/r4ZwggFfsfzzj9Lur6Ap
ZErezYbkFTMLABZCMo12fU5zSdo8fbkzfXY/4LSmmMPbrfj0zADuuZNPyiQ2kQpKJreKrrZiK7TT
X67Lb14lGQ0kj2CGVEe5x5OrtgWj4huI6Phs2/x2Hudbhy8Ycgd4UsNWb2iRKB1iYVqmEfNJnyVP
kqZqCxOnzWv1+rogM7p/t3B0QgfG6KrakScOYDS5X0TEYz2Cec2OLrLcOwnSYEcb7+tLg6WHnCzN
nkc8EesDPcGaTpBkSrgTjbNtqCAaKLt5MypNm8pr3vNxaGmBA+Vn8TwDh0Rz6Z4cgzUKhZsGch9o
grhrKX15BfYYBxWis0t7Evf2VOJ4DojciIuRZ7qGZivCWpNY8IsEernwE7V99OB6sIQC+S2lPsPL
7mjX7LJdiehON7SLcd5AjbMfzuuKGLbHyibMIvx99BdXTNikyPhkuk3PYlmeW2qUmFAqBI/l6O+x
PiekTAKPYyZ9u4Bqq8XaT72ehOsYW0fIysDTU1du/N53Ba12ul5+lMKn9JJovKs6z28krG/FlULb
BoNJZMLswsgAy5jkxksqnbaK3XOfKyqYNCa+H31m68owgosHfxrWvKA80LXAHbj/GHOwa4TFnDeC
Q+/QQ4fcBmRZhsaLlpvWu2PZYsGYDuzfM7PH2yYoKGQsOkTlNjQNeho2Xpuqv0dJcxe0qVNAPqep
jJFg9frBuBywyrCXVh/U2s1L70Npved2H9/c3SP5vITmcE/CHAdzCMFO4qk9DFMXuJAEpqeb9ymN
7yC+SjMY3o5g8x+lP4znn6WoQLNn5+4kPz7b8hfDvKgI5Hzqnq87kwEjjVswUqZ/uJ+eqdJnsH5H
0tCPLT6JZ2i14ugd0l34okOcNYeCKuCqLUdJkNZjYxtuzFS85DlazxewblLd24cKA/ylRoFqrtan
1hlza3unnoAgUqdAuxvg/c6gNY0BP+6DQdH+XzjpKdJoKjq1j0NnyaRZbLzgH3L7Do5aEWfUrCNe
FFghzu1QdetRjXSF2/vq6Vzr4smQVPBPvieMEtOAaR/fvV//xlGdkHzk+91dNlMEx0Sh1qBX7aTr
I7joEqT4NjJecvTHHxexaq/dwWHQVfB/2dcxM6pTAURDEvEG3+giKq2ZSJ4+fvnvVqcJpOa5G/KG
l1SqtKNs2UWqUKtfajnJ5LpG7VZ3n0OtumpnXVlpuVTMU+xBHPUJe4OcYn7kUpYq6aRfS5UEcyFt
NLg9BiFSn2+lTyDpO0Lz9pmPuJXzUL0vodTSN7YAEhjP2more1uM8EC/EiFewrjAu8Hx3gICELig
zYGE8c1WWUFjKtJ5HMGwrSUQfPGLJtxpF0ogPLZSZsE7ihiBN5i9JlYwcxoLmT+8weqZmt0v1ooC
cPfHWZ3+bV7z019XnnbHB+iUnVJLQGj/wmx/ZUsKz1LlrcVXdmUc4aRe7Zj6yXwtHOxTgPJ1RIz3
DhvidcoESWiYZbSa6qHM89TuEe6nRv7APaq8HOKip7EjDAMQ1D0ZK55UEzj1H57d5I1NRlaMMUbO
AhuKUFYI4ca93AsTPyi6BkTlnDqF5EFfxNLasm+O8JHmX0+pDmfsrjlDA+tI/HrTdDNdR2fxPGSc
PXu1r2Ah697+suX6VL9H39QhswG5GmpX/wPGQvsomhrmSsArSsg2eF2K48RrCU6mf+DAiPnEKZqY
Ip7cg+Y2jKekVKKIgdY5adxGKZc/055bemGvwk6MFdtvzw/hXTkYdasq0pgcF4tCWaTADTdzc8nA
YtjyZWH9DtaHlcqiJiTvean/sCh4T9Ba3obboKjsK+Ln8IQnTCkArH2EAwTR6QEW1VufNY4VjCWR
vv48vFO2uRPzfvy1dNfs0Es3J6GVb9qcYZstTIte4UX9Noxhncg2XS8DT0puZmiIew3ybNwyvK9H
x5DUniU9As+U/znRK812RfB4+EUK8ZA3m102UTxs+qzZfxCKhSaJZ8N5Vwql07gM+y0TS9o0cI1d
sbw/PV9Vui3qZHz7XUB3IcJDHJa3Epr3WLXJvhT3fiL2iMIP1geYQl1zdYvwnAAGzkwzqOjf6U7j
B+IUE8gfN9vPooRrvcpbBTrAyvUlYXXl+T/D7SQ0QvAyku+mcJz1p0E8+b6izWXaT8UR5GyqVnYG
Gt1macs4Gw+ohbp/IGNnKtB7MzqxT3I+djIs9ZXtrSDidgByxdJ5A9nyb5joxPs3pUg5sBGFtvSH
TxBinP0bpb9gSGewvfxgCG4bfqOiyQzHKYIlGaNgmRPCawOvu9faTYihnlNl/kUbmOgcGTkY32LP
0ZfqxX+ZH4YWants2Si9oTsWV0Ktdx6+FgeF366AncJYzxO5SkTvQ2wt7J+Zu3ueNyPab2w5YNwU
stfV/zcZ89VW3D6Hp9pvomithkJE7PkioTyIZYOLd24hAX9701fEpWiQfdusnwT4xzHY9zBc+AbK
v97bqB0vDrwVpda0onc9uS2J9yRSEHvqwh92pl+pVFw2tvyY7v2feG1/Rtjqr90f/hWPhlelyGWb
4epdsTFo1ZNa5GCyfW9saPhMN8uETuyKdBgzzpaJsLNdSebMl+pQLhCG8rAUX9Hlvpc52NQjIpo3
D4haoFOsZ78TAKeLcE3deCTr3vYnO2iJaVzEnH/Gic5iARwHVqqgvDsCFmnzdqQiOJIBImNoKujA
4EfvGcwh8dT95rZ55tKZFehODituo2/sLYkCz4eHGnplPqlbIffhR+Lh4/bXzhGV1BIiQZYvMgqY
3gQnBei26YOEcAot5xt+rIDl2cuMHjUBkDedLubke5WSqEVS4aSfNNVvVJld1sAyhnMUhFTqQRlu
aUaCms5sq+J//n2hh1ZoznG3JgHj5G8MqR/B3VsrM2JYyp7Hw9EBSykrQjJ+TyO3Ya0sZfst5k8i
zw4INN+uCkVLszRt/lEGzAsSkC8OpuHeViydKPowSAFS4izFMLdtTOyRLmexberkHmvmtTM4WDWG
EPxDuRQKtl50CDHSCdmhzChrUrfUAfKu/o149+ir4tWfbdr93N8KCRK8tE/pmR7DPnMJ3M+ql9gX
qxdfGYFS6dXAneYIVghndG/uPBKg5UKSF8gDAWPVmfidyU4Ryj2s4QHcK40TAGOhMJNimqaZU39J
aFX5qjif0lkPJpxgr33UIXYlpr9zVQLXLljXoPhcOpA0+Q9adFr2Z6AgEIIlKLH9UnzUpyMVvYie
IN4KpaaDxERtgPbXzeFt2fYL4fjss7tjAg3J8LiPS/4iF0ATo/1lk4pCSXiKUoigc9YiCOpwQ+Fy
aiBFVhOXu4JVbXUIlE16o7X5C2aKQ06yAZafD7i9/+VtGi9Pl2gPdseSVI+A+D4ggdMHYUuUjvTw
EB06JgCxtMLTnaG2piCIXhvBGyiEz4EOu+8hcSk4bNnV7E0taADhUo751HYSPG+VcxAbNe2VGdMQ
ZoE9nFNj5KFOG3e5xXBU1KRA9K9yBL3hhSvcH5pMBtgXENxypChVkRAnxDFghMitDeXuIDtOM0K3
RT6zjfLnjFFKBb3bja4OyPMafEBx3rRRdZ6sqcT3puvaLMZavy5WmM2n/sBTdXpPTubnxoLqqZJP
JfvPQFPhSAu4IlAcRlOFGtehRWq5pM+b19KW2hZNHtAmR1DnJsBgSl2a9Nu2UWzfik9WuECd7Yhs
1a3rxzKaDfTcq5qfv2SqG9SXxzaLrQMW1ym8oQnRb8t16GoROt/zm4TeNM8pleDOpGqfXeVvPzzi
Phs9S/zMdDN2BtvZHklEHL73s1AtXtr7ZwIZCRpNWJHYXv9K1OOBYNXNZH21EiJwC6Qhkb9qRRJY
quvkG//QoD/mdGcjv4PYYkcfIe36XW29M7tVR9N+L8h3E9HYxbPTF5F3Myg0nW3uB+jEG8lkLg3n
vqVfuoTvAmpYhem76hdiRkyZ7spY/mYuFVXNT/NYPfceDKGIP20oewXA0epCbGB7HLJY1DY+I5n4
X8bMnTwptUMyzFZHjCAsY6DYqaHSiU04e0p2Bimh7zKoAbGIwjuMeTrvBc2baPlq6bzP9+GfyhrJ
2jeL6FTTJwrG9bNmp84zDm62pldcyqPvrj8GsIpsy/sxG8E05fvnVBgVwXwkH4Z0kfEdokKYEc1T
tDN331oX864i852V78wrhxeASuJx9p7A7fdJadrV6XOy6Y3MzaaCEOcdGzGJIpFYgisHdTUgLq/q
e5etcY+QescBfVehtUBQgctZUauVmiKJ8ZnMk3ASZ2kl9tf+OzDiN64LpRUazGax4Y7Z8xPz5qU8
bBwhnbPIDPI0py04vwToD9K+gdrUULL4yAuWp2i4cW9kGFuO0xDioNTEUvJbSJQEnu2Dmocb26Jc
dYdbKNTS4bWg0NZeX8BpRnltOB7WAXvjaUFZDHlBLV2lLaraOh/SKizGYyTI0pr1cUcIZ24RmJyW
j6ZoBWzeaSDYbPhx0EvgP3xJAuvJQEOYpk7CAQ7LiPa5D+8c/HeUXDMspBkrrvMwMb+5/gSVx2MG
tSwtyykxmPWnNcecsCKbPETN+LCcxKIhDZ5VkX5Y+aOpUYGj7vdAOBaPEJqPkr54AcZBkDvw0r4o
rYi7JcE+Lo88wX/8ZEnhiZg+hnJ5i8TPYx49L+GHnpjOLWRRBPsUszIq6WHIyxYTtbKxn+9II0iI
Fo8EnNcl5Nd9L/Amwn1ME3yEdY9n4Fx2p3UK3NK0l2yeY8ZtRZJvBapoSGUkCkCObx0feKLsF6+9
Riht9L6UgW8hQG+9OnZwyzs6juMqI/BAdFjQoXOa9AGd7NtcGFXYlWJE4Yq5Sp8K1bNXc4TFLReT
wIaSa1+QRQ2yVhNwiP/54L09OScahK6taAtWLLWNKqJtAYt/wjYO9lx8JtUqFlmQUPAiRi7bS5pL
az8QnD0hHT77ls052lXI3qOduGquLHxTsoo9ahJsTfxrIyRQj+K6hjB9aRCYd0vyMnsaemPZn6OV
DqkSmpMCvUEX8UnCz3vkPOOOvVQgeSSk9pZefpaSbkjp8FU5v28iQSmMcHfrJ62Taq4udmwRjWDv
2Z5/jDbKgU6npGBzqGGOXWEqXZp/Pv2+e+dKs1O3w+qwNQGdB8c05rf1OLVllfDyAMc5a39qF32y
EseyZl71RE91JN3BSRlyVnbF0a6KPtC2SB9uq5uPtRp4vU/lNNjQjzewzFmE6b68/0UsPtem9Eri
MEAszL2RYsuveyt80SPgzrF2LagS81A3ltkv0R/u7ZzCAgyt9J2xJTcWC1brVi58ALNg9ofdCK0o
dF4apcMimWx9RR14U1i5WYKOIE1iWatGUesyW2EzsCbBnagWqIpqijp51OGO9uNreBCjIRU335AD
bRsIqfxRLJjducqzOVp4PGDXI9boqzwQ17+glAP5AKD8h/51Fq+cvKWz+OugVCElBCLyZ2JoIsat
frdQPwKyiGrdGN0WcvpnA1AsvIc1Q7jcnDTPKBE+dm45fxOxQieuCT+aXC1E9UDyJ9xVeLPE4LMh
pDe75EVXFiFhIYKWf/L46YOOAZskrqBMe7T+whdmMeR2tGllGjkDRjoZSxzXbUDoTNwYp9cIpzh4
fFIrSzMrQYNZFZ5qZwMCHSmjUfuj+C1dwBbzCgyVo4RyxoQpftSjvDZxRZvaly7yjdG6IXxEhqWW
bG34Siirs+QYGutkdi2Mx36BxKkfnQ9poIERsTYwWmMcnqlYyxS/w1r/G8/BIbM/c9hZUqEc6G0s
8LbNqE+u74DzfGyXzqdIwZfyrVj9xVGBmsAVB03uKA0Ew4zUgCEmD1cgjeVcEldlxSVZyCCfg4b6
98+PJpb7iU7Jsyd2G2vouGnmsilFCcWubWHJ8lEFixVlCbNxjbwTkCSFHdY+xbFnOt29l0bUj3Iu
Pek1SDI7sFDimAvpksaCNWqgHevwaurjlVd6k3xcptjMXGYpqRJ6xpRMrcisTeSoVRDUNl64AK8i
fcz8itB0Fr9/nAd3hEbIszhaUfRtzJ6ZaWLEpCniVdeuZW46ZucKKqzQwzAWpEiTPFpGq2KCs3lo
h3/pJUbjbP9J46KDXp/DaZAvflZPKh6alxkDGG8nWCPM4cKhzBD/U6iE2p/NoEE2uq2M4khCgfU3
U0hVxy0ULrC6enUqxF0DJBn2Hd66svQ1KS/axC6GOWOo+wbEZfKJLpE2Fo0v8/FQdQNo8KlJF/VC
EYckXd8Hvd9rV19u6kZfC7+YdSrfSx2mUUmEbZ1aI2b7JaTwp3G6SUkpPADcmXs0hbIggG8raoLY
iyLLnALkj6Hao6VKl2mLMR8q6YzT6inFBxXnMmn4kp/4QvsszNs6Rm7C4z87ihZfAWT9+AN1PrHC
nbPKCEaxZaEBn/llK4+cYz9prL2t9esGs8zxD53Qnwm6hHd/KnIC6xsIMLZMU1sohio6wCZTku7W
al3/LP3mZtQji9RlnGgqdXif0gi2oY0BoFplwW5rylPuTveIHdb4mt4UQyIrRqFFFDNcmw4OaPGT
OLpGvqiTHPNiQ6UcA5wAlNv+DD4Cq2YJMH/yGJlilcyIR7BZ/0taNsYm5Qf/YxWW2bHWkFuNVwIp
M8v3oozS5nuV8gMaqa1QB3nigpf5R8Q0CL69+KHW9KpVFZJzekBpxlusaiLpeeqXREf3nfa/Fr50
rAT9nMq9L9rXWBskWGH6gCWCOMJBqeZMUBqnlS+/FQO3KwdDHdj6i4MEnV7QZau3udW/Yvr2vtn+
g+qCj+YDzeRopeWa9dLKeyi1Df2C3SS/USNGmbyp0ZK1bZeSjIdg5ciEMttgZEoKLOIujj7BuyXW
c5iBws9guZOKudWfGQZTWJ1YCVJN3Le6FWUE9/qVCdUOSL6ODYsCsaLKv6RfoaCsUvy9Q34pg3wb
M0/0BGBGTXYUI2/QltQG+SNhVdndN26Hj7lg/34qv4YCEjut2HTbOkRk/Fc3KDlth5yFHQ7ftduc
gviEoGOMbAPF9nDkpFSOyfEkCFvX7BOjcSXYLS/BFXrV3+LSF2F6HcKU1pTfvhRb2FZwB1s58mFo
bOQv2+MHQ4Z2Q10mLn23kr7knPWfVgGmjoju5XWRQy+fPNUGUTpPMTuMn23IOpEc9T3coi41Rw06
qN/tV1t1JFFh90oQJgeOJzpm1QYhqwlVPReFaStuZuVVCSiUqAWjjl6KzcaiAFprLV9jPkdAet9K
hf1qY+B4GTuh4IiqApWI/OC1wqi/yIxk+/fLzQx7BQ3GE7Nk3k7D5gESdBfn9cgcMjLjGylP4v8E
dO5uwI2xjp5TB6W0a04T1b7c2ww5KRUKIar/KvQzAKXhvJQi6xVIxKqdB/Tnr0cBUDzHFgBPLA2x
YYMFD4Bjs5ME7xKHNV8ht/xQJ53e7fbpiU9FWqPnVfGltmjY++mSBMcZxL7WOTdfigNNR5t0/A+7
A6Iag1RTkKhHX2cNCJBkYiyu4Tz07KEAWEGHCqLIHk/UmeVsbT+sKqiAaTh00WIQSOOgicS0qaag
jlrHI952NDtNl1jGn8k1YCsyjlKNZIZaCy2G05OIkIAaUPoYV5Rec/kvVuQ/fEfmed+wlpPExAyx
pgIrGn6/W8NcdurzYhMATT77qll0oUcMamn7HXw0KIp6C74E1I6Ua/kY6fIKzk+suCKbh1VPRKwp
wC8hn8OxB/s2QMjq3WQEIxT8r3WvdZrYZwLdW50wqbknA8ShTht3O2sCl74Y4jDVxP4etGK1oCI5
sJVCmWATS+DqyGiUAlRsHdySq0B4yY9MTCb74G1Bh+oh4W5ejAxdYZ6+riB4+Mw2XdVRaKf6/98q
zsmb0K1PxJO2fNDOoESudagpP8+UcRkp7u0xaKComCb1ABXgm3DBQ/W8R6O8Epo12DF8DeDBN3zz
wtKJYtuoh9t6OjQvZYNdwmH7vApMwzGIcp/zFCkkogCw3gwO8jz1v5GXf6hTo2lj0tO1xl6O0+60
2j0QerOojvu139PdqOAD0WyoiH9Z4WGP4xsJMjlK8EoZFMenorJ2UEk58kAIlgvVXDai0/NYjSqF
xLG6kSyguPdveZaZb+tN8ZCbNHDkt4vwtfuljNay+yuMymS1f5ieAgPoMAgPM2pNUM2srIKYXneS
kdO+fGe5myS2MJwYeDoWzBC2oZuSoGT9123mjnJR334xxpIo+wZ4SXAEBBcn/gJZe0A5LY/ud1vR
UqP9Ck5sa2Y+17s4zmLzi8KfznYbBZ/2bGjW19hXrjy0isLj/M3Ubh5pXlxtVlSR6S1YAZCUM0pL
tuHEbFzO/fcs8R/pY8V9wXDRrvEcx14Fg884OFQhAh2JCi/uq2aR4vf48IWGNW7Y/GhwRBZhjarR
tF2p93HQ/WcWpmT4vwqKsIbfOY80A9RRqF/2hiGRa3a502r+/K8R6oeqK45yZ1L3QGvR/Nin8kWF
3oLKa+fCSYmT1waj83V/yLZ201PVLIAl7QRr3eVuqYscmENVrJLqMI5Pvogbfgm7GZYu5ODzaZq5
P3YroZaSkklk9C7RY3j0twI4PWX4DYkYmKM9Da6VATICW7APbw9kVqSAbmLTvkPPkceU3X8HTgJN
2X2F+bkl4akrWL374XrWCgt5nmG/5ACzruQDORK9AzfijPIgfhlArSRsIsnzrrQ86iVC/tZ6PEAt
/z5BWtxTpovYL/afpegMSJ5beDxyCGhnk7pnlDsR/gL2RBBniJQFdGTLJzZHk+4zEA6kB+828IWG
0ZrbgI+LyhZFqdf7iHXVghGiaS90SGp/EKQqPQzaEo4L3N7v1OpK1OhMfUKV/uLUoxmbu6cC1So4
AMircSq+/vLydYWUx2OtbkY89RUbw0O80VvN4dbXhYMk3TzMxrMizaeAP21O0sAvKdV2heFTobok
+rEDv6R7xE1C4acRqocU89ZlOABbw3ys/hgdorMqvBkLRmnhWohmLlJNYvNSbTSHmUR8Zjn6lATL
1dXiMlykyOrZKW2fwRh3yIo+I55HKtt1XYa4erIb0XzE5xem3W90GzXAQxkyBQaPPDBIJHL2PivX
JLYE39EQQYBB1KrPFj9SGJP3eiEh80YQpKWsRXkZUWkUxBNnelrMld+lqK2E9se2D7SXaCtkc2PK
TbL1WI7Lv5Bmse+UyUSlNv/h6WsSSxGOQK0X4BH9nOQXM7g0UbzUWgFQVQTt5Ix58O5wlkhEA9xE
A006TLYoHDbdo5tbNH+Jbb8g7v7FMsjlg9khY97xfvGPk1Ibrrh4/6CbhBeISZ6OM5c3uKzWChq3
rBq57Y9HhXGiD24g8kMEOY7aY64Z9DqRiM8c2YxKlXROrsKr+9Ywm9oHZd4mhtPDkS2vXU77YVs1
P/F1Wa+8xoLTlkvVIvqZzHIAgwiWhiz4EcNoEa0vt9fJE2fgtScsuVn6IEIvEmETgBGwNnKr4yjV
GaVN1E5aMoTtWNPGL1lkKvdjtXbJfKPmFic163QI8W+/Ao0U0p4JL5Nxc0XfYTzUBBAv7tD8ZG2x
HKNpnhd1PXxYToLiTmDLGSeThq9ZATqie2Vr25gqVHBepx4tVyVcpdaMIrXVCfLLiAmklx40C9kW
xNyAIbo32cmxMnAVZqRXF9fTm4U/6ysFxZlI64drU4fVgplhtX9MWN1MfEBIED32RagLqOB8P4zY
nvpPdGP4NL+IYzFWE50xCDnt0rjtCSIHn9abU8agIhoYwtFMOUAy1DHH8Cg0vDWzVO53Q2S+qqhu
SDYghCSE8Y/tupqMFaQtGAFyBHD5t1hHg8QhIarbsZuTi491Pg0ym3BmSr5kGITWeZo7tybrlHD6
Ea5FSHJcbNCPGvV+zqBE3a0IUjHcJ147P3MFxFy/g5l/eIMOhoOY8mdheu2F/EbWtH8mJmIBDxmQ
FJyn1zp9GK9yTDuUUUppTVLUBMcSsgVsAp2ftkO6x1PFKFvuroCCQq1Zi8sDjBVdUN0eH12edFWz
MSwFbfUbm92MM9+X8t2BwKdfvGzmNnA6cNspcIAEPzStiEqSW9JXrrmFKx1cBr3vHqnSoVNskIdD
ZdEhYHl9zLcv3y+iplBepVIdVoptoHcIFZe9+VGRRED2QV8BrT2Xl4UoGVE/e/B5t9SFUPncBwCv
EjQNQ3qqdGXyoe+Qu7lUa25+6BKqvLC/15pNWy+3pCOaHMkb/KFXzWeUn2q3wiDyMGKwo2uRUNam
Db3CTgRddmInLzfbqjUXlvl8dBv0fdsOAlE1AfqpGMc3HE2nCkBtnLkmbTbCgcWjPhw/Bhl8bwGD
4SPZU3FJeDhp6W1u2Lc4NnOvwgBMhQsWwsqj5x7zis7Fe4hdBlc7uxMlXFJfw8gJwRcjU/XokWsD
lNAR58nNfbOBSaQjQva6P1IPAkwGS4oEmMqJdn9OVyuIz0q7vdCJDrxfSLs5NVc76PR1Z34v2vjS
cziqxZhLi+q351kJwlUzFfekXUf6tuOmNLRnhfxgCXAGZ23iEU0dXTm6yDPqvFnI7ue+5Y6nQAVv
+OstwRe9l0Ywe/xUQZKyu07yXMfQ2zFl6G/SISHfONR3wxjEz+wUD1ZROKsZ4+5OB6a7uFnZBbVd
orZBd86aqFmNGTTa7M9SMcjV5Boj04k9GQQtdbf3eu3yP5EO934WTg3TJECHKhG6OLWZ3EE0B2lS
RJfE0KPed7wSf8ngTLFCqAptosz89olWeDQ2GX3Yz+X0xvlwNk7DAQ+SwSQz2R39T7gMxKTahqRc
czLjfFpcrn6hnLQAiwPw/UjiF3LrEwpbvJwcSVt7FPKZjzmfmkHkzfBvjBTfyCx6EQ2JgDgza4s0
EiM0Nqj82/Gu6nOwfzkPVolYHAooBxq7CcOluN4VPyxob2BMpCUrH+vn/fyrH/RBZQ74LLRT+ruB
P/2WCRHC0G3yUGYwhb7GIjRsmGM5AxFSOkmymEuoOC/N0jTGLzSCWbrawBoZwXcFrJK4NC/vFfNd
s9BUpcRNM+q7SglMZKo1U4culI1Ejw3AHDZyLR76trKAcSfAqFZT2cHA/ZlWpii+No92P1nsRX7s
xETl3EZS7ljqXDVUCecjqSc1kWj7JtWQCirj1Yo9b3+KxyEcOYsi818wlGG1Hyv0gzjOccc8/OQS
q7EQmZLFfeRlgup7WMO/VzTTPeGwiUDk4f5edJ/QlNr/cHzZYxjPF8YAP4fRhMQZ7SmfwjXthUfu
9HOAGAxX/OJIbrydjZ8ErFRmK0BLNIixGWb7ZhY5BWclMSip8uVzuYUz2DJQQQLqKl6foMaE4HaU
m4DgSxPV6JZZwcOYBLVveTy8iKy6M1Qeq8T8kfTHTO1HSlaS/rVE+k4FjCWDyNFYfyrio3qJdQQE
Uf/I2i6HjSdZc/uFzrYX4dq4m2xZtmr99kZDHrjNFrjfluK4wJN5XGoI72YFAHwAfveGWyuaDrkl
6xVJOpi+NlZtUyipeWrGDVn5Tua0VRUtvZ+M98DO1SP6AVnuyk/CRpXYOhJGDHle+tWuU591hqvq
pWjto07rzfLctvuVwAsEHAAw4JixJu8AKb8YW4U+r+AfpwNZ/Xr/jGG8WmO+KQIQOUvJW1s79VUA
3P91BMmUCRXqndFM9llQFcPVzZ6exYBO4+lUQA4IpHHexA/wkq3ap60p1MqyOxF/1SOkML4YiQPU
Gu9YaJelZIx5bTrqRVJ7j7EpQSLHRw+ko8ihep2Q8zaycF1YSIQ/FhmQaHSvwQbKtNFvYOvk9tpV
Iwq1aI46hf83XW4i54GPCnKGo4J/m8yyfzDjH/yLYZ5eJtCxLZPTN22pTVxJMSovuD6rD6hXIwlM
83K7xWBIGVRlI5Ide9rCejdjHv7vP+7acbeTPxX0MCu0x7pPRX5NxrFFAn3WE1lNHWHokNIp5WcV
IAp//+8ZGrZzOmPYv/RtZfeFrPdtQZNMcjcD9R/v+4Stfh1+3Wv43g//rJZZZLwM7QyZJLXdrZ6u
n0e42ZULem8eikd72V0SUYlkEYdYnkiULJMESYBzbjx0T8ozO6BgiXkH7cYqiyV1fJ9BPMl0G53T
sitLAwr3UOxNsqpIrOZDKqkVT6RFj+Ht6Gt7aXQEoISXHGs3ne+/WJLPHIJRmYyk58dWuvtvEoyS
+ES+IOm+Mwyl72Sf3qr3MlT/KuAa2gdTGNmGxLOpKGgPhNzMlHMFZe1mBX4a0lb3D3cYhz/UkCcp
Kz0FdQJQFjJ9bMgIKVyPA5rJ28RSgql1hIkd/NSpRTgvsLup2n9sj6LUK+4sNeIhfKWz+9y6Eb15
tTQPsM7I1HqNVTb9rjy0ABP3mbk0orhKGx+Ra4D1D/4dUNO2BTfVI9aQd9qtU3jSAfJnS4ZOJdaG
bHDkPLwGIY6CR94Ws7kIKQwEGWJQgvw8DoUhiKUjHhFpxTbWQxiocTBgT9CAlL5f2Lbw0huphdOq
db1Yi2JJ9ZRYSBeW5+U6+bg7+lCQ0un4VUtnxBkuQAGuWe369F7B0Oo6W7shl4gT9fd2WFPbUS8y
ct/1C50q4yWkkZAYK71TaB6KsHoBo2FCdZ9TRIWJy5DsasFslimLfTDb8/dj/qOJb/8OAFydvs13
/HdFMLp+JeQWvm64sxE3gAY/VTBhzEuZvo76AjLzqWU2sYx70lJ4Epb2mZwJKkbOt6SWvrR1Od8p
Nq1NDVmeNQ8apehb2pligABi8CAGgwMSOakmf+jLWtNm4YE1bn27vPSCRPIo3/oJG8DCOY3DfTSt
WcKJz6T4nqEetGdz5Wx6VJqrRP4quGbmc/bEKKK4B0P6UMZHAuMblW28YBFUtRjPN28hIrPbByY3
2FLJtoiWhwoQ86tSYFXRgDYsOHnI3fsQ9xmBGgEwW9u/epRpaCqum2SAqRlbTfMzvnursGF6QqHA
2CJN9YHLEspscJ4TVJcZfw4QNBguzbhT7wynFPwdjubjsBfsBvLBGBxT5RS++7EyGyhO7dAbmWRz
6+Kv1uetwdRiuWNXnUvHQnAQWmpxYrHAM2AIEozy8vZZdWSp2X22PhgnF7W2JaYF7QNSjS9G+MII
+nBaH9YicyhElgaZ6/eNy4Icio44H1Dp/I76cZLv8GAy8hU+pLSOC0zPVVCjz9djpwQcH/aKUHU0
Xbuu7uJw/e3Sd9usFm7o5lPo4q0pXvA4SMygRQCdesz+3ZlCY1dI3+yO225hpm10DXKZUOYWGAIn
ivIgsLASJDew2WByDDK1/dQcvGldYcLed7au3Zn1T9mBqPMxitRPOxjhHsjqWRHnymIiAJ5aicqO
A2QpHZ55CUZ3i1Mdrm/KNNDuwGKErXW8IeJHFkFUKDGiVcJPjepgC8QXePFF+Fey4fh1LngTLRa4
zBB9CTAaYKEXJZALnC/JPCnxowlpGcWlvSLb8tCTL+Sz9R+fm2WP/NBa8srdLIe8EccObS1Q60HB
hrqUNFy/oS8Ywi7NO/imQebx53nDSK2tovUpvTckAJJh55n23LoK85zlD96IiOFMCXT9Uj13u+Pi
Dn3nVmKQwjLsPzvTzCH6N9jf3TL6+34+yingETrI1kQbh8+3NCAH8yb3ehcHFTEFFK5+Amq1Kk+Q
n6+9f/UeKwmv21jdFNoNfEt5xty37gCZqdS6TORei8kh+QEgX4mGRHOr95Crnjo9kWG8Gz+gqtqK
PRusuQKYktJ5gT98RqiX3MGVyEJ3/GpdIvKbAiqzkQ+n7/nms3xCkFxnEGMI2WABAG4YEUGNFqtR
FIx91i5+0BfJw1gi9b6N1TyxIna/wt2XYHP0wmtYm8cpPF3nmcRyXL5mLh7qpl0Ln/QHN0su0b3m
8SqffXCm0LksVxzVLOFR5dihS8jONzKoLvdeXnTCDBONg8mh4TizzECXcC5Q38C2bqLReSaWvQFj
MZBeODZX93lSDgmY2PWtmvDVWBP3uYDqE4PTZkMynCLjHubvGRzFIFgo4oOvqP69fGNxfUx64sw2
vJ1w7DIlfKubL+j2fPkjlKntQdAuJj0UhctuKYAI1rtDBG64vqm3sy0LM2MgjRYWp2LRlmcuxlWP
+/aWGzqSX9PikT1KrC0CDo+TbqkAiuI0eS/tiQjMgJ+JUKp/wDN+5Y/dfKRGHIoH/yw2TuVvIxdd
E2Zryp/phkHiBgOeN4nnA+26cdgXdo7+1UvXjB5iX+z5XdORBmmo96Fd82+EQKeQf4AwNP62l/sU
JGn8Hlsap5KOO+Ut3Afh+w7RoXzOk3P/+3IgPNBKUMccgbduODKahzm0xey7FmDrXynWJhPGD6Fl
oCBo5ybNq0GnsQyWMb9W5rFYuDj52v165Y3PuAnapDvw0aP49E9RAqeV7IgEX8xWeL16v+z9QSCQ
53NB16lnDnghbCogw68PZ3We1y7XPanfuQB/va/cpY5nqMOP81EeD3CaqDtW8ojmpoP95QwhTSir
uQP+5b03Nxj/M/FxMsA6rw87oO+32nx5W4LwaGvnxQYqT1TbieXLEjfD1lokMUvriP51bYw1ObUl
bMXBWokxrGBp//Cs0/GddJFsi4m7lGO3fLxzJLGRAJT2HNaoCzAeocAGBVDB8abf/x6m/MXYlTK1
DHtBb9EnZxhJmE37to3SiO/PjfhCnK6PgjFtR3MqmvDhsjzhu3Egme1U8MudKfX5kZusopjEIERm
S1xmuqp/7QUknTLQj1GvJL+lzBpDgRCwulmQA5c2fOq3i53291bWBy8p+G3ukjOWWS0CpF5JXLWx
UnaPGBIGDa2L59MDZR2XJUBjYkdUlld+Bpo14t4bY4KUrm59UwHW4R7HxATJizC8CyJ7BleW1yvX
JsCiaQILOryORfIa9nyESS+paMD4XEXl4FmZ8/CGLpLM9Y2dBv7IKIiFVcBTPK6mIsV3kv4STFyC
/lrdtPalWpifNxDZtqfFZMAYOcKa2J5iFwFPY1JWC+IfpNjlbXXAKGeDNoc25cNWxxC0X0Z7is0R
4nWedqaKlB8QWzHgA5piH2MBQ977yl0YMHiCbZlKcCMjUAQ0WaRl0KLPs34KdN+CmOMuCu9EheQS
Iu5tI8YXO+oSqACoVkifojbte2RLP1hD9jkrEw13zVat4c12PCv5RQjFwCbnGS+UHmmSLsJqFc6H
rZC6kdrRGiYNXKcmkaXP/gh9boqMYiwQmJbqAGhPV0/UwHoVXGq17awRK47YoHCXZFUJFT+3Lq2p
U71hT28CSa/6gbPjfPm3PobWubiVZxq304NWzTS64bkDXs2Fq5hnSBc2aGtaybL9G9tCc9X0sqOm
5+3Z0Ru9emEs9lxOZDx0bWbLHgRcJ2HVJJbQmm18HORxrXyY2agNYsKNoIqxCTjP93NzLceK8H0h
pR9z4EbIlXvzxJvYNP3eGjSiVd34jr0FllSjtNCvQimnncD6JWy2kjSuyQXydOjDS7CNv+9g13kB
hT/ZHWETo9sbr/N5WznXTGCPVVeZAmwuV0UgavInBrloZ/Cw30BDUjYyj21Y/JQbsLHADitYt1JU
QLIdzzypzCqCBotdPZLtmK4BuYCUu3s3C2EK4UDq3KVCWX3fq7VQitYfbXYsA1nNPo9YGWCx3Or/
jQF4CxG/A4ZH8/EoCMeLNZr3v9NtC2vBb4WA2YJjj6zPx90XhFLl+0pXtFtzF/b2AFgToJlYGnvW
g2b5kqRMUHPgnHHiVKyJ8AgIQxk7FB2ejo3WW/l8HBhLQHsjYizcbwaagFqJBlBOelEZP2B2Sa4z
D6/BBwnUijzxJFfUsie5lpfy+bj1A2siftyFwd1vdESZLR19oLm9hEHG/cPnDKrAR/LCfuJN2OAu
ARTJJ5vuei77qGb7ShSM4Yez0JFsuC6iSqJ4cN8kgTvdxppO94uNtQFGCGDKTVuB3+hokcIA7XFl
ZTXe2SaB7hbo24azkqlMJ8Gb4yAxNo2QTAqTtgEfYdhfguznQyKcS/3R+5oAwu6mbdzn3hucFOOe
4SOgEJeGIO2BiikRDQkX0hFRLbDTGegGUezLanG7ILpNWxubNl73UTaf82Yo1ZDBlA9/sksBVZlx
yYJ4Eo5wpYatVMuAVPcUN+clwDYdwNyU+AiW87Ya4H/0uiqCR8qPz555rqT1dbpgoARGF1l0lGkC
7Ip7puoIKy415EiBLkO3boGr4ZZXr7ZbgDIsQaQ0/54ydxyzmIm/0+wDR/xMrVuaIXM3Vblpmys+
mrX26BkZBdOBzaZV8ZPpLJIprjVeg0l77xREiWPTZkAWPUkFZKGSGsChSVFZVUV8RBe6MfVKcDGA
6AaC1DP/zvQot9/zJkoJ/Ohyh5LxvRZ0enbm03s8sj+Y1/TVcuS18gATrbX793X2KSpCDPdg68Jr
uYYskHQKUzt+qWDvShY7/vfPoZqcGec1ReMi3jcTT8qccO2WtGeFvH7az/Y9n5ILHSkjr7jFLWw5
PyHtpbVdjYR8VR8m/1KonOnZ/ws51OPPN544f6+y/lmwjqYlvFmf34gB2JoZxO21EJqCCVPj5CYK
wUsbYqtDuQWzYqxXd4G1Fcb8s/FWyqN5BsYCe6Hfbbbe/hQSo/m65ynAjqgi0MxPvP+xA2DHT4SO
nCvtjnJ8+dHrOIUDFnjdO1Q9/pSFNyMewhpADeF+Aq8MlMqIlYhuKuSwOfjIQlBFwik7OpRjZp4e
gUAMOew0i0IL5dwJlG+pbi4Hi5ndUt96RKTHkmuHNWh7amtZa1X08H5UjTRXZ3GSYgDNARiuCv7g
/4N298xBYnI4AxzH75VQywhd3xb3PjQR2DfK6J8dSN8h1Pq6HSNg5ir+xKEUFlc6HO/6PL9kGMXF
rb2twbkcXnyOG1azghArgX3eS5eO1AtGxmG/B2LFpJU1+Oa4mQa/fmLe9ENTCQFMxmpwX/w2ES+t
sBBfSMaGvCx2qGW4s11Xz13eDid4q42RJv6V6nM7BPB3Up575BtOCZ5gDWmX9NIE2xujS/yUj4rI
LT2gfJdc5soeAukl+hz1kACUIQS6MqvK8+iArvgsCaC6FIp38ZfOZFI2RNhCNLJzfWKR0e7eQV1A
yr0VlfsRzohng3LL6SOf8u6XWr+9GfqIWHkcRBGEYJtBxciS2mmJkHQojwAK9k5K33Psz54Jtr6T
3tqfuIM3YVr/9Y3mlEMh4qmmjwxuy0ztpT7v3R6pTrDMW2I2P+vYOQY8Z/48fiDJ+llCnNUMRojE
aIJaWHOEgWiV69u9HQvi78PAJ3dpZMGoFqptb5M3Ur3CWTGD6FAIo9YodS/nwGNYzmf7eirsZZjQ
90iWToNjYKs7wZ093Pfa6sk2XMCH463h4LnqbNw3e/GvAsZ3wykyrOejMh2yl1Drdz+E/Cpn74H3
SkwPoXvd6VGNjnxpj/g3j9FrjJv2vX8xqM7exp0Fb3ZgVwSL7YyTrQPexwfvWpW2yJMNs8v0VRXw
RSfTfgmi6M8KJgJmARXnAFOZeLg3Rp6aAaQJT7Iop9dOTP9Djc+jhi94JqUc+Kd5PYChkSQ6IqFj
PLum4snRvE8v1A/i5D6V2ZFyApRAehX2MWMdHhXlQWMBVAU0FgoGaxM/nB+RnQmSHdqQBp0ljn1o
JlfbBr76m1CTmnPN8p7NtU1fwCBjDPN7dAmtU/rQ3BdHmY75bxNK97A2p1g0B2VwES2dpMMHsFYZ
10PljSp1+6Y06yroW4FpGVkvIh3lDV2wM3s9AVXFCHt9k4/BjMJxXwvw6g6ZX+xq7TRU5ucKD12c
xT0xkIGSj2YDjShmpjWBEfmt/L278yNe08dbcspDRfB+stxzvdkUnNzXpsF2Ae7qoVP9m4duyyOU
oQgM9TkoZ2ur5InkmWNS4dvsxZQFPWUbhn08sLqM+hpEb/DUhp2R8+33kHEEBtfXCLz25YaEv+ba
jFhZ/y68UCnLNanLs0FR2nMdEN8dW3Cn5XhCy04k7LaQDOr0tAhbEvY427MIKDmvFNbcZAobMR2R
MrB9oxt4NlWjOa1I1qXeqDA1uvw2tByFKh3BP/iR2QeYr5KAEEjfilHJG0OR0zWoYq0R4xk2gftI
CazgVVDtZV1fvf0cx0wBxCI+Y14J/+Dmr4EeV6squ7gJtx1GkDdaeyqvDkvg8TotJTzMMWZrRK+I
UM3St6qX/PoudlorCXrROdx09JR7xZwJJgeTq84xQzWTweGZd0v1TEJDRgEByrdc/ncv/LOAPqvj
BL8SpgJXclSYA1XoscJw2RvlmMWIidU/sIg/FAU490AAtT9W4g+Wv8RUsxSPAkEF4iyeabzBQXC8
IjkMaFN3fFnalOEyOZRWPPObfnKnLbtDsAZVpsn/ZktV12IMv+MsUxUa+5AFfWAPPWypPKotvRgH
Tkx1YvxrEJmViPqvqyTp7Ydydj1OkuvaU4YP8ayvBtVJobgEdSFvNfmfqOerrHgSnx4ZGSVO1hPP
YpFSZMvjYjKpOyaIZ8LRUziu6Y6zBP6CpFgdmws4IC3PbzYPRvomOSuiQG60fiHrJUK3Ix1iZJd4
lKfToc6ePxDpeFK2mBDtc5L7pt7KWwvEgI2ebREO6PMeXhrvPKHba1SwMD50Pssw6dHwPF+Uoacx
gUfREYeT96TlhCU/P1i3Hy0LzEMp9kw8EMRcl2vaSpqz8C1vHDIxMQeVEUvB4Q/G5BqjJe73acVs
Nwisa3JDuwNHKt+nTcWZ96spbzKJdHXL+tTneR7GAWz/w7ozsyET9ymS5GTcll6JpDYO+y8yUoSQ
fVrtA9fK/HN5vWLaO3T3EXS36jtOXDQou80y2fXJair2JpTjlp+ZzPth5QrrepHhvnL2eXBQwEZD
uLiUt14MbqLWaVyxVPS8oC6HzJGaq5vgkeF2B77YC0ClIidaGedcRddeYKnCYKdQwwwHep/C81XQ
TYxyKPY8n0cfq/znQ2DMVEimA1dq0gj1O/buAqhFKL26VZs5w9GD0/euIxacByGZ6YAp17O1vY/a
3tadpq4ComBZD7e6wnxBIR5YN0bscYcfapjWDJFDwN8VMZ2o8rMjRUlDg6Gwc+o5/gghsjK7fTcj
90t15vrZXg+/WU6JKIdq+ydB3kFOyIgOfL/icC4JeYWe8l1n+s7dnBDvc+nrENmo7oQidR3fQt2R
Gti4a6C15dtRDKgoEE9MTRRjCpHU6TGeuPHoKJFggJatZXN9PnZ3bHMQm/A329ZEPkdy/DX3QxBz
Y8p6gB+E3hQ86hqqwFtt55qdvCmc5/mGAERH3z+gQroeCpO3Sx6RnPAjWP2j8Qx7b1iOTlADQw6R
nLqSCyznZpzxqg81ZUXIwUqvlEyG1w984bmKgDh+vXD5nYus7AhBL2ts4d5WOzbtOveO3fgqeM7s
STye6pZedS5o4NksYwOe2jQdioPum6Ekhfd+4QVhu2YIywje1ccNbQaW4hTkvQrlZGjs/AvSR0bo
1FHxwswpa5tCuY6eVuCgs+Nl39adK5E8VDhvn6G37rHwjzZgIdbWvr4UfJ3u6xkjtMmldEdFhjuR
HfD9q+ZriYdAlMkDrlTnJjG1yWnRzx92QFrWPVtSR09Yqd14w14UvYtPCdQdQRRPLxyNHTW3URi4
sZ8yEWuAR8By8E9IOhamy0AgQl3M4l0NuLHbiMiFsNZuEUxGn5QYp4OSd3U8s1YWAFx3qOfIrgrr
UoCEISs1KE3Ple/7YQyftN0rXPXmnKEfi/mAA3csVVSECYIqpZNWeTB2JWKEx3rIgqndwAwOfSQV
e12Bpm2cW6UjOqtjePPIwLpD3PH2VYFnha+TrmdZjkjeRfGT/sZoem3hHAcc5Ok7vZY/Uu6FE4Cs
GWnaMt1JweyF4GwOLtKX4Bk7/TuQOMKYXMoKfUltnKR4zoh+W5m1jdZrAdPXfWWQ56Chh/2C+IE1
GSyKSAk1pr0J/PwGt2cTNJqjExyPjc509vQMqur4PR4X4J8dBTUlt9+KMvC95+1aynKqFfnctFHN
xG8iPML1ayUh52fD7duk4ZqidIPFTREPyrF7XjI4jz55F7Tp1MLNlRfLONc6UlGxwiG/cZVZc1k5
gT/n64rt/fZ3auUwKkx1i9mDrkk61krkbdT3oiZzoS4L65R3+jh0Xqdx604sVCsdd5zZhtHLDMMo
RIwN4uzsv99HEHr3oaFdITLcfeUePMwQAu8LEeBnLQsvPBPl5YkNR12tT/e6Ay08nSQZuxpnZ341
8maFbAa/8A16VNNVEanoIQMh33fs8VZm3ytAlM2twLK+xaHirGnbxQOn3+cYHsQ2S8R/9GbP7Yf/
VNkkjQ90rLlhY0xjmTIFGeyg+vrQOR51pBG1mcbqaJH3LM/4uERmYcfInaAEzCzy1l5l5KNbb+Fv
x0v2me5j9q+ftGv/znJ/UOscPFQAMAg5HVhuW0mHYvYFsmRX/Z7n7z3aLhoJOVYVA/ldW5zYXKSh
F2Q1QBcz6E/R20OPs/df2X0B1oX9vQYkuZZVZDWeu6PCW0wBObjadkR/JE01iu0fQDchxfpUGR8o
QyU9tVcR7KLk/8BjM+JM2wKsWW2R4O3h6uWkB/PJDh+vGGpyJxCHWt9JdR161Xv88F/HlwvFTkA7
Z4RvluSA1xzdobHb8bJxUjKm5Hz1nrTAeJpuktENBGSOe0p+MeNqW2b+qDA+P5nOq/U2f5+TPNIa
VgoCax1HudDb05ffw17MfmnmUuETGpSfFfV3xorghAjYF+934dA7KDqLkUQgiaZGGOya3DG2cD+m
QUhvzT7cnGkB6r259ozQUUImC6YUZW6e/DvrG4NqQdwLD4q9SCZqcRBaemSMvs9Kqgo54Xz2ZjVp
okCteOYPB/EPvItHPxQ8lGr22gAG8lWVdTCLOsvGXVCMLHp7k+BtdRkEttw3NWboI+4BfTnRP1AJ
qUbdk9LdYobFVSGZFRf+ydwWXk6LY7Cwc0e4N1CIxpjAx2hW39AC5/mm8R0KYAAIRXeelMTUvelr
6cbeKX1NR4AwvHYTVyap5viRGMk+SG0CfxBwayjJeb357HrzHd31SyQyOPF8C4e79yM5iqtP4D+C
ubTVUXJKPDuwQDnEFzD57LrYYzjD2iiNjyeAv7r8dF2drzUiM4xmEzCEgkKzVi+RfmqsHtePONln
ogj2lSSSXro3jytiYHcOsdalPWxlDIbKoYzVOstzCwAtm5chCVOizcyLITv4by75hQNllG7w2Ugh
boOZLmKVVVboj96Jl/QEybrdqLzVUOyVkZLcpCtHilnLxhXcdxXVRANN7ULn/UH/f8lDgf5YH3N9
CTQfYW1Y4n47UMS0x62zKRi3/aPwL5AcKlSoGgiy/unFusJkO5E2b/jucnySLSH4Fycvz5JYna8E
1ZFsP7iZ7VPilyqc9RRjGbjqy6wK6xpV1g86xFWYoJiPRYwZNZHaUFDzHaUmmFqr/wGKiWhtcHTz
yBHG6CQBSMza+HRModlDR/1AlVcltVc4oiDRUwiCbKGrkOR9WfjLWqIHGOcggiJwugk6hj2P9cUE
jg/3pxw9Jfso9tv2YTKeZW0gT11N+rtQ38/kmsta/N/BevrdWo3/EKnCXlK1Zy8wpTu+cJnFG2ie
tp86zLbbosa+VF2sGgbytYDD/8LAladg/CJn0rC79ZsyPUMq65M9OYP80uIH/rAkQvJbu9mxZZ3T
870cCFLbcYE1V9khprJokz4ZYz3QUUwXi0UukgfL+mu/qK4JqgLJdpN35N++7fbaXWWmnpSnDZH6
DI55rSgPmCEs7tCB3SFlicl7XhD5EkHEi9//ugiu9Wl28vGdGpJH4E3HOkCIsteL7NzBIkrpfPp9
2r+iwzcIG1+WaxndoOxipu/1p6BedsRFwyxlN445wV16aTrHdER5Cwg3VFM0pl+M+iDc4J94xCyK
OIjxXbTk5lhTbGY1nJP7xlzg8TU5coLR7/WapByFBFGa94V8kguKV0hO5O+bSZeEtUB2Ys64Snw3
Ai7Ih2un6+ptSpaUbYgTbA/hGjYCzg9cacD/dC0GRzgMtLOchPRdSqiaWYaczNKppcagaB3lw3bO
j5fZlt45WzJX0RzXATEKr9q5XtgEB3vKQbFhaBXjupWx8skCuTcZ4fiBQTdnnVMhJFt6sfBE8l48
2maz3O/GO0fjG9JoLYoWcXCYZIA+VwkXi2ORoC5VEvSExI5pMJtCm0YUBp+3bmikeh9oZN/tydNa
We18Kz+r+PhcGzJYRRIuJFH0donWtualscv3Vkg/ywBX+8CZyLcXNzt5gCuFTXB4NQ4K4fiVK8D9
Pl6eTwPDed5CkeTOTGnQu7qn6tDETQQ5nIUTHHiIxWxBdrfQ5o1+nQHle1Um3CKvjDl0IcDrbpid
R1k2gjPj36Z/iB/qd4GUS4ADa3uJvEE/trf4M5AiQDXiE+LbaUDll051HVuj724YchU7kBoOJq1N
OQ+Ve1xGZeI4/bkqY7+RkJoxmFs25LTViOTwO6UW5g6z8uYXcXli/PeSsLWDo8nzP1jIl15eaEzQ
zB6Q+1XQX8f1KwzWJhOh44rxVj+Cyghmpdac4VkTHGPjayJPQoGlGCG/W8K/TOeaT993nAdCUVkd
22m91MwGXoKZBwZvouQ+Bb1yJZz+B5koU5W3Cn8z2tffcBDWgjCURXxrhbZkrkrWjZgRfdGqTVSB
rg8MZlOTbTOtD7c8h1XgyeO2DrjLRzzXhhYkIcOQYorL4dtTRHe5f0uObf2ul+dGclQg7qilB3bT
slWl1ZJ52Ww8sc0iMF+ls8rZ6ibBz4NHwsCWkMFz+Vrbg8lAcyNszz1rGqvQj2JmsG8vAVnkmqG4
Kx97tpPQ3m1difvJU0dvzE0bVnRdnx2oMy1zFBmTA7AjQB2WJ0Lysu80nrVUTAb4Dcs9QyuzODVz
XMCbZGBLnILFc3Gx8I75vM3Y3QxqZz0jDF/cRR/zNXkPD/XZr4BWxQdBF5sv9tYZXQ7r830gPG+J
Ho2gC/zRdDi7rUF2T4lYzGSbf1gyy+XQtP1Fim1bPJSK0UTHNzj3Pbe/Jft0xyIPpcVVYPMwrE6f
V8whoJRW3zBuPB3prJIzbSibwL2lfND88ja85GiWOWk0b/CTP2GJWLBkvLM18sHbFq2tEtB2sRXM
yv02uy921SyZQG14hi72UYh9D3HYxyo7fVfujcE5bExu0+mi6gb1D4e1eOJMQZgnjsFCIIjcx5mJ
9im7iAU2zR4E0GFQkxjk++fR91bnOu+42yORSZ9C3clL04xnwFgZmbOZ0qtmOnjeR5wEPS9M5Xz+
cciAgOHifzgoKpkoxpJ58MbvuH/Vvvx9Zzm6bAtkLBdde2T1ccqEoDdRfzJSij4hats7Zo/0LoOj
mhjzYtpZ8SkUdxlcGB/MxflKIfFtvSi05+m8jttKGtco3aSTLGkJ4f0h7BGPcRX1YXnc3xU/H3uG
8qM8XPZNPLD3y79VuPdukmRo/uGx1INXC3QDo1DgowYXoST667HXcg5sGHgFQ/8ul5LMJ66vH1xS
Gom23yWT0Fy5NFRL+1AIKhHZ9dl+TXZrbs8CGJgJiJlIwxLnezk+4r9pT6fJo0H/yyG+uVFMCVaR
KBTa4o2guEUYbJiJ7uz5R3trFpBETc2bLy3f3Acr/Z9O524Q54yvu8JGmulBi6sQUV0Ibavc4wpb
CF3FGTnf8QGD6MCCXXfVW5o4bSsuYFBBANwm19uGf2MKfOW+DPkq1+10TLFi9VUkfWl6xJ824S/v
d+mo4rs5oHBq+YjCvk1W+u+P7lDFjQVZU1dhEWkI2FLwHMQOeacGvaopuhHTGPhHxESz1U/GXUCp
HT2EDmZJa6nhmaSqIdaq+GVZUkowF6Xlo9gk0F9+UMspFlhTKlSYwBKcudjR4JvYNvbWbNFA7TCm
bqW1i2aT1ytxQLFyGUMbrmV0JLXEXJb/SeKHcD7QOf3Zj56fwLsxibPaoOgFWgP3zitmdv5WWAqc
uLkCtBkkTgOtFrzBxRFjRm733O8w5wyadV7V/b9b92pcB21qK79J4/P/sUuGFe5Xq4kGccH9aS9I
hMF7mkRRB0TzOWdMy3bOtDNZP8x5Kw1p2GzHL1T32fRwd6k/BU3A02xzafJhd3e10AKReIYwXAfQ
ohyoifKHJXiehQDw3id/rtQwapBxIIakSvjQBSFWOjYObaUPt+aYbsS70Sq8BeoMYk/AEAS/E1bQ
qKNWJp1x/LlyqJYIekOgqjKAb7YsGw5P7oyO5sHG9oEr9z6MrS2N8trDYxN+41/lfd+uu0J1jMBb
T9cZ2jntyrumizd84j4VgOtNbJT60J3QJcIAdREvvYnpsmsfTtmh0zvh2XKqPmmisOKUVGa5oYBJ
TS5hFokErXg9tdP8G0XiItD1CRkVR8d1Qb/AfA0vXeT+cfDRRV+TqKewwENMa6sYSTIWqn+wY8i2
JIuRzdhjvJ5G9nLA4ptyIEI+14Sg6suIi+sRDliYY2NHcOaQBXyHBeYvHtN8JY73Fot7sYtjk2Zq
u7EIIsrvrQZeD5abXYd+lJ3/7fLCnXbLfn78oWGPwr73ItcPvrmYMAjkOsRIu5UvOuVaMYbVEkjp
MOxrSa6VLghtlPSyjUKrtf6VKp2lgEmYEQdvHIHwo0E/9t9w5zMg9nkQR62sfKnUnbY8lxVE8yjm
nBgVsEQV3UKVT4wAHzdgJVvVFnLNXe42ffNt3h9qg2zLY1DCH0LkOXGN0yT4GVTg9rjf5lRDXIIl
juH2hjLChrr4QX83tSQBVvGXzFnSpY1jbQlzd3qxo1x7tqsntoL4SoSm2183TdDRv410MvH5wLQO
iU7fY6bW3A9Y1a3fZRGmSlq+1O6Ut2mubF94MV1yZuOs1MZqlEBG4keIFzLVR8j3yEFqPhd+eQbC
+tCLISbpMMeuX2tyRPBQanBj31pfe/s/xuYJjknuIleoIHGKoQrVo1UvrUXKjxlnI9+W5B4bq5nY
7pQ/sju57xrs3w/PvAZ2jYERQT6hl3ouUNkKXZLk+bvvt0yzx+1ySLnho2ZG9nMmQFgPgNakz7Yc
iXioawaM4FXAGqfuN2L/E6Gac38V6YaaWR7QgQGfLpXBNQVNU62fHgGE7w8FqczhoX9cNiWwho8p
8UWruAhKxWjnYr6FDebcH03qthoXS38tznWoMBTvnmbneHEzg4Saggt14HtEnEiSokzEGBfk0k9Q
o8Uw1cqOVVABcl+XAm8vPS307/+robIN1G6rpmWoqUhNNCcErmkz5W0FMWLzx7idO/EH0W1Inzld
KbE51gZE+lDBwK+isu3fxFXYASLl0cNe8IuYIiqdh1ZbR1nwf15GuIgtbf7BFebl79Tp4EdMiyII
9GJlCQtoXRBy9bVIqYHwdZeZ3IMk2fiHDkyxTcXokwvu7Xq/WnFcK9CODmjazbRI1rNY2RVuhRpL
1pDWWu5HhWKrBOlR1uXx7Ds06AO+jaHUIUObpJgOK6GKMw8U+Cv7Jx0Ds5yZDZDO1RCL1cA/iVoX
sjC81evGDec9WXtV6uhvoR/oPM9ethgjRjNDKvTbLAw/8eNZt0p24O9ZHp0aWDXe7URbmhfdJWA4
GB/jcihlkM5+ShNPaUCa+wQIx1bugR+eluKoywIjUYueq/fmCGgjgjFqcyHN7SZvN4uZrcf4c2ff
Jkq1kkijjuAU/JEfIAc/K8lguGn3trPMnAadiCoga10rHAKLnHjBqaSnmiBkNLi4V6uTmjM+a0zL
Sd+UQev0+bJMM8BhtfQ1c0Cdmgp75Kpr+7gT2H5BaOJSQeGIF43W8lnrMlges60PZwYdC23/iBI6
mmULz2kRkdzLP1iIrrqr615jWPUFPz0DQkTaG96tbGJMFUKnqLP5PlRst3Fpf3v8SdVFZkG94mLf
wUdo0CNRz8kHlh3PD9Oj26KUNklNOyFOvlmmnsXwOZhIPVAA9SqehtK+mJ0ak/Ibugr/tc3LZUtD
nr2kUGzXennqwe1rqnYNd8VcABYw2u58AstfSEz5S0mPGLU45/vXBJa8DqOAgiFOvDmh+s0tpZ0t
6XMDnosDZ1T+TMpIp4i8XBuqYZvUvo8PqaSO5qgbhEcEUHDEB9Rgc33yNeknTHa/nXgacWIk9FJ3
HS9R//uVHOqLjRPCkroexDweASFjDubLX4jU7bDSyRQ+iFMCX5q8oIn2sM+4Iucb7TKasmHKsDNQ
ndHRC9GCfPrVWZBai9M3kPRubTBO33HGZ2235UC5H2eekYbIOYAbkU+idvqkuJjAzrbD90o6Gun6
JbPw/wKLjecGiJdXfHo0PIF4UnDf7Y5NmYe0HykPEhdhhtv/8eofA/SJx7klTXSPjqNwFHdG+rLb
g8m0zw/qorNgx3Ra+YcxMuTwlluIeyx1W4PB9plGOQMKyXRKLRe9eGp4e9csIyJ71/n3NrggD4yi
baCnQNhbJ+UE9k/RKDojv4gjMKcRirb+Y6O4HJez6ioSUfYVGLjnw4rE/9mYOtOmSbyaWTFuh/L3
vur2TP8nsAeLwbHul+gkLyWctUGr/XNiFOUfQGwdz1uUZ0VOpjOrsM4zI9wp0dXaR6j2neU0d323
NSvtKrVQHlylROWFCi8wGpzkKgGQzkQot2tk18L/51oGN+lY2XSXU8fymlV1PJHqw0tCDSkDHOU8
wrKuvoDGWoO5g1OjOrez1YFxsKDyVlh72qC3etnFfMrVS1nTvhUyllPNF1YD9TOHSo6rcDJWfgqA
iggU2iNOlupqKKIbNiU0198+/8Loux5APT9nqPgV9T4BNLunQAnh9+KI0ylnfgQLZZpE3TvdOswr
8biAK1hcGe7fXSy015pTEuMP/oFdZCfcFcQvUs/5ALiRtjUnn32DaQNrLLfTLiS7HDSsmpQPKHDf
nHTL3tGhRmI20PSuDPTVpq5vWws9PEgSGnSiZXgFDPyaKlQK3kP+iSJ13OGm659vH2n6dMI20B6b
FHmxZgF1PCJSC08DvhwnUskh1E59K98miWLTZSiec+/84Pf73x+E1Yv6OtQGJ9tNw0wWLScLPqLm
fKyLBCuw4sCL5wMLU5GDkbu9tX3YmP23ort/3a2g7TtZrWjgQuwdLjXnTLK/qtokTImb77j5OV6z
Ihbccq3vTBYFsMa8iG2iiIUNqG80nxM7QajzD9QJVujbAWrGOg4lI2W5VBo0Gx1SQVcDjuAcxVED
Umaq+74BDOy4wSpbNKdOYYjPgTKAD30CAIcb+tVbSzZj2pOA5d1UYEKtwJxhwXkRdjhJsnFJ0Z2V
jtTFJWm/xXIcXFQbJhDo83rmZUkybdNoLmlgsoaDFA2QdI3gt6Ri2B8JJcr3WduIkM4YXoYtd0FQ
+8V+Zw3i4Gw8DL9lNZpgldKhg4Lji12jNau9BJ/dTXVCBbqd03ipbJQKBYjYfj5njpI6wQbRQYV9
y9o8bnkvXWpvhlxW+/Y0jHDJ4H6lRjL2hFYYjCjXlzGwv5ETKGnZzQYx5h7zwxTpj0GFIHjJFXgm
LtN+YP9I37GRBdYQTEH8w64KCzydZD0z1F1i5WznjpbpyoCNt2+eAiDomTamNoOoaEB95xrmgHj6
nHu/9flvKiQW1a7blOTARMq0aRqrrBv4KTitY32PeyLTGU4HAQBBTh05Hmz8I2leLiNyjWvjPTtq
sn3SEpzy09CPGOmOsc7Z3hTw0C5r8yK3O3xi8kDhROj/MfFU1Fno+f7pzyJLY0UnEp9rqAS1BP0q
1gOiNWvmvypgRrD2hnCr2Kb3K/So2HFH0M6h+PkjhEe6NAebyjL9aQ+hJ3aojz81ugxRVlx9s2xu
5n6tkV8RZS08oH3YfWs1sR2WKlOo9o11Anwa6ZA6zJl36QdlXzh9kE4qWnTWAZmUcdSUPL30APUN
lJtUw06jSSjdxUFJ0qVpkdV/utPGw9p9pW9kJzAiH3kNJh8u6kUQ3TQYj/hQSxRkhZuSse46jzKj
WLm17z35Jr50Ol7ZUaFOk++CmTg136xN8z6RMdEKrMzPQm3D8uLGNmPMkQEzwobjPLVzZk0Q9n7Z
MLohw4lu3QQHW1MIBeFhlwuE7citA5kbaCOvJAxhTizEJlJp07OBCF3nHMRt6jpA40bxpEm4GAdw
f2kOEHKyVdv2n41tEb6Vzb/oywkRyKiaLe4uzacgj1W/EaHqI2GyVCYGQrc7UVsBWCTPUpLDyrRD
XoTi+H/ZcQeMiJRzRU2l/hk+2iNmkSjqMKKwFetbt8WFLluUMccNy5E7qG9dPKId+NTbjISAN6UZ
absO1ri1+tUuPJEbyNxddjLpcnGnRzDpapoPuOfYQc34dXmUDSKMeuewj0Lo7HqRfAxdYJHN4WrM
hEUcPF59HJVK9n6PgUu/3MikcqgX5MWW2Jm0gpmLgTfiO9wc5/VsqOQeEu4yjJSHbPRt+J8VXhzJ
ZKY/C1iBpMsZllk+Jyf0FH/KDXz0dkg7p68lvWGEaAAZXH2asMtxq79kkRlCE9ihsRH913cU5KuX
V8W/voxiIZd4foLI2DHEdY1J2X+hwRolO7LATZsft+LCRaHdXVOBiTw6kuAPTdTkhyEfwHkLHM75
HR/gOZTJIcuQtFvlxpUJ3jeK1ipJCKBwTt8Yw7c6ggruM71dJJQfvlou7zvi/0qiGPLtbIDw7qLk
hC+3AWawxKPfcx8XeK9IAiyKvous0NUYB5b71wEOxtLW0cBBZPxslrXYAfg05CbnHA7vWtzRI9mC
8WL5/gr5qOJiFOmn/gaLsSKo4ewy1dohzD7LrubZzNCK59pXlMC/SZK/+DW8iieQr3mftxgtC1Vh
d6YiKMUofIf6YFXuHb2W0hNrbmsxK0G4p/geF94VqPU+rRahSBGtt0e4VHZwkkiUoGZf9/YMHpR/
c8KG0Is9RZyEOeivR+ZeF4E/jvbqciHdIB7JGfUl2SGZxHpNcaTNEwcLy4fmccYLM8oW3eb3KDvT
InYtyroB39MBY2I6PWpf478v1sZtHhiY4mU5OGGQHDTKYSyFFnhOOqQMTkQrOKEZfAp/XoYEV479
5oHS4rcA5Y1w0g3OJqfkMh/tQzO+69vYvUWObeQR96u5F8tdi0/ctSJezEjMqjKJsX9aw4N+tkN5
FrhXG3EZI735KbKJWvj+h6HPpq5APcLUQJj2InwO4iWVB+cKw9AWpgao97l0Nd6sNcg0Kf8r6I2Q
Ng2XNwYi8DP17djaNMSTaZKn257/KjytJkqF1VrDksNfXYgB5TN0OG8xw82CDg5TyeHmUZ/9SRxJ
tT48pFEsX43YSo4oNJc5Rrfq+iJWrG4YcjNPJ6fy3UuzLpeb1x1dHDhg/ZsD6RDEr6mT7sKeg0qO
oAqPxesEn3NLZEvEpYEDMadu/12guxWEHkCTbNk1rJ9mMY58GT+HGsdclX1oh73ivWqX/32hApo1
KNBcj/v3WfrQCzxJ9ZOBiud6ylVdByFSyKcxy6YZST88/j/e4L//pRd9mRI4dVIX8h7ilMuwaJK6
NVyY+i7XcCKre9MjbCLKQbVUKdPyJKxuULVcp7+kKY9PGcaTv40F8zCqwbPPv4jxanlkh376bzvc
5IqKUjmXf1sNWdlkswwkL2IDA5DtT/CEOzhMMFecUho5FhWmL5mPAbIQ87p9Uji0ZXzr4YpDqZeI
mUYtQlNkDefx8ZXaE//wJNM7uibj17yYqrOHuGgWlqz5UAIoT+XjgyWNc8RhFPAtly8w1AWdlOej
gx6ObsYhWf4JHFY7eSTcIMMuUnv6iqqNVHRThrtoaQ86t/KzK7kgaTw9xhxbM0JMUvefAG35EoDY
e728B8ySZfG+EBHrT2CJvzErf1FjePfbEo6e+B91o386fn48RjGpLVy+RhqE5mJtf/iYbKE9LjYp
3HxbWKFVpYmtDgovVjQs032WSd1pPFg2wfRFVBT4STyPgh8ObFtuVdUa1th+dG9eJXS1onWBUf+R
FqpwZAUpu0UxFLZ32lcXJaFXiUctsYQE+HHYA7rSwCtgU5fH2RMJOuFjAaFYHGGsSlJRDpD23F4t
1b89V456M63XUxIFJkSQMnSswG89UjbUJ9TpHqHqf1p8Vf7ZQQf79q8oqFHm6uTt+ZlqfryuQqXN
6zn2pFk8Zz94Rw6JkEi1siUZ13oeSjKxsJaI7oZRWJ0ZbQHV4cnMhGGwoTL7G5CxZqmPXTDjIzhU
Sw9dn4JC1Wg/5u36uDbAzO4dy+XiM7OJCqIhJFn6v/Ed+Fkyz8j1+lvGZhdebxiH1wkABrIuWXCX
jv62fQSE6tcQuNIkYJbEu6dFFdR8K8L3iZqvpZx8b/8Cq8+Jh1ASviGz7e8yD+/x4pEXjGiHKktU
FuLxvUV+pSJYSU7vXIy52c9UkiBulBReWcYGz5M/Arfx5V1qoH6eUUHINZ0aQMtUQ0/Kn3rjEbyi
rEgcTHgv82NgMpJgpdgCt/woVtrjcNhJjGq32R1A3l//VXLMENpGuybCh2iD3oGYFpMK7PogcduR
Luh3aVNmdjJmdNmjZtKyonAP+Ahb/Umqh9s8xzKIDqVSJTWDO0jRPwqq39Kr+NrO5rhqQUkd81Gr
IB9V8gEJABKQzr1fgNGPxiqgFPb01rBF8ufqbssUOXmFXq0X0LBWo3+CvBijsGpFmA49mlLo+xt9
EMcqsPtOpEUPTwJ5Z5wDuZtYIs9P59sLrF3SQvA0rbCUFrelAiTVBmwn4KallwoKDQe+n4ysuZ+2
siMMdlUHItkC25/HyylGQnK3a+rO/IPp+IPt+miW/T6CAcNzwN3RsovM2sxIyuVN24qyhteVXala
bw7MPhCIPeKoWs5+XbkCDFFJW6EaUqXMdWrSVWb5ACjnlzW65lKCAL5LJ3zws0vwNlhR5rrj5dPj
0/V9YlTk59a80hKQNm7ipC7nZD1MJy+xXvNVnD8ccJsbbKCJOBclY34M52DBJj2nsk7wDbOscJp+
AnEi0uRWxKMPe3tHfNEbd0EX4de9aMMSlVzL49ntIvWxEIzhrCA+dLvygjommlkbUNJPqAs295rC
9Qzlvh+97Gm1uLZboy0CY1uojV91ijjoTv19gprPcQLVLW7OJ6TVzVPeih42WpCXZMQW/xEbdgc1
Ary/yDFSnmzC2jbWRJSRm82DPdMxpD5p9nRB4EQnEUnFUo35JnlcV928kiSLwxp/p2IF6Aveko+c
F12nQaWNykdc4gR4BKJoEgcA25DK1VmWbtvnaiIsEUTnXDlpJQnfzElKPCMSjWcBLI3v5kBa63k9
AqBEyfDuLwCmqwkayi6i9MwBsKoJgSZyrsid7MrZVR2zSkMvvtB+VYCZBBnWT6Fe/rEuB7FS6ZFn
XXgWlJ1gVuoplZBmbgpLkARJ9uNXIpwGnngCvF/nS69NcYrQUSM7A2gFjlKiya6mE/k722FDhrqa
spXylxHIR1NsVA4PyFthaMzsCO1zbUXPX9gRHF86ItkjwRE6H8+o42mUsPuvYLCwDMl3N6t1rrkL
9Xk99IVDS3aoCHgN/y9F/4+prPHhUDkc5D4v28MpjkDYhvXjCCIVkqQslzPge8j2/fRfW+Jjyky8
pQLHWGeFXEnFAe+uUuxGfoVhRmf7kNiEGrkSkTsBb3bYSz/9q6gdzjPLXQOLsRtlY4srn2Ao783V
IP2t0DHe1HuB185X/LPDtfY8aRSXnTyHhV1Ns3v4Retku17ixCTg3Ef+kyEjyMm1dMOAbDbfN8fp
3QgQv7zCQuxtnionp5+EqZRgyh7REtk2eObmw26d4UCDjt8b1yUIgh7pkH3yAIHmnHIEcSDrSwkH
gFI4s4ENU7HK2UOE6fbqMIpEcFznfKFSq2+wUeT2hFKbrwsMG+6YMrlTt4EwR5n9jhTgG3ClHJyM
7DfwZMeuLypdupduv1WBvofakDlYzntAkc7jcWkeYJUyrQq/Q3B95dJJQQq/lqV71lbTt17R7LFi
NCrVleEzW71pcjXICpLjjxcAkIr8W23H6+yFpPpa/I/kVSOcvgv8wMtVAykVSHoop+xTStzNFBp4
fJgDkaNw/FTgLqHc5QdN4PSTdni8p4VlrQ5mMsB2HyzneJA7SMoKJ0IeR8EO5wZqEvaAWCLzdl4h
vYCX/8iNijB6AIIyTmB7nVPAxHWQzvKP8QvQSHl9UFUY0pcpvxSqVq2W8vTWcVMxX+fHHeH6waNQ
FXlXx4gJ8mUfxxn8DzM9kXC67K3SxGsweRcue0j/daZPRH6Ob2sdYQOkUBxxQUQQDeuguqOmlnAO
7ta6wYdH0ZJjwK67DlS3kGwqQLWarahwzYpcaB3YoX6Tq1piLXx9g6y7MXPSyean7EUdyIgiAT+Q
Krjw0Ip5wIQIKsqfNVt9rtuIigR28KS1wSK8hGl+DFnqan148CX0TA9QXKxl+k7ShtYdQIv2h3ns
7ChJ2VxDj22S73Q3xr87s66S3/uhjPUVePpWJP34yA5xKIEiuU/HaGLyRcbH7ikqxhuXzBMHciRm
t7CkEMUOHGcPbBvLVaU8ZFk1wSKCixX0icYJijeaMqGeEsb+p4SnuO4/F7ItE26nQgvHKU0TmZf7
nBgSMFJfPzakhHYHvvaFW0WB2C7/hCHnyRQORYM1eI1PRAWBOj7Z9Bbcju5sPvtS/4Noq/FQnC9Z
BOagZf8ir6R0m9+I6mmMKbHyHJf4RKWxI6LiLmC0Lq8nfZZhu5Xo+Lnsh22lGuMKWCC3fbC9h2ju
nfT5MbaHJVcyi5fTaeko3bd8V/n4uGTBh+dRmenyf8W2tUdnqdQNgt0arNO8sW3POTnAC5DoGSRP
pN1xoLlQBZHGJTTLbA4uydcfYgdT2WRM5s3tq5ncVmnpHxACMAUlrJo0WgYlKj/9f3+JWd4kDw3/
aop3RJxF5h28T5rIB2Kj2Jal5NFkMnlg3VvLUaahYDuovyxX6AbbdnrwNXGuGegglooiYiExDEgp
J5IF6QXQ7qnnH9oDiO288m1sB/yRLs4FiiUSWTza5TZezoTLwBAdDjSFI644bQDZKQi5kD/jB6bO
y7WhsExmd+q8EQiv03SZTxnnGlMyhbXOYqH5n0Sgi/duiwcFMN4TgF4ePjjuvWUD4cSCjBezs3Si
zsK3NZMhq0ixOs7M6Z47+p0zcJLD6nhBBIKufX8XzIz5VG3VeUWKWjKLDgpy2uNlzf5UT0jAowZ4
YUKhPcqGLQpLnIMFeL9WlZLQWICcT9FGWv3go/u4rnQISDrwFV4+hegenbo01Ejw5WZK2RUoX3sf
0JXHvNAYoqvv8sK2eKRI19IQgPiuLwlx3zkRMlnE5NWZoE88wU+PLvbWHa5kpYaDBaccs73WZCa7
6lxQOyWKZXqYQc8WN5fFvw+Na7UeUmCXGRidkMmb05dLaHM+69HMNN9ZxGwtImDGi7F8FgAKtbp6
32zgs4o+Fqe2x601HIhQNvPEZXAVvYNvKFYHTe7In5uJuE2FCYc3iWVdWX22qcnUVuXLU9EfjI3+
UYOtzod/YsaknDPqaDcqQPi33ZQ4101pTfGow6+NJr8WlijgyLM+oiiCpe7W7mLsqbm0RyFSYRp+
wxq58RljJ2ZDFsWeU1DU2j9hyr/DEp30qNrtYJPZ/bj9I6YrJ0/VIYC+amvqFHc3CZsQ1NDdCj8b
W+Uvkk/MdeAKXdj3UMtmFBdHEy7tOYZz/idgOUNhg0eAxRg11pM8k5CrC729PuhI9pV0qYDKs/9t
HC7pRYZpb9/l/5zGW2E7PGmFOKwVQgqTtv4yGJyqGdV4TEp1eD1+puwmPeRAeGFWKGxGw8Any/D9
I0LT3j9a1T6cmFI2GWdaVAY5oCy9WUk/i8eRXpCl0IndFsFTm7B1Gni9ib1Qv0oIcr4yMDbCpnYR
Z/QQniYFUPvBvWwvzs1uaNdqNKb0YDpW7IKaEJegryjqVhImJAuVHhKDhZds8bu3PUQ0eIqotT4m
Hu4aDW9nsRzlJ2yi7zMmMbVlUZcHuYaWBUe0J6fNAu6kSwxVeZlZGRJWnVt8tQiESheXqMecumiy
qdwkaWHiw2jpv92WR1L8HEinXjS33wU4a6M+lFWV8rbfbMXuBCUDp3NbJBSs8lolY0GijBULGKX2
Th7KrfxXse+xtQRByn0daCHp6GwYXUHxgFyQFzwxbX1IHVom1SYg3g501np1inHfCY3qlyi1YHNh
fNykDW256wFAKhXdJwUsKeXYHi2B8mhN8V2vFc9xvoIvAc5sY2j4qIB0ORibzbd/p7ZwR4xzLRTp
TH3CH+IdUp7ZLfyLMUOpsA4zoWjYP4Kffwr2OKJGmuw3MAfAKEEwao2U+6aqlbOyyPvIrHfYACPw
bwyiMZ3cg4HArGzmDA5IL5lwaJkKqQXn42yWGo74KX2ACSXhXX7JyYgqi8zkwOG8s6xzQXnKS3Gu
StFCPELiuae96dBk+mUAL6MF3xK7V6nQ7Jpd1HyM1KR/odfn3wZLNk/IkLk5MS67AceidYWQBF0C
0X2Rfiq5PK0cdfq5THXFtHGGXfhsWn6cVZ0xK6a4fS5ib1go1vfQfZFOsuvinmDpbm6bSODDEb0p
VW6Bl+1Rq9KJu9e/qFhDCU7DhDVPMHfyRpe2gxYmheRzMJ+kyVwMHNOd2XgcuRmk41hKFk2QwKKs
TBax3B1mevL6m5oYjYuGEC1YZ1LOu/V3rKomRw3g0fEguHr6frMsZ5ySjDyLCD0xoRR6OAX9f/7q
h7ANDZCpOTErY0tCGzF9BC31khPNQLsSMFvuQ/BucMDQ/E9vX2EI3RjBQID7QQ/2mtJjYY/zw2+5
BAsqEW67N11C+yHsbFDlUwVhEVf7gxHxuju9WURMEuVpEV7YqT/ExveHCuW4SCkJcDoGav3JZxWT
VeyMzdY+7j0HQjBI3dofVu8jg3zYggUZXziB91xVNegw1KBjIfFSjCylT060owkePdSIZsRXJU7v
NZj5r7pRHva9SPrTM7NWZaUnZV0avx9ZaWbL4kBPFfuFCiGJIa48joiBKQxBnqpgcNKS/vTEu7gS
9qM+qZ0jOdPjmKkKHUKrBktIkwmznWOgNfJz9WqMP7aHapZUXDTCZKUC58PBhrX7Ggo+rEsm+7/D
ZmVrQqsOyD+Q6OeCruZG9mQQulGIn99vlkIG/TmLDvRDNCwlaTcZDqAIma1Og2d1CldEA8QjpHOd
wCHLhjVcyzpvMdtV3MHlOwFtvedq+pwi/5jeTQNKUes8w83KcWs5RPmtpU91zPPKSvoH+pfxHWXq
uyzGgxTA+Hb0S2PPTGHg5oSrSi0Ba/171b1xOtCeKzXUgXRF6IvGZBquE/oJVRqocfNKKHQX222u
quxfuPSsFKgs/Lr/Yvs1UL44cNHZN9+d/mm+PqSM+az6eBczj1HBmyu207gucZvcNaGcrf0Aj9XO
3WjqQ9ZykOy15gv6HFuVwSJrhLEZoNotkmap5wIFMO0KCw5Sqohwwe/NkO9c92pWYo63wzcWwjiR
Rvy64qqzjJ56r9vNw0SVTecXBa2QAp2RLDyppbBM8NuRq9SnMvwnjBQ3Psu4eNbSu2WuX6pH5TrC
Tp1cROhQRrQaUTMm3kVrJAQbhdlPhPaNY74ijWoBnCioMwrq6vO2qQnXODdzJxrSeVtZowsDFMki
Fnnz/ApXipuN57PDY4ySWYProQ7yv+7xr0SRLDby3jrw6S0vrXw7mlrKCsxZFEyhlTVWDGUsBWrT
UayKAQI5++7hQfqVDzVX40TkesYTZmb3ApfNqGZvMyegEwZ1fEfOm5gVOmobX+m3iWnXosZf0ofN
O/0DkvjGp9ihp9r/76dJNjHRWBHVOUDZmq92zL+gURD/Nq/Ya71umsMhBsu8LtjPHe3sLDzAyX5R
moBsmgi8F1Bz30O5eTOt1KJrZuEHejt7uhzIyK+wAyVQ4BCuX83RpgsgDofwjQvAUxJAHBwcDMPG
LkTTBHnraIfWeZgz1s+eUcfZBwE30Ya81voqDSPAgflnZ4VyoTho8vCHDgDW+KFeB21Rqu6tKCGM
GjkfXxarTZlsMR/9WhYefeb+1c/bOwkFHd2sfZP6YG7wnxp1Wd/+TwLe2KiacFReZkF+4SA00ohW
Wko2bAl8DEv5DGnDJjp+JRSbQGo7dPSkPLIOmRjneGqy7iR/JajAqQ0/fpPTyY++sZtjqa/m4U8h
QNZ73iiobi0eQ7KTkqep0TEPPnn2X+rgN4Cm8GNhfd+7xy0nyHLCqOVIJNGZvNrfiCD3oJQE8U5t
qfJ6i5nROjv8uiFw6ZrZCj+qa566EJvEHk8E5NwSKPeEAdHnAqFKPT6j7gOeUAjEWdIkKV3s1Gzu
UJ0dnY+uk1GHs8vZXvFxD665HBvDXZkSZzg83EjvmOwS4L23wM2zAgfMOsAzdl61ONsggvcb3BpY
x3tWkT50rDc9Ky8nXV9CL/QpQkv7Th3oGC3Z5TN2TKG99ZCE8VZTYCQ/zyfgBMJSPLN0YJ+nnrC0
B8J55TFzMDmAQxPT4kDZtfCmahMiJU7t3EWwVD9lZTTrIfmt6sdOrWnjr7QS964mo6RTCVzKF/MU
YEAgVb5EYMhqcJHV0cwDrmsXrgli/rhcjsGxcnsnPCa+qg9NgXR6Rhb9yZgeknJXyiGzQpskM8fY
a1mTFLpbJIvjviGA38umvqQiBM9K99XE6dDXZVRmddpngXBoGjiJo2oyXfXi5zJypKs/n1dJ8k8T
vapa/rHwzuePleNX2Ok5oNzlV1s//DuS32cMKx1dn9QeSh3GbSGgMl0CALlleHzaZcT8aAjsAfdz
ejJ0l09PgeIdNV/DqPmSPSn6nFUwOkluSSPPbnhMx/QoyeeS4UG4Xiaup3M90ALhghRKlkDLf3wF
Eoyrdb1Z32sWH0nwUyi4SO6hjYtNU/hgQmNQUaAspd2slWx40+VODJk1SwIGPj7CINxtaV6TT//7
CE4J9RIYEC2bQHRHVM2XWV8qOnpMkGO6aBHsz24DmYODhfBAtOi6vSGNkCH3xTwqOiayukYtKX9D
sBoiAPDjiqn7lqupQI/xYbZVhHREeYpiez8lkTOamea2ArAKNdBxCCSTHlDQpUp93qtDGVMOmNGp
lmOoFxmBbckB2mY8uBae1ebGjAp6lE+W3DQbg1n1YO24p+QSnplr4Jip1qAZWCQ7hy08yKKCJzNm
Xem6x/F7IMOKJsxDqP/zw9llJ3RDhEf2Nq1moGWTi3fr1r/XzfEdjpV1eHT2dT0K5m1ENDfysr5f
ftMXwASgXQYttURv7Zecnsw93i5rHGKA6oB3nx4+zH52/ajsKsUOiKOyBIT2G+yuS5bJPj9ejoRP
kBC5dThmqx2NB3byK5E5RXkF+ihYL85i553LjrsVBVLpQRg8mplqvf6XQypEEyB5n+Rg6m4Bsyos
Pz2O01KESnbdveiFV9vHU26HUI6kVdWz2rEvxU25PkOMXMAtV7L3d1G50itJgT2E4Aca+RzBfUC4
qFGgHa8822SMN4tYwubDnw5FbcPpIBo9Kdq5hxBP7QWdqR/HTVxX9e1y+wxbSMakLX3BuI0XTuRf
xRyixAUj2eVSvd5nTqR8AJuTamHIidmfgwojg+mIGwiIeKfOH82fCW1eDYG1s9xfOSJLBIWZELCn
5zUkQwWv1EmaSMlGn5h3YNL6lunAG8lk8s8SlbLWxuEKgB4isS65r/M1Rnwt8YEYLzkHeEmr0soF
AJHnkw2XLpixwIpQV/9/9Y+YiwM+DDD8IGB/cs9aUgDdn9JrFZYs7TCpsHHq5Vfa9C94tNK2+NMX
2yUuzAAr2IYMOxbf9mlV0N4cauYtVARG4ODOppO+eg5PHT9zkD8kaCL+3+t6LcvC9VKzhj5LFzUf
ZkFG/uJmEHx/2koyh9/2dGZk0WtrjkLFqNlvjp6GCTXxXhkpnQBGS2aFJ1QdWqZyke+8V9qIzxq3
OMhgIcuQ9iXz7Wl5WSX4Be70/U4klaKmiKiHfr+ZUE8MBV9JAIo6k78LrLdYKu9D3F7uJIS1fHAf
Q6JPQEaQjDY8JeHC5nC3Q6PVQ1YmQB+ems/FEyRTHHOgnaIe9EwXOSKxtwYzmQwnBKq94VX5i7XR
tH7TZpfaPnd9cRKP7yZq0kCLMG2BM5p09q2y+RQt7AW9W8oPzt7d17bEbq/+Vt7KrFCOzSDY26EM
RZoUV2VjhM3Yjj99PkJBdUYKGybLrTA719Mwsf2rhKHpAGak1EOsslzWYLI7y6x68OudqtIShbOB
PwTgQnvHK1ULJW1M/c71932V7pS4KiGXVYgXcZKXBRjhGJCFPoWmylxBLD22EE9eWYVZcEA9RXua
FHlAa5BLkn908FGxybXS88WdwkSvXLECQSSN0c6MWCZc+svmVcdvTjaBP10it9LxqAVNgvIt1C6s
zt7/mIrXFwqDZQmy/e2Lzslznm+hNlJb21kM27KC12YTF6Ii0GudnuFzyHWQZSrDalKIY4nIFT64
jgV6kLbNCGNLtHS9qIyVA75md8uoBDq+RJab1wD8yhtYL5ZdI8i+fItKyUnnozkPOG0PUIFH63mU
lZiEX2UKEbSYlBxXuurBy8ZNREwJT4jclE8GroARP/vZC984LsRpRs+k5imt9XgoJ/dn/EQtrr8P
x02KlpkKrMZ/EsYMsLrpdpQ9fQMzjb8ntb1I95zt4c9VGYDRnTqckLQk4eptiyewTPV8I010KU4X
hmhb83ebKMjtO6tw57wHpDJLhtJ1X5s6KMUkEPGCdE0bi/3ijLh6abC6Q7PNIWCIG6kdZYDWzPmA
TjjE6whJBSugnqfY+7EakscNBvZ2WT+f/7HBeRSnepEvk3K4MVxv13fe9ZcR9ZjuhYTznEI3G7be
ajbhSfhK7Pyxf+tAB+QJY2CLLXsFxay7koeIkkdx4ZG6o/o4QYZQatCSIDUcq8CNPxWKVFQKekaA
D2OgNhnIp46VW76Zz825GzvVZZnbo+/WRkVCugtgoPt76eIexVhHY4zQYtdoHSm684EXFaoHpW5C
M6jEO2pcA/jlT4tHvehDMIBSlcMQxCiRRMHqYtKL6Tnpf3yOQipu7J2uAVeMMZncUkWQ5OVIZz8G
pxV6o4GD+rrLYTx8cEmtU9fVvPeUbJiS0TQR9LlQ60t2n4RHAxYX72ekrHUlD+4qKJlo08kL+iSc
ELat+6AHDaWwz2J4AAsGFJ7JxCLeGcRmFRbSTJUWxVrZy0PY7BKM/A/y58Avo/FoQQ/nHMru6qT3
WyQBkesMaKO2SWCrbVmZyJ/SvzLOEBoT8hBre9Ldop+T2CGQsNSZsqCRt72bZKNYPq5p/Wzs/pxi
5/hib+EADyC0AoTMpvhH5jY0Lo7yQj2IwVeS+ye+HkP9d4aj/R1GVTjpDGkcFAYnlKC4pS2kemgF
U38KuCh9Vvc+AUJk7vDcR9W0e9ZaQ3vrbulW2R3K85GZ4U9KBfT8hC4sZsvCTpNwETOlypCksJCG
TjmpNrTN8l2urSxdw17uARdMalfb/h7Ym3EKH39PPDCGuGtj1OxxmCWKqiYcibOVySN3ijXaol/+
dFlW2GDsTIGNrNGn2OFZK9yJQC7j46ZNTsYlYzOg4UiWN3Ocusn9KrSw618/1g9bw5+jq8SAKwxK
4Pg8xfxi+sqNOuaMV0gc1SrJY28I26W5gIZ1VO3b2cDQvoj31dDTdeGn6h/yXe+lSGS62qY1YCao
6Gv55cK8vJzl0ie3pxtFNxMdMjRJRFlpXtr8kbfOHK/UISpYmf9xnPeiNDxknguQbIWLBMYCqFCV
hMIZzHblMGY9tGBGgucK+49LMPMQdnybmoSIyT7jjuvMEMZVxhf7uQt3MmeIx8HQ7To0fgJEIgU7
XCq2CByWuYu/ltocCa2VZKtPwj0R8AKne1Y6GHDurtUs6o0bGnjRs7b0D6VGAc2T+FIVC+juBO6S
UfRTbXYNWenYRbvCkgzajjeXvFFDGxtOjCyz/6DCExWvJSZG/bFAhWMpdZvW+JNv+HQh1OCpFNMM
tfb2quWghwWwxAhQZBpEiIGQYRiZFDk/NZ/ouVzq56dJFQEr5gTSb+hkqRseNE3C4SuRf1NSeIe6
ol/LkQS/X0haclngjN8mbW/BHBNDdnRaTFj2AkZPezc6BH3W7Owna6kPnnwx1ZW5A0Y7oWhj2YLD
/jqZF8W7T+MqtKJurS+kLFEn1E5EPvg96qdY3aSbiZoa7luJYmpKIJ9wlGaeG6/0eECxxFXxEjFP
sxSfUUH6j6awPZ4IOu+fq1Vkjm0YRf5RJb+19amabd4+LDxDsTkgFidraMr0JerkVQCofh612GgG
CnwOmDHHYHpD4us00iVjbUq3D5ONNQpA5IzhWW1uAXcIs+PZi+rsw4c444na7Y7s7lPgRFOYrArM
FGbndSlK+25kUpRXoWDUpaMM3YeH1JatU5CrNiiMca/pRkNuth1kX6NvAtekOIBum6j950m9djun
vHlgIfxh7OEDQ+MTe2hkoRLOrXjWgKt+pn/TzkmXIXCM4ng2r83oVFLyydOUhLOq9Dh21iviIn/P
1eFa68KyXhQ0g4UMhUeCmAM6wLSLxS8IHsyktCWlX1gm+MgeWsSjxH9tSLINkED16ZfsaC47yTGu
satUbTqef8Z+VwhtWeATAMRz/uRk/1Zf0YSNmUCsemFPG13IR0xA2t8QHPHjAiOStIu4qA0PV5gh
wXRRsH0oWiMVFoPTkx/9yIpr9xCFZs9R055INsmt0jbewiGK8GvouuRi4Qtltu8mCRlZqfFroEFa
i546t06ebHuhiqL2G/D7DrYFKH5LshVu2cuUKUv+AEOhOuHQw06eC7HZplkTRDV22JyMq0zH0nZu
TmuWziTTvnso4kAw4sgoPcz9t6rJc7NN8nHhA1NP/QQViEbkPMQQJlUpRyTDGzu3esqf4rcU0iC4
Us2PDJsHULyyngn2uTYyHuoMl7UFn3vugWkELQ14mAu5Szl+DM4MFGcpWQKcs6BEz9icE/agaY3V
FdwBH8XOEJAOxrMDRHjtj1j+q6GN7JAQzbuiAyaERp23mlcDodUAU7WHW4FbXWcrN4oY39oRwDAD
h/JDLIc04xXiL9S5MYJAYBVd6o0iOKiu/T5/tD0Y2EywtiLZu/2zBH3TLIA3zIyeJSy+c89CkDKt
F9lwh8K02wXegqPvKaaulrOXh7m0exlmEn+In/1NtHPr95RlpPXHZbMjmDX4w9T65u/ds0DnUFmy
PU6b8ERFvPEYXYdmBv4c/MBIz69A4Ndt/y9Pw3X0+lO8EdPdsXPddoosxQVAU4xBZqnBVov9WYuE
5ddW4f/6Bkbvf1b0Nt9iTO2oIzMRW+9aUdkt3w9ExypP/lQzuhVK08oxoTurt3FlNonnhNhDDBCj
D3xbXtT0jWnS9bhM+vDpCEWup4xvtmydVIKRIs28xDk5YU4iuMcYGsS/Bpnm33lFiwdb6dwBSdnC
wjnx77XvVDGQVQLf7E5odQhEQqPNc8OnxG+wK4+WoGEoxHAvdWlMvkdwArycBZgTehGlfXciq2gs
8e3SlZOL0nKBVSbihoeQSPb3VYtWvbOpuickuYI7vGZWPpa8qSPwJCNn+R5nVwUoooHMG9DFrVBX
ViekSVxirb3llH9McyzSZRad8/CA3BTv1/pw8GQHzS7dGKhwkqszUuoiPdo3eaV8LvqeDBqrmM9X
T8uRsY3Y4UidLILu40tMOJ1KXdGc/RKjp8o2Ij85qkcRyHFkKA9LKhhO2irxHvzpgpQ4iINU4jBI
FZ3BThzXZUZvLPauqgg7y8xQq/eOLY0oXgXea9lHCvfDd/RD+gxln+nh36n0ts9vTSnSgBwJP+N4
d0uKO7eeIgBXwvuduQuGC2ZjqUjgg3B0VUoo5aRXwxjMacSFEZ4Y2vCNP4QYl4R6QisQKQCtef8z
ujQJv4alvogKJZatyKGNldjvZJnLChwTPQGFARryYXNfUoeULSbXwXiGtmBvxvC8lsnnfSO+QrVA
AbywQP2g2gizXPjiB8IZgf6QJlCDEHFLhXJu3cvvpCyqBfZPKCiX1pPktBqyA6jCo1zzoRmnGLex
vn1KoWo7TsrJSmkdFLtBje7ssVfZzbet64A7b3JXT+YuZjwXiMUfCbZNC5gpEjuVDnrAA4zJveF5
ZDyySo44gcpBER+xlSpALgrFjOvyGGOYF23XpuHH1UZLFRR8L584WJNvfzQZaGBWid37AMo8Xqgy
zVSJgvttGF19zdVU1ZGhC5aYSGYCxOAP2rDYtCk01NTm8wkvWlIA/CCVGF1aK/xTwnvSurhOhkZu
vE8YlenpPn/4gyoBoOPYIFpHMCNWFOR9BZGCdMg4HX32pvIJ9zZD614towkR/wDMReUD7qydtl1n
L6GXIXir1RJ34rcjrQocy97T1fQof+Ydg4ZbMFgzm76oFqzzLVBR8WYHqgQx68AQHxhE/EigfoQk
S2dCYX5mnKjCmXjJMiSbL/DSiwZlY0LJDNiopKeg3gfr9yfn3CW0P/CDiFWEpl9xk/C9JVVFGc7N
zyTwAb7Y32oU33lmZlV/gqLd7+gHhlJttSll6n+OEKzNmd1pqpcdbBSloKQxheFTjvNPjDEl1cL4
GvNnzMw3WoO1WUmVCjan3aZ/zGeBDWNUwEmtOpPFEiwD2e4L79oUfXfddgc1x/NfLDA1ZprUqeg0
4w4I/aQYZR/+4u82kV9eUK+Cv1vGXHJAPWarwnvMePcqqsk9yKInJc+60TqX8TXSZ9kdmMpbsU4I
EBxeecdZIzKVoR0XMpORXFUdfRgirfmYxjWIX3Rkfiesaaw+e9t9syIg7EDvM/Sjkz7E44a15b7p
WcifOWMhhokCZJp1pO//Fa/5whE02JGyzrZg7rn2TKncEa5OM6HdnP9cPpFCIJtcKjKhzOdbAnpW
8d3tMlg9Duj9npyGeXcCQ2R+LXk7d3OM9vR448gORYCC8OBqm7sitZaB+TqhWJVFyA5U6NQmLaE3
XfL+zCcjM+g3QUw2QbBtV0fwliG6M/gBsgeE5r3ALOCVZ4rmJTtoF2bK2iA0KkWJizDS8xMx9qg4
ccJUVEcBYIYDDL5Iv2IMMmzDeOxjUJND1CQMYsWGZUmoFXZo26Y/2w9GYfD18Fzaj4rS8x8qGIVC
rg/qW0t7fr709kbpJrm98wzlE0Pnk1jikZV4R2iWIjT+4zDbpxbmftbhYTo+dTznbubMW1RgLXMS
lHHJGv9fKvN3VFd1BP/tDZAv00HNcdc4hFRYfqivgiMEN3qmc4QCewqHmSNa0ZnKDL8BiBoNSl6k
MKHUB1hIzXKy8/IwawW47ARcqcUL9YRYpvs7LW6uAUoarGtdhbcW4i+vD2a31SE42GkE/h7gizXp
3o5RecbObf2HGKVf8D26ceC/cfCGI0aOfB37l5uajfqvQCvRv3GTT0XuZ5b2v/K27OpAt1CqxWnq
DhoPB9HT8arD794jw/0GymgPvAkrxfPt8WUicrQBjfTFT56FhdbVwOBeuI0prlt/9KdX4CA38b0j
lbIw/hofZ3B5UiBMQz2399tdBH9J6hMbNGoiek/I6dms3SHNPXOzJqj4Z73lROPb0xg/hPYtE/YT
KP/g9Lx/8hK6tTBImipapLhtSKVBfL4qv8HgRn+RpVmjvpXasGSBOf1RVRzX0GvxsTCKPHPJ4FLI
4AzWgl66QbyrqVo3vM3mjYJXRS8uZoq7pEazn7Fu+G8q84n2szP2qP+d8aEoS1JG9pjBTThsK21L
XIPIqmgFnirxg1tPoHU1X8puBVFDZcCl3bzL5fH4Fi+cYx8f2VJP5Wjciq6sI7SG4ji6bhVa5WXO
gpRJXZ2hrRD6+Z0u222tJrvkBROQHFgZKEsfiqAZQpbXoLAmYdRTm0dxWQdOcBLKBZMDAu02bm8O
fXQL76uZaIiQbXAiEb+TeQjeCjniG2eGe24nbipc/AbHWsOSDXffRnGJAdGNQ2JmU7EsBTf1rKXi
3bSez627KCMuo5ys8+U8Cs56/4iPl1uCaFhpcTpKYsyhfsGbbmdJv8gEKA5FB2Y70KadmikHWKY2
I23rbkMb3KHo2eh+F1Xk91TiCNM9G4TL89DifgZFPlJg1WaMWQcHUc4yxwjB+CGiVmPwpL/jrV0/
jYXHzBo8rZMR1gbGiTztWyFXvXPL8Ib99HiCdayD/hwyRQppbyYtw2JWYdKR4JojgtSU6Zmidtef
aPMsR+JxqHatmqbTxmeX413TtSlwck/6DFksCsGFrC0u5c1wBsXzXUpjorOQ+lyQ8vCdtWPVv90e
Q7GdqPOraM5KaIQTbM5Q5DCZZifnsak0t97WEmTMEFvCKNAi5dPPczsgyZpW1SoivKPo+hTIHiDF
6wd3X/ub9FORHbk5lvD2kjLwqaEzHHwv6ck5eR2iW0cn4oD5XrlDhJfCMSRSiCZKN2gpPzMLpHjX
aSonm3yyX9v/Beyltp28G49zYU2zL8taXQJ9RfH6bdvmaneYb7xssMce9isliBaEM9eKAB5ITBPs
qixlV/3WyL6aQzSdO65x2Sa3LUteXS+wxP7MMPB3/ckY0vpduVuHBqhT9pxL3wW8n/QZUzlFwmE8
BABZ0l/C8MJTXHzLZVLaXhrvCCkLyxiuTX0ID7lkP9V42h77pBuRewo2teAQKqO34y7Q3hBtMsxH
uFJphVbZv7UK3Puwd6NPhkGKaL4jmN7RCtlaYChPUhJLknu7meXLOLB47RwZhZtX4p4VxHVJduG2
MpEAMz5sJMQ11k5Nnb2OYUCVVNPglXtMTsA6BoSev9ifkoiCEe5ll1+6SGZBH2ZNQdedOgRysXg5
MzHlOza0KE7QxrLBG2oxwgom9Grt9sQI+3Hp3DRjHSIQHd/mckLY7VPEq1ZCjOugJBHl8VCN8ATM
M/RBHwiMKJgGNDh3/hSyKP2A3kI8pLGUG9iveO9ld6fnvsWJqrhH76yQX6KhdKuMq6TgIFUprwSf
NKHG/a3sjhT6sG5PSq0m+cWRkyCGYjuHtMWgfKSeKHmJP6Bte+dXr5KFp62zxR8yLQFAxVZog8aX
6hjf+6J6OS14MNlb5iat0Y2PkGIYAVQbuf1t6K7SkoENphEDueYJh82jS2CrkhbBks2uM80hMtLp
hif88ZwktzySay3TzCpzlDNkXtUifzvJwNtf4YqI1fTPCkcqVEPTYloOG3tLjzPIFWdVWSdmIV6N
J9PzKYsPN27qBI3BWWbUxn7GPkZy3TnGL1mpKs5r5nNz1HPZ7FpXXCKaKpY4Czj6aVhrdQMgqQgO
mZoNZWUdfJO75yl+0G67vIKr2egOB3X2hwXualpJmhrDSxtalvAGVGL+axRPwPZZbSdKNxpuTGHi
aBK7jWnJ6exCRJ+s/ZXOqlcdwKuMA9bik6dWaqcE8iZYsv3l4tSazilI+UebRd0jPs0li7YbxV3W
eKdpTUtO5StJsckFgWypObXyPyDuRzSE2J5CCaWUeS+mv6aG4FU4dc20khT6Yh6TnBqkbFNWO9VW
LrkV/Bfa2jw7jxfH0SibU87oIWdjxqxxO7TqDhvLMYnhIAieYkrfH53srNTF86LjCImAy2s7FjDA
YiwL7AOnzWiEdyxXXflLTVgcgTrYyNOgS3h+LZASMp80lrfQo2LbuDPG26a6rp7TSoVX2whf/fan
7YCfKHSbx8RLwoc7Tn2tYaR76j1VgmjPQ7oKS5F6eM0sJ9AXh7Vm0k5jSuPO/hyDNyP3DFXR+eHl
tiD9SJv9ha/ZhbSPPr961l+paVHFzkOpwdlgjR2/yMKzHTTwd5nsiibyzpOBCGoUKNWGTcSGjyR3
twitxIsTDmgFwfLrlnzwDprq5FlYDyBgJprhxH8rWW14QfmxJZy3/BIHnCKtoKB2O129ImdfPPBw
QLogqtwwA3ajiAjx7DN9F4KBhz6WOAWqWMOms0Z0jaCQjy8gLmUhkPj8SBRbiWkiGO/ZTuAK1JoF
PJ4fh3BI4/LPp1dQOY3iXjVWvg0O0aHKm3Fmr1DxrWWpxiqt9VN7JfUske+xvKx0wujtYB/lE7yk
tw7/EwQrTSLZYMeA6uZhwu2l1pIS7nzcXvZ0Pjc0yI9l0XB7Cn58CQMO/+uRq8D5NapOPWaKY1D/
IpJVuPdoEbDEalQp9ioXRMO17Y+I8IQWYhH0bNPQIdfUVUtblHdJT2OpWYwQmr+Mn7kr3SyYmijc
UYwPqWsQuXfl8Ldec75cBwu6Yk1oQJV/gDT1fMY242iULV1NAp+MLf5+ESgCJGDkcsYVFJPU7gZ7
1UD2rNGBlgj8cUOaxCP8KTQOMOjMa6jvff/2vcWuH67bL+zNSfn1hqlJ2fTORPpkIG/vutIousqF
5j/WbtN/4Cog2/jxSmL1YSheDqKouZBEuzZUUNEA+NTN161VHoiDFxMVQRi4lMpvntjiaVZw68tM
5U9AQltflPCLW8LkGqGa3Im5SlArPnN7LeL1dzafJA5ydMbGku0I5jsnmsAoYDFgKNcWuZA6tm3f
AeWAOAWnJEhVq6fKrA8cBQ3CzXzOuT4Hdibw+GiNKQqjOHNn8JrZI41mGDGfSc8pM6zFUY9KQjhe
CG0Ep5AroqFA+OAlXjgeTsTUfH7CNnhBlyuVXlPBb311b1H1B7ijjqFbcZMMxx4Ulq0b5/CeFkyI
OMmR8WbTAsJzKOm77GJp4WKh6n2uK9OqehxKl8aLa0VyA4CY+qwzv0iqGHHYqgOk0ChPsSJC2qwJ
gGCLRB+fV9xY/pRCJZkimo10Fgm99gARV7yjU56RQqAg+OOqPCjZvYViz9ikfyF62W+PYKOXwJZd
PSVwcIKP3BFKL15TVumjjpo6tef8lgAflYRhhbbBri8LWwlF3BGXBbovb+q5p+YUjecSYzhuE0Px
cDjZlL9WYp2zTNwfzxdKYErTWHTuuTSI2dCibdp0pCBhUTJP5DSPnLeVCA3947hbXr9p6GlZeqXK
uC96rMivy0tJfDwk3zgxyUk5Esrf2LlJ2kUOtqZxSjqPnb7aytA2jUsDXwjRNEvbDKE8+pFl+T0L
TmIAkNAxhh22KTiD6812/ndrYcrC9stmUgYxiJP92DU97sjgaAGAAzueA+aiWH+ZFg90n1zWAQfn
SrESZEAo2/OwqKlbR+vlg+ieu2LC+vds9TUULVQShkQzO3nKj0iH9Mjzq7Yntdr1LQw3J6duD7So
LyDHtX1HvQU27eExlZmyLvrU7mviqlThujYNRWTBqXmws+QXM2tjc2YgoVmVTRUIUGNTNfgsZIV3
FWHOKdZ/wkN3qGXjUXHvTAzbBKUSn61iZs05OKfQerKZtYruM99tK/HBafu80/B1q4BT+7c+ED9z
7u5oJufeHuaAKMXeDzGD2be17fQfHbWR/MXUFoi6I6oxkFOK7/FgDPoto9XVgMXQ9Kqmi4bTYHds
rHGXbfH7nh7GlQXECOf415cTfkgHEPqBvV4HORsZf9D8/RQJXPrtIRtt//MUaZMNLgTG7y72L6jm
4m2vvg05Wt/Osf/x3HkZbNRvpanUT0+DwQu3Db9I4SA82CeZBBIVbYynYcZ5zr2yjSIm20CNmqdJ
jaLy9g3TbHp2I9QqHRuc3FleT/iCIezqnjmsvO15ZXVIw7eREdyohKRe03aG4qmj0h/zYc8o9PJk
GuMeIz4FUNbLGG/LCmw94q5Bgp61CLGeI5soLR+JEy8LE4EzMv9Kic4898x96WZ6JJaVCoKQH9aQ
J0Sg8pQsNVKp1gYDuj3jbYtbT894ATfHGq2m2rxOBodVGUlUTX8em82LVjNJuGTjrSU9BEecFgud
5XFJyJ5ong9Ko8ZVK/ahKp2KkljKh5CGVue9UkxapsKI3grR5FcVUhqDH0KoBQnFz7r0IkjEUo45
WtUOiFrz5aejma59C2GJof0++OwdWKCPj/PtaK/1Tebrq9pVifgzHUqntYJthnuSLukij+GgDyvG
3Z3DUWbA3WNMFnwSKyJmrxmDaRLN3MLAuXC6YX77Sw2qEZz9K/Z8o64U0Fm1RGxkzRdXueL2LVK4
mfBBSfmkoZtRLh7LCDud9/hkvB5NJN7nogcXakIdRklJL4HeFtdVNVgAVSBOjAi+SCuuXTdXxu9u
tHcHGrmY65slBfd3qTvZiZwO5RUjt00pGRLEblxj6vds99ef3YNbIiXSDxrIWmNBmIr6cCm4Hjga
FWp2gzVH9Agfd5TMOGBBFFkymKHbE0gMO4ILRt/QZELZL73EBPczdWv1XhdqmxM6vP2AcB07zOLZ
pVuRcYQzPvk4QNZEcvTtWf0E2QXIW4Fmbu2kvtSDztcwaxzbGacDijxc6bTMwA/poYQI/FtTFODy
KrpFavVTsIsLV7fHEycnVmnw+3aMPEASMEJ/WtwFbS6mXGrkef/0c7IR46Ikg+E5ObZV0rtXxrco
pnBG/I0MiOX7sdhWQUOAnu38hgXDP+Rq6ADePfAmPkrUwOOgbLIWUd5OELeJhcMTEgVJsLBJrgtN
3WibeAxd2WoahGF0la+ecxnHRShbEeucxtQAma8ABZa0y4daBpJoRuYIZPb1gL1Yr2OUpyR6WmRh
oiqmpuqfNv5T3Nm3IYfBkCKB4KgjpBY9+6RY6QGBvMg6BQ5+LvlknjYOiJAqTeMlZxvVg74SaWTg
4GH8ZV3eFRMNIPN2P5Fv059i0/O5V+KioXYQkgPNxYCvt/EhS2d/5I/IzBi8aV8d9Wr06yl03Sj7
5ahKTOmG0G/hFRPN2wOr0Rq4sFMTqeTHN8qgzg0okCRjgcgNr8l/iKVVsgpfIlWAnTjOii8BBXTm
j2YGv4tUFbGXPGufyU23tDqJgbga/bV1C5eY1uqom7wO0bx3EOqjJoLG1t/VlUZKgpXzo5mcTNzO
bNWDvX1BSLuzbqZuUxgTaKZfRj/8zIswER8HjkUhmEgQ8ie/tAU/lPqXkzJVoktTnimGlxm8niYD
x2QGjt4aNqiyMwJ8Za5RynoZBcIQ4s0pirZT0bCqtMi+deoZT49mSbFfKEeG2T2YQ7rWCVFkKC1G
Gbx8D808+uKGR9XjYPDLrXOEwfm6hDSJWCFFf0rtHQ359xNpj9olrZLos8hSLjCGAeN0l+AQ5Uwn
Ce5qImmEE0ilkE5JZl7QsHSclWbGvnn8B0fJ2eDTAD+rfiDfjSg32T1UW0Ni/HkQiOJpubNoXEEG
uebuLDoAKHqTocx0cjhFRIO3LubmgpJmlzqG135L3vfd86DGg/cxSdsrKlIYTo2rWGNIcSLQVWfL
a1tcjiEgIioAthUQXLJq55y14+gexCVCl96u9MaCxZ7tU2dTdB2BHsZLQLIuWc/p1fkrw2AgNfpT
0uaEjxDSsw4UQQTlxe7LBWFBcuibu+CDqMclM/jCmQO2vhWO58pqcw/A5y6fUOzQMYKlERSDQabn
LmVIyvlOueMcftE3gHvDajlHorabRgCNY46AlKaMMtFbdRZouiChExUvVE0NVr/M9G3eosMI4TPj
RYk+KPvt3Vd0QpqOVDop2S5LK2sApTRCSfujkiRG8FU9IQ2Mbbkn/DQ9J71IjxAHZchkgQfg1TZu
Y7nCzFDLZks+2yGMa/+P22HIxnCYHuelZTZWWS2tNXvWXIC9iJPc+wNgmwVtoMMEQSbJEtweTVO/
FS7FLqP/CDAyj786qM0SkjjdPBtvRjlo2ozbuv0Js3B3eS7oE8Ag7CcA/pl/3xzA5B9FaNdeTaW6
l/kpwd1/srT08pk6Wb2LErUCCbhrFTNLwgRxW4xq2XWUHEj1evqlOGseC8D4vMepZXC5Rbhm858d
9Pfp8Ud61b+FyROZClmPRc6OttkgJGFWQcAArQngaTEPDg8zOXIJ5tTbqFiVB+b1ijbCYmtwHfYT
gH++Cj0Vf4/JMFdYqy5S+lsLH/ybBfd8UmntVH0lKik5JCD5h8valLegqxwso5nY0NWgQYcd54Nt
9mffzTUHoj3rW5PeHcaP/UYdM446BY9wF7TEbqqjCfRitRwJ/Erww4vZ+ZeyTKPMVH5VCcRL5vEz
oOyu/XD4etU0/c3HvRlWzKzh8OrCmHjA9YkseTZQtAtEH8cFvobg3HwQFS0m+/uZIF8pW3szUUTD
LX+kWHzsSpZ4eCzlOkb9Pj7TR7F04BsZGcLKtdkv9RW2ggA3nPplWpbGfJqXF5DY7dt17Aa/JlXK
HRmxXyC8uyoI+1zdSmv6WZFzlTwqBAhdMyy06X5cQqYV/S9eDWtD0Pc1LIFf5Zpy7DgWR7FPZN6S
C47+VeTBb8M5E/ZhpYIdPDAn5v6+LApALeYB+eGT4wuISFjDZg9AK9t+yLQRL3Ht4MGw/343Xnh9
C0RfMDrnosF1T6Y/bl4RVLnsQTmEKcFo2ZN1hjnEeeU9efSWOSWG+IQgKxbMrRQdT1WDZoJlENy2
ceXC0/KF06ZqLIWH6x5G5acHqGClv7w3j1sOWUJkDO/fdQ9E6UDQACW+13w1oredevOf1ElgMHnz
lKkoHk/0LBG/f517D9ymbxOESonKqO0+vlxydiC68nz3BBzX8sKI+Y4Jij0wscaGOwxvSSnfasUU
QHuyMyZVFyR4BZ++TugLjRCG7PwJzOWyYMxE1HK1fNIonioqiB161Mf0omXjZLdGY/6e+liQgFLR
aJ2BQ5HuIwz38vHFB8c9DJiQsN7snVXb2VteWhWaeP6JDrICJWqSxIsD4yvifrpr8UT23VB2Wtz1
q2DJZK8Fo/1AW+aSZyT/9HhvEKOJYMEkpntNzxnQBEktB3UcA6K/Qrq7I7kTmGrUJdo/yuAG/KkM
W731vsUIM7Y7WbH0PoCOrvIA7vrkT/H0P2j/EuFs6CruRVgWgfP6V3JXA0xZVTcyOWXBldMgM1aE
05zvV76x1hpt9nXhOd7fAqcSf3nrZ9i9JA7soqf17RQf3coFeUSXu8iq9LpXdtxXgiOkbx+Bw6c2
4ZfmuHZDoP1/OiVKQH3ybfb4nDTOTSN5/96GOo/ehMhcME7dRegWF6kKKLmnJJZvSnBKdsVXz2LZ
gXO0S8/1R+TJrY16ft2VfaXWiE4QvhUfEpJiAMJBVoQbCxWxzuDgQqhKerLLq+qOZfZLoduwnXnI
2LHkbe4voeqzqROtMOqQ5U5FUfkte11Pl5rcWMrLd2N0Q20jFCmjeCfhm+1/KvqA4i4InDMOVuXC
fg+ygcB3hHO07CrXm+rCB7RrQbBpSjZqxFZHLPBkATScbQ88Gk31d3nJxAjH9uqgJ1y5wfJGtl3N
VUiuFwkNE+0JwTjjB2M3rwUuzn7DIqzwrmeY/AkmrfNuTvuQRcoI1X9CgUXtyE/uYyIntA0Dce/b
KnL/YBpyb7nodAEhR1ZX30Cwu7+ZIypBRCzIOOLEmLVU3eudyPqRRDKGp8kH+CQXG/rYI/eei13u
Zr1jPdcOZ5N7Swbf9rYAvnnXSt8ndTIJ3yilgqKLFMzw2FNjHvJGUk+7DEabFwjU2PA98TGD1jNR
OXZinVj0Q+gME7wwVdmmWyDyFqAHgrE5eeJnOpawd/6lO2/IVJUIWNxL7dUCH0fj62hhkpqpczAy
HA4Xyt8sFKp4QdvOKzqRCf9l/ejiF9tnOWTPqsBizC8NnuFZpJ9Y0wQcUu0cduLxTRz7UXrc5E3+
qTQqMwWy5/X49dBEsIGPU2engLeePn8B3pcLrnlHv8EKmPu2VX16cqRLZgLp6nVSqD9JEasCXJu6
theE7Zg5rLiupaz3aesQCr//VzdySWFfXshpWvgm+/ttNCRUVu5NcEFPdyvPaKWomPw2KtQUXKS8
YGsPIy5TSwM9zhQqbGFwQFnCLdqJRkT0tSvZDV9P1R71HyV26yH1roaeub6Lo0pUUoHV0al80lYt
u0wWxVa4o0BpDCbBItB38a8BQ6sbTeaZAGnNDUywsbB5jddGHESSXjHEL2Iy5toBZLugJOeKjFGw
1EFowCSBmCWk8CD/eeLO8/iPmK+cFs+ehV0h2Wfp5bDui5OHoeKER8BZDde5+ZprFmsZYwiIshDq
q4mjJg0hd51rFbLSNXj53PlvuYQkibz+Iy0XmKS3iuBMKOANA8KBpXRV7BR6kQ9meu+tgVSJ4mDp
UlmfpvY5S69ZeJD7UOZP5otua18FDttDLFEROOK4GwFqWW6Wd/iNeXp9mYxbB1ildkLd4BOp/J3Z
06WhTqdz6kSmJGjCpp8gpIIGijQ7IVMaXEvwIaETFGE3c7jJDFIpGt8l1owMaY/y4rF/iFYWAtqE
oUNIESitbjZaAMR6d9Q2Dns1DPCCK3/vuKCb1nq/gABBaetBjF7mkcNYE/O71cmSYOT8/MxUMPQH
03BL97IybaRkT9tHXKH7UTkdW7UkC7nWiAECOJfq0EuWNcQzzGO1v3bwHAgtiEy1qNy803oR9L21
0pVwlsRAt9eHo0XPcA1CZ2U3R6bYco8MTdse+SDqtwWgToZm6BkRki0oOLq440fkv7jVK0CV3cYL
hwYVE5agVh7swg5JYi8Lzf6ItFVSrRO3nUi5KZTDPvu+KLPMEdBxi9MmSTPfSIYjMycyxBwQ7bxu
SDtSLdCtf60EMox096ssUffwHOX+O+SMpXYRBe3nujfiQwoMqOmYgLtQnVCDiBVTchbqwakM24Sp
54eHy+AMuOPv2TOeBgi9FkEBY/c4HQXZZG//OE/53uuNNGiyKwfqdRiQRAEcZEKrr1uSUnGzRinb
azpDZal/YUh7yAu2SGMGSIgStWr0OUDwdP/5JCbLUZs2lhkWil+eTGvrgCiJKaX1QYMWcN6uiAmM
CN8bfUJ+7rs2EYIzrb+46ZuGvygIlom+CM2XAFR1JVFT2YnqKWYBtwt049xUnC7BVZgv8F9OiqYA
zUZV14DIyAeO98EG7qoQn/ALJIV6GHdqCNu65jVczX7k39wHusTbCJBn6DRGmfeZehimUNTlHydN
9nDdJjVqFpjqid7lLGfn9Z/bAFzeAT6nNNqIrcmBvD4UuA+X9Uo342Z+MqeaBMCFQkWxilv3y5sq
sNgfNIZkeWNc61i46YFFFzVUL8WpOkt3AxkDToXZkLvd4YskFzswCm6+1/pmJo5qCvlYn4gASuvX
RZPXQ6TYGyP/QP5kb9Q3vWe4jMw31nYJ8Fb1iuOO9OOvVus9eWIPDb0f8G0FAh5GqAVCU/7CEOy2
lAfEXP14+1VqemDpzX9Y9QLvynIumTBttt6DjGykFZqgYKBfijejJ4MJ8fv75IiRL01qqgf1u64C
nwvsqOAiU7qiZ/GaEV3j/tWBdeQtwgI5AqXWgA9pDzjOBJOKpV90wWCZo+nQdnslbBrGcq5nxKWq
xnRHFLTsQdhE3TO5jY8WQf5pM/52X2K7LGw3qz7EJ0FpjRLSX5EHPTGP2tuI/Mf3f5tweDFaSJxA
F8gbCCJNC0uoetQ9z8OasZ1xXKSNNvVydM5ryNakXQnLWTD1O5QDHPmgw7cL0kNbb1SC4uMunnfM
YkzdODjGOimw19w8sPDgA5O0Xz/hgELW91TsuQsCIHVkGC3erKIshzmZ47jxkEWqwDRz8Rvt6AyD
DANNpvevtYofX16OnyMJR+5IcFi1AYenOGJvFSMkVtyHi249zV0LlNVEaW1JjKUEQc6qVHtJ2X8L
BA36CX6x4D4QpILbAmqWVg98X0lshnqzqpmmkle4WCkkN/TEvSWzmDqN88S8DCNV5kKvz5TL4Kba
wnzDSElWhcL5lcoukhKpJ2f8Zv+AF2ZdG0SfTPRkkNBryg0Ua54Risn8M+9cwsdCLYa4D5JnunK+
LEwWX1RsEqj9G43kEgv6sKvfOANOUmlotIp/FT/XdXfK9SV6ueNGE9yPhdKy0sc2AQQTx+pzLdCf
eRvgFQGonmXVuOKPXKxW0OpixIDgNuMXtBmjdHB1k5uVF2wzKUtW/5W/yxnL3VzpO+JcrJRL47bx
JScYYNmFLmSSLZqzdRMBdMFEetyes+9fB1EYj0DSM30AN4N/+CaVGP3cVkq3JrbCgODzK4PeOSzr
I8tkgqKqsN35da0orIGMRlT1Hxul4bTiWJhFJfAjzmYzetDJzVQeXgAF3ESGnwThK0WNvHUaUUpg
XkCsjLNGqhfW/blwNvfo74m6PwNGU8BbfV5gOWtWKxFkH8Z5/0xkJlBpc4xGIwjNPvmzV7gnCLkM
D6OiFrFwKSei9Qg6qQz1ZIjStq07QyOY1ySfz318eBeXT7pn3fG1Fh1+IsF5wYpy217RamLw9bGd
zYE6dnQz8Xts9+tWJuQIsDwKR0Ka194iO9zRvreQKA9PStc0ZUDiH1kGMgnJ1RJiO2wfYHnkMQup
zn8wEtLx8tHdHSWYr3YWufRpRJtOlwnLKIuORdFdOl1xABQ7A1Jtz6bUF2S9RafXt4yKl2VIuXGp
fvoNffWufU8RAFl5Nhc8yvMHVG1lmnZdMAEcD62yMqWYU6qi4+ALze3yw5b5O/ubpKIdkln2pGtI
ebGjr34sn9fzoc4CH/tAqs3z8/U/HUM0x0Te9n8vY/TwrcDOuChckBqLu8STYCuVEzrGYCT8n32E
Uyd5ZGIrs3OrVStvQOvvjOaFZ3q2Xe1IziaFO6464lE00PER6eXqo+DAr4DQjYiouitCJOOYCYcZ
5fYT2n6wtqWrgTN+GyaZO5yoeeYc3XCImljbxnnGz3clmikUNZoatv+B27iSJyosRTXAc//za4zR
A4LKwOLShetZr5N1HWD4ODe5nff7hlHIcKXfTBh8eHl1wRPUg2hYm3IXZf9NLKslRs17G72O5gvM
K4Ec0QFwBxTqKh32Bl7Z4fdOhUD3JwphSI4mmvT4ChkwNfD4OpFprnZmxtQ1AvSYBJD2OlnRlcPX
f6KqPxMBMel+DPxeF9zNyH9/6060fKyy5SRV41VO8SZ7jqeboAtu/+eehfE0TZqNOfpQt87hUQoJ
f5fyBQZtv5+AmQPapMkobSJI5NecHCQmWw0SD36p/wDOXtToIKv4TwpzEimiWsvsKUkuYy6/dY+M
j/+DM+myF3G0l8gmF9JgiIqWZ96vxajOvUrdBjaPG6R4nDAhniBngoIvT4sPE3DNcZRo7V33XTva
X+1Y7wM2ZP1qcXbzPcsjhk7XDLG7gOuwiTSgoiVVbjS53cO7+tln/JxpNkWE3YDmgWmaGAK6USFj
keGykOI+KxjxF2HqEs3TDy73kuTbVfterqrfdxtsMi5f8BZ6ThQTaqly6AE2kcIfpBTJJ5p2xbG6
jSsbxsUmEyLwpZQwCc1sM/MVj8/OARhq1nXiheLhqDZnfla53J8FlkO2R1R60Ipy1ASJKf4mr8K0
ye40W6eO9asOe0HifDKoz3JA4X+ZlS0+vY3fCxS3znHxxueK7DIiX+ZKpyFwTpIshhQPxiFbzq/9
O9LA6vNj0SkhkAU5DZ04SXTEZzOLmSEQWtft1VqVBZkRdm203jN5jO3VkRiQGLvn3UDvnguKcdkB
qLd8JjQE3SvqLuVQH9AOMwvlf01YqLbCEwyUkkR0ONusBR+mjxfmvPpo+dHsX9Tl/Y5ANhajW3kT
JZF0YjWVCPtcUNf/PMArzxyLnHLTlABk7lVBaMpo0q/gLemQ5Fcsory7ZlBhouN4NUzmFolkDN+e
UWuLn7kQDvpeDHnQFBAVKSX9052t9GhtSoK9dAmqGr7hDxawoUag54f5jtl4a/2UjStT2mrU1Cmn
y2OnKIIndHGA3LxKwiHCuyasiew1JKbw1g81p+G8mO6v2up0nTMajUP4uXnEkrmAmVmgc0pthh1X
AwDTGakjj2JwsE8YU06XvuFUuJl/1o9gmACfZkAsOJ6HZaZOSuvX35xc15p4cVrBDMjS4iViE2b1
/tzco10lp51NNRhZT6IKwxGtdamHvjrW+PUTfXhiigC6KiAz6OKOai44JoryMdLDskepiVB3Negd
Fa84M5tzqji6vaV0XFkuN3qIaf1NLYHifAzmXqRlk56nh1ahmZnEm+y9Q3Uh3Di+g3gpM6v5qNz3
eJ4AeLvB66pnDX7Ph5J+y/WR99mHQFRT91gFTCrHcD4HSutG63rrAqZ9pigPEFebLN4QlT56bSs+
uh5z40of3z7gHTT+UYVlHq9tdU3YE1CbP36zeJDg2ubvL6zjfMNQTStM6aHd9uXDDo2Qe3SpV7wj
96GiWKAfg+jRH3gSzkNxG5OafQ0lYSdeRNoXluRtvELBCqBQ/j/edw8rbzRwETrPLc8Me8eafsh4
7N/gupmw8Aab9jfbYSwfvPCpm3VJlcUEbeYgNMaIrRyyic6c4pT40cgSKrKSc8icZVB7gnv/ySqy
KNtNlyRRBipp3YdHU2pGar6iU5hHtnFYwkh9WhTN1w+WGzgk+lLRouj2nM2DnCs2WHzWAyTx2kJ3
5a4VMyA3XzpVTIMPyoxHGjBU6lbknBN9GsQrb2AABqTqVdavuGHE0Pa2zlyObzZYLyrlu5mXM+qb
AYuJxExCV4NqJXgwJZA5ufuMbFJmJ3aEWgQaKXcuyojPKswiTfiwPTZLYSeEBgAwNSwlSu1sN9PO
j4uU0EA7CckSq/MAIxRf4BeQET/5Hyl6Nj9EjhUpwjkj7Hp1+j4znL+4EgeQ/KbONM8FDodOXbFM
Fgpv7jzJy92Q9D350EL2fu9fKhCbCeHE2CWsDTk7X0yyu41IDDmil8JBYcGXnk2FWmR9iamMKj5K
JevbdBCbO5s0eMOglLIjMwhUpkpS9Lz2APgkRP1myjdAF+tJWB7OzBZQbgkbvU/Fwq2cAW3wAbEN
4zX3xFYbhKaCEGZRDaH66JEdjIAqAo481MTRNjLlE8Fr0wd1EAl5X5E2nbLS3SBJvsMOGSxA8yNK
BKWiUFk977knqaqV53sWhjpDNKzwqoY702ZqXz4JSxXNG6TCVsMvBceChfvUp1JCjUmO84LvWH4I
jMlko1ct43+ZlEFO4Smth4pU3TCUmZiSrYn0PuGLNaXTG48Hpzs9ymw7WxsjDPjfMcvs6g46BfWc
wW7CSGNsHKJWGZoVlr9/jdIrJCr96uW1EqsmrPJp+4wnyfPpa1aYLm/omJ6TTY4GiOWEqchb2Jky
iaDaU0r+yWKVuSVh263QtiaZB04EeRAqQKnXZI52FXcrjPrJyXsurUDCpLSxMA7aycKScg+UQC+r
pXmbxiNzjhLw91fPccBu0bQzH71bTLhONxOBkOtKxqiJogOOHHZJaeu2uxoDleaz3tc1daDjJ9gR
5dh0bH330vkpO4etyq2liXtOYylPn2s87ez0BxYMSr1PYOmVTKMMLLm9T/V5a8cCaG/T7GwJ/LIs
mRSewJVcV0XZs2bM1JDcR2rp6OGGxmbRKItfo6Yxtq9hR3V/hfLC9pdYoxOHVfmjUKhn8aOrr+N7
2g45MnAiWkkQBRjAl0pt1Wva/qFOvcDfJdYM+vnTj/bO/7mt9wAY09GXEqjbGZc8SDUdTBALwpXo
faqj7Kv/h8HKYMhicmWNUbMY9Fu81RDwJmqPJt1f42rWkrhbW2Kyuw+cCScfNnkkZTNP5aaeMpMr
XzY2oiLohwXOJ6M6grBnC4BpvJnXUhyjEtuzrJqWWQJV09dDTkeAHHPREbho0lfy4OjaVjmgEcSL
InX4VJZNTmIa9kvevSw3BLOz2vxoPpU8Mwq1uipF7rMXEXS9d/Uh7k3Pfqho0QfHBdPqVB1TM6YN
sHbBt23AkAWXumbRVsx4uYmpBnpUk7YQdu50kydvE+0KSdlsJi7AP/pAxhytAhT49r+JiB7w1NUb
+s6t2H5E+YojaTvOHSH9Bcp6Ne8GzlVTt6vPX78bsERzd/EK3MY18wYEaVVWZNDT+rhSDqKBMqNZ
tJjpMVamhzdfgKFbzC7/vxBKz0HK8uOt39JvK+4ss1Ico2uxuFghT7xx4r8WdGGsdto7R+0R0agj
gEBsV3Kh+Qrnp+GcN3p6tccPab0EYlq13eqkgyO1vE0iQMfDXXrDsEHKYZJZG5diTbMUdyuvxMeI
LbXPuBL7SDAN8GuqzosPDjB+LmDYQI/oOFAOYGt5QdAgGel9GAYQBXETHtBgTv71aiU13Oya97HF
lHLTZ+wy4JjmkfBjekvTCj/vVIbkmO2Iozx8EWthCdJa1zDY7ZginLc8ToxyS0f4aSsVn5EGmnRp
dNZLRkrfHn8PW9lIj/ronUF4WI7kt1S4V5j5Dx4zwdqxtxAkWOjnTMSyBiExWIm/wyR0BMqdPGJZ
04z4uX+NL9lnwsYhqdTmw/jzWY/EchoP7V2duQq16l/+c8KRyxAWgsvUEf64Jb2rXFjHCH5Z+8gP
hZTF6AfhuQJyw0TztLIQXT/Gx383mxi8HBAoiZE275GdTtl0WCSe86lFeAYPY9ktG/JHprLVZzFc
9kd+e0D+bevC3wIW23D7jhUnho94KEKrnx8axBM/hCtIUbkD/sZcmFAirkpUPSfsJw4PpNFW076+
McofkkZg0ltQiW6VAvsUfI9NBPQrxObMWZeEZXFSgBy8E+32KwTUzl7f6cP58dsEwBVnxMcBKFe6
lYay1uHTd0cGe5cDFKPI4hidej7fUg0zr6lWYNtZP4FSPs+SsFmwtfmvg5QXHdZZ5CxpCox5uEtn
cF1S73PTFe8YGx8c/gGYGL+22Eeq1GBpoxr+8mNxjPyXt+B7Fa26UjpxnevfaZZeOC/0AHojE7pQ
qqiB5t9//CA1g7ObDbjGfIor0/mdE6HGmV1gllE6A+OYKarSTJ1pa+DP1n/iMNskRY4676f4EU2U
ysUL0laxc/oqnC24MjXu/8PaytRU4jOt1d1KtBIcOwB/lpAHn46Yx8MiGt2M+uAewcNWNoOAx+g2
qin+ZuDHHw81qj43IDP+NnrFtYc7s7ov9ro1nO32PFIAcCMuW9levKu05uCz6YOlu3HRRlHrEr23
2RH6Q9yYpE/0MakQa0qDxjSvJ7L/dyCgayO6mFQZNRs6CMnlzSJgVoSAq1Q5GQmI77hwM2J7M5Xc
7dFp3jDwcDlT35cVRmVxBsfHrq2sv+9RHLcla0NKGJPMmSyb9N8K0mmSAfDTOiqRZOai+HRDHxbB
NTILlPcuU7JbAW8GNFmsMakr3149wNkni+UJ7CjLGyXt9rxZSRdPXya8dOX5hs9KrpjUQM3OzfxW
0QWYIpAwaZTJjZ/0Xrwjtw183o8QoTvtsXSYk3fk755EPeoXNcGqJ+jBFmxl9YptHSHmorPfTtaa
5tfxj6IzhegoVFGy8nWfccTH5q4Z9l0CXJ10FLhGRUVxDeaxVYn1mgNBUQeWliCNKRPao7Mz5dnS
lTVIt6Ck1238Yi8bmxeHSHN19s5LrTtXjqC7NxOUrSsI4atqECl628XhwkEAQ1KX7JmQUdhwB1+F
qvlv4CNrKiFBYy3mFHRw9Yiohi0KkdsB4N4npuORqyOmfPm/bxlLAema/sTUOaYaBmaxnMC2xtnN
ZbCqNprNV+TOT+Tk1PDCRSgmNgI73rQMpxm4hmT987/WSKnBgvhMuG3tWcjs2mNgj7lxzY7boZAL
SdoZS8d0Y1QETBcXykagzE5qI7LcSM2sL6ewQWoEiR10eQamI/qHh1Fd7IWR4ek0I5f0Sddogg36
DGhXOfJ3lhgrpkZYwbPPYjoHEZg8P+slGjzGlEvU8acWTrlkdjO3ZIf5dTbPJ8U3WSKHjb2PUvNb
tcgEPRKeU/+XviuQQLuPwhDl72kAEmBIeNZkL984qVihDPPTv6JsKYcpZ2VtM9JstrEdR6szqUEG
1DfzZhA6hghPAoLdcHJjPit3U1t5uWs/4/+lehDP7lLeWVyaCWtQlazjG5aU1NgCdtPS4b/faB8A
LpNLeSYx66rcaYCnaI5DOcOV8L9xmmSsxN7C/EySrA5Ec0aRV5b3ixCZynjC3NM4rSBwtAZZnVlE
nCr0bWIebdNgVgLzwUW2vWhfBNs2s8a1E5CoQKx/YyNh/S7qfR/Mibxne838fbGNCNgDZGIKGIOK
04ffL4BsYjJuSgqQYWlzVGlDAcS6FF5xWwItn8eBs5sPX5iYfkylG2Dmh8M8OMSqj3KGR477YlSb
yqXq/zLd523W5gvm+/0dl7ck/ryrjPgY0Pwht6/UJ0JB9GRzX63rb2V/qLthVkRAcCHhQ8rY36uw
b+170m+K3Xnbe76gpGqXyLW6V33fZ8iXRPRXsf+gUB4pag+/1veG+vosH6lJE7RINjvx5p/YLECN
RNJezj2EyLmNPHL/WS1S28No/bg3nERO/J+tMOdehVbTxoY4Qz70Kx3OcgAeuf9g3qf+Oj98v8//
iGkipr1MbGhsZ1Au6AMxppow6Uoz3Nkw79F5X1Xp46j4Pv5qDh4LZ2u3y+DBRsFcO/QzV2TlvRQA
ii5TH1zobXouWlbDevmk/0nKfxkEtZ4SC3+mm7lTYxuNWnP84hNoJKwMuRE87JKtmV9sjgyGYRJs
HqESZztEDrTgw7c3c5KP+TMvjLt352Dmm06CZfx5jGmCoOFPQMb1B4y/0XdkUPJzf9TfHWbq/VoM
VPK1wE1YwExMamnxw14wg2C+X6WJQKscNlzQhaclbCW+V2mVqyKJDjHQBuGIKUKSHuNCPdrqEtRU
q16elKyUyIRRJjnuy7RcI8S3OyG/JFOrQYVAV6mmNSNkpI/jtUJXeaee5QLx/sNZamMJbc9mDCdt
QNSanawkQrr0ym90mauW/LJebq0LPvAULLE9Zy3VJPilA+fc1QDtU3SEsPSUXAFmuh49BpoCvJuE
SVoFZxWSGv9Smmxmt+KZlIeDznZvy/JHVU0qAnwJzwF71OZGdyvw7SXsDGvCRFocB+eZLrt6YfnM
nkuKvBLHMZyOPvB4dOuGrzu8/uuf5hPU8uvnDSpiQ+SPv8uuVbr141H3d0uBX74FSUUKeezgGycF
tpIxhhmdI5ype66QhetzvAbs7AF9RkZP6EhqnuhlWCBvzB+D0jULKZAoKlETVtVILsh/xI+2D/X2
muZXpuolMeZPYTxb1IvPhTGZsdm9gPyKjGXJ6n5SBiivfV7cjLd7SIM7+bdEo29ovz+E29rYdD9S
3fCTR5TlQwZw7+wgffZ+oYMC6YyOrD1qWn1fZsEAanb8LG7+dy7Lg768yfFgXkcDuOP4jjjYqGXc
cXclvsI6FfFi3nszQNHoOqoyNygKBDusW69jqrR3kjpP0Mw1sVJoidC4gq0gdKlaWmOBPDL0ct0b
A90q4u3FrqwOPdNZUwog/IJUC8uhlQ1B0YvQt5FlClPFVKLv4xufkbg1Ulqp8g/J2c300nguD7Jz
61TBRbmJfUmcwpUhlDAdSpVQE6y5MvOQsrVq2J7v9q2x+omEg1OodVKBkpoK/MxkNC/XXhCxgJEe
djjCP+X5DTgPctU+EigBvs5AvcdVX6sKRV9im4woOKmwDPS5FN59jLHMCyW715NnNtSlaD/7xxiU
kBi/nAbT1H+GNVWhd/vygTL/FyNlvfvrNV9tovwW6kWsUq3o1rTZrZ7Xvtj4TNgg/T1MRoBFVYvq
ouvhi/mQJakWJY6aEv2TSUOQqxPNlp9hHUSJQlU6bIcNqjra8CaCneYh2kXoJAl0wCxgApK7vUwn
Gf792A1F6jbiO9XvBvZevs7ryZjSkuGe49kEjwm7IqqMFpf1upBuVIyAAtWa/F7Ap1FGJBq1aHb2
iUAHwNWD2rKMShU/T6GaGucDCqwjnHDzjFxjTVzub+Ph4bn2Au9l8pM0sc0u73+9cYJD0kwhL1a8
v4puzotXE+QMihjXGxFM0NmJWeAIVPzfhODwhUVEBrqOdYryP06c6sZ95djX8RwPUzSOHylpwPE1
njgSCtiw4SGIgqvzvQ9y16i86DClPfV6p3WCw2qrnF3s4AiI9va3MoH4KJpARd+NQ90rdKfw5RW/
K8mCRqDGa1576h+OmHywqD0iO5MlXFqlFG6iqRsadobjcqdN/CQBRF+Bu7Ap4hxgiHGJ71kTgebm
rDaiEfaF+wQd9N/OiUgMQ9so4RRy0jcfcb1z1n+kX0uYzIoaRm8reuGMsiHv5Pca0FnGfyCuxc8d
VVeUube5uIEjnzBzUqlgkb9xsHr/3+nZqLAfC4N53X4ZS5W0gOU0LbbVpflbRE+vW3heSn+Ldwre
wcefqzT/KjLxiKTxuzzZc9reKUT7hy+xFNI4E3ryzWK3ZP3cmCmu9mNlH37ABiNjVCmcdEvQ3h33
CRLPYDtTCu8DP3x6LLPo45N0j2iwUSwj+AM5ELr6U6qRpBU9NOS9bmlsSWHa2AfVDNJbUZxBmg4s
K61fYhy6cRTt6/cXrfFGui836v5oT1e/DFY9FGyu8rAZ1ZbXZXuzm3J+dgLBM2jre811Oy4IvyrL
VUglnUwI3FPTKVywDbXrq5BpgSmcB2240xwXeJWTXMmW6aXNVZ5CLGPtvqQPXVyfo6WnaYevACG9
ckQL5KsDkKCqHsAS5ccWjTgdA8tnsL9pdnrO0TpyN6ZOSmeZnkXWxNHXibNitEnwGDy83AdW/Ok/
8IAV+g21FTxedqQ2d5YYHB5i7G5EwqHMHFKVVIjfGbcJvAVff+ilJgnalgTtedBLfVAZLFQi5rXl
R1CdPw+NzylTgvfH8dspy26bh+xEt7vOFvLcB61/mBEJCYUutCh6rTIcwszy3XnMUu0eKjc2Z6zA
+YkNyhYJbOCIW8EvJqAcQ4DF3kpqeP6IH8LGkGJ9sLdnbfrN82quWUk8qGlwBPrBmPunLQo9czjg
MP1nakAyyOYDhF2CPX5nILut5fJHmbmKoFSRVy8k6CF25npHagPVkoTnSlEgO5xlil+X7cE2V2pA
+opwft1c8iLJDrft2n8/RbkyNV3MgTm6q6Nj+x7CPDyG2c/ljv5xYViQS+t5FnSB7nvkvEMpGJju
BHsuyyXgJICkrj/66RCpKJqaC0aP0u3G4TglGvBxJQVNmaHk7e4DVShldE9enlpcDect3jo29k/q
bdVp3Ai7RzPgox5wX3ooVM/MEtUOX0ApOC/HpzE2t6+bG64x6Z748/4BwCiOXWHb79kKKAUxLbm5
knt+g5br63uExaI1YhrvjZs4yNTLNkX0VzVop4eZiW8DrCRpfr+gWqiPE7rwI0IgWMQuvzooXhBX
wklIKRlgBVob2KMfFUiODBMncO5Y+yA0U/6qMUFy3sH+IypauCC6fmuhzQNGk7RwQUSi7nH4Evr9
8Jtm/80Vef2FbHgS37lDCpFWqtcTqrJw10lYFifoYP8b/3S7pCwgj3AYYS/48ODZYsJ/G98hT/iV
llNtazQwMBUrbiMmHYpfJTo0fgl2w+0llIpP209om0kvcZi3i+rpBy03BHgrycuoDdHlOQ1XfGav
QcWEZNzJpnce/vVYRS3ZvTcFUPHzDOhLJBSEEHOEETEYy9v1sd0HAeTAH8lhWjvqhLWEamyiDN8+
w3aZ5DwfqhPYe2I2VAUMyTz8ixFBcMU9+oYzYDFcFl7A5NcxSVG9u9czghnEzmWzmHaFgjPO+Ouh
l3g9WV6FMQujZTrzteTvsSQsBvbsUo7gSKGF9qvMbQ4Imf/MIF/ddzP7UCPnL8sYEwyi/ixKHFOB
dd/FstDnWlxL8ZkcTNqroujOP8B+5/Vpa91qUVrEB1hZ/3x8y4Dme1plPBZLAti1tZ7vqbbt+qjT
hFbXEZIVulLpH4ZYQ0mMHF9UeHb43Z8O+Fsx3gr0vpRAub4ihxe+qCEmYJwLs6uD2SVyH6d80mxp
Xl5wMyXE2jN0B+phC4JM2ulYjP4hdUfqnVTkBbsQr3OCgOEfVj6QGcJLqswqTPCGoSQ9YUbWQ/M+
/17OXsyxCbHwUHjwJ02+pTjKf0IkOZjlJl4t5iITZaRKPpw3LnrtX6MH4dgkefq1eXA2OMksSvqu
0RLBc5Wl39iHnZpUtXZBsbLB0e6wRyML2gOVlJbeqsKRPzZLsdRKXvPyjerfYuEmYU7SzN8unK6z
rld0hn/JsglVadw2+WXCK35/VICFeCqmFU37z57MQYxIvs/WeYe1hjQeHiEkAll1DyU9E04Bl0y0
Z7S1r54Iw35FKIykQ3Tcxfdl8b1sZAWqD5G6urT0mBIaHPjF9/6/4Xww7YPR42fSjJXbWfir/3FY
HgDCvP2fLEvr91i4LTOYiQdWxz5a1x6d1uJMRq6Xr/+HMU5usAE7KpbkD/DzBLC/oIvLPITxrAR7
rd57YWnWFXWPwLmku183GLjpJNnShRCendT0qjj242dC5HNuRFVRUlvyMbPkKvvwoULn75pC0NBY
dl/oi2lxUI5d13xfS3jYk6qQ2hK5PAdXItP07nM0amqv42e2akPyeSEkfmtAPNkIyge6e4HkJZHJ
QX5M0Hkxp+za3v0kOqjz7AFRI3evs4ApO2XCiC67a4DHpfpsT/BnOdJN8FifyOlC8KmWypNuLnml
Kuf6zifIFDqqbPSdhcYv54GpbYkNIt3J6WL1bjen2fKD2tuBCZOUn94qT+G9oDek04owYllpxwnY
pQ4v1WAT9AryP+yBRaciDXeBTTUe8UuOYRz2TX4v/1FfV5NQmTbGR/m04sQusgCZgyGk8NxDG2DJ
BoJjkZHzFE7BcyTHErnAGiFFS6Eg7rx+LpKqQt7MFeoQY/JEEdcQNNnIBSp8wvB2D/TUk6tIwmht
rao16vDDaxjToFSG7QY+il+Bv1AW0hBcxixDpPQQlUwkmNOHE0vNL5+zOIAxzxuGJQDKQUmW0Z6e
n5BCZDvNbzSDudcJdwOlF6oEZpKnZA7rC8wXxM9we97H2I7XPryltlmSCQYBiVpDw73qR8lmYvbi
gBfOxR4UJ6EV/ziLKVeUtx91BzScoL+wN/2MWzSUEdrVGGGIFEWMjgqUWSvQ27OrdueKqQw2nkD8
ETNAVrhmOFZzZsjdgzeV5CihDn9KkXwO3IIp8o40L9t83TCOhzZzzVzs75NDUpJ99YDlAXAwiIIX
eTZLmbdiPSQYt4kD6x6NNmytW6LGCSzkojjconTbCAAm8CyCmQhhW6JtkJdsF52nPORiPdBOEJqt
PMrpvEWa1jXxsZnFLq9SMeXJZDXoaXnuLM6+kB7haI+2BUH60td+PoNCFQqv8GcuRFLLeVwFrtIR
MLaPhCQkVPzk7iT8h7LkjkxHWhNryM3JKJ0vv6LnT/4p17klkvqMj2BElIsyzF3VrrhMaPfAxn9f
32RF84m3Dg7gD7nDoC6HHk1Ig7u4DfFqevnuAZUSPLrpo5IW8C7XmQqWCJKSzNBIATva/anrkQLx
6E+JrJQEUpq5apiFuxlPCL/tX7+3NegtIzADZdSF8iFt43FMguGF1RaV59SAPxx7Hqw8Z68HEUI7
BqBxD9sy4b2h7mRCQWfmW6ERzWSxcJ8b9DMVrUbr6U8pxdUGNJn51n1H3tMku5XFLxUcItg9fze/
lPNzgKjRVHGs9nP0XRHj8q6xn0DYsYK0X8AkP9xfGpLWqV11oJYE45Iay0h8/+FU1Ir5q7Hirf+R
G7tPuVQZ+QdKHeOOpwaAjmpKResP2oVjGxUY6HVJet7auMcH/LwSPV27hhOiHYO1i8PvGgz5JGs+
yw59ffdcwhpjVvP6C6l5sNRopQW0PQBjkP/a1Pl1147bHJxy5YBADigRf0vTTuvLCNqMPkT5wVW2
k2MGBjL3p2195jS5CiWY8qBgBK02PsLqR3ghxCq6Jr4Xkl/AY93X7gIwVVwS8J3p/LGmVmG7O03Q
G57mmhnM+zKaw2hiVJBXu8ka5c/KmovU2tUPD3V0Qt4ZZHYQxfqYEoDzUxz1HrH6OHPxRYiG2j9B
NNt4rf6cKVZ3r3b+FtLHhJn05fUt+lJXOkO6IRq8FrdtNPuNwftl9cRqOTeRUdrhkqpEeFNI5QXh
xuGhHl6Iogz+sCiOWU7h7oEg0/yL6dSF1UTks3WaEUB4F+Bk8zui9zSNY90YkW5n6vKgk45NSkaB
iE20t3ddShuYYnnFs5yCxnLUMKJ1UDm25+kQ25IPKS7lrJln2g89g1e6C0hQEiOdVPTj3rBRSWxu
8hlk2cyiACCyCVQ4KEiH23U8Bt599cNOSkcv9AlwiiC1XgHZKz27qcA58kJoCJ1I1AB+AYDCV/vh
N0g/ifNsYd/CVxMreCZFbbtnChyFcE5ZxAjEuJFYCoRQzUqD8iae2AKz8wfB36r2HFpu/wr8oXFS
GdTT37jD2TljyZc+pYPqmEUPdG3aLEoGZomRngNijetxIjzqq6G4yYxJw7S1qkZ1S6SX/1AcDlmv
obNL6EmGFY3ObVlv0/dJRbS6OLMvZUizLBqTO8FWOCIFEB9FrQQguP6fkcIpfTb4T8Qgi1Svm2Mi
AP1vqSa6PGz0MLYVlM5HCRLKTTwHR0oLiYHlo8TWEUWTMJ3oK171ggloOas4g9TPBnNkyRWuQ9g6
GpuSLRs1z2YH29uSupvNqxmkKobOUzU6IIBoa012UqsGQn2EiSdvRairQFTTScmeDRvO5MTkzD0C
2olzu+4Gep+JE7K8dtvD+3IX6E/Bpfd8eCWgclMDG7JMdvxY04JFJOGfRjNRleXTSYBRheJ14wFi
pXc39LMU9cOKoXMgf8arXCNg/XLeZIHKMY/OjnHt7nmEPDVEZF5whIUd9+VnYkByu9iuLn9M8Z7D
+eIZB5coJ/9N/Nw7cQoYxtP9xfSMzg34GKGLcAqoRayYA6vM6NZNlMk3ADt9ohFstWJsojeIkA3y
0YBKpslnJWgbotS14EfhfmjLM0mUveiS0Nnnu6b1mKIeddMoSpIGi9gfXNmRcPO3zyLsJGeGGFCs
kZdbdPmfKNBbAOL2LokXFNYglFM2LK2sQOFIZOYoqLR0Z8HxKp+UU00fWeqBGCGTgKwPXgMvhYMe
n48d5snMktwvhO5pOZsFGu+1TZ3hrLwGU7u6FETBBYL4HxcYY2jiHYLOKRardh029YIV+ldjOUvI
UDG0IopvMLb7B6sduJTIk2L6vWm79vbt+z4jYb+rLjQ6ccSrn56GQYk5FFWDNJddjwddks710c9W
7hE6MwaU5JmXsCNz8V09hRJiU8hjxiT1eftVk3/ZaE2Ab21igmvZydN5fQ4uAxK76esZN3HEGGrP
q04QlYvmJJJhMuX8hSkLnZlfgvL7EorQaAm4ASyIhKwZJCGGSiqo4AB4Gq/XiJ0emMHThOEd8oR6
0TcRXYD8/zzDWQhmvGfpnmgwFUU9vnK5o/d5EAaC0Yf/Lro0gTGKMvxDBEOgIPzkw99pSgO9Vrmi
iHsr3al6KTHyr2PmDfIYKiSa+DEkHjMJHTKSSoq9z7h31a783hy+IZ0X8H2qf1zf4Dnz8fgVVl26
AKkPltSTvvpaK9mc5WfcgdCAGEo2Nxll4/9A1KRTkhjKuslAUn9AJCiZa8F4PugOZaX+DURABnRg
9xV1CO7H5uVnbfgMJC2cHaES5oO4aRVctiTsY2m8eKc/7cl8OypFTr2hXpB78cxzlt5y9SXVZjfs
lkAgZeC/eaQ9wLbDUaLL/2D+EMuwjbTueBhdrtj+7M6kWCdDpIoEuz7zF0xHh81j0Gr+DblD1svq
dpwKHiiGikPPf7bMmaIoBqnmAlFoG9T2ZHC+Az5y4FiuS/m/ml6a0VK3SYUMPYm7BXdTe0I0DQiQ
O6pBdHbn3esGdpm+pKvmJwvI4oUHGLvacwrTkEGPWKtO3ry6dzk/KwNAQbQ9UFbhGud2PTEHsBZF
DWSjYV9ZzO/hBc0uiD49i4DXX715DmKMG45sP8mwu5AMA9pyo5Yi/tnab5xRknoiMChd1pPff25/
NI5Qu7HzgF2BJnqUs5/8/xb2oxe2aKXGHVfe2+kkDC9FT63QM8J9Kkraj0sNlEBWEXvNPrKg8Dwe
Mt70/Vg9e9JtxMcvOsD5rk+l0mxNNN8Q3pmFTE3V1m9efCEwtRqnn5gsXDTlFRaTqaqyj0rXX+rx
1X0jOXgaeqOW9tvluyBp1P+hliO9OsvB3FAQXh9gX3z21k1ovoGpfd9FHQdJfWBR+jlliV3d0W9E
sgY3PGdheK09nqyzWdRXhl0SVO6FxGo9Roe9ZVjbO8CKh08pHRe2sEsZOMvJmLmE3+mAI+6rqwPt
P+jqo7B1cnPWOeEaiQ1Jb/fHF2TzZNL8Q8LUIoE0wTT9LspASVtCD6n4vqro9MoU/Opl+iEb6+L+
diYs00FkNUDNPTp+bXZnchn7wr/3t6K5thunN3XvvrfYTF0JSKmb4t0A9lVir3i3nkLcFbn08wDL
4Dmfsdj/BxAf8NL/GkSbh5v10VcrLQGzxtrVNRx1IaX3tVrfX4dYKyI4yfXQiuC6gCDTGNZ4wNxz
/fMfo2jgKs4+4xlU9KGfvULawJaH9g6nhxKgQX7Dm/sTK7wkfQF41JiOOqKcHLTSvPD3yMJ63l9G
uoPqy68GUGMhVZKDQ/TDEL/TrNvJI43GHYRbPJyL4UZXKPNPkRsG/zfjV3BULrHOAwgby+VtsveD
OgAlbXKcjIxWzTK6ddwSwTc5uJs8ceKQzUD/h5IfjjC2WJtc7rGsUks92SZp04gzsajPKsmfMRAB
Mx0ZhLTzgtgbV6sgBQnI6FXaZ9yjzwFQh5ypEa0KSHwYgNKHQv1hrWxzJoM8mcoO7qWXcVGXqAdy
WdN/YDVrzguBsVBQbvb1rNuVmaOASTY1gAIQG9sGjryV7BpBSdsp/vsyWgfr8INiqIAzkuGVG6RG
d7kLRXIcKTB+UdaSZY7rrDj4ZPAZeHC9fu0SYYHv7WxnBib/wpetj+vo5hoanVaT1xCTvk8xJunT
p9Fv8PCqGq36EGa57YkbPQ7vHiyIr/cor0iEHZjt7UyKqNn6K/OyK3BWv5ggk7mlUm6YmrUFzfd6
b8kqlkib4K9rvSIaSiGQqwEzGgTtukdeQ/W8TtQoXI5MV7E/0ZVUccPz6k10EkIuYMxDqu+ePX/Y
ZjjDpvKa9lzv9Mc/g+OP3CCFGjvz6fDZdyqnhvn96V77Q5LndBcSrOqpDHFcozUarKLkTvVApMai
+Rn05l05ayv+aig1sJuZxVZ93axWEicbQjhQR1MG5p6ZaUvDmuQ/a+WbmdJvCxpyU07JCb1QA0i1
BNVxZpRJz3k58m0rghzQ8EeJKB5EIrgzck3ovf5Daiocx/iAz1nlf9vB2RIX8k3t6d1JK/JW0F13
SmYy2yRY5TOnl97lrzWV1pM6j2glEYSWKEuxg3IW2g/z3Z0xZDlJQiXHSVWcW1vvL7HY6BRf0SPX
Bzf77/BWil9u+/n/n7zsdiG/FkVR44KVd0cYYwXz5ASEFY9YyvY0kgY1OgimZnv2FmuT1BneL+QT
rubBg4RoSjaHofGfl4pUnXYXzQfwyphuiGL3CtqTnh8VgtbokIJ0wozAkd9Z97nNAsZlm3qBORxJ
XUUiK+Hx+56CuFDbJVJSd9Iui5hYdqEV0PkPGgRYADSyRgy6LKy904Hd6HiofGlbwaNNllnuqtE3
bBnnK8UT9qUSxOOMdQC3bcJqEPiDrq6zyb8lP4Vzcuu41PVRac8wsYRbtsUKvqKb/dHfXUk9uP27
L3sa4ETmypJ9AN64VDDfZkpFChSKW1yh4jKUmXswGBD4ek23CFQVCPBIfNvbL7QRv/R8VFYk1YKO
ZlTvlURGQbaMuDSZu2JybndwlDNU7GQvJKzBCcL0bKCx6iEaUAR1X3xt8dTiePRQ6LzkGGFqscgO
+VRpO1wbbSq1gcM1X7zoqJHoyBEOrZcJN3UHADkZKcD3wM20flDl94rlNMXaf934rOBfkBWCuEVE
PtCYvmEheRAdr5LGdb1MnTs+ygWhCewpCMxGI7xnoSCkAkB9+bRdQMLedV/EGENbb3vXBf90Y+8L
h3OyrOaucDfGKAhclVdrbA1HDo6rgFIDenT4bUVNoDqXPii35yyDHkCL/QEEbAwQZxczKnzAQF+5
tZT212/J0pSG+Y9vpdgKoGyylQSQ7tXwVRpQIK8b57aI3dgWTd8VDd6vQ3opA+gUXrOvIHGJEZrk
IKLBM/vgc91VidVrnS/ebuajqblFZDiRPjq8GbwXsqm8XWC5RFrwPfDocJ0GpVmKMc6jEMXV28uT
wAayBefQVv4Cps49WHkGO/YHN+v5lW1f3QwD1Ctf0hv2iw0v6nic4HSgGlxm44LMxyPgfvLeDc2d
B3tILJlHnYf4MMZi9l+bWeaFmhGnvKJkxmBh6uNWm3EFIuMBWV8Qg1Kfhv4xRCqqEPmCyt9qdQqL
6JzJNPvZHq1qWRpAl0N8drwB8iCQfuM862Q2G2Ps1V/i6JXfiixlYovmtdnuX8h+rmyy5WaPV+Jm
fjvTxZav+VqTYmVd6jECuaH2ElfXIEovNKnQCtGfFQA7WMTMaJ3yrnkVoY0vWVTxImGZWmVHy/wC
2MNYQFsbOQGpPwjX3ltAe5cSZyJUoa8j47fZ4Dqj5gvYYFnZ10A5sH1AiqQcesPVA14qnsSfp5ey
ho4LciiadWxZxUOk7iwA5PHHYEQ72a+Bo/s73or+caxuv6x521MThuvMg2g3LxlFRm6WKSOiS5Df
g/k+298L24sY0YA6cs33KJwmOhEzN6ZazzVDNTYN507glJYWdlM4nkapdbIc9cLw/P72Lj2YHerT
0+7XRU6DdtN3A1SV8dCYVSOJfUCZSji82aL+VKknKrWeSLzu+AeN++Bv6HblSAmEyzVURPAlYUNR
bpp220jXg7vMEBVE1hWPqcD9wQd6hbb+fpP20Be0ihvng/2TRx6Zad/ZaUmuQuNmS7oIC7K7/Xnp
fFVslXaoRJ7Lor0rcwOEZlSnclCg6LzMFNExPc33/Xqa50V315QPFzZRMLwGvZFoyu1xym0obZYJ
/dzrwB64A2OnmyYwnJZJDdZgD370SxvOEcLp7dvodE2JEzRpY0fus0XeUjpCi9naiMfrbTBT4l5X
HsZasxqsoz5R2t8yA2NOtb5q7RRN6EatPXkP2QmNbReXvEJlGC4hS9zmeouAIc1ozeHrFXRwKRAe
lTuz3BaTNDurMWjKqQUtGPOxZDAngbUOYXso85b2WT2Qvlv0BtgGRn6AUa4+annsfQFYj83/gGt+
n/0xhljiJj5vbfgS6RfPGYYJ8dh8wIf3JBEzHKJcf4/2eIwAY0vvp/D1W9uPZjxYzkdVYPQTb06c
eOut6Slr/fsNlj1d4RgJTaf1HbFG4wdDY8Clh7PiSeDsG6o8cd0q2nVVPm/LyucUSjlnvExvgyaX
dWz3KLBCIiAzTAr/v7RyZ7amxVjUeRNCpZs3nSUcRk+rShr3GI53/Pw1P15bLhSnoRQlOL+UAVU8
bmsWOei/V1puXsW1bKfAREKMrmYPM8KRyfxeXWqmvf1Qg8SQszPdpqKQCSqLFYa+uIlve3gEAjaf
RmQ+gbnewCUoqNtz7qNixmO9JXn9zkTcry7abyf+AxJ9qDjq1Z1Htfh5Z881ns+GGFFvMnsUfSFh
hePOBaQTvu8za6IGzh1pF6zpW33DlMixlnKa3Kd3phQxeClTwoHz57+/XzNZS9c9IcP4foOi/XGy
AIadoBXVmSXQgfZy+OH35lOS8Q/glDUXO2yN3Gtq4Wyc6t5SQYEKBoXlGJHJuRYh845E4Y+mUIuw
I3fzJrbt/EtouUhsZAW2jeD36pPVGH5SrwTCYJw9UJrbgPEG7yK7Y76s/5FhvP9IRFbAAHN+0+ME
VHo7Y+eCVjerY/P3ze1nRZs9nQaoB4k5/THKarb+LzGJFYnQbZwCt71qFVZjEkvn1V8q2K+LG+Ht
ekz6Z5LIzvcS2dmkwV+GGATFDe7FH0N0tnVJPmu0275/Y0TELdkMYbdFdmJAdX2rZZjqk3MDzIpb
QNLvODzgzpMbq697rNZ4SFdbaZmGqGpSsfX9+To/N0Alls3OhsIL8now79jOpMJtoZ1I5rsE620F
Q8cE8YQsY0sNTyh4krKbqyw1IBk66YlZiAf+tblqv6maATlRMXkrFxQtG4XLD8ZqRyXhTZw6o2Ds
pCwroqKm9U/3Vyx5vDHvXy1Ebt5571SOiKoRxagkGqaVD2rDH7+jUdZstQHUFv4m5d6MHvsYo/sV
CVksPoS1EKJukeXMUKcrJwVZZb0HHHasAVn+TDFRiF5QgbkDptXVrPr/86u3ot1P1Z6atpypnfUW
+GZALRp7zX9ZcNVU4QXPpF+f/w9CBmFOQ9R0m1cpREG8ZmZdu2acwKEbtxTXZ1Dmngaz3TYpRfip
7SrkJVSVqz8Q6m8HgRgRfiseIjP91fVznWuElaPm/RpXWTlgSqlVo7r9XrhtNsIlo1WjrFEcSHf1
DmJ8xleecEpU56rCAxskNw667u3E4gpuU69W5yvYrPtqQgBfsvKQq2aYxktUdjfjMsNDb2zc4Zoi
nFqOUQkeVUBnfAorQypE3JDTAIAXBXuhKGEG7skZKoRBq4jbjXJEq0eNcReuo1joREJvnj0xfAwF
1MZZEv7PRO/IvFPvJWZbI1y0Nle4jZT2Dm7eikO3T2cbfraMoVLvom4ElwXbmHcC+ZXYbXcAIt70
vCJeCnlTDBQw0lzHRAJRpIHy33/S3VzyzdoK4f3FCaq5M+aNfYPjjmq/dhgibQSMQA9SrdtuUk+i
4FOYO+KGIRl9DcbOuay7hYViQeDUWJiBT3RXDprojo5lzy+bPj4fnIiW23wSQ6UgAQY5PF++adGr
v+A7xuurNeYc27qOxweu4iUsadI8V+r8ILRk54Ktt22fCf4ZZSf7mfUTbmcKhu/VJqup17YTOuyO
eIYGUZ+V4xEjkUjT+U3b6EpZWpR9ey/LuC3IixkOeRszQu7EsD6X6vP2NzLyeQ86eNuRf57thM0N
QBH0qv9ASviEFHzGlycQtv28K2vsleZhyZkb3eyeJmcn6dJ7oQvYFSXgGMk4G39RCZqqPKLJ3Za/
mTXLN607kg+uTmbCj7/GSNbl7fxcM8msNvD8rhNo8qFwExgH3A/F1Wdl5GSdlJmLZ9vAzXfYjMO+
Qp7jZ2D3/cOY6wz9vTMKPotJ5bh8RBnajTkRdvnBe9ViC6qajbuDHt4QtYKAq4VuVgbNSsvS3mw/
zW/mHd6hV1M20NllmhBfwA3ojqb8mEjmk64A8LRgdUNsamjCk9fVzvyVj7CyE1wJf2nzjl4N5TkD
jrxrLQh0D2glzyiBOX/VCoM+CHQboCBKKVeZGXCK7FaKeLc/RNr1qjbv0VE+vDcXWJBfxCK+dxgA
vUHA0XK6m9bMpW4QVVvdLtOIbT0w18H+tXeYYMoKvMeDOdozLqlzDoTpGPeqUP16pwdaeaDbZM/h
SeCHXuYgRUDgNpCla6bs84xct5fCBxR3iXKdCjtvCTMXOAEj8Ie4cJJZum8H1D8awLZmPPbplrhL
bbNZMz/UxFFmYZKzPPlvVEWLS2OWzeFXHLZ0JFNpoGzmv7RtIK13P8gkewVqqT0PANhGDOf9adSr
MkaJuZDay2lsKpAc2S+VfIF05fa6HQrBWh629JDCyoNvn9qK+vh+EKPQ+gCxSYQUFnsIsm608c/t
FhB9YrRXd+i5OQmF5KGIXWG5MEPp9tbwbjLX2EH0LJ5Oqd9RVRm0tmqiC+LFcWWSTh/Fr0BYBxs6
eC+6Wgzn5E3EyGeVUysmGNRxjSDU0tPLpUDU8T4/fA0smowTGyc1HlJq1MLz2Lq2KQLvajfaoJRv
hJK2hFdgIdH+KjBejq4aVQrsUkrM9iRwDXbuZvOt1MnIs1KJZr6zFqAJesVe6I67iE498jWrHzLI
bN8ssFC3qYYFloL6Ja/rxhf76w3iF0ysRic4Fs7Oit0fj6iNRj2kl+jtMQY3sJB97Z2cr3LxUw3B
Z4dTVi79OxNmsJ2l1sJEIy58WgZS28uLDTvRI6ii4jq5ZxpfzheR/FiouBj0oKWX4qrExdAMnFIV
u2N1z8fNG7NXNxUpBJnkoDQ2PiUR+BSP3uYWGfMW4HKlrGOHewd8MJP/PZ83VrD5CMGAjr9XSKC2
srW5sqcrlf+dA9v11RHWioJ64QwabfcYYsTnV7C8+1VGUgYsVCXqRkvU1wbzEKP4j9FGL6poXPmx
Mk9wMiGw7+XGBB74Gd6bxGBZDBeOi0PlvjxzEx8dNcrFGmKLaJk5wyMKJD9P+hn4UvrEC9hhV64O
ViAFSk8rvoEL678KdywH60WzhQeTda6vQ6b7QHicDe5QNQ2BXcChCtQ/5urhXRGGk0GFVxFIdgJL
HqAfqq1Im1nhV2cygEmMfK08MDlGFf7GKH1Xv/qT2t6OOLJw3MD7DBLJOR4IZIq0unpuTDmZ94zI
Cg213/bOyWW7Ti3IZ1rvxlnpwQADW86g5sTgGRRw1KFIvew8BB/pn/vcAXaLOf3zd6dYQkhuxH2T
HoEoxULpQb8TQZ0uMkZ2WAW9y0CgzjD0pJbNeDFfrkdWVWDf6IllxFVg3EfcP5Cifgtyt6WpjEQF
EqsNHuMHftO34/DnJmY4c3uyzI63Ajl4Y2UzWMFnZfmKhbqxyDBfYOEIgpt8JaGkKv6Ajmvq4zC0
oETkPoxhGfLQ7twgAfi9sDwPf7K5TaTRZUyk6ooXTDekfiGmHLgNyuorRk2iW93I1z477i3h0wZq
fT3Krc9Zlc3inkG4LSWNDjY7fS7/gwMQOeJdVI3kS383qhJDc1NZCdiPFTH9b1ibg/NM56CXeeyD
bVCIVCG9HvyVGwaBwwp6DzSlGamP9/zXw9j79krUy7DFcDoa4ndHAli+XZr434ReHKvTpWNrVj9t
Cea3b+Z8n1MhFvurKOIKZWAMHmVGIBsz8knpgaSHiQPwcYMn2TwQ6nThlp//UkEzRtGK7JrfA+Qn
7Wq1fRiakWcr4/WzTciY9fi1LoleRYjI8sejNgWoTpJlbV5PV29A5M2e6aJaQhT+KuQe5Lo5tLeK
J9jGdyGu3J13csMZkwHZiZTGJWoQsr0riqtbxsjmTYKMT0vhNVWKzOWagH7nPx4sHYytgiggCNVV
R5nxE0tvqyAenIUP5qWCCsHtXKFz33LtIq/QGE8y7M6Nm++Uu8Qu83FG8WyLaV5ZF61CQYsEr2B/
1KJCn5nQNyqRH1qKvBnIR0/ItriAp7een6H1tLd0xfVpIVQ2d7h0MBxGvICsIm2bawCERN4/cr7n
PGTclxfBkaleDry/mroOfC7VIYD36AsAYnvW+6J32jlcU1XqSaCMbUFqm1UgFgF8JWs3WflgzNB4
cwfwi4CLxyqTT8u3ywB8fU0oC+msMY43eyPol2TAcQv+jyOXrzAE802+0ufFF6LigvDpSB9oEnCQ
W9I6iQPD/ACBHSf1//DjsVQAOOxqMydlaWfcICiV9lF+n/wibjhB8Gg2XbnW713zAvQFH1Dv695y
VUrYrkyp2ysdqEgoFNrsE+5xhwBepOVC/SP5Ilfx0KGN2sBbQUFQVZ8nEBn6JVmhwiqMYX+yITHt
yS8Fz5MnTkbs/dbu8gMg9oXkUBImMSGOQjozKJBH1Qw/kl9v7iAu7/tCUvKgn3eMq+Ise9BQM7zF
gnMnB6J1hL0s/DASZ0HImKMpbsauJV7dG2INFfpIN0CMXkEBBCrtVW1RuszGZ9TnIal0Ybu3y47B
ywkiu3gXm648u+LFNTsLchVhAtTo1lFWpe6jKjFlDBkbxEZ8m7/DcD3grcz5j0et9NJDT0BwbUa2
wxQyDNwsjidBLn6TaN1hnbS+fJb/IXjfZ/6DBoX1P7i8LZoGArIfnb6SpcRcYZ0o6n8QUKuNHcRx
cQqolGwyJr9ScthWiqmQ2t6q8Eu+7pBmbVCswoqx/dzBlDHdfQXAu8EFQMVy2nIGPUutzZ2rDe6O
4GioEfHGJJEEebwb2NRdeRkEXHIP+UskAoRgGUuaYgRoGySaOmNCJdsjaXvaHBaXy/Mo3g0hMK2x
g9DttR5lWLayRaNlw+u0mpEmmI4D/M3VxqtcxodwINh4tyC3PXRMdSvlZZvMqgxYpxIY5LXUj4FQ
jx79fQbmOCyQELjcmx8Ew/hJ7iTyJJVPWKlRUcBxSxZHpI7G8VGKvrztdxM+vZRG/Elra82m+C8u
cPglGPl5dfAfHDBVEBeVJEhyNg7E06rnsDrnvfZQVyH/TjQpLQB7EBusnIHd9yN81od6v7GtRyKP
Gq8nCCjq6G9qtExniYm8Isu9hJZjIy7hstt9OQwRyFfaTZoyQF+5kyF33u+IxQGNax2P9J7gWm/T
u2jzoNomc0CBePNg4k26pQRyes/bJ5CA5CraMnl1qdVCNoy7GQj3+ZTePAKZS0hRZhmI9ra2WQG2
cqRVlhTNDIORD8TJJi73SeCFmJ2LaKesa47BSVSa5jUsFs2OgjV0A/b21xe1KrmLByG7U3Qv3SwS
t8xxSA+FH1PT+qufahngTb5iUSQ4Il/qhdK2WNMtUUIRS1AjcLBPVwQwjEisAajJ1GchnVKqOrQt
mEYNhhReKCn3Er2U6Nm7pEH0uzB0WTpbHbuf6sEQxjc46iBNtWZQm3beERowu7dlc8v9xd6eF4k8
1J5AbeGx+bRJPi1LJX4XFweqLRCrh1OA0+B4OoFaI2+4GVhrRl4srVI0Cffy/rkd3gu0vmwHk8NM
poTMNN9Tbr+t4G71z5R/2koXuHBpxHmAcJ8tZEFhUWiIdoWYOrxVnx2jNolxH51/VvJ9tSJcD8Ay
ZDWaXHy96SbOUSxI0+MdyGJIiIAOpsMv3MHD9qyu9dpLtgOUh66G9mkI/3sP6qGNMwRd4o0RtlGn
MUolTCu56W5uiL8kthhmn0nw6HIJsOhDE/FgYacK75YE31kX02DhCGWRMpXfQHND2SA8QmSvgqwr
5rJfIu5CmmXm+W2ZIOnp6Fz76cbIPqVFU5Ki669n7iwcGE5aeDwq4HuHC2Ex7AJlPMqPCySA4LD4
O2wD9wUdTPKQPteLlOoMbYOmWmqYsrUtVDg+AEnfkyMqmB3Svpc1t26+cnhAyVyj7henp8i0Mr9Z
//zgZvi5wECuLPcbceJ6H2zmMXt2ViJZZQlqEXIC89iUduH1RtmR2DBPswbgzlaetYyFOCSGabZx
+a/1uWrRSBc8wMK+CMzXS9LpuLcr8p/CNCGvh1BGIgwyBEOYg/3bT3yLCd3y/MpfdPEx6JbBITOC
C3haRMImO6uW+RQ5+MslPzS6c28hpMbr03pdcL8GwfgmgyUs3+Kt94X73svSqXWvjKPthCFZ0Ai3
nrD7Fe8NO7YzEmAFnJGrSig5bRGCs33Dnf5GdNAc9RLRE0U1hWHXnfQQYtNo2UblpA5osMn77O3f
OR3D/bgnhH9VSnlLqepOvuj+qVcyBEsknARKjdsZAcSTwDhBtM/hbz6jaTm3bz5sgQrI5Epv4/R+
3aNci21NKA9p5x7hqCwaZ1e2dn/TqfkW6obY2UGoOTv+uEUyIyGB98JmmXe3Sma3wO/R2Dl9Jn2S
K/ersVkCxegCdkFB0sInMACY1gC/YlFC7st6SAXt0XvN3rqUADuqVGfLXPmHhIo1czSmS0Z4nx/Y
FYoXfla1TmPvYXXs1wW6gUOpNUreMKIu9WiH47c64cJfM7uZv6+e6gN2YRwjFHFangTKifDs+gVL
DI002t7qwXxE0L8YxJ97idhRfY6awhx6tYuNIj1OcrJizPR1cUYlc95r3RWT2Uu6xKD6fEGl4+Yv
yziIdKRvGHdqbALYZj+WLT8hipe6b0ZCApfudsGsz3crNXA6+OW9zv8p/5/pcI95dWsWkheusVo5
8uPvtiilNSJ+3j3DaQwAiU/HAx8wjFugTAGjtvKU3IDvWTuwhqe+xhzZz4gsnd22afBqqeTBp2LS
hSpqRQlp5GWIr1bLwvG9qzVSTW1R+q7iZPwdC35ax9YFhGZTk04NWgxc3kBdOXXAvZRS51sejYGe
CJbuk6p1AinEElJ86KvmWhEHgiAEIqb8E+e5T00TjSDRez2908U6D/Tvz1IucZw4Cv+y9ZHs51H8
T2iTgNxcot9e0+Dot3kdp/g68sUqUufK10zFgFFe9ZU1pmZDVJczXIhCwRO+s5s8WaTCMcjjLQcW
ZshpFVjFV0VCWhbjXZd8mH9pzVzuZAtzo4Dht0QB57gbE4v22B44hSC6IcQO9q3CfdWt5ZuXJ6Nm
JJXNY3J4AkKEbFf793KUjrEcJ2ttwrIwfFZbYt7B3uWhhC/UHuHt2AcnOu0EAIlKwqnd0+W2wPQL
hQFBALcKXjTEL7H6RWw9dWarVN+H9vP2i06dNcEsQi/AwIdAOpmnNdVuEA6Dru8zL5gzWOIJGyAY
nh60KUd3jvdgn1lnpqBRH16VrZ5gq4z6z9bM2UIt87mruedEwEaKX40cZvOY0EbkEmBvyC+xYydA
EuLd1ODhFAt43kX9qAg2grfJWLGIFQDpiWv47oJxz+8Vx6fI6j2ozZzhwUoELegyhx9VdcZAC1FD
yiPeX6Fu+Ms260kdZ6UXlmm6ELa+0CXFHKWowyJTF+IxqbFhzbAZP7aF8lKtpYWv3OXZVXZae8+u
P9xboiSlpPsq9O1qP7iMjnfe/SwTdA7GZSSLJjY1NpDCs3ozWmMoxrzS/kHQGJvv5dNyfyF0YySa
WukahXgneTV+MguRFsPx99XwMMISndv2sFbJ7eG0Urcc+vzc2HNfmkT5xocwUpqdCKA+7/AcrgNp
hwFUFoZszxR8gRVTsA0qL3M97M2vG1UqiJIUmojIeCxyXAfUxjv8uoZMgq7isCSPVwE3/UFpxA4n
4xOBg3X57i7r6o9j/btYvSVA5mYrNBXwYhX48MxhcGmXsPEI3vnp3GV4a3To+UW+Rg7rVRY6BvAd
KII0qpbRPUMA5FF94JhNmX0j0v2tz5FGzBDl/pmBLjIjYAFV7QPOCbioBn/O6SAwWSdopZnJsQ9d
dBZIJKUBRzekk+JTnNuSNIyWKEgYteqLU5m0ifoJQcklFfQ5I7DXYkUVuVh+7GNqKDO7dHIdcqcv
HzxOZNF1gZkuxCUy3eop3nEe8rkW0lv0gPyKmwoR9Gb2PJwglg8LnV/1JKmvK++Poz/mU3zg/U23
+QTjWMggEgVU8bffyK1TtVz3tNVRt+hqP8ZF8i4TffQGAfR2dCKnsFpqzpvbw5RoDwnSd/7VAh7/
3gZCZgSBeTB1TQ5EnKTufi/nkW/TAm4/ipjpSAj0E+JR8acLa4g4/zwyz8Dj0QZIJMGL74oK7g+r
4ZSTzGuH3ocSLDhwMwu5eeVdnkBCOmvybFyIjZA+TlctfGn03tlgUVdHadoMWmbeFE9Yr0oxNjqq
ULxLD9NANsFpHLew5WOyUqQ30Ajc6TX5kJamjkwn9ASNIBPTzGsFbor8MTuct2BWaehKdxyKqrpe
CbZObCRiDWQowrooksCyLbVq2J3wmwqUOosdMMQxMo8R/tMEVYyBZ1gd0WSkdMmGlWBUB+wAzq65
ulpefI0Ji6dzWG8sqdHkva3sViX91lNquILHsFoHAq1CId8KB9DHFTOQVypclJMNO5cM9i2cCK8t
8HD7KkGwRQ+/De0BZtgkj0UwnjXPCSx1EmDCHuelsPUtjk30wLrlwMYJIt59nl0w9I8gYmFNn13P
8l7HS0wacTAJNO+LQYOEnss/T1iF5iN3xD6mBMqEu00/pMG7LTF2q+IKWQDQCWHx+GlQZAOhLcQy
1h9qRDbxITnecYxk5W0Kk2p88IwoaTqi20oPlelICfxkOFNynW5XFXoviy8mSQ36tTyofzqRnXd+
s+wo4cWQROx8MdWCQL7sryp7rLUCFaO7OPFH+e38zMq54EohywQiMmka2D3j3shwdI+mLZ7UsOvG
woDsAX8pp7Chp4E7PfeY/dHpmNII33+E6l0mxstYpnULKIHqRVjPGdqSnK8HLlUlLirGzdtu0mzz
xJRyEEyytqAtlt8d+w9NmjtX14ZjlaG+tKFO/6PkIHhTV9DsIhi6tsstpgTxcvH3PQvBZV7yuJub
qk06GQXUNzR7OW45erCQtz4t4Uaol9Ickhn8FLTYzjydBpP1lNkWVhe+UnI4zp5wwb/XmJtRbfty
YACFClT+m/ZMXAHWAZ1FpmRGaL8NroDLqCAiuGpsWDgxVCvLrBy/qcXxsmQjCTyQVYTob9mrbcPO
xGlvbdn470xua2WGq/C9HWwy7znGX+BNzoj/MGO02UyxP+clIcPTFNlUcx8VQrMO2mo50STMa8st
Aor+3Wv/tL7vEhY/g2jv8oEMqgYTy4EqBkBHrHQyVs6vZXjV6XcEF6xGfv0UdoySctfUZEIASniX
/Vbrzl/KQ+4utK58LtVFElBxn1FJdhjcCmQSkXzS66b0VxObZLurU3AdQaKCGP8JeEjVrMYpaMkO
0o/i33exo9107LxP3VGzlzhpxf0fLc+QpAuLx4a4L+EAA6nOIJOpPWTt0yrDw2bprVr8yk0dwowt
usvTSUDMjFkdwb+sYgORlkZS2RfCedoEdySN28PSAvt5VfDajKXQPW2NIhncd9sbBvrSC7N2TvWF
QeBTFXVv0+dmNaLg1Z6QZrHUQgj8NxLEbPoxjyj9uwMaih9w/lWy81CDDmdEoXPItgGINvpOtAgi
okp1Rj4Iht8Ge7Abi7+1tweq1PiTuZm/myJYRdj54sBgXvpV5uv68RA+5KfU1zRMEA9knX6gyYk3
HtsupFhieRSi6GGTcOVEO+gORSC4F89F/IECsW7a3WD2eZO0Zs2XGpCe5rVA3eJ2Pamur+9p3SZH
EiIHkdGEZQmea+xrtV+LPgvJFWegZ1uukstFgHeeV8g8CcHRc4y8dzeHutzaxSzhwHh2bjWkuiSl
o75k2irvI3nBfy1fNTp6iAlbG4pkIK8ZGEJsK53+4plraoRMSJsqQYEI7C2YQJ06HXQUbvG87azJ
GkmQ18n25VXCi9yhxKWb77LpuI+VB+q2Yp5uknMlWiahsw3v1B2UCiXt1eXVhPEK11Ca9QzhQE4O
XBOPCJKA9HPPgnD+HIrq51N/5Ki7IQUuUxve4OjGS2IhISY+drwDrg7xDZtSonCa1wYkPb1pMGA5
l4MXEhw+WpWGJFrJHr1j4ppx4hMASpWZi1EwKihAv9fbqGMP8C7ehujKCqimTRBDBx51AeP2IIsT
S84im74UYGcYQtuujijHmvmE3BseDv/VOoegnl8qnDOwSZmpUMGzGS+RaGr1a8RYA5A8KNgbCfTu
79qEHOBkkIhi6gW+8ilWJFkwuVkbn9ykb2otEklppDZ3DuAG2n5Mi2fI7J0eG8B88gkJg35bgrEk
UPwDzHcldL1AnFJau66SJztGAp1D/qTgSfRdjjo540Tk7wbzHurxVG5mZlKip524B7gfXWL5IEl5
LeRLAcu6yJfGRWdyJsW5vVsRnJDhyHlGfB34+reZidCJfZsaFLgQhVkOVR4SZvbaEdYRpIInMxGX
SJ8j+XnOYlPN7c6ipHp6wm7rdMWpxgdbFOuLlKkxzxiDnhc+y5+Q3MB3Rwq6VLSZoOL6CGTkGWjI
qLFxt8M5wHX/IsMPMbdxpyp52Bi8HchsJn1kvKzX+cGBwt17x7gsKwvTAJdWhKLaTZZCiRrgMlo/
YXPQn5w776UGoBkmLDUv8j3YVg65Xbn2CLRpkC8Upa20oINbXsG9AuqwsALmyT/M2xYJMQ9M3I65
MetP/9CKamqaZSuLKrJ3p0cSzdmxEn2ircmDeMAUNMs9PYXrzet73RKtLIoxe78IEMdnzPmz3KAJ
3nf9otGFcpEPcZeuyLHgs35vYp2tXz2zGfUZDoi2yIMhg/CwhWJOXKN4m8e02b0RcZ0kfL3/QXAH
anHMMC6uKSo+UXWJcvTYKVpyguYYixJzUfawUrEnzKqZs1tazwmZqIjeHTQ/ZN1MHgr+i98cEsez
/+X3Zrb4NFILvCctT6UWQcJXyMnZolsL1Mlj/ovFO/lsvXwNzojjk+4W9UsKCTMyEyzDa9Qh9Mng
UhnbrScj10vUqA8jF5NTbWEzBnwpI+vGvS9LA4oWcVtpVs60MdlySz1Bak/yc4++QgeFCupu/+HT
xUV3OPc43FCode7khTlLUP5fHaZ1SjHE8XrRtiTIr972ey9q1WC0Nfecj8L4J01tdDlhWbcxsG90
KzsdQUO8e9csXB4LSMKxV5ta7S/moIHdthv8fvDCH4kR2UmFvaVg4nAnphT2WMH95IGQ6xPowv1N
74t+NJr4deufLPOpiPq8tel/EEg1uF0h9ODpawxLDQynw7yeb88FXhmEmY2OdqW5iECb5zKcBWhx
SIHyMOnoZ3NOCywUPkVzN099zO+RnR6+nwyaQ/IloHr9omUJ5/pTXwXhw8d7QXbydXudyor/8Ipp
8o1JcnI2vximMUlSCdVtL9aZWmAJ2A9CApEz9DrcUSwbiDo4LMz1FKQMOlTdsK7DrykbNeXcu6RQ
KSJAFGYbsWazuiFI1BNYh6nHi5I9BIay1HOz5z2G6ufEjJLzkWL0ixTmjcrmpJHDshIOZ/k7am4j
nywr0jX9x8vv8xnr2XSiLyn4OczbbVMTGT70YSrVyN3zHjypQt3tATdcjdDUz810HYQCyJ/ktNgx
37CeSADZzzUqx3kagUZ42ukggnJZBn+mycsFcAGod/FGxqOWB6VBxxtIsFS1QoftU60Eva/CKbU/
bdvBtWxe0//OeLEqJYvO8QFDCQQ2wqil5l+gsG56WajMK2ar+I2ynw+z91Ch9M7c680pK7INkK40
+yDKBVgUaIUqIarruzonl4k8wMpNReVd/hPPc7STK+VE6BqwXJiNzRvaW9FO+VkGmbuKjg8hFOCu
k6IY3Yx9i5DKhybJQ0thpHrZpiwns0S4ZmQi+j/FBVwJ7uWo5vA9gE8m17bEuInAFZrueIsyKnOl
4wzmw9ghDq59Sb0nyhtQmj+Y7U2ir99B14t/94y/YFsbfwAejbuAHKnHvADrcPsckYXzhWxcXr5y
GRYepuSnBZGVVmkcoJmYK+NwMkOilAxTGvD+hYZgGcChgdmYbvGSB3j3j/A5DfNmh8fO9S2w8CpE
0LzQUai+aEu6ZsdBu6SupdB5r2JpnkIarVP94mPFmrIX1wdMa8n2DqYauotZcdrbH4sihgTOlPQO
Jcb8OuMFN0LYQFWvJXr2YTVv7rz+7rooCCYCviebnD5NOcS3A/lJysR/5jmEBl7tLS/w6nkrveZt
0mSVQylP3UMCdUkpoX7rLj2gD0UJR46nIX9by846E5UDRUXYVcsSr03fYcqYjJuqHpMN8KhE33hS
UDo1U4BIwiwwo6i0IuIfovhDHWy+WjZ+eFoKXVj+a6VTYO8/Ic1w85Ml2SBj62lJJwsh3fH8OR8s
isVNKR3lz4LeRgJFvYqCr0t1oCrfwG4No9Vf8g/W3J+gVE2yIIz4R9vyaucLwPjExdPXB9Uvl3t4
shq2oLzEZOnpfiZkgVjs9jMBhDgsqJPjUbt9z9cCas8zdByvwDrbk41c6g1pMT/Outo/+nzGmMET
nGdrwi1lJuhzKbRTWXbURI3PtK1k5bLyJT++OiugHZQs1FWNwGbGHG2/dRMCi3HtAc5ffeT4miLu
hQJpdOn3qA6vOZJgOxa4neYgdjg4RotEhH548XwIXYbbOUy/S/oq4j8HyWPYqwTzN6Ommdcf6bYG
8yLOpWEoccWk5ce5/gRnI6ulDYBkRnoOHxRRsTI4ZzPvLtN8dHUkiAug7S6SpVpMpfc9JSj/803W
tiIPSEM9fQXlu6SF76FiI4yMV0aQqfTlnoCme1NapoKh1xikEj6rGE6kyTddMXt5xjiBG/hD3fOY
vYRs++V/xEo06yGd1sf11nd/Gxp2+vwgF6xCWeI383Js8UAxE+kZsX9pl4h5o65psxVPOAEqhnIE
s/g5UwJdXoLje0J6+YoDue7MLfFls1TIU0uFvQABK5ZUM7nNl+DPk/7wluuF6bw6P+zdLiJTjCKY
rsdha9Ws1u/a600ECy+DYjetXGgQH+xhTBb5p94c0yUIIl3tFCdcNMvbtnIcW9d7sU3TzwSE2yqc
gd94ek3Y/d4PC9GImrhcP58O9HKr9J39ys/wjwcDT9QoSsrIR5KcvTuc+4hTWBmk5ejXVXjOKI9g
voXtOwf9mE+ODVuLhzCcU6TFFt+4eg+oyChsxTQbrbgmf92LE59BQ/nRR0Xrb7NOGC1ruqKOFKjs
L08LYJesoEmCh+mG3+YkwHrxH0SK9ifJwJEX4r7ZqgHfh0RgKiGmBx/TbJF2XH4D6+0uK0ZaCcxk
usnAho0y7YqLYSnSl6Cg4VAVqjautFkktlNHZXhuKr7AxKXGSERDLVsS6ChZVsa786rZTi4pK89F
AX5wNUTDAj+E54WDN1qoTBwM3PfE6+Sp/z2KEJ68lnQYl9Huz5Ac9oEUAqfpvxuZglv/evGi2AYo
+F4pGWzBM8BErv3oE2OBIkcRzCwseCfY81P+mZGIAyaEPtS+gI1S0uEuvqs6OSzFOMqRtU2bTCNc
gwqwUFmnog2Jog2Ct5AqQvaXMMcts/wrbFxV29bCpVQCL0DwgjkqH3n1XLSGFRfW/0CyqjFY0RZW
7vMzi3NhMe77MxvW3Y5DXvOLfwiT4d8GWT67o8YLrQqcUZwNCrcOgzHOZ7+51zSidP/bZgaPFtie
MSaL0IcBcXZCQPrJp8O9hvRGoAjMqCL48La6zcmJWLHmi6ZZrwsqoYwr+WOt54SlAh7pmyKXZkcq
HimOKMyR8nd3QVTYRYHnBPEogmosb4iC8uA17mVqdyFs9xwkvnH0k81qjyvB+E6EBke+lNjpAW3L
qvf+hhYr9ZhvIT54wahte7oALcwPQSnN9SD3Dj8BjxolZ9J3U+VXeWUp7AmfxBaUJV+jLvZoLYsx
jJ500yvwB1BeyZriZAMXtRvBDLFvqaMN/WXEZFmHXZA1/SxZJI4KuT8sCur7UQjH6rbXykT9dUr+
fKHcwFjjo8e7C2Jj6W1guk8CBzB6XhpM8dljxBU8VbphwefyB20tvbrXJAtSdSNuMZxhIJFs3deE
RmKzeWNQQLcU9+YxgaTfD4TJSJ4ROVo8XJH2lwe9+FHOm6ghcG00dmXgKqmroC0oc9iC0jT6/Xha
i755prCK0Vh9vufEfG+SfN3HQYErb+dbtakXmsX6J3CENrJJB7vUMgU7JjbptW+fYdiP1JCN/ID8
0vlK6/HZ+wpXZinSD0bbWkZj0MkNhmVSsmmQMbRIHcJz24zhuQI1tFCB7OZxcbgbQ/222MjzJwmN
tl2r4RSk93pyGSBRJCK0kwF8MhWyGv1ng+xJa9WAfRADBrAg0LRnn5+/6kCVR0gPzU1clRrEeT/Y
j0fi84e2yL6ra/c2u8hc4nNTD34lwx0Os8hyL/CcsYmln+g/xt55w/ZDds2fKR1fj+CM4Q2xOhj4
onbWqTH7LUXXtCGjLuNmw+GZYBdq9bgJH6zKlnA7YOHkJnbD1v2FVyo1EsK0IY03fOK3fIXpPnSb
WIhic7OzFLSa5aYKZFQ58GCDSxD+/KUoJbheiF15FEw0YZ6i5+4zlT8Ax++82cFHWvWeKqeWVknt
YLmxqHOB+ozsdPbfKHsUlnFoewWt7vXPIUhevUdDwloMvriEDPJCUKICIuvnP/dnIkKjWerXYfEs
dsCo+4g/75sftQ2hqNJkcLevDgn00Kc1eXg2XW4Cr4T/MFxIOneZL23utQ/7BPqTFqfmsKeFOnhe
7inukDc1uom7T1DimKGwNhw9gWsimkjBsw6gR+Z9t6Af41muFiVCdz5nN8Y+YLwuaaZUYZDeyGsT
KXO6vQ68pEVXZLEY5gHMqJY3YknD9eQsK0fXCMtJyEreDgSjnT9XESPm0Mv5GfXmVJ7CANXh5EXA
8OSy2hfCYs1s07soZedhy5PI9QwDBborNXOWTruFpl8PqkI+1d6BKYiliqiYz7R2rQO5BVMBMXFE
FsxznBCCoJEX9783h/ybijwmWsA2qS9T6eSIpQnzOT86GNFSvKG5aVUyTBrkBqll6tPr34oPWLAQ
XGj/FlXYXXYfNcwFNfJxsB8o99unn9hgH8CqMoH38vPAi98VbMAnpd3L2FKtV3RB2h4D5U5LyN7V
Ajbrou3wUov/lL8xzmWU+a+/Q5cFFWYpf1X2CbD0bVgAaE3VHjuVgDp6fg3mVKG5At9khdQPBmTf
QGBrFw/PEwN4nUDM18K6zBtFuXmdI3abh2677s142tvEeEej0tKllK0ILiaRRaSd7kr8EpjtwF9l
lrGARLpuq9Obq1WWDbaDEXa22m5wpWTGLEw3HmTnjt2jgY+mhQCvLpwjqlHqnNwqBaazhc32KrAI
GLQJqtxCMEDvkJ34rLyWu38oheOj/luN79r6Nqh5VdNZkQRYfXa4UoKz17+Y7kO9FtzGNKAM7UHf
Lw1V2pcJCdnb0fAuP2kxfvMJK9wVNsYa8SYDAP4Ga24/JQF93G+AMBPgY8JXQrCUxtJiFxg6c6Sy
C9OtWD/Qx5wqgI5BQ5HdYjiBHuzcMXXxjxegm5H3NlwppoyA1mGsreALDNT8nsgPoO/o5hPU1VL1
mJ4erFtalECtCUC2TMBzAPcV/0vk5mQws6tdQYb557Gqg2grlzB4OWVYDqk4m5awI7ijovraz8CN
q8CF5mP+FeQ6K+sO0uKb/D3iN6yKFzGuO7iZ/lyJFvzlbJktSzmwXSkj20vqDATOql0Zk1gu0/W3
fk6lxiARJCpawfdcPn+0AYonRfPnAQQR9vyqwDBJcyvp8+cwk8vA4RwRkHgUJegW1YAMv69SSwu9
CrQfWKWR3J8qc6muNxle3dVRqZaUmznyqB9LQdaIXwCmISam4986MLmEg/FsG7i8Lc2m8VMYnIUB
lcGNfSoN1cfT9qx57LkJB4RTdC9aaGXaWczJl9D3Y0QgukxTrlTwznPrmhqCqjJNIT8JuHfO0nMh
ZZQcDW6P6PxujXRXpctzsEIq0vMnQTcpyGdi7hoRne1W80t5HvUfv60p6DM/mTp7bn8pe5YttI1J
yNMycDeylUneUWN6/iWKoOpolD9LaVEPyCr7Au6UPtEyeRKFgaZG0mPcFXZt02pH0SFR2dhkimR2
wia++Mxi1pTfD3mGTnjQolr7fic0hRSrKf2swZIa+/AheIZqpep93oy+Ex7DHKLDqqL0YBZ/SZEm
UUyg2m+9oXsFmk7AXQPRmrdb36dreg1x2utaYRn+Gz1CxBAq6hXozo1yZJL/d7CKS4pgz3+T25Wr
yFkTN4DRXuK+GLcw7SzMESHND+mTIFYrZ4pAuBB5US/FlkCk8/n9DJEijNPbR11rYFnd2fzSDGce
WgNctwJLAT6+hXohMIGRBANSqaZaGprKFupxtBhZByrX/C3adr8t87mUKFLvbEkBvJykvd44OAva
tUmMmyyZyp4qY1LkKzbVQVYyLGK86Cxh5EV2MGD6nMgO5/GihQIQ5i8mDKBuLgF9MVoRGEUd1wly
XyWQCEcCQJyXorlU8M55I/qEcdU5bzLBImApdDC9bW1Ib9t9QKAiDZMS1/UwwGM+Ma0l7g94N8Zz
yK1U3yXxWSsPLInwXV1ffRs0a3ZvXdW4YOnRXT5Til4G93LZPdmqqCIx4ZesG6fYKym3L+Ue7P4a
Jui+ZfiAQ2TLa8meLKYJW5kVqLFIPbN+Fur9MjlfVaKTT+6izU0R8B9l3QKPV50rLgc/3GICH8w1
KY6sF/p3uo/Zx/CmBpb/Ytm8PqyNl9mX14I2/petMbMvTs/mr8QQNuOj4ridPd1Dj6WtkF3VNAnN
pbTeTv/oh0QmCckjPcgNzSVX6ndd6EFi76bHIfiKN0Xglbcc6eSWg2IISUIOzF+fJx7Nt38PxurJ
dbOQMLYFTSP8FioFSttMT0OI3emi00VodxCH/DXwK21mbApdma2CQDcD5TDPXY+gBhRpADFBi1Y8
6/5cnplMSavh9at0RYgO8wMY0BwMUHdVJzdFfaoMm/kWGEVcFTcjtRgNc/iLWh2m7RkxvwYXRl+n
Ra0Ag3lPJAm0ngdhqsUyMEcMGwRph+jsXBFTt5+i/DYLAJVkGAEDszKKTv6RZ1VJrgnoVA2GFlGd
+8+TTNDfSdv01WabDfqGje5rmmDDDvNSxTMnwFBVa5O2u4JzFPeng1yp1euu3YjVKfKBPqPVA385
wLy0T9OGLTxVE3YvpL6L7MLmM5/zbexkf+npudlojlqdxqWUjds9Grs4Tq0D0VoxrrwgTgT+B32y
yzE8YHVqDADrdMfq5jB4Hl+DEjUNh6N4b+R/Fc4C/T3gb1GUvFJg0X5VhRwKKKEASvh28mF72ZCa
ueasRuT8bWJEEJetvxHqn4puwuaheT42El+rmdicm/s3fKVC9vyHPN36+wJHNQCWQL24cY/1FQs5
EZUa0KjEtAyC1Eqiw+PyLXwCwuuQZ6srsPTuZapkt5G5xy5hEZxkXRJz2ggFMLxIbYdaR3jaipWX
ezjj/GeREw9nlw5K//bIs798OK5v1l9KSkwxeq+Wk1k7GEeKH6rz8zcXPUie3nzXKXFwhat9GR8p
/NOYzHnmpp/i3XsV3205MvRTvdXz8NCoSxwC1Yx3QcfDogAd7lxe6tYJ+GMOHy0uvcvjuO6Obj4D
Wysv2Nc3FpdyuhjNzhyDqrl+cz+iVjFjDCLIaTT6rfX8Kk2PLUx/XpKW3wzeRJj89PXo4nF9g3oZ
cCeOMlCr7TiIq/nz50aMSoDrQGhsIw+QpV8QzovcdjzIWZBPgLRTtvqXmEwR0IbqpN0buKEILiTb
EWvMImYv6D+6c2cf9gRwcMZypUQze5QUGft62CRk7TPRC7f9woGgkWHATz/6ZX/LvWX5cSLqAIpK
JXa1U9LUwLuSPFPSwxub1zqqzQUwJma7Mmwf3pYk2CyhHxdFSKrqU+MMliorKvWxG/z2SDcHGrG/
3bTuYxldw8hU3/p/hXIn4psaY/P76KSnnz59JaHehWSLgvQ5m2048FVX6LqYyENLTr9PkvVXujbF
MYLBt9VblXBDxylnGJxc+wrGnwk8ajFuIw3WGy0HdfqVMYV/sqWP8RocsdbuHlIp9bmeuHwkelEp
2FGdlER5F9R3YWXNWwlq/pAJwcj0DGlaDJGi1Mgs7UUw8rrzpkc9Wbvc3VenzsA1QTcAhsNWPJYK
n3BzTGFNJ14v+WbL0mhd6liOhld0/9y9CvSuHz/Cg2QjqRRKvcQM+33QDuY81d86x9SyUG6GK8+7
k9VSFXfOPDHKqxxTxE5nTKHDkOXogxmKgkox+/umDFXJCs9LKx1oUCrMXKFkFm4yjzopb8q7kJwC
oAwVStvL1Cvnst063ppTbSQ5RVrxkZRhpy8DVoJwvg38vKTUKhP31t5P2zJc35aJi5EdlN5hNx5D
U2EMAcONB8q3DhagI2+k0x85YN3CeQT5+ik0fYPSj6syTzCayxo3Sc41v+HiWo4LFGNlajuUnuK6
Hcx9k1Xybt2/7dz13J6IsrllTDeAD8cyv4dyi8+Ffsh6KhMXFhNGhMlgoW9rDoUR+x+2wm3uwQbT
dR8OJm3GSDdi0EKJ/fM/jGZ9uSMSd9SqJDjtE8a1aZrqmL/MnbN4CmwIojsWVtcjsiIUnxod2ArD
oEcBkbnGjOBLpLTmZe0iZvn6bC9r5T7fb57OEjyf/i8f4mQ60OPB0Lce7nd3iQvUF+u8MiVHVjXX
aa70daA04kZTzTBwfolCgjspQ8OsJK7lbsvZLDrP/omCrIrNawPJpuS8zrtio3kB2ZRhWlg43IIY
tNmFIKEPgOn8VEyl8c5j+qYI83vCVM3EOz/vX81SJBSc8Afa3P225uonVB26woBV0NEepIi6+766
aVPEqczaYW8sxZhCmg4ggW+aUC2oEHX5RSyKi9HSKEmBTJ4q03xxjgxfgfFFl9hgDR34Hg5Cv40R
V9G1LbL2+Dljoe5C8gOCkzjapJL6vWvhfIcTF1BiBGP0gEhR5hNS+/AH6U8jiqSVDB1jeRA+NaSW
6WVfzJWKZWxwoCQunElQt61hrb8oxH7UlwI6s+GSFMFhzC8RMTPddCgQO4Gg93keYvvvNUTMzqpO
6bcfs/WK+s9oCbJVdbJnEshPKbiTlzMsPZ1WeWVSmd88m7RVdOrNdH7Z6R5ubXLmcA7PedCBhNKe
ONcLS8vH9jTbhjm+OIbb3nYEDvdgftS9BrOhZ8Qj1KKNBLPr1gc52Hh/qwMrUMh0gFrvCpXZi+Ol
yA5RDBw2NCybXgKABFReWsdX+uNz+2KNUV+t3y+2qGTT3e4OKoWhoYH3BRUC3hHu7Bkfix1vWBA0
nbheyPwyt+15MzP8AqKTL4clSjc9hOPq0o8Jx6HMh8Xk99rHZ5r4q4rXKd02gp+XBOM28g9dv4In
zKoBGY3Y7qN0LRfmnYSwCJ457bissWUbUKm1945wlm6bQSJycv7UIeAKztuoiJ2aOko14xjW6gPo
TKE0qCPSPP2sxW5xa8ItfMcDdIhRta0zWM8xjcuHVNEPSqlcQBww6Hcp2A+eGOxbu1liN8Ik8gBp
Pb6pS1Tg1rvNQuJtfc5m/vcPLy2SVKSFMUxc/vW8IdoER1MoDcr4ppVzgvHezkeWeTl6ChzsHNfN
gtOLgn4OYQQI6l2bACCgJMRzSdtfv5uOaMZ98wSk6peN9F+cPpybB6QL2P8q2ja56bTDU3wNndqZ
Ix5eiZEyWOqX8QkwcMWkQkqo9pYU3x1zX6Z97z4Dkfvc6HK7WjTqzuYT4pS9REu1K2mzjmW/lm8P
EOmseDG4haCMVoi8/WV+7+SuZwV9fgGXCAkzJYpeZuOkd569w6AjOI8APGj5XWIglRrltR7/+ndU
28aB4CgecBeWHam8VbkjtrHWH5Bf+nx0tClXtcN/SBNdYNnPZ+kC7M4OzTBnKgTHZHOKBRk1jc8v
TjiqLv2Zlf+fobLgAEtx0uwWYMD5lTVA8bZX2RpMEw6fndEIqjzhCpaxCjMcNXCjhoRmnzWCXaeL
Hrye1zfKYq65fGIUcyr/XG9lsImVtaBx+LysmASDs/rLf9gjJozwbQVvmwy8CUqmz4dWQ4rGJIC2
CtXJOXc5fywvqaEwFVd8XyFHsLZJ7Ga92K+RMFQ8lGh19EQl4bKZCe4ErG+w2LG8/P2xS8UhvwZE
FIjDAI8jlNZ/mBCvgtFhNJI8xfEhBG9jEFY13GzZshiHQYCdTJ8k2It6ilpDJ/bGfpR/iJvsC3Tx
3hcaP/OEGxbRDtSro9xwE2TJBPXh/4HrlJskCGz/8Qm9tetOquelASWvYZ1XT07nv4aZIi2/bvY5
FiIb3+dwVCF80Js3YGgeqz/5vFJaw+tp5nOxfiMBxChtd28usFO/hsuytLW3dE36/RXVgVMtgz8V
+pAbyItQq/7S9vTpnLC7Dd48az2oH96aDO7e0gtjUE1Zu6uAm0ftfpc5ydAMhCtRblgmXcn2YtDu
fBuGjdnUZ+qZ7wk2dnc2gV8OZJUv/zb+V4CpBAfD/TmV4Q9bBLAH5c/GPvd0sIHDeocJ12JGwoGv
zhy1WGyMj0Me2lvLwu0lPSUR0U6u1Mzuj7QEWGYwVuCPnaKDM/1qyEH4DJbg50JD7HkBQcupxEL6
B+FAOj1jjXzSdVtCnza3e8vttFE5Z9icRx/0bz50/Fo34MzaSA4YtER5gPsYVykeEAnkkKqqemQG
kP/HxEJbF2gdNhS1Cdk6ngvkCOl0yK13maOusZBpXLlubWQ1IiVnYAU5g5AMBBBhbIN0zIQPxmgt
sB+tlvmlBRZ1x6lbNOnVyzBIy6rgIME+HQdVOb2OMtH0GihAeCCsPZKPWM8z8natanP3hDWy2pRT
+DQdZ/wD+upTrdNJRUjVkYAO3tEPATVT7168oU3O0YWcY2pDc2j0DFnvJ2bAOo187U7oxUE+B1wt
PnZCboxnJDI2x/k3lpOGnL/kPRHHFPa+PeB0NY7EhwqW3GyQKXXf+zxlmpn6dKSy5O5mdfbhOauZ
YeIxdCrG/LiM/m74/iEi3UJqmz17P78KgNBOyQ8iBWM5XjjThy/HxC4zSH8u1nrA5kSwE3U554vf
7YV1rO+2azdFt0b5O3KEe/bd7JlfQ1o//v88IiTC7p3c/qdtn0INGGvWwOD9CYZlgmBFMm+SL/Bi
br0CYdvYpCn6NR+3HbEh50o4q2vg04cFkorQ91TIHErLVI1imzrziLuq83tRuOyzSxyAEt1URUaw
aDmtyyTLmhSe6Do+8fp5oSdnafBu4Rynwz26Og0LWqSj2ITEW36KmDK5nPjfbybmewcfqwv0IiED
KGZroD/i/oXcvZELmQz43kDTkbBbzFYI6B2hdfshqqAo3zgBfjL6w3VJgGNWyqkEEpYlgpT9sVxb
h64asn40qJVkG8ACIUD1Ipc3OQkD1P5ou2Mh3flIu7OwQpCxi8hN7asGVHdsYqP14/kD9je47Qil
GtF2KatSqj8AS1m79VCesFlRxXb36+vvDpKGnA7hmAgdv8hflVNAipK6Yq/KTfcAKB4G5KL0cZ98
qJDTEpre0e/Lj22+pr7W7BVFVlCzFkSxGBvjotm/dQG2S5+h6SC9kUK59IWGijGCeT0MnvXQ73uD
yCDJg31IkEIQcNF3L2AOCvqVmBqZqav/s1j7JlaSGCUPqgrkpRRBEDrvrHXN23umwKEiDwgvRY6t
ERdb8VzzTM+FC0WCT/XOlzxj3CYaXcyUGIwS0oornMMUUt5zQ6IgH1zpp6wKpVOAv/00FCGoqScE
YSi+r7wDrIXURtDwiLuHh2wNNmTl8Gi8tJXbj8c/amQIaGdwAJJmajZMrFKxcNXxuwxiYzyaVbkQ
I7fe3EdABbc63tEbKXcTtF89nUlI7b9wN2ShKByVfrNJ4NuOJpNDC6+06wERo4f+S1tAO3ziAKXr
vD50p+0iwTxWHMR78Pik4rLufpcl6AfigYueAuqtRels2ozVMoYWtnOKR4LEoydtj6e7QL/ewbvq
Q60DvJaW1/opck4k3dn3gXdrFmfVhP7yk7hBCSRIztlKI1BKr+yKl4PDgw6BGWGbBcSvZE2fpviQ
UDQuHTHIYt3604akbXiBbhfb2yFxUSOj0nETFmUKoDx/fa0MdBPEQ0iWYAqcDwrrLaT94IHh1Ggu
8F75YY7/kkpHCdUmpM4zidWwcjK2wGgoy6oQmFr2uZ53L1PCxMTp9qUg0g2r4817NMc5/6C9Mv6W
cQgE65XHVPePA7N5pDpmtNrYt3c7IH1kBIrqj3ABLcu6WdRux9+1AW4PgoKhNNrQEiG9nbxjIrot
BbFR7ZRR1Y0f5h6Cv15/eHZmq8v2qB+Z/CBZEgRRIcdn6t3g2S95bEE1kzQGbtURR1p1r6V9gyKM
zn9co0yQO3VmU21GCo/OkofAkH94ma+q/QH0Y88G3EvtdvZ/NN+TEYFvHoQeWQ0VrdK5g3kta4jU
CY8ucR6YmlyV36XNAtM/7F1sS1l5K2KHB+PypIp1c6DXHrT5tXELMPDbznRxrD0h/ihcjYaHfmpI
eK/Z4C6+60ms7DoXDuKe8cjdkAoQRRyyxJEJXpK4HcPxu4DM/PLIdzWDYRvA5kGQIvWFLlh6q9qI
wD6rLzJsuLMLl7vHH/jRJ06s1gxCYKSxeKmMNv/iIK30i2/jAibWDYs5MSz44dynG5OmuMP7G5Hn
n9uvZ7Snq4KDF4kgXSoq274GL/bsgZyN883xd6GTgi3pHhymb9yf1qdstAcsV0gJ66Bxj4JbMvuh
RCofHCkd8VzZr7oFq9KpuIB0J5rn04fNh1BiVtpcz6mKM1ye5sxNtt8G39fGxLu450UYGPPCmwdD
5BzeQB44qiEnAtmgc+coUHU39oxmZuIwQ51DgbM5Zf6Uou0wCs53cVqc8/GTQ2bWB6SMZ1zTvcDi
rgbfUCYyna8rS1sf3QDszUyLe9Jm95N+2UdqrjghnBSsXzRgAg/bVfrgVrElfGRAYKsvPoU6L1jj
8JFv/pt02loRM4KMoH+obDaGCoGRAHZ7Ho1qnskxJbfxoJEGpkQHKCNCPfaXA9C6/Z9cNAwU949N
/KFDDVP+5+V7XGzuEPhrKjbkD/YSX5pDCsxSYHriysuW7PbLJojRFe53qbZbGzziSqZ0/CECXzIT
1nVVga39XzN04whGqNC9wz0QrYq8bBYHN7sf2u1mKiGkYR5XQ+kZkO30YL4Drj4dzjGT8cfJhNSL
axZp91SnmH6wzu9U4xaS2ujStnba9mtLJoH+GDBRGSSVaxAJJDx64KYSwg5uEJW3I3D92HBFJZJ3
3iwP1M09xoPzFhPBbh31+li5EIsfSXboAULsp01CFDPjz1GL0BNMC6ZTrCdc2J4XcgdlYOuvN9SE
izjKhl81OQbLo2uw+n26H/xpP1G/BJun8XHk/RzAC71iI9pUxG/zLLNVNWaqz3SMOIwdzWyAIOmE
azjL4go6WkhEQ50Yru67nmyPXY+eeGOS9rJ4I8Inz2MLLSWvKjP/RBno1hJttoJnjk9ZHRa3NPWL
s7z+Nov8b2X9lg9bNRgAlVjeYxDpu3vUEBe/8ISCkUQeoS/Msh0DbbSCuXBwA7l2iI0YAOpkGOVz
1Ru4giVVY58DDMlhMB3d5Vml33ENRb5vHBlZA1x3UCzpaJIfLUCxh17sULcnWX1Ob6mL9HPTOgfx
EVC9FsYCFLLytCWOlQL6uMX4l34gtV0ZOpYvJMxo7DLH/SUt5uPF3gahAcFxrKJFGi7tSPvaxpjK
9yEF3C16zJt+BAG0DIJMbmge1VMP0OeO92UhYj0z0a/0Fa/otGUhxEz9pjsxuzdf7/3gGTn9kW7/
Pdz8GyTHfOsG0OqQZRGPle4OocLJPywQ2DqtvF6es8u+FPvyA7iB9D7kf9XFE0cTXLjn5/Wcmsr/
VJrgFq5xlA8hLg8qCBBmmyRRFOePqSKz+M8NH6gDkT/O/4FJ2znGsmq1q5mtw3H4oGSEV1kGBG3m
WgWw2vb22nxV/I9wyt4s8OW9AbgHCbu5J5LD5B6etcAkpnyHdxNuFZ+CYITnxWbBq1mVmpyeYVsk
f4xC4NXWodHFoo53a+9j2AhTByU/8KBcaN+0NYMXiOWK7gnRSPoulakK84xZfDtMmtGQ/I1nATiW
kA+031u20GukhTzo+EiKXa354Lg8RXEDmj78AjU3zjdxkd6Pc4EfXSK1h/uNR/lvh9u3j1+GhR97
03hFZRjabllvEJjMUmr8BIlkt06znvvjNDlydEzcg1ggk/QQ9D+NoyFxmXZ+BQzI0QWu6h6ihdfN
ZtRGip3XIWp2wtt4WRfF05HPDA/3lMr1MUkk38cwI26VT4ZKfpJqjTfVvbFDqy4UrIPK53v1swEZ
9P33dCbM/N9iHQAHkoqUfr4PMIvPgpa6rBtSGUwFFjZutw5y4uMDya4WrMe0Luw/YqD0XsI/V7Jl
fMussHrh8nz0ggp6u7D8c/hAQOQBHrS1PEvEleUzhOUEt8DifaNFi4SS2K9OfiyI9xHM9EkT6Kk7
xFc3bCmMrsP0PTOW47dK2xuy4+uTYpPTmspqa2b+g85rM00MeFTG6OPRPCnLxjGT+T0pQFPWU3N2
7v/J6+kBMdUqdJni5F2pDPQepz/kZrozT54zCF+dw00cVpfcn+C6sFGB5Rr06SPK4xzLWdtwKXdE
brvogqxssQZUksEsBx6sKynLvu9eKECcxMpM2wH33sy6abFnIa3iQXGtMgCi4UhIm/MznYWC1Fdy
YviNRzLfoN/w0MOS0+uelgMdLPDkon6WHmSFGorvEthlOJ145/LUqt7ihjZjqX4e7/OpZAfEjYL1
xlUquZChUusdTvd3sRcfDad6iO2T6EM4MrEM1yBJh13I5H1UkSZzPs/CdjuXEqeFSJ50Jnhfe0YH
UOTuYKtoyASOcYRzMdRMgC0qoMlVxEEqe2qLuMYfiVzss8FlmKmxJbfBe09zp+XNHj9+GfSXaOAW
eocnDHgLpnIa/c8mqZGoL3jutQRcE6q55OhtgxXh5WLAiTwi8jApwL82LWedMRwEzbrk5WxTy/0s
Ygi5apj9uojfQM68c9TcjQHrdB5DuQAFpCdyZMcFLMgylkA5pjk2TRZ1VRwcyHMri/Oa16k98qos
shDm2FXoVyduTRo1WMo7I4BwjPyV9045rCrxiE18wdWWXa0bSTSdfJQSVQtJsxaTqYz3wxUQUSXp
BH4fdJGBEX+BWLcEcQEGIOeOeRB6JTC9IJyl6SO1clxecqjfSZ0PTJZf2fvZgPOw/NpO82qahuNn
Hg3qxH65o0PNXmY6ch6PhRixHpycd2ArMB9ouLl0RUHuKkGcaBmtS3XoPDV1YtumQ8R/GtsmnrMC
Dnu0xe8BI+98ABB2OY4J8UXousW/tPXPzdXB0SmADq00F9fSRp92FixbY7nxDFd4bmZBDheTSxmP
3KTRmxTsAuHyh979bdKeB822NCizHxRs+j0SvzyuVJj2qLt8xo7bSTlkl5D0vLuWkZJ3S1DO3GMF
MhmzLTUBNcdtKEhZ3iZZyFGSHSun4dFatkra8ja8GkmXZ5DzZESmSqtnHAI1IvFcw8L/gN4TcW8u
JP0Z5ne/0p/OScgxrGSgTmPp83C+h0mzQYHZRG8/dPE+zyJSitGJl5kdJzJZHhr8ppZE6PwoR4PP
6TMhKp5/WikhLlMIJWsz8KtaTv2yTVMF8TFnUcrAlKuFY+wAZiLt5xbJDu4wf78OeKW/OmfFWyoV
EIXDf0ihXPPyq7cd3D0t91f0bqD4IPt0lA5vJ8oGRRIK+wU5fG4iSJ70DXCbTX77h85MC7fztliv
JHjOhtRzhEJjgqwz5ndL7vdOLGr5JVWP579Kvwiix7ODf9pMV50QMrk+ZBB94lV56QbdCK0YyFpi
aifshfOrk2NiuB6pvYF0sC1taQy8v9eZY1o1oVCl+xXEZM+4+TJ9jX6IfpgjZ6pDefatDDeWI+FF
TTPm8ukGTlV8R850a9jvSMt/zZlxAw9UTW7WUgZdNosfUYoS/36oaN9FJLzMtwo632TyqFZymDy7
9YKOB9htZPoZaNQCfXWSnWop+u53W6aBBTz2UmWtgcjNMI8e3lu016EEIan1DZyhHtX23AA9Dd9+
6qsW4+9U+KQKE39VFly1uLBfnGGDdnFI44udf33Wh8dfFQm4Lx6/T6aFeDKQVwWlUjihbdYfAG5w
XeTf0W719cVyPUcSh6UXlB5i6jvYhsI7CgFZ/oFjapygeRvXm3JE7cqRGGXkobT2+iUZCdZZVgK8
ugu8oajcnlEQ0By/zS65T26aH1miCc7ShxI4fHhk8eYBfkYxZeZS/dYi0gPeZ3PMhsccG1RX00ZM
n20AHm0iK5csKjAfCvLBOij4wYtiIdqi0zSiIacd1ZYTNgwwQul7n5sjKeT4kf4wNcy50no+0YaV
8V+AkP4YX5B8Pe2A4F+jphjuYHCSjEWecFu51t9DqbhfZ9TDcteF4+AyzShf/7jyuJLC5PqRv/QA
8jgE/ADyonZ1vbXSj25ZRc1XNhviWLch5iVNmudT/P0bETatzcYUPjl3dBa5ok9kSWAigNckUChf
ehBwGNb5MamWK82CuX3Tac1xpl13FI+WhBewNFlyPgncux8w9fgP+txnIHQUtsPg7kohAruYKRTH
RcbJGL7lXNpsdtVh8K55NooLpm45UF6lZG8z8qHXUqCmzYc2hlaI6woB+8SZweB1aoHbY+2pfJGe
jmz/qgZ8VQbvBlWqHIuMjmUmoCVRl8vWsFNFT8xeKoZMs+pUOj4HmDslITrgmgVXCVvFOOou2CDu
OCqqQKMFQLLCoF1n5bUMxJ8ZKfWH7zOMMbGTaQcyvwyoavTallUiqHB5QZMcotiWc+VHJHE8cv1d
10dgYjaLFYVJWw9PV5kbZPMoUub7piKMXsmKC/fsUNh8uzZ7Hr5iCWuGqOoPJwdIPwgeo+HIoaR0
djuwdsXaA1uzQzzgGgh4mXoCZuQ93mAjRw/ohHNjAoyI0dsT2ubkxRnSTG7fHsKOwa5irovC7TEd
H2FmQKTFBz17/3RhmpkUrSE0kWkajQTFRPblOvcOagzlHMmMFWmwfYkiyzt83PQ0pzDe3QVy36W8
RU+mag+7yLY6Mpk+vP71JzDlC1Vs/b0Ak/PtOFtXTz0Na0iLmA6P2Azt3CBuF7zcKhi9mIyOdHm2
K//vazbp+ZTFe1BeeOUxnXzZ8SCgzwNlGRuXcrBiGzdOCRqwTZrZ4w2xPUC8U2ntI99A+NHqQiUw
0ZtiXr8FmeQemv/VijXWngVMo+tdUEiS/rjzSgOFoESGyx9t08h9rwVGZ06lp5zZOkkj6lTFPnck
nXiThK8QYR2gljmwSfV/+7zNX/tLZamVGwjaG5h2dLOYYqVMZtcxia8r1Rk7ueEyzg95T4IkF+TC
Qu/QoFuC4G8YZuvTACCK/9wEN3D5pXBoeN64Jlk+d2zjSRybb0jjC0cOG1+PbYpeqsOs/1Fh4noa
/CnZ9TOHPnB8MbBHAqsgffIyrpYz0SFRdLI+ZxYLbiFDGpxKC2Kk6vVZi1Ue1ASUjK1yiEAZKKFb
NyeAPYR0WHvGJsEsSfyglKU+3Iu6R+YyzHQ/kTBmF20lKR2LaLBKhKkCq9bzl9rr0TDOEgx6RH7k
4iQ4EdpJeZb6GvjCcaDBzbfuHn/aKf1NIbFk0nuXU8BbAVN0NkClhyTiegFN7ilYBPY1EplGwXN0
cu3/91YWnqlMCbsOdhKLb6ZxQ98vXGyrAPwz3K/+Gsh40bn3AaQdAtrOX/FpGdZrmTylCoDjzMVO
s5yCtMIKmxcg+FO+rNPhC6zui09mCltKWq7iRnH9YikGJlvjSX4ek+I1VKCduQ2jzIIn9iIX1ktq
CPHE2ZDAPUfVMcIcvadu4YXBg2cRfyXnUzTSJgNGBH9M2TRlYAX/w6zYYcyut2wGjuT/UXb7t9hh
oOOdiQ9EGi5IunvYuVppiq0Qcz83iKJxwx9cbzrNO2tzNsL9l/EWKuMgCHDMt8yNarrUZ3IKvJvl
4zFUrdzyIJopahbOXxp+ciOktBBXjJR5BirKS9HG/GbC/tMVz/o/J6zZUB+hf2iEGb9SWmKmrD4z
9zySXi4IEDSwRUCWyVWRZjtsuPkQXR1JFTmWhErACEhHo+mlfBj5acCRXhc5ASkGRjG9D+NHrpRY
pQ43iEk0aEJgA8Aa58Eh+O66xJ/TTtNnk58JL5hv7VBZkrWPVEEp858hX2hlL5zpa/PPoJTrDdAS
6saQvUVDV8JAoE9fZdtiumjA1pDaF/aw3PjxQDIApb04Loqiu8Hw1OTfGpPpXsCJjfzDygpevT8j
U1ST7XDHsvoO15Ll8rKQxk+U/4BgsJeVjgdSjuTaApmK7GsIfw/LVAgRnFhzq1UuAr5t5pXf1aKe
GHvVVw6KQ6bMOIY82BEXJfftXI41MXPm9v94o0uGe6iBkN+O+8xHU6iaU0eKA5VR9ZwCdz0/ffH6
bCf+t7+Z6bkIghaWcqcnAYcX73LJa1AAAe6arZYMtLZLjiDw5y5t7Yn068vVJU6nKPDJ4yJhVg4d
Nx8FTUAq3CLHMirwiiOO9N1CnwmW8jL7ooJ5IFrCayMTeMXMvgbtAocNwVpW7hlF5N1COGNk5WbF
CvmrVqoT51AfPE4zC64uTZV5cZ3mXtJAylGQ+39MkfGyEmsiDEYdQi82vehnUAA5gpvFu8Z8PN5F
eh5LzW8H4ZanFX8jb1HJJtlW50lMyc4O5+i/xUp56GX19kgiqCmeXoc9zVoJrHKcER2wAbO8N8Wy
r+oeawI2VFkspWwuOe1+1M1QE3FX9CTDjCtWp3wKYYj0fOo+caql5MGug/f6tK6ojc/sUAgSbH3K
B7dipt4jQ4qqU4IR37cBFmx7TyC2icfBazRnTcnGw3S8onsBzJ1tJqPcIRB23ms6e3+G8YbDFTcP
f8rk/oMVW1KxviirZbUst3exNZBWQZY5uyIg0pvYe+LWG25RYll0JqCdThjS4uEb98AcnjCl+bMW
t7IzNmpCTsO8I6LrUvW9d6TN3NpoW2dCAJnCE0/Lo4RAcPugIxvySew3yuh4NI9FCZTPFOLg6kwR
J4a1Q5XUjUX8Q68jN9PhrNtHA79IY6emu/5idmzZ1gSx74/tVWvQvGsbGXLnkmJ3MNLtDVoQ7ePQ
anVroK4I5Y5NXYVvljLJBLmvlmQfipPzJNWbZFrsJJE3qDO7Erd6bRf4o9TTEJqquPG0SJ+JhQhK
HhJqD7HCw+CkbeZeIeZueHneEkmW57OGeOy1TgVMA/GV5vdw1NQUEEY555bVPJcMG5jpGEGTf8vN
Ryf1CLcD1C8TIpt2K9sN0ZIho10+iTjpM0pbCUucvIIq1/Ykk+czKL1R0CjqtQaQ2Kxt3H+N4hgc
fsbOu2YTlwR/PdCN9Xm+JfAMykhJMEN7aFXNC6/QOi2+lF6ClHT6e5cj2axEMxtsuE+gH7mrx2AR
G7RPq3wlEAuYMpIb6paqjVom2MLcllFyZInqedBil0dUA8TkMvPoIZJZY+zEPj3+q3c7rb+OCPj4
aImh0I7/Qf2v5HmuC9HHUKm7/V5cbp1kP7g8HkZN6WXV+Yr48Thbl9xC3nuqGyLKYhuJ841QPQkx
+DLQXYgeCWwBclP2sErgODcu+J6hmDhxus+OSwPHnG/fCaAG3j1pUmwIIFRgzlLDCC/Y0ueOusnV
AEqLW2EJJtR806dWxaF+9hIe+RQ4dOOfhWMymputwvB011SPxX1OndxU/Wl4yZtPi1mp4DEdxNzF
rgNI60dDHAsVWsXOgDu6zIFys4m2miFfTFf1fyJS/0pMB8P9uAEP77qKH5FoUSImlH2UqkxPLjwI
Tba4TyDfULcshSPNfqlNDnBmfYo59cDIg3aD6mo4AxlwyAWLJ8vQQJH2XRcsPRoaBjU/7T8x1c94
N77erIiO6Gpg9d+d7VVrKb3O/wjHAnLFVGOVQK21XzlY5vspqr0U5P18XHjLrzOPGDh46AAN1Dhn
8IQ462LWkbHzZkMaVLpS5/AFZiusbPkDWN/i8gHqLN0OCptH8PclFcbKM+zyjk+vCX+qJ290T501
F3LSCoshTf8XCreFziG5/lWYAGbvx7lUPH+nfhUijqVbC72YKksoXJHECf3mW+fT5TmDS0vpdy5X
I02Lc9ukkfdpSk4ffhP7htamc/8McMr/n0ZhjnNQQN7bbChlp5TT3m+iRqNaqpkHeTmzauHITY1J
GJX30eK0k0+VMHVfvKwk/UNtmKMUU1vaqjxDghxgAyPAmUBZn0pAOdTZKYY/a6usk7E+4nQh4s/p
3l/IFsmBbfOjQOKEZROFT3CoRQ3VpMsfTqQ/Yq2m8ooQB7rYrnPlwjFPbY0PWWokdj/8djdBmLNh
vxhLQLcUVQ0qmIJtbuESWTXn93gmwqC2eloCnUD8/dHg8/pIR/9ad2LAsV/hRaO4JNYT5gWmQHj0
IWJjA8hYPFaJP83D9M3LQP13WX+9leBGZNZZ2UmXd8/KQev8bUrp0TZVmt+JJD6LL8gT9qClI4nt
g9GYRURumkkuHwXnVdCFhhhDo1ftre6tS0jgoEZKnxDBEz6v5Fhl3RIOzVv0ZwFDSvlkqfeZAlcA
GO0y25p6Is5p93I1S8pbCB3vqu48wtXBW9x15gcuBeLDisOFpUezM6QypCgO6jX4dXJX2mCrFjMY
Nxzy2JgYWmI0+zkJHO8vN8qRoW2wuVuSGDQsi9YX5/SLnuAT9u/unauIsRkySH2hRjn+/DlXkorC
c3s4nn9W2y695Y93aOVCClCXqitR0DU1f8yyuUGadOvwNl01Ga+ePAXO6gy/Myh52dyj2LgidL/K
KeddZVZeZoVHI84UvlaSeTKMqNrravYomgKcPIzLeX+kOMk6POvQ2MZp/GfaC0uNrR89BUZ7s66v
+a44j4bypbHD2FbQm/Ntr8zPRZFwYJxlkX8/ohAMNdT1i2ha27kF2rsj8kDpQ0iKUdt/vo+zEfLZ
GlDeLzAS5ER4IPmFNBCbrHrXef0NqUO1dgvlIqaqp1tR0OLeDoAeVI2MqldVuDBt1DKHDtUUNpHZ
2w9nmipXO1XEjjJ5QD8D70VQ2efiDCZz0rWrO/kOZRxKdZ4MZ9JGIYfJ9JjNmAO9fkGsI3sDAE9H
BQ6gqDYY2mUPEPepceosDH7Hro/8m1agn0Lz8N4zndNFkLMHy2qj4QqvMRn5wcYJx254cC/es3e/
gPQKjfchppW5nVfU1RhGYPx0vN1uhhG2pJYntHYeIlBTIZSoetfDybqdoVaojub0zJKVhCAZWWxT
yFKC7kiUnKTov2ereomsBJmMmWaHD+gCLWUSPDPsWI7M2P69BOcK1SX8E3QHgORBF4tRMSq+EVGY
kfC31npTtWfZJXQEBLTxY9L6fsa31CzVZxxocARwcPMKQ+bMdaBiYR+skeHDwT10AU+npqwCEWcT
lQ0hP7bPF9Ia2EqQFxJFloFg5fS0PeeBaBLQtvH+IiPEezTlRp6mW49l3pY5+RDqaC8fWDO8wLpA
TVkopyiOzCEPXhh1RRKfDAoEZM2jX5GvEk9JDqFoM2nZinSFSHVsZoWjA8QKN8E/wsNCzvTYCsjU
pFEI2kwD6vWWSYXhxvghUrbV54eaqPtkVyfAOLwH/tsvE1DgbgAZkniN8WTJGvb+X/9EhZGF4zfl
8V5xIYRPJP2QHuS07OMDasxQCuv7Juavzs7HgDckOPwUzZq7SYAV6FOWxKHL79yQNM9kRQ2V6NJj
THqcvbQ8zmLPaK1933DQq/M6hp/qR4pGfJLmVMtNjMfYdjb5TYqkSP9c898oKBc/8223X5MExXRD
5LCz1mDs/9FkXDZ6vU4P3so00aKBOXMdG0A+1CfyyuItTxSlMtCJtUf3HMBbjLNeK9GP98G7PFQy
SQ5V1mTAq/rSvWXDWvwjEle6rpT+1J/ILZRH/dtyznQswIeSws4LwD1dKp9gWPYQHkl+VLkBhDfs
m4pD3f3yYk1U94xYzEgypje9xnNEekj3tfn7M9ImS6Co2EucQaIw+yeekWlMG27rc9jCOd5AyDSk
fo18Wj3QZgbhpk0/oLkz3L4HU1s8g8LHERJmcNJ3oj7BDfGqsPeVOKvoTwBUV7bVg5xB3ITMMGw1
beDjiUdm6tsny+523OxL+j80pqBS/cLwXt7534nCSDA1SOXs3+jt4sxPTma92V5hdnYzQAK3fBaU
qzWSZCNOXC770T05E9+GOyVLQBpJB/TaTwMOr9bjfQXCng890gvLickGBRCxeyrYZPHE1VaiFgn3
WDVMQ8GV0XcaizBaTdtCXwOBXOTPT1EzhPFs6m8ttKEM4tlMJ036hA0RLJFYCO8TztR8+1tDZ2ty
5i0Z0s9YDrKkhyYzd0ekLrt03crBFre06nkSFXY7/L4gah3nhFWgfiY7uBSLS5miCBNJ/Rx9wfgB
Ss/PYWSwkkyoycBaGxlImmDNlnuiLZOErV4idoA+HI+h4nXN2BAojOQzqJvY+H0WbMrgsMy85s7I
KUZpa18POKH3XYnjvrWRCrNW/xcGxfJP6Jkv4YbZISTcREb+m5/jSMfgbS1aYSGZnj5PV94jMNO6
k1nBNSaantdzcCOQQp1P6Gej1voGnELRc+zsZQqlbuaNQEl3N14OT6Bw+3l6O/bL6TA4bwFnP6k6
DbiVQis79uP1cWslkQGxaOi4Atuz6boLRGm1t8XA8FQ4zwyk4cDu5/1+hV1/YReWZM2oVUF7HA+K
044jKCetsJv5j1+AGkBPqnDRqsxI7lCF40XxcgoyjMxQyM/ZU9ToShrz42ejcqWszrqfvQ+Y10qK
xjXdYDS7xI8EI6NMqif/f6kMVRmotzsOdmFkSij0rcT5dOzwbu+ZlaIOeHdTh+3HUbD00e9QaLh8
c0w7L0BA8yMunIiTKEJ2sEssewcw+NVSM2A9/HFOAIUwDae0Io2zZkNPyD4ODYaKG7E2meOhJ88G
ICtV9MMKc5IY5W2I3vmn4Mfvnc5vNtqUWltZ+57YloDlsP2JowoE/3SXNbA2IVYJZUdqRiyUSnxT
Gd2J5pSYknUJteyRkivvLS3al+E/IcVuI9wHaCN/YXbtx3r2xJE+NKDZAgMiYySAZJMDnRN3r8bD
uexfEKDIht8Vt38kzHEtWJUVGSTlEgsnntzz4COZLc/TCnxRnk12hkvtot5aStSQJ89ne+/unnQD
BnY03WG/UotuisJPbjQyxdr0JaKQNHHIcG2giEr0HlVHcBPPGU5e7pWet8CulpZghBjTyOu0wcha
aBYN4oOjb+lMRBRCkwgE/0zT1DOpn84MlQNrL0ejghKLYNfkvwMg3PouaekMGFAMRE5Yck63MI26
qwx88292ZYS2awGABwk7iKD4lt835PuTI8QSLu9om9imBjBN91BJfK/9UMYYTEK2DcHbD7o/BTtl
EeioOhoczd3jVdWXo4lNvXsxkRpRbkDzMObjrx7SCbakC8RoCGoSY5/z62oIAsdodfT5fdByWMd4
gJQR/xKwTkrjlhTliMfzuKvuBV/v8cT94qVvjHj53SjVAktMXFxIpKMjhfXp92aNFkRahVGbBcMd
CPtDthV/BMqz1XJF41lKVFJR1chq3yI1/VLYP+o/FL5ZmMPA1zRUuJaVWvaM4CUZHzzBLHqMAMys
/N3CBkMGMpqM99G/xXpklj+Lr7bATdW/A/8G/KbFLnquX2dodaA2hy0kFWaePWdflZdi6HiGA4hx
SPQnhu+8Ea2gzWN12cQVs23J+c25o1LFoR7Z7ODIzZ2EU8HKFp/zfdvZWm/YsCn5Gma5HmRCzmAq
a2nVie2bJSzAbzNlySf5f8OhD2W2p5oh5mMStXpR2GzWR4kJycMNhFe67xnlWWZcAAWHsnqwltGp
dIPwJAwagsLwT36jTMmNo8QfPI9WpzcixjpwmqxTkJgKssMtCq3K/290osv/yyNfNBoekPSpbDmF
VG0iLx2ZOAjqrfdYuG8BIaBf9f2HLgqm2gymm7UZCXky719/BRxalEDNQOETzR3HOsUl3udOQwaR
cZ0jAPziGpgoFIYeZ6Vyuxl6Yv6UhMtmsevNLquQqiirl74Auaug2pmOAZg0sMt1MjiWGTGiWG2t
cNRtrifAXUAnkSQiFf33oPnusoM96XqUN+Jk06jZ1HDH3m5S1JID1kvTPK8ZHrULKdbBdRYc4dPf
V019uH3FznmIYsxSHlp+M7x0iSeaHGkzldeNpoCvreRF0ucMa/zdnNGZRY2/BbP5anIwN/RtCWeC
O0CxxeDNrHIqE3WtL3bI4lWI2DSJBNxtgMsn8ztyljdcYoP/mtgtf5LzWxPEKewDqvQGjPncxykW
qCu7xbmo6xKQYR/XXd9UR7ZL2QN1x8CHHGV+htEwjBphzpUN+oPhmJr2OAPsu90wZRBc9T4Ho2bE
vdGnpqaSJVyGU18ipZqi2r63OVIRY4YGNQ9H8pmfCQoMpFm9fYbq0KETGEmoSBwyFoj4HpyQVnL6
w5sjE3W0/TQvFheVqoR1f6l6XNwmHCMAe8a3mzouGLefzTijVo0UIbWpCPbBDRqNyghe22V8iFsK
WutzQaN3l9I2/ApxTbubDAUM/SZhgeUgR1WY+x1tUxbfA+ngihbg+De6CUgCjU16phU8mQvNP282
qhvrlw+lJRBk/MCMTZ47UUK6Tg2M9NIooZnsmQI3oVS4UC39+9fti6jf9/E8b3TnbbLIqSppAl5R
V/ur5m/rmyMcqBi8znoRsC9hDoPHqYVf52iDjJhLpQ4xeLBzOwrdKdAHO7zPiyX+YSNMSvQ1SpTr
Rv35FqwdzfNHTSN6UW9jpgELRQXIIc3v3F+F4d2GPLiLO8CNKvsNCNncjcotJaOQNAyuKkqqdNoU
1COoCtCdjSiNKLerCLS5LZeqi8qgr5GIXfGeI+MYtPG6/tt4JK+Q7h2S8r+qO7I/UTLWsqcDIDf5
j32zi6wvQQ6V+cfzHwojeO9tg8MMpQLTlW0PjgJW9w0aww0rlE5kzKlicwjtAnFegH9Qt99XtxVX
eb/a3W4aRCjmc8BNN5blktOFsUoZdQiRMU0OoGz6KniycItBBlOgLftYv0dLXk/x+CZDkB76atD6
5CBHJyQSHL1OcUIcnAphs+gSYap/aOK8Vk4b7nlS8dvUsqRTMkJRblcUZugS95uNF02zKZP/hUuJ
LsLk3NjSwPK3BMizZbK+8Ar1S3SVKip07h2WvsexlHs+yz8UzRgDenXlkZfLq9I7J6zdQYNeQGLi
FAZXUgHw7KYMrw9PryTi+nonlxIR9skm1tnO7fo9MWE5DUP6xYsQohrjdaZOp+9dpa8Yq3ZKeVW4
ePN/QcggZZ/0vnAZILvCqsvbv9M2+li1tg2x96B1YRzaGfqOMDztbzYtdmFOIiyqNfrw6EVUbDMo
xtHo50DwAxGNzCHmOLs0niSo+EvcrF+mg23m3037+RyJ9OwX7bGSy/vVGqXi3tDiaLfZ6RuH2l8C
PqaDByAI8tZnFj1EZQnMij2rtOdXFmOq6cFNy8x91XoPr2qbzJFFzgq9S7O5vgBEmBeIYIPGi8NR
rKOrOLwx5KpFaK+6xxGjumBpJbIEd/DK3KSZqdaOx3uLzFHmetR61PsAgBe12W0JWeqqIkgpslKz
nP8xJz+4EayM9YbOA7aYL2zy4rmzyVUA6Ew7GskepRO6Fm/UwVQWSsZroZJcSLGYaIESNr2EjpwJ
tQGtjtA2WGvpUWrtfHe5g8JU+MZrcOS4R8wX5Z7hgk3jdwaI99MDImay8LPprRRRQVvPYh+dR0bu
74tbhwZJb8hJCa3uwRlEXBdJqg4M8mh9S6SrEy2HMGjmWVCdYAYo85BdVgSv5VeVSXJp9n1fzJty
78j01O5XCuM3DzC727okHBHf+MaNTnz99QIjZzWPJLlwEbhUpdXVWRkQJUTy6xlj5UsCJ4i+FM3J
r+S3aIdTBFdqRVOycIhRmHpxe8IrW0J6/eM12ID/9ulO/D6sxAwxo91cZ7tgaJXZ7KTtXY14gPj6
HU7mcQ8PB++9O0cqOJpVQo7u2gbAOBgW/BlxNFSxivj8iZgqY/PmnexvpK4qi9pY3NJGdGU1ygeG
jOj0MxeoNe+0JEbh28eze5O2/2pgim8kTViShlqknglvuEhMBPvTfGtlbbiXVRtDt2UyXjeiRXlf
+ag574arTH1o9rRiTsW/Hm9zsKeiHOE0XvyLedBAaVCq0pQC3oX0B45TmzhnKeKymflu36S3REgt
YIf2v+U1Hm95brg+cyWec+bh45qMljjMDcIfLsM0qf2UaRL/mrAsZyUcGT3EbnQLE4YePplTf05e
9etBMvJmiMqoMSR7J34GA8OStYY+B8zkyAXvVSIv0e4wkbCPt/boit/cR9T14rkv/1GzlnHR15Jn
PFMBg0gBnKM7wWbG1tXfkE/H0yfVWg7S9wHheyUCDMHz3e2o7sCqKujN2ZGvOyHwIm9r4dhgL6Ze
BGOHP/xJod6XNXZbLyXWQnLp1eLG29EYHQJI1micPf7PtilfiE04PQJnlVCXwlFjvZGe0ttwNXEQ
NPgy2u5/xMOX1XhMOmtHYx/OX++GmSHGgWGnGrHcDQLIx4nM2aP+pJxsnqUi3FMyThRvlBX7CcDb
1+3FwCmWJRUlH9lLug2obVTKucMQ8c1ukq505QyBk4H3WSuIApUWzF4dBAIC1gd1+brivqmcijmO
20u4qDP22z+77IjPTkGKyL1e606qxwYzDlorQBrAXzlsTQlUCknVELMYRYFRnUL+XcOW8f5ATrqi
SYhPGFeDtGxDfOgejXXWf4oMQOc1/ahnAPEh4n0TBaccjk3QJ2tlrei/lJEXYTtNIj+JF9RwBES+
VvLGLm+ldQgQXGEEzk+A0oufQ0mdHDxq+uWDpmjNXCqhz7u5IeF3d3Zvd/C6injsgcwgWrHm4b/v
quCylYtBVVzs4ClgVcNdJQ6SeUaR2jI/CG0+sqgCSfbVdOv958jM5ftfzP3SWNAMWQm06ezK/+vy
yw1ENrA1qxtRky98HLZoqdtx0yLw6obR+krtQAKq9nucp+EkBWFMyZd7fv4d1xfDGmlO94SUaBC6
VeBJM+sjvyCcWXm4X/5fyhJXC6VSVX/ZPYkyqgPY7lgNkHkk+mBXdIANn5XkdtPfPI8pbSYzTrEM
IbEoa/+NkVjYE5kpRhO+nUE9gQIxroQEZHFxuEz1zI3RODtiAyAQ++LcO6tdkaLraa+0nUIqFBxI
5NQDs1AY9mnmAnKAjXk7lFlYIeObplluCGaLHbQzjy2G6d37X/LitUOaIUoZ7BeRm+CXNj/Ve1FL
mjM+wLlP0oZrAtA3tf3ftJtDkMpQiYU76ThatwHDcewMNKTHp6y+3/uFshdtaOIyAF5vXm0ypDGp
8dszxLht0E9N1HEqfABztbJcd3FpFmDyM/z8Pjw31gx2lUOd7LUvU+UTNFzsl+CWobLYhjuGMvNn
ME0UWUS1BE7liq/uh7mowD/aXAWsSQwTChWYnZnIzX/HXJKLZAdEeQOFZDclVcLYKPdJqlbCgjfi
u+iGEYcCI3VfPiUvi07teRHZZ8i5DKMRn2UNfPUKlYV7AoUGzOEfDXDXKf+5tOmI+sxWV80rCClb
WFxqACwGq8VLZAgwfXIYgCL4dkVCJ1u4DLcKcwqgk9Jjp3wjM2C+vfobfdGgADO2U7pTxkIruwk2
kojIHZc997SxOUjvQnxEqlicaskkS3MC0rSe27nhMxkuo7H5WXdLz7srQyxQTCtNmpULIvLGyTuc
F+fvU0knsIPRHiLc1RFiX9DnpysvwUU+67gm12xt7novMWOA6vsu/3WrwoFKw66WQTXeF2/qtwoG
CCBAsEKRphFH8VHYbakFWrmunHcUdut2odfhS56Pob546Fe1s2Jj7eTJgYgPXToAnzWzeFPXnFoo
Bb4uSxcU3KPToRWQ+zPpxVTv3+I0f4xmVpRjYH2VSzeetmHzW2i6D1w4Y7tZNn4lz2pfdu4ysoT7
8MuRvV8Eb03wFNNxDiKhr+IFPADla9WC6xJFAtSml/jb4KBSrxo7W472PMBbKdTHfpAWjtQ7vljD
7OV2mqamoaAFiEQEomPwztzwiEEMjaw44Yq1kUE3uaJOnRvlXNVsads+6756YxqDAGq9qyj4m8lk
vQDY7f/OgYqdUhk+MKBphDeuCaPUc8QafBFQ92Gaq6hdlW1aJ0Mabm3xZN4pjEJqCcUAMTM3ANb1
hBrsjDhTJAJZ1kp+p5YbFPryQ9h1ISopKQ+gcXjT9IiGMWAcwz3FbiWoLTMkaoc/yKWwnD/mWSQb
klCL7zelzm+w/jsukv3ViBJo48i0PcaoR6dakbMNrYBjAJk2FfuuhugjXgMT2iBTDb3oGzsL+6TP
dIlf0glNAm7aUIWmbahKP7Wek2/rIKQdHRyeBcRws7k7jpSkvRqwCBBrOefJAgxpIdj317T4B/Vp
TLCOmID9qrrUAVgMFSjhTnJLlGy3cNTcTTfCFk+cc/eRmFCln6+iKLeH4kU8uW71N5yl1XA4SqX7
TDknef1Ss1JGaDZZcGaOjg5GrEaZoIBMRjj0RXvVXmWuOE6V6iqkp4apzLgruJhMXE4OxNIkSoBb
KnvzkL+lsEABpIn4LB4G4nhuXuLyxZ2sfUShqkLC8iE97m3yXzirQhQxnk484znOG+5YcIdPag+W
Fy25NZMRRit5XeBGWkJx0tO9BT7NiIbQhHWN9EziSyUN4hQf3qgDLp00B8Wbh9lJqYZ0236hV6xL
ZSH2DBn4rqUWyjZx2R0lHhi362X+gdSATGjKvUurJD00ip9bbteLzxGl4QCec7NXNeUlTPhwR1Gf
YsJ1+f4ghWp6CQH/JnJHrdfsawSZ+8qEySH+OBAM9nsJHcZTlf7GyCdOJyFZLhAhA6XSRfiTMfpJ
8ok1kowdHPFUe7tHx6iePSa3nOQlkq5qnUeIp3y4Sj1tGarp+PN2mXvoYm15xkEvHhn1XlzSLU82
L1s5ATFwr61t/B72YvDg4qPAtWC5mlzj48wPFEw82krSiUZO6heWjR8awyurd3LeVyMOCPPQUFj4
JGE++51IpF8+q4MtKjfexKugBgFKGwnDqSFxLaAqA5DPMkh5UUGFp29Df3u5vJAAfZYTd1/9OrrG
v73LF5JTL23uOn8D+TWf6VZjCvuQSYW90clwBG5LWxTk1i+OD1YJdb9GHtL/85l1N6ccBb9RXaD5
TuMet8M8+BBZJLr6dU0UIbHnRCXxOuhp+VXrDcSKcmbsPO77kV6ihoAaro9qXcn2Reb4VHnAQoE4
nxYLhjyc5VAr//NIXzhON6zR5j9p5CzHTsxEsEDcSrM6s/z2gfZ906PUNALsH0vms9qVvXY9ERTm
4DBZs8Skxiv76IF4ZdLOBZJ/qyML1lBRq5m9xoMQng7uo1pZ3ktVAE8myVjx5ShS79cQ0hJcxoT/
qqZxNbGr16WhNCwkzX2fr2WJ2gSGDEhcQDRHdv76I+lDoKgk6Eyo6iuwt5/Q9Usnr1jkZPVATYDf
tHetD6jeMayk7joTJevZKWzNmJ3DuR4figKSeorENaIEbD9vJyn7SA/HO9OZNj05nCCxhfTzyzmS
rW+BKZeAgVVg3HRuBsxh17pIG3sGPxTsMspio2g4aYRdV0DfL9fBusI7k0O9Fm8fM5HTVGc4EWyE
uwMJ1+Yi1nGaiMbVr7/S6d/OuhFWbs7jqYcXmE5htxw5mA0BaMT0AgYnCP1Qj5VPFbouHYhCLLBE
V/URoxxTnE5rev0H4wBj/gTL9lWjJiudm/7C10td+QK+f/jt6o9onV+PMd8E9XYE08I8Zj2DD9Zc
9MMOw0xVe64VMFnD8BtnD3ltp5MViQDOWtMGJhTfRQAASfKeMjj0YvROUf85rRLIvrrbQ83dN1TV
jedRU4vSeoPaT/uXFxhlPPu41b/tf/7n2Q6uyCZHoqvMSUAqM5Uz8ZEaNeOr77/JQy4mw2ogaO0t
Wenxm2e1sKZlR8YVFdvejbDodripCl21KIAHHhoelqvRPFauuc7awsUO3L/WFe8+OfizoUQRRRNt
Hl/cDRSyiuYK5LHsh6+x//nzPZECOU/g3y+xnB+1najuRVtwuGmhV3ZHh+FtRoS47gsWEUKnBQkx
gWTNBLBbjYrqK8kzMJFQU1F9yoHcWDtn1B5Uri2BjEe2ugIZaG0iTEMkr0bgiKG4uhSaPuevexQL
znmxOM2gOFYjFF5vle4O/8A8WV6fJUiK5YI2EpsCtt2h/1blwjef9BI3Q5b4TnC246QIm/zWFJWw
nU7/HMiA0F6FAG4/eSgq24VoQskUHMy9clf0nHzRORxBEziwmPuv+POiVfB3E6GbVZXw5VIAMa6V
l4ICWhZRpANxlJm7u3GTdFXrDHQb7hc+W/Dd0QLI4UAC0MeAm/14UNDd2k/V7uQbJq0pgPK1VuZC
frDGXiggNRGZBl3/3gGjU8Ud9Jz+10J3B7URGaT1uigcpq7bf8km8NLVE9+fDDVm/CqJXX3syppY
MJcyYi5wUMEAhL82Ih2mETbk3Z+j44bNMjiL60fplnbIGrvjg9/Ry+BG9L9AJSmzPDqYf1IuLF6F
x1/xFo3ZBGCjShvnxad8WqccD7KLKXaTGwbaepW7OWGZOadNUzGGhUMbpmdo0t8kbCVDNWo/Do2u
pZA7ynfDs5q6029+F2H2VRacuir+q1boaofhmkl4CKwDF7RyuUO5XdweAh6JJDt+xyXAwXGoR+mg
3MY+nKTYjuaHNXV2q2Nnc0IJwazfGsr4LYVvNTcVhrcAZ+yKCgHsbPoCllfuWZu5HNUtrdWGNyrh
M3HRCE8Ng/heuxFx98U6KglxigFa6sIh4EfQ8rgtsLbBbtLPtbP2TZCXGCruDka1HP6uJ8d+2PqS
9kKpNYw3xW4qHGI9dkSPxIgFpc0oqNpYMYXPRhPq9X5oRNIyZ3vAj/ZFClQBUXA7A6eQzqrI18pt
h2thL9pJhShkdD9G4ZwJkP375MyTr51UcAp0zjBJwBSCPSoQcgmE07sSU3XyGrJ6GfcXotTqnE1h
Qyu52d7Y0pMw+wxxyQ0WY8xTQ3a1xRQKLFyNmtDcqEXbhRE1fiZ0NX4KU4zT2bZDJbxi2iIUFJW8
WD73E9eIjzxZt3WqFKDLK3DiflkkwdVBLRaiiPG+jSEXdbDa9Dco+IuiqenGpzo71TBerJEQjxaw
PW4WxRmlLmeh55+xSk1w9TzBc4wmHsHyL/p8SvHc9hi3MVH8LRXfsZNoyj3rLMeIeSJw/PW4jXtP
s57oBvGp2KN/PRJV5H874yuO1MAVIKg7Vmjil8nnH7fe5e7Rve6fvKiRagoVOzGYhZ9lZcuZkksE
DURTe7lkq6u49AT9JMzOmqVAupQmrYP3S2tTnaJwHKPdP2rxEcmlXumVK1Bapu2o4hNqfD9mVtPF
F7Ohh9E2Gt5ZMe0gS+MkLFa9bc2DUengIov2SHJUBxV0xMTXSdtIVLdtyK7TWqXZRsUm/DXqF6Q8
b3KyIEHICoTzLA3ISYQ2royuQszFDvvs67VUzDnGG5FkiK8opGA/NUBml/piAfn+dKDV+iCDKiFP
5RgKl0SYq0FisHsQxiIRB6PyIbNsV7nBRJODuIGLljTGsc7Fa5fnq8OLMhWFP24WyeBdxxL7Wa46
STymzISpFB5YIHHFoJ7m/O5Q/opjAl/0xf0kDGag6s+rY90ffcjTbBxYCvA2ZmG53aPEfN8ekz25
Jil7uq8hNx5ARMC+q6loiJKqnlBN9RLZeJ71sBl2TFqZpaYxAhlNHQvWJOZ8SWHJu302lUt7CkcU
v37PAkI2wpTugnhnIAeBXw2wK2v5Gd4Obfw84pEdeeXAMmE3qH5HRKzE2pwJNotyPrfbM8dUCWqj
eUrno1v8+EdvfxodhiqMm5NUXXD01xhb85TCrb9jNRscByzK2coubyyQEHtQGD43i96duSSu0l1H
dg1VoVitbNM/PxHwYEZ2vlLzeApmqBRnOExJcRhJe5KHxWMRS4b7UrMBHxphsZD72K9+lZ8dp1Bs
9KhEfFuRSL9qJWFaqXE1EybEmhlzu97kSaF1xVJV1BI31ov9rVxhOf3d0SiI3hfMgRGZ8zHfztGs
m5sYXXUP45CczcvG5t5H/rLSAV/EWOSTMo7wvupfWC7YVhRei3l8a/f2dx1CMNj3TUTXCepGMKp7
aNXH+FhQlFNZrgCU4jLNkdmdxryKqOLuz5ZP9ERkkZidYjfpc/ONmVwyK42fkF73OQmsmuDzcGVR
C8LKTHrr/8Gi55EWeinSMs+1NZ1FmPOqPCLH9Cy7ZlbDQMfkGJDMb8K4Jwc0maaNifwgwntpFHcc
+vh8JRQTGm7IRhJwtoqSF3DeRgtzvf4XjOQ8U4kEBGni8tty89rg1UjCeWFmOizHFFaN2F+0s7Rm
M4Mw0kfN45cV7Ti9ZbWK4ywypufVfFIvTjOESuh46UF7SWu7bmbQ/+Rr4ALoYC62d/Mkqq4LyhVr
hFjnsZ3I3NLTEvZMtNWVf2d/hp53Kvr269yVbtNxyMXGYaO9AnuZXo7ghwJPPJCikIHYRU7lwiHx
ndQLwXqEA+qyiNo4lZE2w4/NhSYaSuV5DLCUqXgv8OCC5mFKsdni7u9aEN7FkkOZfAUmlxhAVzPj
UWMeHlFzaKsR7T5exga/txsWZWKLYTr51eO9LSttBe9858hJ4LGutBV5oQChJ/CyCkAZzKwvJNln
UDOnklHMXGHGxFPgGPohCCiNj+4M14SbpXWTl/X/uf2FugougADrWl0iUCswaYXgmbKnaBCddq2c
4nRRm5qEnC/pAVvZkLcHi013eS+9wxqX0LxAvMonPCbjBRGm4jk/x0jMCM28sk7YZN0UOhHQjwo3
HR2VyWpmrfr4jheoueHWiHDGlWrMUL/9dsD6C5k+y+7entfLFG9SBkT3YhvKfdDL5K2TsmwDQTIi
q7mlEoCMeSdGbiGlu57XKeNi1V6NMBp0HvyiVp6v250Q3UXMbySem1lnmIlV64BG9YM1dcM3A8V+
dZCzW5PoTKAF6GgCWRzN5bpLIhfV7UHiGbOmtHz4m5vccySo/YETh3ptFPtycxMsR7xLvYD6mD/6
spXQHYc+mh1BpBclktR8EYH0DqNgiFGNJARwXkvqENSyQsxtmOLa51FUCSIjT4Dlspkm1SNWtEAf
MdLQb0MBoUxrM5gMok+5Qgv9Rzfy95kAJvDnSq+z41FyeJWO26FBLpRx4U5tx7rtUmM121NRrbHK
3yNJNXyz7J3aO5agFSvzdwWfwiZcL2g9KWj9clofmXH8jfn4zERCWT8Le1cyh69WYezYC1lFTugz
0M1k+MvSujArhtKpNvg/cO4xgnUrhNESp9Uw7fJOUOUg6KuptBP461kPHSiPnktthbpJpPiWlC2g
sXVWPs4JOkj48S+tSSYlYv5FBMQQBZ/kw2uTlgcNlP5f2JBMV+H9dFii5w10Z5gBXvdfiUTleWz8
x4r6XbZAFJfzhxbeyRpz8QxUqmybRnDHl/jozaCfuystZFRhOKMXXcKvIe96WNy+ZVmD+GrndNgy
CWtNmCpKXocW7cb4LKHZ51SmABv5rNRcavzc1yLAZsB+HzV7L3Dj75NuuW+mqkpBDXVL+F66XTq+
id1FMA111DFjBkhX3ofMnG+3KJ+9vlMh+oQbBVDY3vb3LElEkHu4k2mGJBgh/80T9F9Nz5y9YTjZ
+KMshJl+CFSbwR97H6Er/t6FTZbI/sH7GlUzY3vO2SeMqYLAWaN2arzEYXJPIaVU9mMuxDwFCZyj
UWWi/NaZa8vCyALuzGSti21YSb0LojwMpIoGPtPoJglnnHmpBZtMT9A0UbYVlrpvuC9Uo7kTjePK
ot2BMbjrW1TRHqreOM/MlIefkGoW0cnaq13B2xNTz6Aq9nR8mzeFQmvo9PL1wDKwguHQrADFVJn8
qpIn6BIeLXY1N9MZMrYvMUrkgrleksY758dRAqDYd55pl4EjyVBwGZQVw9uK7lVOzPHsiAyoAgXS
Fm56j1vM/9a/+fhJE/N+d0/y6Sc37LAXPDgU5TPPdDiqCJO74DdU6dsB46CEb446gEgyeCdUhwvN
GnN/G0RBgyjVFYtUyn6BBaJN+uj+/JS+d29uAd1A7E9Gm43C3grrLYo+l2XrOEEX0FAvif3gCh4R
ixYGgg+kdGd0yFI3L1jhaSRG8T1KTt4fgV2j25e/mO/9wqbxoZEOTMCqdr1NSOEv5Y3PqhWnGZwy
NG+aYG/y3qiVV2NVNKLWwN03Cvq5zFJtUjSjuIZGIuALVZ46i7qumjMla9w0NgKscyVIzH056UYb
Jo/eToG092JfC/wA9Fd9NltWElg7xciwfbwYkg3HBgqBvZ9A6yZel4U4KnWsmJP8W3kjdq7Za/Zg
a/wkEkmEf25dsPkjiUdsiIvWBCBBqFRhzfhUEioMNBrkm1866/u1baEsAzYOx3ID4onmOwdpOWaf
H1C4SKHLS1hdiFjcbM75qIc9dIpF9h7ero2rKQjfmPrBta+/8zX5VZsmHA/dESXuNgsRIqGqc0YL
XofbjYnMAY8NFnqgzC1aCUCwrM2RGcaJr7YhK2+97krl5BGXjMbBeXsIcA0erb67kFDUSAkQKZEc
/7v8WD9bjn+E2lJfxw/UJHJPOnsj2eAmzZIXXAS7PtjciK2ksFHwXDRH/7zgImq0g6SbIqtqt3QK
SJVRLwOImBH9jiyhYBCLYmmtJU8+yLiEanZyDbCDlIjkDv7pWnNzUYbKcNQ+73h6x7r8qD25TEbG
5k4zhkUZEZdrf4tT6UuEy+9F8kaNhr1Me5AVZ9ZLGfWqF1qX8m8E5YuUbNPIYjoLJjLdflwLJU/7
uTwCDEDUWHGolY4By1/xrGLpN4Az1JvvEIzGuZ9p64uAO2z4CTfp/H+yTzXnbi9Yx/pqPINEsUUK
gHebBi2/06e0DTq5D4CTQVuLxHnk1T20PqrkkWtomcZPxK2ad4nO11sxJ0WyQBkeqflrFdbODkad
Ta9okom8JKWsrCTh+GqQRs1PwWz/yjghnkQEGpnOZfOmRQ1YnATNtuEQp9zu7JXNWG3UW2O4FcDu
UnMfcO/R54lh17u1QhFbOoEpzr+OTvd83YrC7pAvO599xHjsjPhPGj2bO5JGLhZv82iEBT7BHZAP
xsLCNVFRXO/5H2apKFYvZc2MhYSkNNJwHxCgS1UPFsZjT3NiZtPyYF9kWCAYV+iE12+0KsJzTenk
4IICGgKJs/vifoxNH6nqmjacD+QlbYbogBv4pVBZsR0W9IQ9njoqHtboAEl8xpMb+kGqx01yA4r8
xTh/z0ZB+rusl1QUwi/hljp8O6Kzi8ZUwjL1JbmEZWjQTJi9Inz40/ZDOIsVq3OPy5cvt6YFEh4M
B/wV5+Z7RzzC+mD2a1gpflAQsjQnh2pU/SjYApUo1QcfvruTJlnnUlujZzSNlePUMWDrUgbaUo19
HOk4bRXTRwKpmHPbu05dOT/e8G3gqlx6+aHWovtbq4Nd3abT5QTuiSgOYVSwHPoeAFLmnZQv82OC
l7mWmKLIuPzHi7zqeunAdIodeabzKRbEyUD3/pnsuHEnTa2gKIILqVYqz9R8KFJjy7Qs/qFN/2Eq
Z4qOjvEkw8g6Aq4VPJjsvEBI/ngHo1AbpmEv9fHSbfejguXD/z3fCWWfGE592cwrB74JiYQ50tgt
Cfdnit/76464t8CalYGN7ZiJITOo8xqCaYxW6b3JSk8fVkbDidRGbXtTwmgoQJWyzxYsujqSeIK5
fvUpccX927zcaAYF9yjo9ADjViwbG12rOZqHff+0Xypd4H7NMGmK6dxz7AkX0ebqSs3hzti02UvD
bUSptE4NE6Y1+Axmjq3tJhZf58iCnM7wdDht8swR5wYSDdYGb0cqVRv67eqC+JwkZZbgf2w9l4QQ
/4KIpJBGiFmcBNw/U5KgEM/yHLt/fVxTeB4qlz8OFV1bFigrPwOEzQcRhZ4iYkKRW8arJHCXjyEO
QGsAL1GKKaP2ernhLY/Ddl1UZlBComZvwa4gMToVa+UcNrmww1SetYHddTaG8R9Jfqp5KH1hvrGS
sKY6zFXFRd9BvtZcgLANduwJpYRJNpqFXN3cFVfaWr63Tv34M0NUmJiNL93AZ09w8p6hSlD6Ovbo
tjj/e3T3O6DYwmHEhOIen+aYoW2MQm6tTnxYLsuQzw0zR5jKzyodXU/SQqfeZQb9o+u9cVCNYrnr
yI5psUklxquozodDNYSuIJljtAhEHA7UQ9EVXACvCyH9F7nnmPimHXqkZCwFtnk8RSAwPnnxA3n7
wlICN2QDJuPf97+3GUdShdsePUjEza5BdAvvp5IU2TXjPcHqWtplvAFcp2Gg1mnz8EWV59fPNu2Y
JUBB3lTFgybJapE0A0UHMtHGHr+7dRzokzWQhKbvOAB+Emi9nSbTq7yEkOqdQjEh3/2OSLLKBo2J
KBLUNa4dFZS2ZLXcYyNnAWeVpGf94pIuwglLE94Ft6O3gcav1hQ/+kW/znV1i9Jloae9rjBkH5u8
e55LTLq7abWkHTvWxvUHW2pEdDjjWPJti3Z8gMsh9XvZA5WRBmWPI+iU9vUtTULJtmm6Uwd2XazP
NdOdt2G3ycsbNMWT81XGGLrDacKgs4Q+8nl/N/qDy6A+Pv/C67sElgINEXOsrXMgM36Wxqn9MYeT
0cMsjJSAOX6fTwuD6t0oBiJ5/d8txrpb3kYiRj4vGhjO+Sb3DoOjEmcUhVZzDSCFVTVHQupFIVtg
xbYUMGjaFFmqxaiAZsY5OWGDHehpuPILundmKyqAm+819otmOnrUMEmn4bFPxNCFJ7Om3DvPuAb5
JZhsczlPu0xmIhcKQTkiGFxwNGpfiBFyqnZiAd740t/z1NqUtpcYhItOUqmeXZkInRuO4rDmbVAU
dlpBee81Z9Uy6YA6au8YMAE2jZQFVDqpyTX29790RAbTMO5mSV37gkKdxG3DL9oQ2yTwxIflgNju
zEvd50/HurRUM20d5bMVqgDsnew9ll56d40+GNEvKNKtRaSwQluQsIHSXnaFr/bK9x0weiHuZ6BD
GRDfaa86oLyumeC09TJOhFziyZZOuCNMdoeTtZ0AWOOWH4u+x4WI+jE8XPAnFOgfdQ3pXZbp2ACp
Fdzw1dCW2qm8S7rfyOu/xpaqvyYCt4NWYo9EzJ2TN4sqmx9/YvMKh3+xlEKDko01JKrkOz8LnW42
wYt3/T+4HFRXH+XP6s72RuNzUEdq2QzsyXhPbPZEEi+HI+75R0iKCyquydsr0cPgx5U7pOqb07ky
si0pNjh1N2HS1+DWgc7ELff5tlQhVTmGbuDR6ofaUKGGZPv4LVQ6BGd5j1DdP7YfNBulurm9duuW
PQ2hRrjPfrI1qbRKmVTqq+UR5x0vBLX957jUe2ZVNm7VEWxe4zsf57Kgt4vOHSCgXBSKlT4FBzga
A4MQTxEEEIq4TOwbWMbBsNL+FO9M7dhwXTlJXkS6zdbYMJl8VMJ5RXGuSeRjydic27Tib1nkMTMT
efRFlyQ4lX7bdfnq0Ss1pq1g8LPhsBTy5D+Jqp2by20qZ+T69lBgPWtJPybFEb5/aBVK6dZnuvyE
HI+aDiPKH50K6dPeMHIGdfi/M5EcmJgVzEUZYr/qx3zQQ42IZ1B3UHuFmGvspNk8gZwcMthhqb51
XCmz0AsH0yCKV52PIsBoaanetMcilveecD0GVtIOYjvzsEoxmBJnXYkbX3g8u00354uQzQWGkWWR
q//UdVDPQeIyCJ2pvGi/IHWv9q7/LQlNwCh3SvyBVA6f89m3dyp9OicSrk2T7l5Od+7CdTgNSJ8V
OK78P2egVIh/P7Nkdly9UeQ97FTCnHjQG2/hNUDir14LFPp8AC+HwaDe9lco/9fRBjjs30gvxCOq
uDSV1AheaLx+KrixGmdHQ6b8yiXYtunYD5sU5Fumn8QEcXKQiGLZPwEJ/yVcvwelSUlLum62rMVK
tGW7L4w77IJiefCdtuWiPKCNXL0clc3mNAnG2aLdtp74dGArfJzrUdp/Q3CCD3cS8BQM8lsw8t8F
2FDUSf+I9D8FpBirikSy9OS8ChkKrVr+z12Sb5+C2DZkDykhaKbW5aWTEF0fzOBDtFv0TPTzDH0U
XhMXALUrmtIRb3EPcuS60QjaTXJ40JlA2Hi91cZsOb5tYczEVpXcRyUrEMxGmuHCwSUOhAEgiGc1
tdTO6tpV/H+FFfbNcbm3F/zd4FZdPHR/yAc7fSTgKYQjkKICodwGAwIohR7CLKxafMlBYuA0uaxw
b/hxxiXU0fZRvr1KDNe+Im1EErWfqdaGEPAN4n/hOR1emhUgxyIithzmnZUhTELrsYzokb6ajOns
MOJpcWs//izg03eT5Jh/Z4EAODOGj0VsaonraQDJt33g+/Lta02IGr6BVUkjNIWrCpMwb3TMFSzR
UGbWZ4Htio+SdTbfpFTVd6JEow6xalbmRNsvRci3BSKaMyzQo4sQ80q2SEJijb6LxcaCk+adMxd3
aAe/A5bji0g8EPRyT65fCsqdzrSCnC/yXmBOY4pI3ghWURxXUTFUyvBuEWXjlauzIQKxcxUS8Elc
HzA65YtNVorHwWAiqvuaArVaAGK5/CRbCDMjNhMo+KW6EfaHIu2NemrT8Oy105T7MvuHW8m2BE/5
n1uYX0BigKf+0dsqlVLkB0nMewNAFlkeeIvU6CdHO6lw+jW/6tkkpilQeoghHZgFCxncTJ94uVaO
JS3J7Jn+4mUZMqFwuWgiP6rMxRmT6Rtx+EayrjzdL95RDUpRzvUY8MZCiqOjGOXueglRNCP4nasY
poHXR0nPlznbkZuhBC0mlDVo2wiUD0YVFfMrzFfbrWgajfdsBhU4vJXzTBRovxwdLfpY8Lhslg/1
UqzpbDtkqLWdLAezwjq1SI0OS8fyqO5hBHSVSnAJ7ILgD/2uGaKP3AUK2M/1smtD2mVTRSgSMWfA
kzilOJlWTKrczxxAJeHg3kZzF940ptwOOBMbYWfoI/YPwNlKtRlYIrP/EetvUmZr8VEDhv0ntuPJ
XarvzDo7u8/fjKOlX3stK6Yaj8IDJe9P6tB6xLgGHPey25jVer5b02edcB/DYGiD6B3/oKifUqqL
UgOlDky3/JXe3AzxHH134hcoEeGjbHAZ+zimc4mymxYvlioIWp5k/jB5ihXjVZfGCMNWUwpBZYyu
yzINVK1q6oABdkmkil9J7kdCzxA9poTzJFe2noZ8N+gRfDdNZJeee2HB2M0NxajMf9smkp6McG2s
+jq5E0wRkcz4hAhTPYbeZeeAAx5DJ6zGLCq8zaER013pBbiYjje8AmUeI+Fc5S+aNKmR4LdbIPdP
1n7OXNzwP7+Wg2depGcGYrQJcqqsU/t02Wog7OTJzcil9FeMiZCKFJWp8jAw/xAtnRcqChfpUUjo
W90gOu6TviX8qGt7PG1kw5KaNCVVaWmj8mSPcfjpDK/6gFYWxgL4I28lv16PwqCBrFidhEthViiO
3IauCLC4Twa4VIq9akaSb6XHV2zpWLaQ+VVl2Yf94E8dSCq6zjZuAFaPF1nk02w/mqDWUyt4oF3I
atLbN6KjvyblJiTQ9XQtOHGeL+W/H2JP4/vj/CUPc4Cmhr5G/ZOqvu2I4Dzq2qAaBxxPOqz3wh0Z
Sr7Bq+X45SSyfAC2wtznyq6E13v9IEgmaXgsXC1Bk+W4Tv/55MiazmJHKc4zupdAVvuGUasFT42c
BC8qIZjdwEFBhcwvx8tJR6nlqub5n97L2ivGCMX2uLQqWAOubIKF6UDIfTJkk2XxDH4x4NknsjcC
G7X0tNYUi6wHzGWfmf48r2fqafyFyNSRTF35PM1k8zzCADd24EwxZH0O6I9qgY4iOhVk9QVF1Ex4
rtQInxXvj/KSXvxdTG8g91bKKsVX+IacUjBUCbL4J8JFaZbXG0y5wAbSNjfvwuwvdhPgE6nNoXoV
SwfYyLj8ZGmWxOzzFDN2uftAUHg1IM2keSywtTWg5S9acNSGoxlbgjmDYZZNKTz9SCOISyZMp9H3
SszjDJ+q2cFgUiAsgh+6tYtd1/x9iK/z7PI2/14kAy44dXy2iRjl61w9QDfsfK2DGswzRy3xktQL
9VpYo6YCeLgwDrtjq/mS0Tv7hFSI886p/jWGhwXVcAgqvrh7YSt8FsQOyWTB4NMhoY/T4A2zHbRd
teEebpCASaEr5EvoJ8NA4o8RhareATKWTvrTFbV23EwtfseCRc8oI1yH/zaCpy7Fb5aHUuk9j650
CnqHn9Am08Nfj21HU7A0acgG+oWJ8ODIgBV+5HbmFuuMqls9sTmd+dT9uAXKUvviheXW9y7SnBXs
2rlQPtDNvsSPHIYzwi//WZyi9ec8QsJuY51tJhQxWFaC8ndNUM//5CZ5XaJn0AEprG992YuQukDp
Y50z3CxqC34rdI0+yB7UBwxGbnM/mxHeH0GzeIOG1Y92Q76vVipoqBBVpr10OqSnZNX0Se7B+MCi
9w3IXsF3G/wt0XjxJ5daR4a/YwF8c72sYrrJfz/QsBC/MWabJIxEaniAfSYGQWInO3YBOqHgoX0l
1DDBFxuLyJUDlA5q2x7bpCtqtCCjoVun1tLyYWGwj80OwJUpoifsiHQ9bCxRAQwSfzmcn0B+q/cT
hB3mCt9mZGpX3bPD4i9xdLUrffCpnW3uQCLK3etJFy5SAczTl4tqWA2wgBYu4sfRI+IO34knHb5Y
R+LFHyGWiLCADNHyEU6k8PyS1kA7SN81v9vaxUpXiFrUqzNNj9feZ2xHmCcXR9UkIQ+ydKOsaFlF
XQH0rOyIZX1fLR+AlTGuX0zrLWh8APyEqnJEZaoIiiz9EUfrSYFS5aOvIUZ64vvwleK3zRFIqoyd
mDQLsG1fZXLvxnTWtEP7YRabCP01i3WfEqGNusAmBbG6fHmdxZjqqzAXwa7zd1kD0wJnJXIcawpj
0AZ4G4nLFwBRxrciNPxJOfJnusoCLpkSzXwVuBig972lrKnl1Fkrpwe1VspoY+1CYgmnpsveYvvM
+3TGfIbIcEM1Bnd2qZHVOx4jJ5Hsx1JyWcYd6OyDsTy+GYihZi2CJawzGvMT7MYL1dJN8H+agOUt
RdAWdqcEDEJCWnYK8NnBm3LvONBdjgD9eNeqWT2g6sYUz7umbvXRrEU0b9j7b6GRoFKIu9aaNj2D
d0VcRkQTzIGBOb2LP/f7iGwzVJyxb/BaIld72Pjn6Fz8hLpby5kQ1i5CtwynG8Cbrfkx7/zpObdm
rMSIufH7f9PAjTNxQr+f2Fw3RgSZ2AQrh2wBJKjdmhxLxvnN+zEQhS/eST1jhgnS2cB39hm07ALb
pNSMj9OTxM+V/dOD62JobTvl2Rd7NMMaYB8j9W0ZAza3j4aydRGDKUO6A8XHmtLAfYWD9o5+UycA
79N41ht45L1jC545++3zBi1pmoE3pB8O25hJ2ZI7MsKDF4WQF3Mu5X1lqsixORnNqONcc9SuI1zr
wGt959ep/rvGsebCX1kiSgUEyVON+2m2OZqEdDDIiXFe2kpu9BFEr3STTGuH1FmU3Lo1p14ACQ0d
BbnsjMozyMpOmrI7bTaNX5qMmj2uN+sk/UKbLRtHX7TqxQC+4tqrABw3g368F95wr1xHyKhnqBU9
73kYSQe1NpDb11PuoMrXaaCWuW6dAMRZ4sy/ijJp13t1YVUtLQp2DbYKZqn8vSG1kAY7Y7IVSZCA
u9XNDboE2w0fHsWd/6Q25f2jbfdvjy1v0cYDa4PSzV7oEG4YZC/AMiAxQUmyZjoQ6UhpgMCIunU3
kD24xh8frYWjxNQ7WDYdYdESGyOJs+pz9OCqXfpLAybt0Xlhc1tucfET8a4ORvGys0ENRxhj9+qI
DB8nei7vxT9kh/0xYN4rWRS1AL65gWL1j/HfVClBGZo5Eo38epXDSSiPFRW1t2oDDS0ay67ZxgM/
0G+Nj8MTFojwqfIOKfs7USOdQXB/dOZi421C8y/fjIQz6QGN12XjDqQq27cvFrW0WAdQx/IpwqIo
hVt+6l5Rb7hJjU4ELrAEPJvcXgmHdgiKlwbQBDC252DUmBICY4MoVo8dHKUZ3p8DjPV4AOIEUwQw
TUi8SV24jZGV4ElcrLj0lMJeyLHb4PzJ5dFaFADQ5XDFO4UXDXp7x3IZ5NMuawDto0FLFp2f7Fs/
2H22Sd50JKWPHS4Q/CFXB+PprmIBIcSJTRrNQInCStPUftPanwttVgE0anG5fXjndzrpS7E9y9Xl
xXehVxRGpAQjgNCiyLwDjv9uaOviTyicP4ObeV5DUyczqRbUzEl9C0VpvQiAYUqT0mCe28HPwKiQ
PPtliNhFe8up7oIfZd9bqahk0/SIZw7FdVECdLpyPlHx6cuiywwE/7J+KNuI9wJbA5hdUlYaXf70
/RL2nG3LFiCwo8/Oh1Ee383gVK6pewpWQqk0tv25esdWyDV2Gs69qGT8UPJ8ujUvvpDdE1W3m1JV
JyYhNIn7fDmfL3VbXBEp5WNLr2ZRaiKdcj9afTI+7gWTyedhwh+VSvEkYBp96nS7jaJws0wLVw5J
oggbA++YRORwqVQfBO98TBtURp5MtxVUSdoDI48+DPNbU0KvX2W9xYxDsKsNXWCXX+5QvPaj6mE7
VVl06fnC6uOFnQVllTGJup4Z19Mv0zeFaJAuH5c2jSO/dpMLUfIoFd7hYAyzg6QEFpmbRw45xL76
dp8ie/i0ngF6ZCyiMZ1UmqMmRpgQD2KtmacLGsl6RsSz1zodWYk9pWHKCAOLZLaaYN3BX0phdeam
GMQ7P0vH6jWXjxs4LI5mHN3TN1xI8llyrIqK0vnoJXuI9SqGTQaLY6ZPP3mZAC4GqoVIQ1hLydsh
iHx0HJGlwBQ0I4jtkoJ4nmbCZzYWTW0hoOQCyYv1FTvDXVqur2L/o2FeyYhDsjcqLgeN4NGWL+JN
zAD5B3pFpS6Um5JG7S5e+XdIn3yO9vYPkeOOM79TJLT/UadBn3vVVWGlLt/J2nK+kr/xtBjEdVQR
VqXUp7Ekyv7WJgRJA456ARW/JRhXIN5Esiu0Lgrcgiac9sNn3LcWBxiyk7EICjDA/O6HfwX+BcPh
j7dCYHjMQAf6maVXKYgq3oh+9UIR/BIH2F1mdlV5Wq6BlY2/JGEiv/Tcx0Qav3MasETsUOSCyKqo
3RxjJBnE3d7R3CDgiDLdR/DWRVfVnvZFNuRMTZUbYxQwWvcXAHWhnM2j3swfZ0KbjXfbSRzJU7yE
BVM0B0oPEmnKZ9uT8FrqzHZIvTWNcPx/m2Zfu/ljESAHu0EOD4SGhp55yGZedf1PxrkRriOQM1VW
poZ+QrDBaeTSnIN5EcqqmRbjJYcj3coNgp+ywgqWsvFezpFQ0yzJnP0HXhrvi3olpEoMTnWAaFsv
9tVfDdseoycw/th1iCtlDmrz11086NvP2OyB0p68KKT4/7kcQsvatcoVeurru9zpmi7V21eQ+Hzb
3crvPWWVQMxHVDwJugcsetDg50yA2JkSu4YC12UMJLM/EiDKU9kQXEwdu5FPUKhe5dKHARA2nTvS
bNFsL4tA5vdggW6maRXESW0wjJMjmC2w6IAL1JxajgYFarl4yUY/0kDcMkrrzj+N8qnjTBMLs52H
O8OISJkiAFGPOeEwNMx/+OyzRmL4GBxvY82JhogWN4Wm1gPy8LEpxwt0hivhjolG+TcWm4XdupLt
h1bBOS1tBvhox6nFewg6knSgqnZ46onDEIfkYakDnXlokGFbvHkwSwo3MW1cJ4UYJbyWYba1inzF
1WXUsyLWcEIJsqhblKqI0A56O0k9uqSTyj/zc6rQUKewi63PoQUSk03ZtaKoAj6E3lAnDki6mxLb
thTZmRk3wmtVN92rgWWniNX9OHfTMxZMqXkdT/7bt1ETKKqihc8qN3jKFVLGgXj3ZUz8Yi0GDAT7
ojynvNSXrVnecNRiwVxYkXIWShCOueDYzqM1qBczjyUtqLMvmfsveDp0i4bsFxruragYhPuBXbx/
m/oMH4YFiV8+RtO3FW2BlhDPdoQU7iGcNlsAK+z2msPo9PSxCAqZJ2Dxv010w9Qj2YUWyaqZycJY
3g1vQy5Hri+3upFAN8IenlCF6TZDJ/YSsp+gEl7G9vwEU4G1JnvClZP62lhoZt+FGOE4ur9RFmPt
YvRQIre0wB0qmPeALq4GrGAErlK5HYV+E2wg8nc50GPHU2pOE565dxSmMVL/3Z323Ax8db8UBSME
F1t2iEJkxZY+yIFEKWQgrRNcMjqkvdeMi1HutrQuxdGYaOF6jKJ5NMrDHIoUiA5QBHLcog93gdo0
p41NT9Apfl8q0BmdJp6kDYUeFibuFKTvqYBQOtuAtSVOjU+M/H5iDtTKLUKSRBF+xju/cA8Pe2iU
YvCvo9AT4I8a8zWdLV+cxsyObE0dA7w6JbfM0XuEm+McrJFoJm2jK9DHygj03kVIcR1hEp1tLnMI
WEBql389sKFuJ4F33ILUq7hXayUAiC6DnN4I/ibVSHmyfh0m99nYyRtY+D+eFwNDNlqm8pxTQeY+
7XUt3n7jPhcOmDjyArTAZzjjCC7rIhLUQykOrZgI2DQAgf8eZg55Zx3Ig7jwSp1BfyxAyn50lyqA
tOfjW43Cg6Jpu7Bbu+AI0wMhiNfDsifU7cObIOWTLYD78FzDgfrakdp+/w6sJFGHyBme8eUgcRH2
bQN6R9AVnXARgokQwxDJka+Civj4wzDdgedCachIUi8Bnnf1tym1fyN9TmPMgPZ6FWvEPUhIu4qB
SsMflUFGziq/BmxqUl+za3V0wHMm076eH5JMrXizMdP8q79eG8Rc/QeNRFcTQsmXZGiPaCY2EHf9
QVLQ2lWqlcJyt9fSI2Rs6Y/cDE6Vn0lR8fVE/W1QKgBoYOcQJepp21IAp9dl02D44zC1rjmL08w4
CLrYd1gfnc5jzWmt7LhZp56Fp2zxBVzwRkSDwB2t9pYJMi7v/RejqW3t+KOQdG1Ue1nYd3pWIko1
+dBbpZWbC5ttWJDOEkVRQtaF407g86G/t8s2GY6yoM+og9pnHy73wOvM1QP8n7ETj6TgCwPyFeZS
SJzjrBkXnOTTQtXSLcIv2WeqN2xdUPOf32jO4c6rquoUTzUo+qmEdu9oJOpyr7RBJjzX7VhiOJrt
hhLVTCEQvmlAiDG3VXsguh74PVBMAkL/qDFtIXLGxq4NdyRU99OVSHsBJ9BoVQxHbwEh7s+o0mNj
wTFdGetdS4ipE+TGUyMFZut1VGVB8AwZynAZnmOEin3WRGYIGiO8cMyB9sMvMIQG/lnMht1C414v
OR7J+3P21mSWv28++K92KaH2kTyNP2jqJSzlOA0dWYAIVzu0CrVz3Ni0m6QNQuOpWSpG6mDTV+rb
JXR+SuLcFnNkT4hx8oAvaeyPpX0OPGoZGP3pbUYAbWegO1WvIwx7ffPzPHRk0uxX1WRKid6Or/ov
59lTTLkBRN/Is5Ta5HiSHMUdWGvO957ANLa9IvQUjmf6l1oT6eS7iOJVCeOUqQJgY/ldiJYqb4jh
eIFxZdy9BFN3zxYJ4bgqbYI7dGS11yROqsUb+sKXKUkZHHOnkcjtyMCwlxBaz7jF1QJvEImel2HS
PpqLf9/s4K5zl01UV6nf4LpnuF565Uk68ZrfgFj4kv4AbWIrwLrf4BwSGaJnEf3uGA9dWNZapheW
6MdcOO5yEEfIj3IJlYkYsz12Z4LV7S//PhxyBh+f/AqYA1ibGCQ1MMvGlNg7BdwnrM9/FdJr9hw8
iCiJpzPlJV41UeuRIKjeLbXOYYgAHsNNLkRk/NKe4tNHOQ+W+wDH+Xo5v58DTPor90HG5DlwKHSn
I75RSHDj1Cvvnv634S8nXvFbg3n2gRUAAwUjmk4G7qlPRX+Sz60QUNcAMaYoPe0uBzbVA6RTiaXM
+ce9KFzPdjrYniMr0hM2Nsuy3LOkkTa5QlfCBXC5DPYn0Oy4YMK5fVamJ+W84xdOCiCJyKp44Rok
diS1Udsqz5AxwTLWHleVak7BYPRvS3He40+vXZwnUKEKSPdvhfSaaSSE7V3U9AsOY917Mn5GZ8uO
yRiAcZRsoAqWAHcLjfuw1hdyTIWFHTFgZx6bfeS/UkYLdljEU7x5Ya84yW9i+18x4WXCpxDQGRwl
9VUQmQNDP+FKJMyvSDR+Dj2Mtq3S3z1nE4OJlS2Hf2wjRltoCXCzULgn5rz6WY5+D5JnJLsE2ZZr
vZIbq+rerdY0NeE8xj7dznzGYKRoiimnOzlJr+aD+SQC0wSiF5/vCWCBaSPXBfwNHlKnabNaPw9n
WOW6IdE/OHEK0PIMpnoVUKFiDlVWwu1PNCt2OpbT737Xx6cNqpjuJhfffCuUBsoPoMKmNhi/Au60
n4lcT5sKNNJDudj/AB2ilTyegmHe9BjCKc8x04k+iewZL0Lsr3G3c2Qvx6yZ2Hj7id4oYvhKuv9E
RdA9MLs9cVHWfAbwVmi1VYkmnMCSLkZrqblWEPQkRh3Xp88Zjt0ZeFRGLK8Ul4A+3rEumybYY7Se
BXxK9Y3MzXgKV47gFF26DaapkG6O/4WDTtdQkBvHDWXk9CLNRuv1KFDRKsFtMruaUjI731yTylaB
XRQiTPtvitNCiRmX7S68SoXzlZ0/50YL3khGWsugjx/76ro8WlNNuKBPBOuORe1/VU7Dr3InBvQ6
3cXK4WTUTGzD+43AuqldAVSPJo0tnXxjIiqscTWtSIFYbN7ne7ipDWplYyP8pin6j7c/UIuLXe3n
7dA6BpsL8Zcr2z0BU/9K6bXdM5eyebG3t11Bzj0ITt7IbIg3yODTxoAsbJdXrJyK5VKTK8UzeiLA
5Tn8GZT8gwyy114d8v25svCv5cfWzbDk0uWnxiiqrJcxa1ng6t71FkoWU7+OGORrfy5cvPBwRsxF
vgYpiHZd/U7BK/9zZBjoF8RTOeBRlprMJOxVMIhVdHnfEQkA3i/uevdVCpVbEuKcNjO35ARxk4x6
DOVLUJgsQBEpptq6VjOUxIS6NFhu8w9WPIBENEUtRPiZxyWTcOoeCNEFwoDOiJdE6vEtht9D3B64
Cy4bNSiiO8foIDm7pYxqB5MaOoRrFjci3eMP+pGCYZ5gMP27KWuKoPKQTX1+2aOzb5d/SBmablwn
oA9hrsh9RjCcCXoa0oRkiEldhBFFCJtw1+oQugMPmJXpVr+YGGBBqCZ07RZxyuQelyzw/U6fTzwq
obRTp5/QxljQpUXnn8yJC1Io8pvlFmwu4liKHGkjybgDSrBCUOywZRzhysC2e0KCNi8qGq4j6Oge
FNfKaVToyX0ipTv8LvQJzMvu43huaTysSrOaWP9jlpVp4eqFY1n/28jgOesa0fY5l5iuu2zqpWOB
cQ76IjIWMdQNTfAxCaM34IvUs7YIcLYsKGJx7Gs+3oel0PXiHfrDMbCqUqnQ1oDMAHgLjzE8eHSe
rhHykBBFCFNhFZLVG1LRAhEo6ZlhxuZ/13t3PCuTVuXiWk5V3ERzJ8Esr0RXKmt2Vsuj7aYv1s75
AwY5TytZKNMUaxS3AOgfC07qjoUlUzlb3KNCB85ilEHh57Rj24UD6l2/c9lhKkIxUA2QGJmuuIij
a17FHpws5XvvQEHPSHhBiFuWYEOfp3DRciIGZRXgC0nh/1pDHhhKp0ahCctxhP+1WpOog6YFF0mG
90Te9LmH0QEOSy9CDL25io3ietV+hJaqCpFdPioSQSyDOT8juS50NVh0dKzDYnt8MsWo2lQgpb/A
kgIrOt8Gls5E2VvzAOoP8IUDfISvGxkVlzkG9XPsXlesTcQuQd+/L8CSM3TYnC3UY3q977cxSoLM
uTVtulYEJ7Dm3Lgji2qUREfcLlg62iE9pO58CnnwiTAY5cH9H3ahCQuvSyl1W0o/VDWvt715V2rE
AMaA/RDva/8TF5zRyBd03z4bUZXwfY/+/AVcLuuEARnOsJ1+Q3W+YpxXeqWWDyQoFC/Lg45+mY//
uqvYWI8hyaTbdQXMQkArZi2HGJKBMmt5ds9WYxhHP10peOS6pFlErcb0yWK07ux7BEO5gpxZ6pHk
m+x8n479fn9N7g/eAgUzrMr6jrXhwlNWjHtA+mYt8kmszXiiJvCHE0xDJzfBqBRo5k/devn5c48n
MnseQlVB36GGQycfK2ACtWX6q4jq2rm7gMwD0NHbIOORotVLrX72xjqOP2Qp9Gsx99vO4ANoH3dA
TMQgGMeY7r/gvFGBClCkeGahUxl0IJcjrCFo9Tj/+bkn0CuToM2nRnt8aOyDprFvo85z65VhANpf
9TmGHTaA72m5o62ANSbt6Mknw4TNSfWKA7G9LRhOryLvw03kJBkc90gmwnE3IxV+NXy8Tx0ATaxa
N+uFRkekzsGqEkAU3uSogi0BL2BfiZyNL6n7LtzXeCtuT2nus4iJyxPbCCHb/sGL6cRlD9M9HKXl
odey4lnZ1uktcmY5yg/JjyoQ8isRlBwju6iEOu6Eqy0MaPhuBIBshegfyeE/SUTbRG0Nxfp2Y2Bf
At/BbHO82VgCUjnYCK4K6Ew9WoM8MfkBFkWx/Ec1bxbuk+C2Z1ip93WsDichQHCWwc7ksTN8C5fh
IzzpZSoj5Dl2EAZgzaA0v4imjFIjK6VSRwLjkcDmlPFecPrvADy/r2AFwSsc0QTUxUAa2qG+Od7i
Yd9k+ZmwTfJLLLry6eD3XU9gyZb4fyxu1wPoP97f2JvWVlsnE2aLxT6YTPj+XA37W+BBFEXu8Tmz
2bu5hOk6fnWdj4nS9xWik2Rj+cjeZzxr/Byfuh1BFIffnprQzxuqB3yLn+Gx9jqeSEhiDFqIthRL
n+a407u1BGrTkAH8NCQcgcMPlfYRde1iVBH1pS9QtzlvcWo3Y5JL8CwhEPfXtCXisPdm3RnTHG2Z
O7mMiUBNm5akLcfkG/YaVUbeazbbIa27UtmIxIQ8yW4/KVQYXzVu0WnviCTkD5iC1WPp41Wp223i
v/aSBlhKFkuuIYxUc7zZmVTkYkJ0JU4YIwy63FwesgTpx9lzepbo1B50mRpEN7JyU512cyLdnU/T
VnDaM1S8EJoz821SVa05AKfp4LlVrVu0fR19ZOu0W4S91q3D4bRZk5Yf/bmv2JSog1x9VJvCwV2Y
HAfF0N+u+/GYQH9k8ro97YGi/bp1CFAtA4Z7W2NQ0Ix/wIOP1wJcX9x+q5ZO9RjGdgHI47cZrVgd
kWtttqpW2rngjWClYUCM5Li2IzjH8p7woBIX6IrCU6PCJd9N4VOJtUPuZMOPC17xACCH6HrL3V0p
4iTfU9sJU9TDIvcdQExVpBODu8U7om0Rxb9bgO7MiIEcHrRF3Ib4Ks5duqbPYrfUOrwdTndxChX2
/r+DEuw8yg7g5F1wmAnxBsxmvxgb3l36JOobtgqf8Yp+uftMrwpEuaLsHIgW2SpV99y3xNvuELdk
5trY85vtLSBWQ8A6QZY5RFrWDUwXkIEsoY5qHfi6FTnUi+orVs7N/LqKoI0ONx35V/MKZyb0YgZB
DBocCqUvHizJYQJ+rGNWHZDwqP0yJkycqJhO1fJQJu3Z5itu6iMgOYX7aZ8TsksfSk8IYKDp9Kmy
TaG3p1EXBjN1YalVJzce7hpuIMow5HcBp8YBtvoRhhM7klDx4oeG1PZ0i/1G6VVD03c98U+XFwAY
Ts3uheCBbO1/7y/6Zec96IvWAddf5tmJwCpvhvozpknC504d6MaVCqwv1spEPYNX+JtJmSUW+EIq
DCIJyJ2PLC4GsX5BBuWe73fOPYsZkQL9tQ4+/rfMqgq45GJfUzSLirjCKdV7TChNRbTtu9sb54Vk
nI2tb2tCzHi1cPNkedLuIEHQ+hi/HKHZoYW932RhxPj7SF69hAuSgyYXGZ+hbgZlSXF2rLiLTprj
Zmqillck/SW/vTt0gn1ZHSnTRLEPJmuTgFwePLwUa02xVsXD6XGFoswwrdyLrF4C/0hrHmXDWqRh
44Pr9fQTyVIpb1xXqOK04nXOW+wzjwLdPrHjMP7l80yWpEeKw8yeAvaQJ2bBBgEKhnUUS7R0Rj+0
V2T1yYFcoYX9RzbZZSL9hfcsghO3D7IA3mRxjjt7+3YqN8Z8UWMIHncS+TGdKAeHwzHidFcawLfn
iyo1RpfXK8QMyntTN4xTKYZITjbcDYkSNhNh31BrWAG9zlRFVYxALoXI5ejWtK/b6u2ets7c5Upc
GBMHwwnKI1AR9WpmUzro5QGIl0EWhLx6K8FCNg6xw29LNQDCTyZ10JwokHgecH8OEEE6yV+BjJRa
fMDCmo0OLsocMoCfDGDM3EJqLhNmwEI986VSRcd4CTM4ixAQP0qWoaYdWc4U4vCozFtCrWZzjCjp
gv6XkZjHiYlZCTTJhU85uLyeTVEjVgKq9++/7ihJDVybW5Gu2WTXXedc2V7tdoGxDC2F4sTUwpNS
p6SpXiNP1dww7CRFfbWbFqYWMGfVJCIFjtRAwd3i+PDGMPh53wD3dh/q88E8HAzVVdNx6UiS+XkG
KORweu3swC51jAeCESunj2laSqAsH26Y1Jy42308TIZvvjuX0Ren44/Jy8ZDYc3N40zPNBHDMNvZ
R0BlUS5k7+SCwfHvi+iQVkLb3Xy9KyH3fXzzWc8I+gOlPUtzjwwVOOrPawP44vChXvmntYmYCwDe
ZB4H22KeFR2L9c4MyXxlHOrFxtJqlD50jNypjYLjiOn47a0agXUjAZA4sUeRywDb8qXmJ+D77KXF
9HGM/aexgLkNQgPi5uJ1bNHe80xK1d0R0nSX0KphPEEea9CvUaiCcVaWnRwfiLURAi9ZeNY4TeEJ
L4cHTKBa3M13SqE4aviMMZu/6y5z3SgfW2XNPt7wDuu/DOW7K57LZAhWf/OF3Nh0HOc34+LVJU5U
39WdGZcUF3zo1Udm48N+oMReiPjvhZOa/YIEiqitiG+2XeskePya6x2oEg4sD+LLKIGyjsjsGk62
rkpzBgxd1TP/d8J6+Ipdbw2Dejz47pOpHfsyL9yRXlR8XKujDxSMR3EkuEZ9VlccBZhvJ2nnufp7
OGIJ/WNpdp9rmpmCKmXSO3b8ZwUeHy7GW/HXcIIMzdselm1ml9dCdPlJ0mWV4/spmxUCorDwcrMN
No90eXZdSN4aLdEb2TzedJ8558QPzfDGKIEOv1NncpvuaZnmRHwMDOuMLM37jqVkz8Lmr/qg67Zp
+2pQLXLElcd+Wf4yqIjtj9o+uXc3wUmHvl69ZHvZF2oADGNWBhNdG+Mdbm3MZTm7rB5fqqgY14vr
Wp3FTYF7DQZZDNK3ShJxkZ6PsFMA+Oc/F+hIV5+dOxuryv5VvT8zZrTWNRw+XU7U3y9sAa+g49JG
h0AIVgx+JWsXFUdUWwqeUThB+KFC+aHsr3HaBah5Pjpww9jdHz2KfnTigGNpoU02B660eM3WxwF2
SVtAJXpN9oBtDDFOrAmNGdEuzMU91e+nHlmIoENGgzPkCRwuAqbcW85qXnDFieREWdy4YCAkfK+C
HOJ17x/lYmHfwpTmofnsTpZE1Tu77AKXHxY8jxh8DzIbhDnHE31Ru8P2v9krMhRizOkDPKxtsRVd
QvGGUx9WSDOlXXaT2On+1YyVG7OSRvO4oLcBDYSg4aHrYDy+LtizBOwg44CYbtkTwSJlFIVC1IVU
k2q8DATFVO5WuGX0MPUairYrQdnfNV2s4D/TrwTD9QgSt8i743QUJ1LqeFNMxEclVOi6lrUz5jNh
yoBu1OepZN+TPaGtgRh7IAY1r/XaGmD5oSls7c9oDjQuh8RXfTIKNM3ncQFiRDCzHFnv9bMwmX8N
XLDaGFB8TlQiJYnnObqrKfEaqFLmmm8LauN5cNG0+3eWATGNqNgBwgrRqCzSUW5OTalB0u8JAMVm
CXQN4NFs7ut3vMM06MxNzbev8UIqwosbkVzWB8FIfLHjg4Hs189u+dzFk0NR76JXKAtKL6ooS6oW
brVPWOg0oYXa0o29dtc1RPvNaXOkcCoFFs/oJ4l+fStcm7SrsFch6Ss2373OBPtSNr+9QZ6+4tfj
61V9RJ30iFB8onC0B3H8VUHi5SMiaETjKnBVWws6wzA0uNXE9WKhwj+CKYUwqRVvot9U1h8VTkw8
BK7WfL4y1feFiQLqvM8IPQIqaWEoAX6EtO9yP9DCRt5V+lbNQDwj9BcwAIVCAxuA6OKn6jpDuZ4U
eVYZFf9M9HqcFHqc4jMzL+fumuJLVa/BFQrVSi/67SkapcTaBZEgjr+dSViRNrqubg8ZjVE/Yp1A
BeuKL6NSgqiKy5bXMHmgIx41ayQ2eLaUflW3zkbRjggB7ejEDAAmOXDL5cf9czD12I3ghaOMFHCs
286nJJI+W6l5oG+nCehCeBLDtEWuXuJv9kmgqr9Q6jBOJAn/G5Xet0zcmYZhIssac6Rk++7UaBf+
OY/Np1rIiJhEOIuU6sCwL5vDDbSoHA3f9xb3/NRq9D616T9dEX9qJ053Cl6Rh/n7/wlT4VnkZ6Hf
IUfZFWIBEfw/dlng2+UJjBOcKyEo/cZDuw4Yj33YrdyGb/cJcUzB2XUS4PCvBmXKGqM5vKYXEMAK
7WrWFJWGMqywY0NPMp1i6ZMJwQFZTOJcd11b21/dV6DG530x7VqJpv6U9k2sZr2gRR/DtSrRMAyM
so/5icTMZ+tVhDuIxAUkY1WKOk1UhcIesoievl8wumiLypCWOPKPrvt1b2fc+cnLwQ2Z5gMO9XYy
1N0jC+nQpcpJ3VNuIce9avlq9xdLw4WXlrWiPmgy8TTpevLHJk2cc4qEMHBBOnp46dA7j+YP/XAR
Of82IZI75TDgNjC4efod8Ej/JrlhBcyYyuwQCt/Km+wDsNfrakbvTZqjVlQYzPTcRnhG4pQXEbEo
7h7zmqbWErTVtGr5paUQ+UqSHyX1PQZeiv//d98Jrz4CrbIcWYwt90El0bRAdamZi0utpNFQgH4K
9IkdDkcR5evdhGoNRgNWB9qqpM/kMk+eQUnbXyrgXAFCfvba9qL0LdC2aC1z7nuSQ++HXsMIFUtx
nP/26EB9ARUuVjqroInhIvoPLy+fq99Vc5B4yjaWNTYudLKniLx3uQJKOH5k1blZ5a3CpLT2Uu0C
y55vdVSVn5gC9zR/DeYClKL1KpiiGblcbEbdw/6XDWyBktcy1ouZGQnaKZh1kkx8gVUUsU2P9RWe
hFG58BPXsVW7YBTiFhDmk069jIFpcWMeIyF0k8Suo8upQjIkj6Bl2VlvNTl37hCRogYk9215ooUW
N4L2ZhHcRfV/nwQz9rkdj0LWnrhybsMKTp8v1A9wL7281z9jHZM8+bWcNKUgMSBCPYXKtMwT/Owp
IVvP5ZB0lrwMIlJ35H/R1/+cA8HeJ95kVD754oPm7WXB+BRVRIR67f1WqW5O88NzhedrVMyZm5az
Id9BnDp0vIqXsB6qgDMtmWnxur/6jpBhFypplPyccmCOshM6InXWh0CHDpGGsNN4/kBlSOzm+7wY
LSXctykPp1HbbYdfLuP7wJLHmVLH7hQIus3eEcScp5IN3Ln8RgjLEbhBGyC6uwXO9gDnBXLElLIB
Ok1BbIeYrIGRt9u3A3sEg0OQOKSs3V8hPqGMdO/xOPcBgqBABDQk02T6DsBjD2lWhtSpm2hR8HVc
f6dYMlEoyBLdW2X8qQQQaZH74ZBztzV2+7JQ4pGH2xH/mrFRAbc1jWPB3KZFWQm7uCJpv5cuSSca
4vZKzf9zFVY8A+Rj0qJKwCsSdWzfeWw8L3EUPUxmtU2C1UeIIvSvitdtELGRWfsGkwZRD3K91inh
B+qMxDStVU28GO1YQNRGUap0/YgopyypLu9Ul1fGEPnd5JfSHDFE/BFkFbgpdzZ9LvvroMt40rS0
NRWc6JKYhGHANR/LrtuETPgmeesrwzcUicr0MwG6IlAutDIsLOo97vfTjZmGWnoI7RvxUUnH+kEj
7lsxVR52gzTKxPZrYW7T6ENCVLu+PyN22f2GIYvCPnZ9MffzHvUX+3bN8HF5i8HgCj9XP17lOvCH
0M8kzaxW933iGbBIevj9dIvkvdBVRrk2oY61DEezwn3Sos2TLutqGxKR7Pro54vi0VeKMvutQgUe
cbVB6Un9lDLfnvDTYr9mY1ZJ0t1daUHQMhu03wotc5S1bz7ex2ylhQ2XIStIahxXa5cO2qBFEYMQ
gGOyqlaD1IFNmDdjqmHzCUGjxGA7nOq0KlB8bbp3tcqleNrTxznsTG+LOw5ZsQyRgOIjr6vU3JsH
l5qh7Of5OBSCALkjjODZc07vyI7xDG84z4mWlNHdocayQu8uL65Iha0KplzzFOo2ZSDcPCTIfw6f
kjoOYyMH/Lmcx4gTAMkPbitGRE/IhfuPmRn8GcL8V3efvEPnuqRuZTzktgdbzN3xstfyBSo4al5c
jfSq6vaeJt8benYF9T3e+Xm+/Aht/Fz6Ot5h4dxSNugC8FVciLvXMkhO7VvGq75mfXYASkmH3dpH
2aT0tae+nyWnBxBUADZxV8mKFoS4PvLgemlgXeO5NCFu9I+djHgaupU33Nqxd2xfazhh8ZAMik2C
9SOe293l6A5fkZFg+v+IlFY/GMW3rWaySrBisC064uvL7dhaeTXRvl9M4dA0jdbcYl+YZQOvFdaW
X2nYYwrIjypH7tFzNOscJuPoBJa+b9oU4t13BScUr5DkQ3CAgs3URv7fJCQE8SAA5JB4cjo81nrf
AaeEoxB23ji3aRoUlNGibQuCjSk/rITRJXzworVlpgGZPjdkvD49pz1PCEoGHLPkRVjQT3LtGyoA
BLTYJGLNA1tBI2YFFklYoWsqIuUaxXy2gfe67kEQ2X1W8/E1ArdLM6f+B12dAZRXe94hb75Kiwsv
QMkplZFi3ivhh/FNA5zkXBhGiWAVnU+ND8FHFD2xQdhZmSrOvZNh/pebGIVekvN8ch2vr1LHxdQ+
NbItoZ3Cjl8bhLyu1nqQOvWiMDc63cs+L5GheiDDp/2m3/1kfp6wJlxTQLh9lfZ3wk1n670NkbS1
GwG/d/w7utmdT51dYS/+D/MfV0ZQvzB1EWtem76ADk8ZzP+3myYITqJArQlESZrU+BWs6gXxIo9R
Pw20hYLjuP/k89jFRiLid2fkSu0wJW5vnGSJmqhaJxOyg1kfm9J8tY0hvN+45tz3vpU89qMwfjEF
hUykNK3YHGoZHbnxcYDT899lBLuPZ3U/LXih8ynI+wx4AytZ61lOHxIqzydEpxOxcJ6y0KAQYe37
44Uk3Rmr7YX2a0HMgqnoTuv0b1ubR6bAEmezZbTZOe0sf3wZeXSg6YcHcQ03Yfym3s/9HaGLppXg
yE8qvd1QTbDzHquMgTdt+FH+bEWE/CIk8GPqFZg9lvK6dkCNQhdJZI556LUrpQDyNVtjzHrIFcms
7sphvHMz01xte81h8YcYN/AXSk1e3R13QhLbs2VbmrmSfWDWuytqsmFmY/M0iL8R/RSSZyfBSEsF
j4ElnIgZlZrxBUbcWSxjQn9hJRfveaXFGC0QP+fGQ7DsKc7uaC2wdM7N2OhxPpo2FdhymvidFf6I
bU674B2f/n4c1d3LBjg5p8c6PekcWNRYiZdBFz0uHYvBiOpfHLkfPm6furL7/GBi9PB9l/ycjAer
P2fRgZcgbFsMbc8RGB+qGrphx/2sVCUK61nx+G7SRxZMppNt+NR80j54bN2HahFJ0HWv4KjY/pDN
VVcq1xnvQqBrbYzEZDMwjtIX4CSrJy04MBoaU4db9FujNvqF7iPfDV+YEEvDqZRwhecNq6E4Vf+J
lHeoiAlBmveLjg/cppahuiBVZBzovUMYRWe9aoZyusulJCpT4id2bN72ibWvO8rlmHd+h2MNzJ4C
CEygok4daTTkHgPaLUFIj5gtxeUaNM5zmSpTAQF6A9cbwoAWBsYdOrYTBJJDAA/6rsZcnX89wBM0
BkWZnHzba7LsnE64VPXj39k3PNLe6IWkKGP2bqcg0qaSCD7/STA3HoIZ+AWVKBssB1+q8BlMl8w1
LSpxIGLPeZ7XdIGxGmZAgVX0exksVJUlxwWPg3Sh+XoaVMwHa9iAkxIPzivVMYJiwCdSudRq6pEB
ZXYg3hleR9TPTQB8np7aQSngQLg0+BlBbyjQ3spNKFVitkHUZ1I3s7tzMQJvT42EsEQz5J4Q7GeD
+nBkRfrEAJs9/5X6+nyVkOwEch/YVvRGby49SUojPDn8obFBmHio55E/CnnYvxFyDSPSrDfkrr4B
suat7yrp8ZS0/2W3ELuxezVWdPVIiJraqepWCO1VZnUWsPwNfn7ajYmCxks4+WjWyZDlRc+c4RSs
fdWm5Gg66oBtD5bCsZYgrshPjM+yAJqUwK9Hs2l+46vbaBgeGyqVtEnJjAJJuSN325YG8ZrvZaWS
Gbz0opnLe7AZdIL06lUguLoOUV1zUbjhl7IlSXZNEoewMq+xDf1rtLk7HjfjYl8PVJVoCvGuxMZO
k4o0WbqUOyLwKqUUNP5MVWTfY3ATFXG8j+wcaCIG7LAzupO0dEkcQQM1hCnN2MyTDJ19sI3s//IL
O4HfD1CaLF48gdLczrMNhVNqSPM44JzMAy/LUhbxwvk9wDKnE9eeb1sxi4kGBWNjlYvH+/rvxk47
LCRToMH+nuQjE3mFJzM72VhHaxp+MByeBjw4JTxFevy5EdnroXIvAv9rvuTwMHgImgJ0SBIA1nZ0
F9aljG5NwA1UhYnoyUJ6wTyJeS8Hg5uaVCMZVIfhNCJUc5YNQ/zg2SIwX9KqSDquE4ExsUtbLWke
A63C8bxxJcnt7dtLmGvQH0+HjQ2haUeMy4TVLKUrwbSQJgmihc9Ke5UcheTVsGx2MRocsSp09iNk
htWc/Q2gdoDe041G0+qIGlLfTY4ojco7aY7uC7b4yg0032S+DVtdazmyhmNk4OJMx30dlUN7xGjE
xNZtvnr++Apo4Vf7T60ojDGuguwM8tqjmU85zyKXSsF4wldZHyIl2qbEF/PWK1KioZDKSljl7pjS
9FnXRHkwqa1Jo87Pl7OVm1rPFVfW4R8lxrlmkPKNRq5FNcB7uCJaNVCi8hLQaPbX/MBDOxVmsb/4
QpxLk+AQrYbQs/GttSJB/EY2mesoC5Y22QKY3BmX5Ch2G9iRu66rIEbA09ot1xPTOZaGFe2dLEMs
EahIHQEUkvND0v2gN+rdrfk4o5PmeEKirGYhhCUI9EiL3HWMEZgz4Tweruf5psbCJzmDTcSzcUfw
1Gn8E2uYZcKjoTM6equvhoX4xJXx18T2cg1jv2zZmVn5jDR7Na3buVoN7mZVU/Mxc1AwaWXBlsKB
tz3JqBLZL+f2iL5iZvOqVsB9NgC9m+RLmPXhSCaSNZwkb040eUkA6hC05VXwiLnhixoZ2AE3xdig
FbURvWN99IytbWC6prrVRJa16CjgN0IDuyGWp6XRNhW8NLlTkUvXOWwCu3s9SziGa23aHK562gGI
TrwscWjFYykr12W5GiQd9kJ6WyD8y3DuV/sqSIdokRExdJL8SygCC5DVa1lilKZqe0A2trXUwqo/
c1Oy5tPfPz+e9J0h9slMGzNN3D/R72nuCDSQyNxvJAOFuWg4QbHR2Z7KVLtnBcbEoQGV8OTWT16P
w2NEyMPywCPK5y1zRtl8sJhMEkXpgkrY9CVwdW9zJ9V6YUqTTie+auknBxfneBNRWwXtEczWVbrt
RGGx1V58dx2bgKgTaHO8ouZJlyH6uuoYoMU6qgc6AjBDrNRRut9nVs50hNQzknGU9kiBevfb69rl
2S3Ptq033CS9rI1dAZkSzg08A1Nhykbk+26qaaouGqxGKzaRe9gRGRighhvCjA/L+BrlT7FE96xE
htNatjMJnOZQg+T3YMuBcKyD5f7FC9i7ALqQAXdLW2qg3cMfmpyfD2R3monKN+LVMJpPQYyCXVrm
wVlAwz1EfiimkzfyUjnV/6JPgkOytiZLwOY0Vsy1tsAJ81rd8HuAETs84TR06KHQWiGeCj+TxRH0
5+3O5LkifOxThEO+9fCDP9em/jQsTKUzesiFRq6nuoC93C+zA8v09lbX9AwevbiuHahX8XHGs/yp
heg1MEvywwBA2ilEfNZ9kzaPj52kqiM0ApNywRACqi4wpgPGyS2I0GPDmyi4WqaGgtVmJYyV+tI9
ZpHQwX0iU8KcjHb19YNNOA4JF8Dv2GaVdS4EC/NIx7PzeyER5+AP4uheIs2PWLcBJcSiuJbA1w2T
A2JXwozBzCkdSQIsFatpuBKHaXNxKSfHtOlsB+VhuC+YfqobMxLfk4NuvhdPNE5m3tXW1Cmsm5mj
scwT4Z+BsLvbtrlfWcVzZ/dEF1cAZaHKi24vElKvLLSig08qQ/2NOMOrHBTDvQC6BtucpUQtOtA0
Nj4S/Rv6pM83lCkJOdJCkUtuL+WzFzcaZ1ajnUpIYCSnbSe/aSOkJsJhfQ7qtC+IdIrvyibyhNmI
tJPNU036rwrHzqPtgOGOvznrLOsoLQW7Q+9j98PWxgANenrFrI8dJ7xJUZJIYCb4zGNCvRsUn6ks
p9g8c8FDMzXumgrr7IHalGAJYVKr25KCfVkpLvRKEF/Qk/1ENxV6J+xmfONeI05M4IXbi/oa6mXL
FVTf8XpaJh70gWUphxYg5vlgxcNT9IWLhAWjkalf++Wz5Pctvb6nuyTvJIbuf4wIcUBRfdvov3WE
r4k1Up9oPGYFuM2XGmYrWVNeHg9D/Rq3mkMQmVEmO3Yde7kaOoJi/wyKEj9UDrMWf7XMo8rhXlDb
YW4zbR4ohkUx1dNUT0dJo1u11QqhcFeqqaUZF1PK5QXClS/n5K1hF8NDp8MUlWZqYeIhzfdXL7Fv
vs0TQviWzR1+voWtCGT3eIsrF7/cLEhsFobzgNGHogSMKwvoeIXv7kGZ0j7XzycC9DSfYpn3ONN3
9RBmGB9i1ZNceKkA5LJRIIyBn0RVBVPGXxM8FND6pz1wAkPE/RgAZu0QSu51kBR/tGpmPh5CsqhQ
VSsu9z842evsF8Uh22zG9cucI/gYIucMZoi7uVnPnvt+XwdVMvvvt7NQUZFDHe8TcC2dVTidE/wz
EMlcpZR/lbclnMT06jBb8bxn9UfvjfcNbmBdQKkN3TFlkZzoD2xTQJ00gVUQsw0i7l15ggEWHdRq
jSLgv3+xJ5ap8Jzl3Um7gp/mTu8Vp/N/m2YI0zMKH/jEp9A47b/0Ikkhnpgk/88liGGU1X8+raW5
Z+MbkEhiGVIAyMydq3NWKLQZpA4yeDikFG1GXi3RMb/vG5olgdPPUCqAf1GfTztKyBWDZnrtHTaY
0VqWrjj82UoI8kLOJfFl2IpaCtZyWmtWiL4uKbqcJW7i8sU3Ybsh8vLYsVoj/EfPCGPQ9fvx4m+U
xthbq7HGJcCkxGQ81xi4cRdauOElDDW/C7NN5KViU/oIYj/ZzTRt+YxHlHI95N5BQwPZHRSZXGjV
adK2NmqC8OgFEAL5hzMqsiZKqv774BwV29a9Hp21rUyXjf27leNatpWcKLaGWm82wzZD0pFwuMNc
ie3B2ab3ehqVT38Jnr7WqQprWTRJAArGv23ZbFkIZqnEjWmFoeHiXOj/wri8qbxfg7eJumA0Ice6
OgBnoH+dH6RWBd+Ua9enG3qZCmx286j5JbuUY2R8MzKb8c/6EWguguNeUTw4RXk1QpjVce3kafgz
8MCygw/qaW1qRf3cgURDAcnTzn+6pb5ev3VfIIZ/zjQzGljrdEpzskYpxBjGavYzlMZpHzrRD5hH
n9/jKAeKfd2OGQ9AZH21tD4+B6+hvEOMfyfAoAG2w9Y9kNF4G8KGeBgJrh1DtwmgxZMMmPtaMjai
SEn6IWiyXe7DXFYEaVwEz2ivhuJd4c7gp4C7S7XMjjX3t4iCpH/IrZz2UAvjt/1mEY6Fr5eo3SsO
sWsFj7bCsoWR/XnLxEVJihWmvHFLciL/coXXi++grGNf3kPZpYojGQ2G+Uiv12xeTr2qGeVFsW/5
iiaJgdJBFTqGpacapZ4IBj7C5QLQO6oAJkhbH7DrWKlsyXXdZbBAfj40dbof0f0tDAWbstkD8Q4O
QILgC/BtHYLv64ruBPVe3XZI1ZRJmV67Lbm1373c3ivu1nV6qz8yjurn4fBB3xThHjolyi8AixXS
MUOLQ0s5OiNoaMO2sRtsdOlwLo3hv2sI6cc5KXGw+6E1w7pRLrjd2H5Yg/bgiju3mIX1YJYhIRdr
7haCijrWaW6gaPgfV9J0QOWQ4zuZHBKqZiEAnlqNN6lxhKEoBAScqF/oX+MTbo8iNPH9zz116K9e
Od1vHcWv5eOhNhonN1crTzQ0GFEAtJwXq2Wl7G5OddhLyy17mLOou4rVeM6NpclVpj6ovTlOsqUH
qnS4pVOjLypI3Xb/feeiikbJ8anbNABlbkhLZkqUKcNNDWJ8xTZTlRFrRiyF2N9e7nlNGTa3ld8m
vUqzHAqZe4ZBUN0Of8AjfBbYRYWjn00Ptcs/JHtCm1a88dT1iXE6ntjGFuY4B8b+2aFBA+lM4PfH
Q2CKbR+BuUjvEQlWxRTXjSMOMW61ur3UBNSkKnSVHW45IOSjBIGeFdXd+OorQc5nAKiLISOCVSBu
0PySH7iYiQs2PKXbPkq3dYHZEvp63Q/CKL+zJMGFJUKzJdlacfolSbfk6NQDcY8Kxxes1PNLhWwT
L/c30TJhljaUfkA6xBDup6wkBwfyVFdv5ho7VFyacpIinkDhEDNWi/5lrvRL4fpCQBqxqCgJP16X
rsTZiVi/FDmvO6FzCI78jVhUeKfq+jQ/nWCKBy+vRVfrpKBd4TI/1avDZPZKyyLlsaaEkF63e3UI
usAyWbMag4LrHjpq1XAW5vCfh8Gq2N6oA7q2LQ3A+G65bhsl6vddMf/lqfuxhCpA613WbOYEq41u
hSpPhLEsAdctnz1QzdxVIhHvht4Th4Q32jwuHVipxd3YVb2Cq5XaR320vERwSdAEeKUXVB0JL+PM
yn5W9Y2Jy6PgXS3z9vfeH1XJNBPVdlAptC/vao0kAJUh4sgXZwineFrDKWuaQwEFF2VMpnn1YKIH
vhrrHGgSBsXuvWi3RcVFnBnU5osAlA4aGKYw8y32DVGXO0fZDTqZsLAAVhdfTP/D4msZEWl/9Uo0
qq/b+pPTmx8uh5npUjpdCNgNOqASMeaM0InD9Vg+TTAAAR+/bXrZvpizIDKjYF2S0oof/J5t2I1Q
ceDrUNYkbhHhE1YQ9VxFZWfwVqYhPS4Eez7nV9I2q7V7QNPhulX/JvYF5PBbXbe+RHNcmRcIuWW3
RAeu2M3VC6FmeCZjJa9iVhmyIUNl4pXrICvtcOxz5wTr8aqdDXjfrFfRW/843vO/9Jm0gzNEsmWz
y6b5nf614OPyqbzo/fZ5Q2i0m33jT/Q/Jl48vPH3Mbb0FPpgCW7O/U7+vZ+CbqJ1CQGy2hRCp34t
1XUd6abwUaIdwi1gj/ZmKp+8TOBrAzcE2wMDkzIUkiOLXqgbyNr368eJ80bI6z/sqO147PCDrwnX
AzHvyelynbfuNkPTG2GuSs4iRb0Qtg1v/ipa1I1Pajr8dfdIXYPp2/Ojx2Lpc8el9rKfyKPiOMQj
6NQf6P8De6Fwpj1E0eIogc8Qcu74Gh3s+eDtkfeIGY7RyhvUNCUIQrWCYq+sr2LZplQ0depGxBki
QCW8k9dTppHw4kKFsL9ixTGJQ4F2cJtS7hhT+UGmyU160qY/dMhXVHkbGOmTe8W2yJPSNFDGLrHr
0o3aJUiOVfu7ios649dzfU7PZIQPpzll14dAj3bh3MRN3A9r8uTmURIFEgm3Ze7pksPypVd5VrcR
/yX68kjP7xQ0CcwJjHAxHaL3BA4+k1BWEoXGe2RWu45MD/Ow689spl5A36Ddrla+Qk/0MhO7akNu
+f3hLuotfm3gIUfzgN4eD1milXkvM1H8TN4+L/fsiIdf8Fl2JkdrSsXMAdxZghIgkBF25Cs0ReBQ
tNaB6iZFzSU6KRFgrEvrMHm9vJFOn9pbLDvD5B5TVZaUY5LSTjWqj0TRYVfdY9sGa4+ZjQdfGenI
3u4gTvEIgsCFUE0Rt5weEdZj6h4mMeCHIx+XwtJFZ2ofnp3ao0Fh/9X6/S+U/Z87TRZbHwo8Hn6d
r3UJ4FqzyGzF1+VBgqt4WvLjyAOJcwTIm7McG8GKa6raJp1KMK0CsIQtuPiOdwxklmYnAxMHaTaZ
1FF0Hv82Au8HbpTgiqcWDWQpc0NYEddG8Df3PUMEmywbFb19X1EEBSmVpt31D05CxfX9WZ5McPM6
xounNoA/bwVVjSEw42TVnRkYVmPN86chxLLfCZr2yrlJIuUbhdLMVn51hqWVtageu7Vt7ldEh2+P
tkIfah0iKTEayRYKPrb0ovyxSD6BfqHQI6in0W/Kvk7i4NKYJdUq6UXK5TWrcAv4aYF745q/0jgJ
fM9bEO8zThsuesID5jIH6xo3olFntlRoxc22WVmZfVDeuNuc6zFKqw/7bb4tftm89XMR0e+hreba
JX/yRscnwTSIBjVpL9Sv1kb4HcJht7VwoPJANIRZ3YNij3LFI33FQclJXy8uXsAV1Zc4xrmqNnJ2
NcZ/4upl+ML5X9rrwHTHOd1+9GXK0xWzJDn6RiJqFYNki8eRNQKWPQuH0J4VsXhQlx+qqFuyP/cU
eB1VgIpKEPv7fKTA7CjFiCqd+4Vj2CYhOf6l6NCWqeEjFrSubxYxRyINVwaf8nX37lx0RbOqnRds
fg//NHfeh0quC065n43Vni/ujv9Oy9NhbWtxMFCyTUjGLYna8hSle7QvfNciLp2jHUn9tVEeT9FB
gQ6A4IxtxJpxvMmwQolWuzt6IVYC+ggzJdsmq3H3oSMyPEnjb4/xGSscXNJJGG5QjYh5k68AXs7z
P6SsnDtQctGp4sfXyL7f8sHKWECGGMVZ9Unxt99iRLJ11NU4v07mVaYg/ULC/hXfehHH1u258TIG
J1ZVQ1NO6S3AjwE2DlJnqWsBAgOi+ewZ42a6eH7gpRi3uQM8fJAXya++IanKILoxijdvYo1o26Fc
kYe571GIHhGDJ1O1gsjNEi3XWh1PZjyLwR3hhZ9ZNemwxv00w0LZr06lIFswlfhiiWjs3j8JuumC
vZkp0lMgp6QRoWjD3WoNJ+Q3ezgDWSwuku3phuS5fwXBBmX8DRnkE47O9/nSKN4PUL5vnOTu22K1
6fYGzei3dHUZOvAd3+SG5YUVOnkCi9nXqhxLnwGqPagnw0RBa2FWOXI488a5JZ8Qcb8dCpacmYFv
dYiBLKOtLiOgSl6c5wJgYuxS0SHkKXMN3J85pFYf8p1TJJR04Wh6f1+3q5FED47Z/tQKrKwpq4vc
ys1e5z/FFDf7IT9dlpdmJrfQGGPvvAffNUP+J+CdZwGDUfsYWhyuDPRRm8C9yX23X7GVm0AdJhfu
E0pItD+Un72DatpEvK++j0mLqIY4es8jky9fK7Vi6MUg4xe7SpSJoD5lclxYkxIY9/4m5jVszyT8
Vub0K/dY2mKf5noJ7ydzMkJddIdIgoJ3E7vDG/76Nu+sP2WVPkl8tEreL8Q4DD3eLYrCZCZ0Gw4c
ww2TLGVpd5Enm5ohZrwqZ82Lg9CIH+/Ebvn6ozZND2bvrPAZ6fagaBFinh4aJxAXItKsbXrdRZEB
p03h4Vy77ZsWi2c5zPnkQRZZsA6dK4eZRXZgqWMDVIlx42TRPF31/MZFkZQbW8Owf4sp0Lw/KLd/
uM6FyUNTNjUbVphUNj3C7jxdrcQfy0lerYptyrT0KGyD2KvvcYtcEZ38QCQFcD+vaTDk1Ao+T0rV
OCCwoy6NgHNvl+unnayAT0P/NxMialkss9wJyItr81T06au935siXKSrwkdX8kMiEsi9uPWRIdVa
WZqTLnZCqZ+ONEb6unfETy0cM7BNoqjGvzzTZXzORdEKcQs3rdNw4gqDdNaLMNne8m4wwnrg65Sw
EVLdbmph7KB0O68R010kX7fO9YtUsLcA6m88zky81JhT/lxVNewgcQzCKkTFXZXyt/XrAJdj4Q/M
0pkIPXK2EQ+J4nN9yA5Zs4RXn6duvcWTUL1VrY6BbhpSOJm19tNUnbFVMCHFUPA19+UtCF3XP73U
xDVHnQb9rG/NoaVBktQtlsPk8dTTen+52qr8I1ookJklZxMqwF+I7Syk0O1qkKwWnSXVRjrA1w5A
JTq2M+uBBlgZ+Sn5ifDGgdyT10DRe8WJF3FvnvRkBlAvK35XE0NknCNASnhPRO7Lk0VOdkDYoGgN
0ock7egv8L8jswkVvqAiODf/rpGuobPWjECdc/BFKMulQvBu0uPqNC/B/r8b2oH1B93UZ9b0m9og
8i4GUp7eB7mUVnpvrLxnLcakbAzHAXtOm02jqsa9KU6jGgXWxHi/AIHhCoU9XHzB2GjH10zomkfj
z8M4eNK7Hlm2iuofsEprq0layrpCg5+KhPjaV12BIYI0E0QWLf9cSYPdf/toiBlwctjwJrdjDkNf
moY7EGqXTJRn0mO9AT/aIfSjpC9Rk2ilEnnTdeSQ8duBDez8tImVUEC4E/lVYR0IUrdeLV6kejRe
EgoG1CcyzcAXSjE5shv8UTR/YFiSyfH7MtKqD58uYxU30AM8G5uBxbtitsmnBFBnUvlwaQuxW61O
eOdp0pZC2+QPKB6aglNmYvJQvR9YspDf1t98KcxWdY1nOV/ETxEcukaDXssSyAZGgLn0tTKFH95B
cC3ySd9gDiYfn70/tEyRIfIuX/v2vyYsTj8xchflCoWOGsdJUVvQ8otBTSD0wg6TsOWavlyLpADY
sPEYw9RFASDGVxeCBKX7jjlSlndSaWxmecP2Peg/2zCZJ3E0cVPlivnFWw/myvv10G1udWOYYwAW
isHkoXbxieWQQxSyKhwZsysWdQ7zAowfa3tlPQE7Lpjmw+3CcG1wg0nr2/jeY68stCWHlR19WIqV
CXS3SQP2kO4VRhxRcPvu9Mml4/lefXZVOjNyHDuuz/Nx06sIYHXiJDRBQLxawr7psAE+L/A59voP
rVEK3fK3eWgsfBJDSdZmn4ChMaLG17sXcgvqIXGyZEXxFg0gbY0BRrFtFltDZO6vNdxXKDILmxBC
wNKGsiaccmP57PY+pj2SHEtAwAJQucRYyqZNO9k/ldoCNyeKeyq7z7iMB0mQBKcHFtJXJmri1kHR
h7axcCSDQwy4jes8IrMjA3fZdEBkwKefiZlqYuHFTaUj+7VyCyYPHnEsV4OgZOLya4jG2JbbqFQc
zmVtr9JwCbje4r42uUWZPnCtFbJR0LLsPz2Nej3n3B2omr7TJCsphzwrz2U1isJchjVs+iUxS2aX
FZe2a//sASm/zDnFuwdGBVGAgjS17L37RPtQ/Lsbubp0UO/6pAoB9E3Px5VGPV21Fhao9Iht3tVr
mxy7LyWq9cGzwUtj7S2cxEqNFDRCQSxoTZwi6Ih5mu1EPOd7gXNysyaAwHEmQK0tolUh9Jvd2Q8e
GK/0aACOXtIIMdorAw91s5tsWSbbu12VhqxRYuKNsS/Yzo8H1r7ztAlvgU51wgQa4x/Sj/pTts7d
SUm4gsWv+4Fex4iq4buRO8EN2Rs22LmXP2XE5x77B19tGQ95KzGsOhYBC1eqeRS1cpqWDztrm7yB
6htsmRFJIldxVGUWh6oZfUDnUBpUtieb5lGx2qK7h/MvdH3g82GnHBYNIx84lfpHazsPQNeRNYoo
LToj/fOldcAyMKVOSYtLNVLmNfWk98rEB4ADQ/XaIhLiLdfwaT/f3K5pVyPS8zO2oruiR7CI7JHW
Nggmo3R54uUNF10g5dsPxcHdt1l9LZHx3MsWxjv7ELGJDeGfDg2xBh6gnjL3ae+1VuWKt013I6D0
Q8x4RcMrBvqFKRzkwrHrVS7jWPpcQqbSsUMf/SkaM/373jaxUbjnx4f+v1dM4oyf6zdSc/Aiyyw8
cZ3kBBgUiyxKh38v+G3tKJSjX5xHapuF/W0+BaUI/xedDKZ02sr/07NgrKQNsRSWgmIeQyemYCzd
hxCYFpwGd5fCQfW0DbQr8gCKPk59NDVxierOaENslqTxEOiQG8NmM1GAZNS0O3mQTAPQWd70Vc1O
Y0OBp3U1PGxkf+lqKOdKKhQyW35UCDi1Y00ROXn4x5vT2c0D+eqgt5bZoTfmPTywVSRh0bwkBD1F
7sgkL1irz3O00DWekqM0R3qs0Kel9Io1O1n2WmbzhNaetoM6q/QMgM/unOErRkoh/TxPlz/ov6/8
VJIoY5wx0Y6zMj7s0qLbmM/fHobg4xbkv+gCIT+7qm2DpCIPIQ5k18X3hexxljudE5EASOgkB0Dk
o03+E6qhZAh7ZbQPYlgDV31x7PhsvAUi6T1Xvw2lzC4GsIrnFsMHdKEeT0pF/fLgUu1t6MbYmRaH
ccgAwtlMpTsTqjFiKACWsHFIPcNcj/nSgNYMU33/0FdG1o5tc/dRSj9aV1c+nUm4j2Emuu/1g5o6
FmQ+w9IcRCcKGztBf2HdV0/qfvBDKKCcQVFNAIrEvmS1z3T0m3JRr9U4C7mltRQENktCEx1w+gN4
JoUr5xLBLrFdttOAsKqMmrmS34OA9ADnpHGcVii+UYktpuo/kaItdgoLmdiIlS4lyJC6SpNa34T4
SScTVarALl7OpnNc69i6hYTdzediOBsy6jxTOkWFEqj2cfzE8NXDnvbk/uYIwmMCdiL4XEhboCIW
iD4fBP6CGinsGvISJ6titnnpnLbhJ5XRqHm6VP9GUmcMDAkgdKvAtFEt8lEVXKUWKCX5jVkpJyo1
eLOl7XyJ8yBh3YV6qkyuXuiokPZaR+sU4uREbpqbxL9ULeg1NloP4YLnm6/xNisWpe+YkPAwXWhE
ieo82l3FhgDzHCRmiRDTy8jx00rtHPixNfySvYeKmhK5ZJ5J0jn5RXE/XTrBq0HEF9LAQNPlyNXH
iWcq4PkuowVPNsabpzS3d+IVqGM2tW5rze3ueaDlX9utT5ItlIZ1ydB+ypd9/YiHvAtYwBLNLM6y
r1Tmgts5Dd4KXlN2eFJYCXSzDekLw3vD6rF9UmXBoUmoYoeqVTv676QKAxraaJ5KbQURDk62i8im
qd0jDF/H0MmneaN0+eKpKR5m2rl7ponO8uk8Qxe17/Nuduf+qgDRjauCfwKq1UIp52Qgjp78DY/G
scxanttoXfhPGphiPMM3Vefw6qIk1Rb2N32REFqEUQ9SBNdGyX/6rxIAZeZnP11MAiD/JUmZi7sE
8OlBIxOg3tHzLiWYwmCfS94oPGPe5nyXAP0S2drmq7r8PDDuGXBi+J+C/L6EHM490rtECUErku/p
sCyElAGhyeMz+eLZtGv3WaHy54zNsvVsPIXOl4HQsLQ+FP710+EsB3HkK8fCmAjHg0+8cC5XIPsm
FF7xjCrYseHzZY9n3TdGXkOB/YyGltpF6eRKpWOkYoDvZh5diA1jtphzXCxhxDJ0LGxIwOa8Ix4x
GJRdwrJV/ZDEoaGNypQGlTndCuUWc5bj25k7smk2769hM4xbpjT0yWJ7FpIG41WhIa2Qh9JaoUCh
BjfbFbpL1LkoYq5tshhqkpqpqq/bweO/ayn2AJvAToIKv01CmSytgE4xKch8NXi9qG7NbW/2kzIM
9hTotIx+6Iq53TtqPeS6oLmlAVGEg1b5josDk0mb66LdcI06S0lmy3QtkPWK2exik2j/6cKPJ1LS
/8WUEUjnjqv1J5njZM/9hc6CyrNgjbbiihv9dPS9ljzLqPBm06Mf/G76VTbEJrqgquffULJxf4E7
cEIPwkGDPIN15mqKb4AYmV/5XEnI8FtEeu73sFIQg7NhFqPAySpvrcRQpqJd4ZWo95j50G8UlPS3
bM2BOPiRgwOTzbbxlUbX24udU/i6H6jd6ETRDMQrpIJbYdFKMvyLifYwOX+l5HtqnL6Vp0flA60g
qv7c5dgHa3NWFfGvqeE9pL/Ok2YvIGOEqYUcuHvcx2QidGQMdg9f8110jxw67RDxNNFQPwaPE26r
dTA/yY31hnJ3hqQOxDXp0dXn9iksX46D3AnZ397Gdph68RtXcj2begS0PU7ZF6tBWYclEsKOc7SY
uP7zVORugg4K17OhBGjhT8oI0ZOxPFO7wVOLgttEKRzQaP8+gpNeh/75I8/zY2AJFp2ewyew9diA
zUVLgZ4P8e8LZFAytufUttvb0DqosB88A2rOznLbdkKhhdpzUKkT3ezjZfu/pQ6tckkdF+otdwuF
/NPCnQ6nXGoIRb+H2nUWha2gYhMzAVj9GGLd/aBsI87DuuMVlIZ9AmFYJdZdisdoy4/5tzMIfFJ3
wfS+zB7FkB/Mfpfd/UlezFicOTMib2MyOKACjSLzPyOhz8ACiKPaVzA1yFLCYH2U+kF03xdCxoov
mYUHlNs7w6iZbqXzvBsGpZnzvPXG59H8hnJCSHRuo31tcgbS2U5azHrjqkiKtOJ6ieAAXudLWnfc
lIi0zyLoUUpCN1EZhxyzEajWawRuLufXR15t+SA04N/xuEbQpbV95hR/MM/FjWjrxB6EOotCe0yH
o0SYTFxdHTInxEWSLWNAxgCe633Nq/3lUfvM+KZ6fa8i1H5iD2LVYdZuj6YXzVDFu2aqEAHsZWBw
Go+DqK6JXKOELI/im3FJ4fnVaW7A6reH1LqsWN6wm3vpHrVWtwjihb6pmvbRwAwlhZ6OOwKYoiDy
3GgeTFyjGTqCxkGOE10CvnSe0yGHlLJ54BKWTWA2Z8gxI5gZ8LvJvPcq4RCTVeRj75nVscH3ZLHb
Nq60RoKiI1k7kvk7ksUSNNf7Hnz44ojPFbWNpwiFz3sPVyHNqrTL8AZud7a4/zq/yGkA/2Xi4wdo
lt8pwq+Czft2F2WmYz5e3AZJTZXZhahZ/bOTzJDJf+QcXtCPBpPdhBbgJBwTwyDMsUkJEqJ9lTzD
nRWe2Scsgp7pSUzd6ssxIhx8fd8/mzpseS5XGXdUzMD5Z7zdhlglITvHWtekkWEwHj1Lxfg1f3dj
jVMH7pp+2dFyyS5yHeUE7I/+jIbR0th1WdScrn3kc9EcejiWxtW8nx0Lu7mpsGmd1JMFbw1KvHh2
TMQAVrPtn4pCUDszgUuT/QjxrHc1vrdir+f1RiKM4qiUEdE3T1Or1vhKjjTYC8ToxfebJlLgS4/D
9ncGao8XUpWndi7nog4+amGD9821/aFlx3gltA8EeEv+N2DMZlkU9yPSAOLGLG4uxbcgHKcw9Iru
EDSCEqsOOX0uPbmQ9SiBHMYHeRF5pOWXpF44uzdZ2aZZmzkYG66PrzQd0vNHOuayGH1DqZmc0BT6
S7CE0VVzHqGTrclW0ke/eaGtaTpCZP7R1WNXHxm8+91Ub/CWeiK+39QuLtsnp2+3odO+1AB1AtPt
fMQtXdjwmkbX2jnlcLfkVnSoJDuzWTuK+UVw8L1FfIivA4ZoEz5ctCYEYtUxZus4VsLs00rpTsZs
ydNTzbgjFOczxO2zzTcJ8wo7zSKEcEfih0CMtvOwgFtRoJtp0SgSqEHdKFA60oZHqckTc+Ua2905
PxwKd1d+N2+ru431IC0EFxX39wTUlaZwOWr6aJdgL/Vi2qIWDnkz3JGhp9inMRklW4wxclrPaGP4
6mqOfA6FwYa9gkbQrVIUFm2+j5eP0pH5LW5v9iEHSPBNeWbv0M2wVRhhWnrTEu7aZCdJusIUCynm
AqXR+JdWBnkZGS+BLcNYR4VKdkv4Bjj2O6gXHdWp0xBhOoJQzoN60HFKTpxTU47PrsuiWGSgZGd4
a2BZ0aFas6l8ugNeJkGD8jiIKuitk7Z2YXYmUbvCkVPGmk4xlR+2WBNni21/VYH2wX0pbOARWJJ7
OBu/nKcU95cT1oxbawWeZmRC9mPY2jzMxMHpQLqMxo1m/Ro9yqsfDDWyHgawmgrdGCh6uHM2nwGC
tUDsa1Dzw7yeeFsylBq6rdTxSioOQQoT1zLtvZrbtLNVtB3Q1CRrxxcwxhesD1J8MLihA23zxzNq
Sv5PSLmV9T/N6vQqGAewzrIgIGi9VXFrNan3VFFgNxBqO3SDIEFhV2Qrr+QNqevt6cImVeZPufeU
ATb1elqEbxrkv0vA4J1oSeMpIRS8JRhxfmQYW2yCVrh9uN2kimfeutcghK1lDfIli3E0ltsVg7om
0mECBqoQ7HQwwXOQ1j4RJaKtU3nBpojbHatAWgCeZABcBzRNbhTvt0BcrQFy8ef6CNGbRO7ZgmBQ
PlKlA4xJbDWihA7KxQZqukHMZkXTBpByJg95Qh8bJN45mFQFSNQHdI3e6vpwdsFUBG0WilSMj63F
076Mputo9IYp5tJGnZIh2x9btsOVB/PqsQ62XS/JJq1O9sXUvN7VSfyiWPXAALDDzjHVigb88Fhj
7FcTj8+bwilWGDxbcITfA2LGAcPWS909mjhOxHJZx4QO+qb0j9MA6lDQ8y3m+bFggHlfo4cOYSNO
GzgKjvhXXuZrw46u5T4B74Yrikg8lI9Nsw/FKMGFzem253vZrMJPhbNTSv9wFma2mZnRhJZcl3X8
gcHbqgf49p+GEr4YdUiawbwOpIS8yD3a3LHVAbyRmqjJtG2PAe1u5nFASMhuuHlq0F8XnUs7gy9K
kUsYl22/DF3tS7vPNRhZYEt5z8RrRzJc58wUz8iqdPwtMcD0m8mO+JUwSVDNOdVzZWHBPVtPWsN1
JQMcYxwCSIdDzJIkixlNstPqRlOL80AYz3rx7YSrtRLse1jwilniTnSr9Te55pnX8qUFsB2BRW0h
bMjlpoXEM4nezhsGaEDruoMXSovAfKTA3i1+LFmPZUVdObtBQE6FXHbr+BVmPNNzKNnbfP1Qq4DW
ZVTWHEyc2Fm6x/lLLQdsYkfWZnxnmvI+umBShR7Yf8D2spm5Lb8Qln6+g1LC7EGK5ndc6UH35nID
y4fPhB87Ows3AY3kMqBKkpgwaomjKsieO22TKmsXeQiRX7dflSdcdrWOm7sGD9IiK8Kl2ZiwcAHA
EGJhjmxoIdRiykGPD3XS4vjfe4iGKTedCW1IwBEHttwFFZINBqqv51rOGGVA8zfPIVkVfFsJ7hG0
F9sflALW/2ZksE22qHHiXZYz/Zh5kriagb8mhZVv9pBW0QV1EbA45Us6lIIaNpCZXyOeKJsNepZ3
3wuRL6cnbo+ZPASxRnxoExMGu63YJohuzNQ34zXgwIthNe2LBLsKimpFczeLIVkWp3yQIFEg6SA2
MSPyhnK9IZjgz1lQ1SqJ7Q+RsdP2lnjmBpEPzliahgUfj9ggqPO1RVf3xOXj1KJL7LdqnHq/yRBf
XOUFRaKeBv/4zlreLztNpC78pcS6DMF8KXOC7wEwyye7onJVc0luR+KzZJtsyythV2HCAXz7Nvbl
w2usehcfZ1FpUAiMtu5wfxBQ7pxyGWloLHXepvcLf7Wds+JRJttu8M3pBPNZqM2ghcYN6KSlW4ZQ
EP7cUas6KGkDKT15OdPmqMtzaYsdGcRL1meT6xVaU/uLXdK742uAvu5lwvVRG2hg1WnjdyqdtNjC
RXEvmlNKl3G59ybOGtksbFu9UjSqbthO2rXtydzWrxVIQU71IM3LJaX6joybbU1QHi+z2diu2bin
1x4mEt3X32GeuYY+HgjutBEbg6iUHzZ0yYUC7wM9Xj7thRqJi01MduLftL19PjaG0pIlFxHC/fQo
A/vt0HLmakG931vveTzlWToM3cBOUaIWaFs/ycmn2oSaIJS6jRyxPnLz0Va8cBeJWjRrL5cGGtlg
jwZw0jT8KnBGNgS6P3QNCi1v4e0kvwsPGsPUxEwJjp+hO3zRzyNKdWylXMu3i2m8MH/juBCfsuH/
8JmWdwzof5n18X+K8OpUYFvd41MYIIWqW/7SWCm0hqJ2zr9gkr/FPyGr2mxlLXpzC+xpePkxGAdU
EODdu66m/lSOUmswbhv2VtzD9T7/BL/C81hsXglrIDJH7Bi1K4FENbmwaCAxeB3OEb/JYCw+cjyx
bHRixApV7Uz6gTomtds4g5ho38M7j2m2kg1F9g1I19h9NNYCSwgbbTiSC0sF8W3gkI5mD22r5L4X
2ft5NhfsyWmLhWbOmmuMl9qkBLxnhKQC/Z1fGXRoH5MVbs2DC+e/0vNlHZPl2auPUOzViJZGduXO
f1omQPZ8P+CqmV80IOGnv32CAFILPkWwbkqQNp9bF7Ck11hZJs1GWkqJfroYemNIHloOy/uzWStv
VVKzrGfOhB07BHMIrpyysWlrNsxgqYdZdENR32bvc0pNbcFyAakgqc6BI69NAL9dVBg/O3Y0h2t/
ePAMvGORd+GfTObgOfr5s8LYusaAp/C1TQQddKM9QhMKcEK7WByY3mCEaUUwDBwt0JmdBxNnhsyz
z5CXeKal45L0s40PdfKV4uKDMsFwCaXOt5RVuiEH4BRTGT97CvypXmlo4qiKBxqFQK7p3/F5kDBD
awauX1287cB40+WRgU00EHmXwTrTuGfUHNgiFHR8PXU/dLsjd2LCQVYMZzlBvGIuxFEeH19j+GU1
14ZY8drqfJnMBLKnZUkABBgDRLqx4HxbJ1AQSIiwQAgcThhMf2MQTrMQ9QBXG1zAzA+3jXwRe894
oOGoUSV4uQI6hXe57OFthTaHnM20ZPEC0G+gskPrbnU5IRiN5m/ErThmYy9o+yZinzh4c9mCowBF
+pmCKqqaUHtmMFyBH5gTJXSooMFJg1xWH05VihCcsbgLGM1K0jI6MvwHkC3Nx16dWN82mR7FdptE
o5tTOHQxpWwkLwneeKwnNR7PPdPHQPBTY4np0CA/A+QKghuuMzqv5cbgr2nyAfg5oKpPwSxHQnrz
+U2iJ3RgPb6TEXZHqXlE1Ug6U2svmd8FQ5H+STysS51OrlLo8EK77QmXjaIMWIy8h57DJL5tmvh7
3tbdGBUn/xYWNEp1TICo6ZMbiFFQ7j/uOgN+yc6gV3AJhuykkdw4v/9jIhk8IVAqdz4DmvwRRF7R
znkZUbNhzQUErPoGGJc/szmr3LLKt8spYAPL+pCkNOaoHyAivhpXv87LMxa8mlFTpN9YCWiYD1hv
7PKJUrGMEcs5XISGTQZnMaSWG13mvPBCEc5sQWDBkhXPFd9K8S+NTeEjk6Qv3a6DpPnTPjoxhAzZ
BK04j6h5CwZPTmkt2cX7sUD8ruv1cVzoK19NUQirgYH2jb2O5g1qKWJ9sYiveOOzxWXtxcyyX+Fo
nvWX8kFSSQwb2Nmh4DOVyjZQdEIoIa1tQs8yogkbzhC/ehK6sb2jU4p1zFyESLM1U3Cr7q9R2tPS
PdO9FOl/Tg1W5HklDN9w04FOQnXCSkwsFeBi2s1LZnZhAI9w2jB4rJkC35r+YipQcFa856w8qWa1
F8K1am9tGPpITXN5QnCnaem6xgAHRVyIBSoYPA2idIDDDJijRziMMFV/35Py5FJjHn8DGS82D+tC
4/+nkxdljqM9qVjt4hC39CbXwJ2H7lxO1AF5MP4FuV3XrGeo+P7XKv49i8tSgXFPVGfzJIxJ3vLg
z5+RcN+G7SmLCzXYyIBsx4jnRpKBzc2v4Gc+iwXUpwPsfCGKWgI0l9RoiGtWn8rs+UO55Lj1SpvA
yCCEWWtiYUb9P9oI6tMW+NvyumHHR9uEs7tHdmalQMQp9BwQtyqL9Pj3cI/Mt+wKTI4wSm/5Frkb
2nUNHbl9H511YL3ey+mvwUTjwDuxK5FzdE99/wC2UG45/GgKuivY9NQ431p6ZmbIA8GTRI9PB7Od
eMWn/2mh388a/uq0+uUqxF/bEUKlIwbycEp3YITjAPFUZ1Mek7keoniG6SfqVAg+bWcn2CnKA/Qt
+MXt3oEOyAYnwnHXhQWYVx/Qe+bdSCUm9M/7ZAzNELbxdPDFAZFa6g9g89YeV/Favh7TUncKcWDI
NOByNRdF8bYdH1+027NWJT11o7vl+qzjz16iyYBN15Rg1WJs4kMY9L6g+om4NEZj6fRfCgKXhySL
WFWtUkfpkFKQ6DGPzk/ne+k1XGVg+ZKMsZTGl+EaWjJqkiWgqDjmeeb97AGHAZ5AhL2l5mRe0i2O
MaDUCZSRbWMv06rJvwunhhiBMnRs7FpAQyQq+HHVpN8OY3VyqGIhy/3++THywDt40Aic41UFg6L9
HXaXfpxdYJSrzD19FIlsE5a0bxaqnoB+sXJtJ48OsIFsQo62bwIAAQeNTpDxW59XqDLZYSj5czbv
l42bPZXCr0xOF/xFE7hIlmL04+jxIWByGgyuALfRryhHcvaldiIdk3+tSY+Gi9r9wkn/M82MXPrI
NsvJuh3SQ6qTSwwWXQ89SFqCr2GmncQll1fULZJPUTfCsw7TJa3iROLUzXW4UN+wqlvD0cTJPxE+
WJpWqEZ39xCcL92jSW+PfAKFim3rMw0DO34heKln6OhGDNfpXAgbNLX0Gf7A3XylRW+U+RAMZh5b
G7rq/LaSyWMlZgLXhRwM8axptMRN8kb6tu69xXepVpBwKaDkyCNOKHN0MavFgdUqCRYZ66JAQN4W
EOifYcXeJJ8577q/DSkvcAYiG+tZBuJOSJwUgTwZS6YWqGWYDu2m1w7yaG/GzyzQC29v8OiDhz2k
8bCSOUdViAqBZ031tKs6xDzw1s4cUhqSD750ww3bfjR2l2bDdNiCZKQQN8EFmChor6qkTq1iZnjm
gszKIRMH3k0KX+fwMaaHsP1aun2AzXG2Jy2NToaaNHY/okFOwoXumVpVhpvDyaOgDMfh9qIeELHt
tJVeUQFu2xNvw8MVv92AWkbRuNo2cCLcMIcopKPiE2UP7Lsgh6kN8CJGKsig65rkYfi/hknHIFke
SQy2/ejvgF6Dr1+arIyLq9vvCYC1NnF2+JYhRJDPhwvkL7a0zl74LvrnIGBKUnl5/d9HSOtbUfeX
FuIOdRAp1VYy2zLOl5+iPwtxXzw6jkQNh09NUdtEFShQmfgsOq87YaWL/f2XzbQVdGVMmgczDuR7
i5tNxe2RRLP6nKKkpsw6bjz/7sXvqqXKMTPqMVpHgUkoZC+SNTX1qXpw4+pQGHh5+hzxs4eVxuVm
T3BGON5f+hh6D07DRtjItaDU24Tc65rTveg8tGkdlxnjil7SWeCJ9wEzRy9NHNXTp0LFm6PhU/rh
ToTk+UX7iwxF+LtiYvtPGC4Wr0unSM19pb0mJ33XpX0Qxu+WDpbYpKYr+XTWR2GK7IrmmSfm/4ZM
K5v5OzrOqImhAfx/apb5PGDxXQZFl6D7wbKe1DcT3kuM+ipbDmpuYtVE/Ho8e2oGrnPWnPGQYgbc
fCWeM0YefBxEmphNqkRXOSHWlCaokZnhzvEvvqnK1GL51oCOpBfEBX4CD+8uK42MpIdy6cEmUXKQ
gtcom3U94HSeGEVfcxz3ZZwh3bgE4VBvWG7zat453g9OG1cGv/clXopw9StpOZmnxjm+4wFf5n+O
cXUsdRIhy4GFJZ2zjtqpoM4nKrCzD8Sr7XP29bRGKfpkLNcYjqeCBxoeWfuOipGpcdKTadu6tFvV
5JOYSQAzcW9L8C+m5um1yrQ0lSk/kD4flDQbmz8+67IYvgtsRmZHZlyoxrPmPXo9a+Gv9Ts/tP9b
5v3yhN2dZvF7KbKuEY2OaAr9x36HoKSFcVmc7Nv2RGYf0wDd+nDMvvviOjw17QKsQlS3rUdqDrdg
5NfowU9t0mGK8/6/zxQ7yZ9vNUDodvkBo/4rPF4/akdx4gKyOqeWWnRxSxrgYRuVZtmrF8TsIFQf
FAYEOH1VX7QpYbaE7VbgWtTF5diOiFfaO89Bwb5VBF2Kt04YGbwHrvCJsyj9avkOIuDZ1FQEEZ+I
fw8TsNYEoMd8Hrzkg1Br/RDPLf//ob4m+EuMZUiaJc1P5g6/Sk5C56lGyEDU9EooV3/KfC8hk0qb
iNbreoGRD8FanYaQfEtQ5eihTYrnWwkIcbtkaY3inBbe2gapq+5swY+Pk6e77f9fSr36ygytgSqJ
Usf1tKXwf00yl5TIRkdN4xDYmRZkp7Caph2dISUwfnlwScWBwGfi9KWNk/BSQJnJ1sGq69ueIVWO
Ueu7f6Fg7NXy6zyEJL8CyfOcbVVx+s9iyWiZHWrTOGT5MjRZ087bAcxwsx+CL+5WzjEfJ05QqNiE
CNWPzPzVjQAv9DEwx1pcju/2mfGZJybl0rExPt6sT1BC9djazlN1wmwLBx1DwosHRLWhhHyDQmxF
SKdwqJSQO0LgtNCliS2Ln8CqDRA+feroCVafksDQAv2qGs0WBjK4QWz9vMkBEqi7QHWKqpzeK61B
WTBnvjuDedEt6gXfJBYM6QXck8lDtcq1bwAzuP5Gc5ObSJhGiDROMH9AMq2Xe64qHFg0LVtHfr+2
mz4KzxapLw2mwvho5PZ5KyMFRfh1YG2EwX2BWHnQ9SHgWF0Zy1x80qa1UuTEZJLctyzlJLiQkQLz
RSZ5bikORcs50G7fA9rN2UN1TZ8GE+tkV97SGeykx/xuZCBxEuU6+FFydKCF91Dh+6kVga7rpOQk
I+ylPZtF57KCcD2xJbxiIkqLK6GUIz/Qxc0EJnAzjuEVSmuc0FHthsLkoifcDb3eY+sKFCon44n1
EYHM1dlNIPMzDPEwuaG7xtalKyITDdgmwa3Fw8l/pcHNnBDHjWoKtGmhUmke4fwhRqcrWtzO0fh5
Vv6CWYFTz1eVB6/OhnK6iHXT+bhWmKhLAebSEBhGo/f88riVJ3bdsTR4rKnc083D1ssrGWhGZ+XE
2Hmdz61SMdO5jDfAwVueA/IFxksd6PiGls1AhQznW/g26JCSLtcELrQNwJgRLfBKhkY8/knA4pjk
bYQI/Pw3ogR+56xkmIzI24xhnDB0R8nsHdk/W5kbiIHuG0ZGk76ZcHATq2UwNvbd7qD6Ok0B/cKz
yt31en4O0VPtv5U9HAhqXsygWnoTOXmPcG9jm06ELmqmj3RYnHblcxFgExWrYnbSswYCZtX2+YJi
x32E+ictGoOEpNKOtrgX1FGYD5R/b7HxROUnchqq05cfIjYUnjy1ryErh/QVxvV46AP2/gYsv4DV
RXdDQdDBIF3RJOwQF6qFx9dFSar1mdNJcJu6KO5rIFcEVkzsJaCw5ZKD3XYFzOCtCWvu7p+wvfCM
cMcj278bHWKExE184PSMYYSn5+auKSsh4xsidhqamK3wwgk/ubyXnTdvV2VcO3dVNt4iQyVN4DDW
l0HbJAG2Xff/yAAruLFJaSUAUjSSU0wHZ/sigP3vv+O0+yYhy2wFOO8S0GrFReLvSkNm2pYzlrbY
dez/ysPEi6oRYkzMDZDTuXr/csIIvGzyW5ZcHwwVSbtQKzc0i9FlJOVBNrdyRStSwOAQy6498Syy
QhsiAIS0euC3tOgO3G5f0vOB78qwTR9SA8nPTcAMxrtoAR6doObg7AThrgjOM73pIVktNnki9Gsd
h7jna3uL4Jd1IXsk6+kZmTqOg8hWmSQr5orgXvuLnryG3WaVqsNvevPTYFctscn7Wy+Tv/FFyTK1
1vrMJAlbIWnve6mQapZEaieo8FKKlH8IEjcff9W6/8n14XJEfvRpWHcDm9WZOmD8PuyFDIaL4q/d
nSEgrc94dY6ynaPMj7qVL2vm6Cr1+31RGbSzey1phRWwZYPOwdQtBQLTb7X98vpcxkOjnKgd/k3C
oGZdINdkGlONHVpfor5hDI6PZyp3283rKHHypoef/fhSpwS1Id/yoEKVaU5CmXb2v7lBRpj2FWnS
tLmTI62wxOEUxzohXFj1Q0/kI+zyH0Y4zCtuIaRw1xyYhtVbR92Sbncu+jOoolHEYBHN1z0lFGlY
YkvthbG8JDpozkVaSFXIX8PWFJW+QSqBwZv0Yibbv2/+6w9L+w7xfYComt0cSelLCQ7/UNDLHX5X
1NZVE35DGoeyoj1N09zhzOyRQCWm/B00T6b37YhqqyEhMR+rCL4cuB2XqTMung0slC8ICzaCnqvI
z3A2vjyf+NX9ShQGL2kF3hQcF7qCfXvHECD8WdPxhYgoYKgTYhjuXafJqd+PhWhdyIc4jSMobjQ7
YIfvPbq0q0P9NZic5/+YqnEn7hVD7PfF0oWgqxurTYRMfQUnd663ttqj/a8aTFwL0tdSmOSm9L7W
EfIqSxE5b0Lub8ECD29a61DpIra50mqUKnhmUZa7+O1N0YZG22DvP2am4pYQCnaXa0WybFAJRW60
0kwlWwmiu4rZHh77pybuAxqbLpuhj1rz1isaigQGdIwpO71FrUg8tiFydJKgMB01JLCJ5e/FFB2D
Dc1Lhsn/oDI4nNwjwS5twstc6ZQJKIqAG3Y/s1uPqpDjQBDf4cv3Z8pWuiZmR1RLwIDIL9fNCMvn
9xGDAkfrblrMUo0oK5TAAlGF4fYii8K/ipOhgLtOrKpDPGmaZyXVKeRUkyKm6/fCcoVVSTc2Cd12
uZHfavIMctq8Tgf3tXFJefdk+s+6irAc+vfLZpFdh4Ke5fY2l9d0iV2xFMKJl5gbe00MjuNvGFR8
9Vn3ZImhy67auXmneAWRaZ1wRf730dR2CE5Mt3O88lSHSQlQboAgYRC3g1WD6mrrqebKsBmhwqPN
FU7CM+oULwX7/gsGBSo5d7SeR5xfMsioZZBomRGmm0U6T6NhJxcypw7znOMyJkLvS6dxDeKusw7Q
YzhnL+F5WOh2+6ZWqJcPek0QnEmBSwudBPgGLiff+PcbVGNNuaC15PvGgAVdRVqkmUl0nAgSmmJU
5EqN5a+ImwV+1D5XLdNE9Hemla7Fz6QLG7fcTcfDhzjTz8Gmjm/Fl5TiFpuDFDrPxWkqa8MdQmuC
Fz69jhvX85WPD5hsvddBUC6nY+FuyvfxILwM5JdPekmZz+PFS8vgUygldEovhmGk9TxSsuweRy78
zDWwYBWa8XmYyV6/2k730bVu7zmGfTaXuPTfZ56bUyFNXn1tMAAkO4lVImYKsR51/wkGHxSEaWXO
aYG+tg7xQi8vDdmRMHfq9dJOUdUDd36jvnI+QriZn5+LO3QhPHuyvpRsHwMOfdxDrsNO4ymI+UwO
SGzh2A68yzo5n5OrQ26qF/lWnLEF0m9wX5CA0j+Sry8pDmh/rLg1mGPn3dvYZq54bEoTK9kZ8NS9
zjnd4fWCI/4l0l9yUuGSyk0fiB0wMnhWHJj0FtHZC/MrfOPom3q1QImof996lt7kIg4MNL5uvOzk
FsZuoCzCGWjU2F5I2jL8V5JXQD0Ug4+KIMR53We8hYpsYrxfyYFIugyGR+4FwkN29FHrqp3EVAYw
qouNxuwqcWByeMWevz4KTcvxIV62CRP/vNHpSYJk2VThjM/11JcpFSPSe4iwW99CWqoIDehpI7rF
Id7KpaV95TW7LVGVahNPxl9iWct+FqpHxpUI6KVngCILJ+57SwS/ufc5LZueox3UWP4rDpF5aJ/M
nQzuKDImjwLG5bc0xg5QysEuyTgZ+ydaPOUq5YzuF6Gm/gLmhzxCaBqCmYqn0kGMgR0OdjU8colW
pwJQoMlT5qQdnFX3iPM4b0Y8lMxaD7HX4+yjArqrheJryCpmu9FdJi5sAYN1pptbn3EcaaLCssqy
PMaxwdJNJRHX3xnG21T8mY+TQX+OaDjhjJeyllFRu6Z0YvAs++0/NuzZuePXNZ3sQnetfhSVPlnF
hMEZtR9KWDlKtBr+tAtFRb6R31q5adf4AEsch7DCARpib7x2SBli33kQpj0MMU3RmTuM4A6Aa5nl
1acE8moH53/ZVuWTBVmb6qnIAOyXS3p0/wLPpP/uKlCSCPI6RBGFIunbeCOiTkS8fJP0/gdW0+Kp
ZmhfyhUAJgMp1S0mokPwW5hYwH0D09LrXU9WPFfUFbGU3S6DRoP6/M6asZX//izsxBCvDSADqC2I
NRbpfowlm5Wc5wcTE0woigqNQ0Av+mTUhcb1IvpeWuDJTzg3sd3GL0HiKL2aqRnzJ9Qu+2szA0zt
yrBS0RnpMJa9clteWd9qaNxAJvD+9ElBAe779ojKPcwdXRNUWPE/9iCjGyP96O/Y+Go3fEJUAGyB
E2m1AKNfaTXIC3l6QvDR2m8Xng/yBI+KehGoalcPsaTt9kP5Y6S1e6hdrKJ8LURUvfkkmdPHkAvh
x2QRZwdgQWa6KwRy2dMcqynR/auSRDXgcDl9d1yyC+O4BBCHJPyaCNlAYTQROs+hQXK6hzIdMYnn
+O6JerqE6OKigcMDpIRAxaXCZ0Kco8mv68XZls4kd0uLpokaYAktssSaYqfH9hpDPXOIppVcLJHl
4Z1NUamjoRHywKuVbyKjq6MB1fDjs3ee6qa9MROJ+NiudnKeu0XsTjFNbsCXWA45i+7HdRS7pFMn
o7xQ6TVHV3RxpaHK/QkiVIb/wjNMiBMPVwaTnBuWfooUi0Z501vjzbH3BXg4BBJrgosN4aVwpl55
wkfC0sgThzUeEUxZ4VgCLH/A8N/YcbABRNdemXq6tQ7ZuWHrBc2pwHtONuanJZAqsbuvWMW7sorx
dM23cQNckSMR4K97jfhGCh10rduxeT8Xgf46/Ezoohuhl1YjnYZRiFvWpr37/8vCmv0+ILiGIUAz
lh7p2JYrOrPVLzplWYnmZUPNmh20PyFgRVyOswV772EWu99K7GTJWe/FfRiTghl2zitrGsMi31CX
UlhVpm/5a5ICoa9Zxq9zTjsPLx1Evq+BasjF3Clmwie8cxdFgJs5eHinu3sF+QevsJJ4Ia5yH0hw
J6FrFBCXf1zcbiObWs6r/cl1e9XgCxyHb3qJTUZhHfuI1AwLuVDuncoF5Ca5i4tzBwzLYtHqwO3B
LLjiIiVM3X0CTWDloC2ddQ9ipiL0UvBsayQo92C7ZIrRlA1AU1j6x4lxoixHYfF9fa27NqjA4lwj
f/apsZ+5Coz0aZd0SZ+bTdMJm2uvt5Ambj9RsY9Ri9lNpystXyj9qEkozPW8gQ9GBMrdK3fXVELx
k6HbdUw62BEF/PFVaoa1j69/6noQHMNoOy0cb2QxN4lSug8z2+GCfNcQe71FZ3lQs43bt4d0a948
C1/q1DypYMVYcLS8cvYwIVzWHPtOSxozX+ny3ad8PhJrEnF6aJvy7xqmhdzRN98/Ffn96rgOM46j
a91iOrICiKx85kcLhH7l0l4YpH4pzMoouJMBs/ZFojCmb2bSKHcc2LY79WqtBUV8w0WPyf18E5tK
u1uvGBZ1UVXUfAE7ahpOVJz2kmMjQx+l1Ps31auiD0u97daROV/qkugTquOxyRcSggr8k4yu/ppH
a5mEqg8Th1rjiB2d/uOy183e/SO29QAcJyEX8Yx7JT4qYOXlAYsrU01KovGXT3UXCVOPqUWwAAt8
hjThgv0Rz4lfP/v7Qhv+FGuYFdqXVVdy2q4dy2HpzLN3+2jSLJg8oOmi63y5eiopp/v2ItblqL6f
Ir+9Cpmx70nlDC9SRpjcvN39CxNrSVJ3eHT6VRz6jIjdkhx2Hp0aiQcG2renkOzgROqvOaWjS5F0
P6hXvIrYFGk0yp6fHmWFh3lsOD0iUv/adZEGxiBAy1R7hSHOkW1bHT948HSSREd/OMFGQRX1y8H+
YcjLRMN9yw3zc4nOgf/jhBLyCKVvF3A0hYV/ZsCn4MIUYPmnQO13bzoaaAlno/zFazkmKJ74KwXd
tmdY/I+8aWLmMnjLBWVWZEbUtB+VaN6gwiSpToN6BYXtQdmD536uPpuhkdsurbESO1/Wq6Ps3Wiu
yunbUec8mZG/SPa61mSfqbJ8Eh7JOtq1Xsej/Crxmmr70Ev75lon1JVbm95DmX4c49GT3HxUloso
c3mDvDsyvz4jlJEpO5+IVo+IdWjMXJ7R91BkUI9yvvOb/B8MMCnqmm8P7wZ0WxSFgNRz+++2WmM8
TJWf8htPkNq02BTP7lZtCk/dFKgYjYGXYHjgvmwsVqnEBOMi9CHaJjWF5qBfTCW/+3MVu3mEu3Xo
ycdSYD77nGNAUPqc41137wGYRrubCVWCFCQVrLb6mshWbn/Y77Rr3qt7ROpYRu6/efewIvchY33G
X7KN/2Nsh4ZjP/wACJYFzwe5g7j79eDKEV9aNhkj90TUGTB7FFo2D4Clc+VchgmYEQT82xQFFNe/
rNLRvrBKhqcjoRh6nA9bfj30WFSajW4vC/CEcZXN7Vmj6s0rk3gR5bvNUDJaW+VW9iP4MZOlFWTm
3DXsgtSH5xs5HSLXIlWQRkaC501mc86+oi/oayvG1NIPzWwy1fsRwXK5WrJfpC3v3lYeulTKWTzr
1+g1TZwAuv48ba57aocFHCknusktjQze+qk5RyTPDzBLhTr/MAau22ByBh71oxt4kIdGveQ4USKH
SZd60+r7d33/C50/NzlCHZo4IyUmALuElF9XdL3+IzFv9jGSweN0fSSPzmisch4e06nbyRUEIdAx
lCOgRMRp3c7UtTZQvDNXX7V6fuIKRPnJS6uTJv7ESIS67WPuD0zh9l4z+lV4WGT1+i+cLv/12jYE
YD/tz9Bw4Lu/7egCgKxjmMDdhrK+NNsbH+fyAfOzH6db9jcTdOywC25AWPXyJmh+CqfCCQbsIj+R
V3ZkVryW8vLPLvx9a5sFZJjyMgw59iVOyzDfv06BLDBY8cU17cLzFb8jiE697rKrEs8JzjGUpy6U
ulOjp+nuAQDj4b37Ltpk8ePswZCkVi8yPNzyzyzbhsTcn6Qt0xTxXKqQ5TTUKrMZNLkRfUtKs/2C
Evn/RNlKKJpB0A1Adv+h57MBu9zOUuFt9792AbwUnrDpdaaED3HLxU/rvHZSsyCNDgRqyfJOiOL5
xYbYgLPLBaJfRcFwcKBsVIxJ85BMOugQZ9lWVIcwD40LMIMMNPbAP2cktZxZIfxngU2m/7YGMKQn
FpJEu1VUPfGSAmouMAOqQKi8pv6APCvQ3J5WmMWZk9Ld17aXO99B9MIUBCZYHIVO6d8BulhWqpUR
HYclG8ELEk/Ok+/SbKP+pZWmLplZyVbTwt/hFcZzXOmChSN8APs9+S7LQWuk9jrIXRz/6i+A63op
aUkJvZJl9JSAHEJoZS1m30GotGqFwhoGCd9Q27wjdwj5Xs88TtYWME7fXoTUgViYJ4KHgRZm94PC
JaQmwR2wvuo/drRfiHdTrV0/v/9GRsHUsla29xpl1/r7JF9RXQ49Lnk5C+Z2kzkcCLaoc40SDVRP
7DMWyIxvRzVsAduBwooFnLUyK1HCMb0J5GwRKNqu9Jh8ETQzWIukeKRIfSl057w1PdPojP0LMvs0
tuPQOIKuaKQfK/EjwZqPcZOp6kWLH6/XqGkbfRa0vtz4miavFWSWaeW80I4BE5RlKQNwRo0+GN0O
SBPjzJ9eSh7Oer+HfSGrDv1dkk0kALypcgS748yMVJiM2DQFKJgL+nN0x7/mcc0GVMRCtENjrz2P
081nE8Warzh384hyPlS402frj34401X+D/exIHxCvbftQAszd4XIR6XY/IRR34wy4AWPNsZ3MnFr
/S/WZc+MIx5Z5QLCkbRqSwRD3LL43lhxfCr6nNt3QC7ttCYDM3EHjV/ivzYlopOFlDxPLo+KlRvg
2jfy2bKbXUuGw1oAxfHvDd/xoVk5/VHP2xFEbpckuzrwns1S05l1HHRtr6nS8qkwVTM+Jzeua9IT
NnjL4wqL9q3te+OOA5gjDOwfIbyWf7e2v4IIlXkyBZ1LX0VhM1a07j1rZR1kNUn1ilhi2JaA0r8K
9iYNRoRu3dz9a7R2fqZ8PrqkRwEeCllBXiiqOpOHcShBEg1YIj88OgWG+pKcBiqAJbqH/t1gCo/l
yYyOK+nUhVWDAIJU1Dp7Y9bW1zR1O//rthVzTE8mowTDgUUpucLCfJi4axBlqS8hGauUot1LTAT2
jPLePpKv4m0fivprL23cRUh4lKZDNvacM75PBbo3vpbunZMQ/gk4fHj4OFdhg6bXQ0xDzlQdkIPg
JzTE5EB0KHDJhs48uUp21+LFRQ366vwr1VrRQlNg6FlSRnJYXlcG3g0UNHZNZ3ZMAbkiSEO/MyRJ
83qrFu6Rd1NOa1+3yqOZCz91eRUmDCV5vG6ATCi/h/c6DcrdFjzQyLg81Z9gB1TFGHiz8Q4qudLQ
SIbY701BaUKr36/yw9LM1dTOM1BJb8FQa56httYphLkGubKwCgAKQOaQCi/oiIod2I/jXaaATHse
snOzwFt5cs/6Kg98LISFyRtCHKADGz+cryicTFGmM6+A4MxjEyIQz6IexdVc/Zvbbdmcj6YkmaLu
Vm4SJ+G6oYtfcm+uxh7OygceiQrILlWLQfhuNH+nvWP9S0S4w0szIrFj52dV3YrntwMA53hwK6sC
c9QUipZocMVMATZwodrT6cCsz6dzJo/Rc3rnn6wu6IFF9ipEQgO1U2R11SOxveU19iAIZQWQGlIO
HKPGCjWRFY2p9OmNVc7fvHKe3ALIgST53EmsSXM53jJL4wUG1qvSRfyzcNNNQCAgm6KlOt7rBJj8
Zzx4ed96iNhGDYHQm86/6g7+GjGBFpiJKZWW/Zg5aCwwaUBLoXyKutv5eiif9RiNdIyHGkTXunSB
cTdpD6dhX3T6UFs705bAkgR2DrPSfDaRqh9XLKBTSAWkpgBGIduJ0gbOQMJLH5CfShp/Ln8fkEB8
vxei87rJ6EKgk5PV6X4IdO9ZI86VI88B4QvuwD8utr14CFko7n0+1yw23OcfE8W+avHPbsYZaXu1
wKjyBbxxCa04LNoDouLezVjmNeWC10GSsAu3UyFkRgC+vbnZ028QpXF/36PH1ir9+ZYDd6ZSov0A
TrNVO0PG1RfTqX4z2D48n6eQGacJ34wgerE55VLsmR3Tq+Mqt5CKylNLLaL5o8B7ugs6NWajz8lh
UM/DbZeR1nWNIPCyK6q2wiPKhMBR1oHV2kIDTe2OMe+IYH4C5BUo4JB6MxhzaBFYNsgraxEWq7s7
1kB2PCa306Hd1MBvecDSEawTWfJjX6DN+Scsn/aadDI39g2lSnX2lZ125+i453OTpUqnhB2PDdxX
7s1CO4BlmKdIQYjX8d+7q+f785x/N9xZDwt6/7fV81jzt32z0p0eEFno1+JQ2I0qYJEhS7uqGxM2
Ig7dhV8GCWxPl18d+vaZtRMA9SYm42uFYq1TJg5PPPaRRqMZHdxmVoFU+tc+cHQGF9sn9FJr69Ui
PQt0EFVbSApu/FXjH1Ana1xcuIsc8nhPqohXv7hbUJ3IujUBB4SKyC3JwYqgf3AJeipUQkCK5qka
v0BlTOr4HDTNil3uKd5EpHcxjzcSpNjxtdU2M+K9+jpsZ7gS+ow4uv8aNxJeIx10ORfpmlmDG5LZ
KVecXy3oq0k+TgywFgzj6V8Ss6w53MFkew9SqIG+9cVQ8W4betwKOV1KBO8kfO8DnVdfjIee3d6f
6WjSaBl2AGqh7GLxWCWewChqZtOBQoPQeoOVlWuUMZN16mI+m8oaBLR6wmfLNT9BR/61YYy2Y3x3
fLmZXU8K56rr7EmajqJlIade8m4Axp4iBB4VV21KTKqZGicY9Bc62GXa+/bvg3WuMUB4H+sO4rMH
j8PKt1egCU3yEucQ1TT/vqd4GIHYDyojb3j+JEnXQoTKOz+TN3x46Z4VuvLCbaSb0qT16cfX4drg
Rfc3W5lTPnJUwKUweYErdx85A5hjDBoHGCkdrGiNHqCY96hebnCHx/a7ZZxQu5yGFmlaI7Rlx6TP
e6B3ZD0gQdEmYA5jDF8aKwZpj1r3pEkiuUJVWiMhNbEGBycwk3I+ng4A8JoJvC5zXj4r6yfjjq6Q
wvom0fCieC3IDsWJYZXBjwGOEMCfwa1OIJLG4cbhjGIL+YM6FVCe4YgCySk6C6EcBRdBVcCt8CZ6
0FuupSNyl8utqzM36PE+9yb6dah2yZ8UFJojErNZW9PFb/8C+jIOi8i+AzAS0hTOapv1dihG7VhR
s5MmeB8D7dQsURkq9nYo2oTQH4bdZNDWhg0l29sO/kKNIlELEjVmnpntn1RVsSSw55mjnoxPwj+3
Z8yOFH2F40MFmauspd4va3g5BpW19nKNljxoK9SAqh+hHD2lkhMEvOv2abniIJg/dx8c9Td/xFLU
E0dQCaoLwsMGy/Zxo4okJeLA79IEm9IKelu9HoFcYyN1Kfp+Z/vL9YRCjvoHKuka0o4edKIdCi/G
fpA9Rdz1INTx17wtmFuo1QdjOfZhObwpM65xLdBjcafqxx9pMp+bnmK2CAR2Ul+9+0OwNIrRDZ5U
K/sfFTEVRfRdDpjZfvp0ISklvBAUrl4uwz44StxpfaUdAz0tgmqwd68yK2byDR+iJemtI8X3lq9w
165W54u/vD3osI6q9tf3/GedcW0MDLWaOWdTKHozIfQroHeIPILwk4Wu8VxJMmlLorcvsDqAYqEt
HTLBXGRZGxAC3Ck4FBs49eNWFbvj6SNGsMR1KOX3WcAvCGvhOa0LT/Yor43n2fllixAu2sq7KyoN
HeV1NGO+pfyRqT6IghglkkI3jwiFsfVUtzAnjqmuMCDdLgo5iYGogivcee+V9ud2dfZrmTxk1mfS
U3M1dijL29JV5z1YzDUHA6Zh8xmlDmPSRFdR76P/1qzZCqQRIXQCU/DXUsO4wUKQgFa9cO1NOmJ5
TXEeTgdnUK3lMfzTSpZ8Nht+zyECNCCdJFLcOnpQI2DPgnpEQA6swlYHoP9XGJYJXML40EHkk90t
AFjmCD0g6R1oiZPHPiL4E/6HQ9UprohRH+oRSUH3DNI7lqUh5Qz9UcmkDmPwKwf8edR9uvOX/bIV
pyJ4npROLJF92GMt+uj6vNXxF79rXp3mxWF1o/J0WyVWRfoj1RI6kyxzjIzkmZaNAFS9FUO0hjkj
xN/y1L4SP8lI9kB69Cw1WznSxFPlNbLNkFzYcb7m2cqsdjWo2tszElypgzzhbMJJ1NC8YZR9mvlz
Sa0iitFnXeRA2QCWoGUa6CpkLCCO9+O0bHVzjDILkSvisUCQri1iIZ/+BckdfPtDqTClGTxtBR59
I+c5joyYySbB1p5mhSfa1Ryy2mJGACfXJOTFmj4reLuojDLt0h+ED+GAzAqYTdrF3H+feMCaYrTO
Sv5IIA19BcdxlyZcoEWNzSGc0kUKHvnqw9OX6mZL0yFKxgVgfMVceoy4f5gqDmlSluKkGfzWUYfr
tp/s8Y+7JPLPgxWeGASR2t5J9p6hqnD3s3IqYRyKjtpIhmvd3jAAkMJ3S8QpHNW/i0zePjM3nHvZ
DLrynuwloRiCw55weBQektnO60qPWAQchF3NZzF2lwYS/Dna7rshniQXdmKnFbEOhKZcZSu9M0cK
X2C2x7dv3N9K6DCYi8NMYfzgZ6d+UDv4BTN9u2r+PMKJ26zUJYYFx99Q5dMcnUOQWfQwHura6MP9
q7tEYuks1/ibjPA6OlTYG73mFyyxJaqYnj6EkpKP0B6VITen/9mSr74bOQ57nk5OZK+QciMfw5/7
iCVm303Nefwxgufk7RHh/KgNRGeONIAcJUf0xhmHz6F6UUseBz1DK/hX4E6YuU1Q0jeU+5fC6QiL
mIktn7lxcmv7LFett+uGbotIUs6GafJ03u1E4WJWR/eb01XRKVeTz3wxyIcD+NeKBRZNF+/u7bTw
LXCSeV6Hc7Yqfil/ggCQBDQ8EgTlXaPUJyDidAo8asCa0LBRS74AbFpD10hv/D3RX7cxSUiZCZek
mm0z38nKuO5Scp8+ok9N8wnAl1MWCwlGqxlRRLT6G7nZwdsqJKtJXJSTskPhzbMx9n99V5ahfuJV
3jQHO/Pju0j+0HumhB8aVxh5ILmYRFBHZEbbQak/Asy3s0htR4jGkRdGAu9K4Gg84XSrqcJiFSBY
N/eKljfVbex5OOFXcLPVFbbxrgyQO5hywII6A5Gth/O0GiPLmOO+q/UdVcy0rf0QJj3DaaQvdXyk
VJAV6YxMsYI6j00xqsAFYJa/5C9u9+z/ztpXI7qRcAQJFqjyuHZdTkx8oMDX+2KOEbayz8pqN74e
hO/ampDwomh3dyOkUWg2hVB0UdMHKToVEPmzo0e7CtdYZC6wfcol15CKORVBOq9ZhyqQeMvHFEph
InG2lM6Ka+qgVKtYEvXZvFukdRJqleJIuFHB35/LFXmwC4tQIT2Zr7znSbB64ONaORTFWZhQnCY9
09hSyV8UDCZWx7Hi+56CWjCx/6nnztrhGiQzo6sba5zqILP+EWT+A5Qjw4VxsuNhT18kZHWMerp1
cjhrn7gSmmjWc94s3oXNF6pF5G+mXgjRmV34eZZiyPHC/T9GZ9DqVtLB9I6XCp3ZuNGlD+8POfC+
so190Rc0u9DDS7NOtfpZyi7zZNzr9xk/f9PBJRfDdU89I00LHbVc4ls8asEhTLSmHXDEZR6TflrZ
HIcoQIaDfcHIuSsgRe/UcIKK2TSOE2wepaePprzbiQ95nL2jWkZgQBFRI09dCtHYAlnJSpHn/F37
xWXVaCGwu3eTRA3l3AhCoQSoDIli2alYmY2bOfUsNoMjdYTCD9YgLDTsivTXClbCT+OEK1OJMR+w
JaiWXxB5/S7kJJgNvzZgzggVD4Ngg4/e3QfFHJaRWf/81ahjjedjUAh9pgzgiHdMSj+M2oMFEtRu
v4KWsZ+dYGEhSB0Z8fmxe4Diz3LBWNbX/ln2Onc0ZZY4ad1Agvg/5VclzFDwjkCr3dNA7sY4xBhd
j1N2o8GqBx7h2TeBPYjCYwrALyILkhxrKjo9K7ACE2ShmwXQhfFA8I7ih6cyU9/AkSZHWTH46xpH
qrd2ZDKal7l9xxzSht8mtzPWTAxXsKYy9U3Hj7zY6SnX9LMhHu3YcasQCWL8Pbmq8Jp+xubGmVTr
ZwHu5Hpo2kIwlVxUG/ZAQAPfkzAcsvfGkzGoUBhyfgPLyD7/2cIKvnxR5gMsS2Fx5oPeWk+ZqyCu
H8Vv9MVu0z2QebdwxdLHG3xqZGy9cQ+1HGUgAEkEr4VI4kjV/1YV4oIbYDOz0izPYOiibmrKZMzN
t5y6UO7aczZYeOkriWZd1asd6Oab0BKnqeI6f3jxSYlyhdQLTKc4ehOsQIExRhCHYt/HkHNelQJh
Yn/s7vnFT79Z78UxpgiJicFn6XSrR14RS5JSAp0gBLKQpAd8U9FPn8SNxNgF3cCJHKlXiQ6XRjZV
BnxhVyhZEVTSNJnVl4QeET9ygipvxSD5LTwj15+K2pEwqeG0dZbWeT5qMNbnkVDZVtyDTelAbtpl
aw914ku8v0iM52qvh+V6TVjynCVxLrSC7R33JJ9x5EWf4PnUpsMcR7GZCUs/j/8ht0VdVdOjt95a
sb7i9TazjQsdW1BZ+OufEGtL/rynMeN91JDyNd3tiV8UxhdVgyuJ5vxUbUTX6sOVsWvMkfwpRelt
P3EtPlU04rch9VgKm1nTVI7FsvJIULWXgjirLg2eptg5PQJJo01RZ9m4+wxKJcBIwcXDY/NbBia5
kScDyOwHvKEj/rRqY/UGnLo57TGJS1Dqm2Iu3RZMgguEM7Uir2GgHHhP7L5jR1JozCtuX1ILZS8M
3mTdWoWzvFCtUE9X1yH9SgMVl+Lob3sehrmlsqcHCS6efhUdAJKzY61EFHVJ8Sj0lGYjMn2nBHYH
JhOQNLjMeZ9IF6pNN5yoE6FXimYk5R2ylwtjk1c01YHMGxXINTNFdO1GCHTJDhGkteWgLb/q+yRC
qy/+NYB2iMXPxB7SqTT3S4gTQo+mphuWtINQDS3rC/FSA3lJg4xeqXq66TNgaoK2AOZm81yfU83i
asv5Tqfe3wGy1iNPYO2o3iMrULWv2XxRHZo2wlIy2U1S81wkOiRynEAOvWq8GDjbulvdoLOVq9vJ
vPO0iMPSOhoLYj3HDOAr9U2KQz/WBKTNxm/6JPtRcNyLTZ6JRCuxXrbpO+5U6diPQWfqsFFDwU/w
UHkcDw3UExz5CV16DiFMVQQC9QbxAnqFvvujEg/ghztkgUl6rT0CcGD/J180rwj054pp/H2Utzvr
pCRy+ML4F1ibJcTavrcqCCvNVU3ceOBT3/r7As2/JUfwhZV1Is7ggGcQC/yaZ4aOG/atsIqT2QqF
3dsRykWmxd8wuZ48eeDlHN8Y+LGCz8dWqWY2xMPjgNnoO6vyfqEltw/DkN1x1pJ+RqXzi447WTUx
G6LA18IyB8a3uzuxAHurkDW6DIxp8UiMWITr5YHRVPi3KLNERMcB0gx3YGBvzjpQhmgofF3EB4yy
PIfARvtVXy+iopt4cWI20kNxsogqnWiRSv1g06kR1qJLY37rB+tba4sJ8oJ7U2bipLz5MG7nGiVP
Jn6LySE+EgbNDy0obDWGz8SWn1hWR1sDDGypl88h0DHse2HV0isydKAm8eyqrX8GV7hDUD7WUc8m
PufNP/zrdRY5AtsVX2grH3b4ElIOiS4Ga+W0X856fPSN9ddS3OHgbSyDqtSqFu4h1j5ZFkXsk06e
cyoDntEskZdD6wSd41wY7jKSb1NweqOOBGzPiqWjWN/mN3MayI0DE9v/kbtDRXuPsMgfeEFsoRCF
oadFmtFvcN1SpYBkvGFh60X6p1r+zljG0bQwRdrgmcM5l2u1jjQi5ZM49aF29983zrsKyD2i2grL
oeUwou8C1QRORy9jwk6p/ixXLHC2y3+bx9KQEo4+L6QtZb+bXO6lL3a84kpdvvnOR8Mu77sxmjim
HoLwjNl4lnhCkTLdmYkwJrYjx/XcAcmGkG588R24ddoX0awZhKfQ0iFyBlh+wnR3EaM9dWGbav/Z
NfGrkclgWRwI6yYRwmTAclTnGIxMOzB6iLo+KJD4P6gggxKTZHxx9q2ZuCFP9AWcvn2W/v+SbMqD
0MjUJmuL6GdW5rt5hfBdWbgkYeFxSHwacF6HF55qw09RSqvmi9XlHCZ/NYua+dywpdbaqaK5JxqN
sJe6beERY5dupfejCyoNXdVk/Sx4q6PqQ8KX737sxs4KLDZW14y33VvRaAceC6OPem4DPwLTqBqD
VN0UU5JbT4JQf3mfpqlnzVvouIIj5LDi4nzDqZpdn7ZpeCgMW03c+eXAEAvG/akQToKGcZluJ/iC
vatGHPHS2qtI84R+H2yZs+N5We9JhDpEc5j/CR9M5D7D9kJofDCvBbLk/MrT6wdwpkivx63xIlaZ
GktKUxARjuwZ8IlLVuhqpOIPG9BznhyrZ/Xcel8itNcA7WYVv7dcRB0kHEaQ0azluCGk6oHEXJ07
3EVLn/hYnRRnfLNZ9NtJMzZHTDb2pK/VFclIGqcoVls0YbJiWzWt7sFxHQsuYVvQeGIfgBGc5Z6S
Nz0iJc/uyr54TweGdsPYZUVHJbbxBWntL8NwsjpVXdQr0OMkWSPu+W6ux4gauMVwqTH0EmUsSK3T
ZmPSMKSPYQlPZW/xqA112p82PE8bSU5kiIJiC+f5SJRw1VIiAMi4Cxda85RLzGy/86kkYPPG019b
Et6c1jekZ6fq+0XoLluM1wrMo7o26SnREL3ay0+vh31NbQitagckJxZc48rVbtsbnp8sgXRcudPe
s9NmKjvqGANaiUEEKU/BBJAyXfcOaKSnfroxym++k7gbPV60ruu4pRQLFVB6rX3Yy63xL86Yi8q9
anB9ExnuA+Zph+tNKKOpsHmEIBmszwvCG172vWXorRN7ykmKlOVGczhBfaGg7wTqmeKTaWSCrfmJ
ReXOUIsvdWMRpPAzkiZ5ZcE1ojz7xIjdYRNz/pG7jw3Y7yDexqvoUhJHLXq14sJK6wtsH7/YvvXy
E0za7v9QmCRbLimDudlZu7u/xpq+qB0a/bejdid+pWEtQk4DZB3vbNHIPQYxw8613fHTGxSRKGKY
H5JoZ1tOS3B/vME9v3I0ieVJGDBpusa+vNg13CzAA3caIepmdKxopMB1HL9JTDbeVoFnD+5XGHa1
U080KAz+JRyHCWcazrpFzCCSS9IGBMH+tWRfOQVOVdqjFIsU7T9PC6zT9lw4zCgZ6INZxxrVFqlH
ESJUUJaJu7nI8ZdGYivFH3VmYs/AYOavdKadZ7MO1EJsDpSgO/5ZF1Lmm/bRHKtDfmo4svGpkkvv
BAs7cikN5macOvs0ZnsjYxnTAlZVlhQt6BPyKoYNlbzNFE6ManjywEP1wKNpPMfMm2I/Ztal6eCI
P65XPezXCr/l7Fyiy6BYUA/l4fTFoAKuj0MrNXrpeS4e6M5F4cMudBIt/yV0tw9qsE9fKwy2Yiq6
4tYE1O+vF62L3anJlBb3USW9PbR8UkBVvSz8dCGyB74RE0dRJgAjaJzgMLmWeQyYU53+dgxSMHlz
RYEHAf4cyiPJouoq/oolfBVJNLtTSIau654JFqGr/VobGBqX68QGumN5tybotSTuxWS3DU9Qe2K+
RaF617ZdztIH8mgUhyIMOzmPMInjfO7qA7pGkg1vqHWXtzGwlkApLanWnAp+kAfDA0KrERW6hKeS
sE3O9MtAiFVe2iDOFKirc4Y6S+/E69oWN1Jnwz6qLxbD27xZYN1jhwMQfSZ/+p3VOWToLTAd/Vnh
YgEGWZFcdLPYjiX0LfIo/RVv3jrr5t6+M+sYQ6CxfUU7RiMtHTQeiUrT6y2mqJwbxmlYBKd6g3HF
5HykXVYrAfl0IFBRKE63Md/PlGiNmEqqDkHsGX5/P9ZpxBFmBLp26z+bCh/iydBb8SUvEG14Q5tp
2Pt7ot3HNTH1ropUTg0VqyNWE9pxAkMq9wwU5QNooZJvHmwg+yBuPYq9J9nh1BYfIbpVi1BWW/lh
JpcKA9bC3kaHilG5bPkloU9eyGNf3lcIciThLT5CsF6n2qbZpJy9LsHWqQ/+dafjJOIQJDDS4qL3
62WuqNoW19nDuMWoV0E7zcnRjX6qUeR2uFuOMWgHA2XFKOsO45SXW/N2vz6a9gO2Y56O64dt17cO
5wyqAXkRqqcfCTn9YM2P7/nEYKsRsrF16Jw/xv0p/av3MXYdT1ahSsKAJs5FtfDQoDxtYpmbYAjP
Ru/vtrQLXgLkvPTSF/F9FRYO221tlgppcOamg6hmOei85tr6FR5zXQwsHfi7cOoBduxGaEGk2Pnz
tZvFhe7R4gqCf1nrlZLwrQzp1FaotkROFPggFpiOrFu2SH4mq/n1Aptt78XFY1JbSWQoAh/3KdXk
bCw94ZcHBegvzGEHk5e4QXdotS3e3mTUb+IImNdMCFh9REPpA0XPaowjVBQdR2/9dpkXdikoLTZT
0phaZVk1RCOk4g+rqlUBoiHyVv6ES6WjdoXXth+FC5UiUBSuFwJ/9KUEdRrLxzX3GG0/6CySqFKB
8jh0FA6MpwbvPJKsOyoNU5SHfjvSmaTMx+AW6c1j3vxztG2+izrfWMxIscH3fYyf4Q5cujhxBDcK
xUYIEbuKZn9n1RSL0oJHdtO76aOvyU6en84WvHOkrucb/X/8kezh/wCn3gw9/xeF4dSJCwr4IKN4
AjNrZZbPMJMx52eyQ5h0KO4VWlZH6MjCMJUBEPHhjfMECAhliueSPDZvqWhRMkWask+JLggeBJbR
lC4JCF5mxkz/odo7eIGeoUW7WG3VF7ANH3WVSyttLENzognCrZKi0oTLvMDYQ1xn90Lyksz0lDf+
DvHqdjtR93OfbWtnOaM/8KZt3wCsX2iVrDI5JSiLwBbr34vIT8LV1yA3+xJaCghAIbzP8JC9JXZc
yNx2H0QIa0FCS13m4+hCoiHf2TNDcEX03LSFYI20w3Z9y64kvL+3MY+F3bWuA8zwQd4pmGsa0ERM
0tUIXrpoROeyWfoAkkE5KgXkALUeQxTvR/nO87MH8dWrHDmweFup44ZFho5kyEHV0AjPDMuN/tEO
a2V1gZ/bLSD8xx3IM++IeMB3s5TITKycnw3Hf4j1kKKUiFcCsw0T6GQ4oC4sFmH+5YqM7Vd4sMWH
7IxjLcEHxX2sngpvmVSLy6RY0T99w1EnJabdphkVoPWyVnJWSucvdEU8z/vkrPD/CWWynZjjm4EZ
FkX4z3fQYPDKYYePpfIoS3PP/sv5fuU+KG/hbSdgVNTZifoWQJCpNuD53q1gg9srXFBfffhQowB4
6ntGtfphxp1wJkpJRnub7renuK/hFL3B+fgym6T6I55nVyt35J+qIqeoZjRE3CipVpCL2jfh/Fq3
S+NFGou62rxl7ZGFcDFu0u8RIc4ndfxg5BtiSB1EunUuFzDtObudApr0S4JVZvv6uAs14mjOrxjo
lHUiQd3L48qsiVLJvojE38H9KveqH3EQBAXPu1Bt/hdpiwel1AaqEJicyTiPt+Rl0K+Hjdb6aq/D
vNEmqq2bZP3yhOKuEBsJBErhtoz6OMG9Q1E/4HPwDWyhAk70N9RjmwKd+i2DtySUosWTNMu6ysp9
RKoDsj1MXXZclwXt4QZEQTgI17s5ZxasKHX81/099spE06t4Ji3rkBya8MhKR/DAvS8CUC4npS2p
ERj1KNV8WxLTlnYFveAdi92gVUC0NjJM4apzj9PxxxagoY1LcquORatZkoYA8m2HL9AUsBcQSBo3
yvOaC9ta7W2FsgKiRLQ7Tz40PqNgFLjOkCZ4y+dJckhhDZA83jT33zIMWf0LiKxad8zk31FBXnvx
A+UYBHo1txwGjv7QIy7Q/nSK4FFHuBwJerHK48oYpkvY2qWwltD2es/ywbWsG5P1nMrD4EtNvvoJ
B07Oa9GolQee9SiRYBNnc/3Bb4SlCDXO9ZKx4VHXqINQLhSiUmptSXctGKQ9ES8o4OwYJNOZ8Pu5
TZL9s3CNPuvpOAhb2LW1ZC5D4fMeUDVCACJ05J87fSp1Y3x9K6BEhqsPgmyxq5uZpTgH3ZMc8Gm7
7MlhpRl4niO1jG1Q6S5W0JXYXjzy7nbT/kpk+iklqMSKT5CtZ9qIjrCIdLxm9W//NUOEck+ZHiE/
YrX3SWCUPC042WGPZ8OUXdasn0fSW6VF9jtHG8HjI5KrXMCcG54uiQhCjqecZu6GCkTP4ZCKfhfX
wsgQnlBysCuj9ml6FRdzrmQt9BTr6zmmMt9/DP0XKjCDFB/swWK7W4j+DbPoWqyNML4YB1zeD082
1WVsT+nhqHxNzKzhdowRFV2E/jSxPBHWX8mP3ZXtUC3Kf0AfUbP8xDLS3UfZmf04ey6BT78Chva5
/Y7oxXypjE/VvTgZJpDteXWZi9WhmUdNqKivNETtACogUHWbntNA1i92x6+rj3onFkLtsLjFb9ym
Ffe9UARFuPPa2PWi7YFuaWUU9ethO1jivDIn67IMdjWwymDK/MuO7YVbC+mCUCVN9Ut5bkD2s0M1
xKdOKJKbHinZexsN0bifhBWXcw9KMhBuK2K3ajJN28/mgmqMNrX2nt49peaNYl+JG9Vy8yDqQtsF
7OwbOXIU92KvJ6F4lkwH/7RICD2epfaD7O8cV9hHS+GEeKeCV6gg+LrxtldQIeDNtKL6OzZOwK3+
OLS7oV9Vt9mgWP97ZHFXJauLTRicl+65dCgAYt7WcfRH+A4zNXqyJXpS4RwvRE9abxGD57QDy5yl
GI0ZyhgVMCMJXm11MsWZR29EyKgUy7kG42+CPLHvwxsOgOMlNJtqewll4C8PsPYZrZjmPcVYE2BY
Nz4B7z7H9wPvkRQ6hYReJh8Af7ygFwMbwOwf83E0OhSgTPN6oOM4ffJT2uBEYeGIxtiNAmhmjjdh
gNKzOB2rqtD0yW9tCCCZFBY3QETUTmQU3IX3EoX+yRd6J6CBQ0ogqoReJ/UycUVGYQ7deSEWbF6l
9CIH7rwtLVu/85C++aoMgJt+SdBJR5p89hX2baUbibPj7rQ/5vxopICF0suZDZjrDpIJNSvxYUNH
4TYHKgp1JotEHhsimTzA5uyqS7kP6AFMClUzdpiZcTog8Hhd774/Rq94ZG365NfdomITf6dMuzpZ
4C6u6HkIUf2hAurepGy9bPvL/10TKHNZqs08IXEfPDGhIbWJ22o0eoABdIL5yXqnUn4C30JyvF7t
/QryhEb5JMxHk9RVkbkafLPxdfYCuGVhgL4NiFtKWbbK0dDIyipA+fa0yFfdelHZscgJArU9JRp1
wiePaWea6Wk2VlSEbbOHz9LNWOBPAALLJEAF8sWOTPKO9OwIv4vOCv+nKBJlAu95aZ3Z+hJk9r3L
FxqB2w8elkNp/p4z98Fu+CxeC53/hCpn2zEfxBUtM1JvrnanJ98ljswl7xv1HwPppABeRMwZmOtO
Et6+dyU/WmFCQHL9vgiMU0OFVSNKWV+ffirKjAzGvLLae+iMrMZHsMtUFeLSVMLpqAT3nM6AUP89
YDM79WMwunRkOK7iOsbmp88hYXwrribnRIr8Ah68WwNxzzTjz3S6nOIVRj7gSYNJOl46D9QD8U1y
A2QYUxO0jKmcXYXxDuRn0LumH08bZa66laSMc8mTDQAWGXAFlSAl9ESEE2emOfZPJQyeHIN4r306
1LStCWa6B4PRXzVmBxCKp9D+AchmpjLP/SNYiD9qP36DtXgqN6CYwqp4lOP8jqUQma3MlrA5kpS1
yOB5I6uIbwY/QxU2AHJfUgcOgNTmjdJbhZ4RoTm+0bFPG8QNBVWtTBNw8hihmKiZ48CohiZbrjRi
KhiE6xeOx6U9RGAppqlZZ5Rrir6zrAfXCwIl6OyagK3kp3pSZwvUO6/KKkK6jbRGOtuiEa6pYxYC
ZKy1UuVAi33TgvHZsXiPHTv5L5axablmTgBZXKHUzW2KE6osTvmJowL88lAkUyBJsCvLaxQvi4hT
Jd5jda+1wLmDOFALvBLsDNw79TtAdkNKAc2BPnPgyjr+YJcsQT3xxzei8DlV0ufjy4VRg5fnn+U4
q7CGTvhjb+jga8EYn0UI4jo3uj4opPiPZXVTZojMHN+MpA933FfxinxxuUkz+oSjhxEyGR3V225L
4LeunmMMMUYnoSjAnith9h/olqhSVKF62Ngn8Alq+ID5YC8qJsdfCz32j3p3JcbLz4SDza64GdwX
R2e5nsG/bF4mPVHRHe/gjttsXb9PumwHz6ZYlFFEqomJ1dl5Ib569R0W/pl7SjpLPWRK/cNCxTQe
qA15rZLKhP+G1/b+EhYw7WtTRLUEouN1JA+dXoLGip/hiPfo6XUdikJOFfpMgMzLm0aR0RI6m9ek
lBHdpXTQZHhTs69G7ZxKwyVt6Lk9XKGqCgaIs58RlbeJ9IXBA+VWZ13Qm1qucD58k9EJRUJ0Pv9Z
mEA5UV8WUJnt3W0bgaEI0Zdu5GC7xWml8W2BG5vNCng4A+PFuA1uY1W08bgKEIRhEWecogyf3nT7
5In761AOhQRJ6JgdJ34EN+aO1LWPwl4bYxqiuoCf3YNmJ3e/8qv5RQb5VRXJjgrZPoGaunQIb3qR
mqxfN2hLSdiQvy3FwsKzwXTfXIJ4X8bioQg8xY2ktfIJa0ufEQHrX4oWLeJb6iXqE4QYx7E1Af9g
URND4BpEd5s0aDyg1QLIE+Baf4DBjHZCbLFhe/51VjPIZx9oxa5pC4lFsTZOmb46qRZSFG9MG87r
0PgGhMV1S+nJQI9Wbc0t0Duj2qLlC8ckG7voyqGjMk42xUzT7CqZ6inX7PrRnTsqLiGPJ3W56tpO
U2E2P9WWr2VaNoX4wLegVL0t9a+2gAHeJxl6t/04Kjm7R8w+hrDUMU5LEWKcZe8mcsg0tSKq+DbV
7tAm1McoRlsayW4Gknl8RmIlE8hlt/QO519OQbfINbrj5KSQSDeaswBAZrk0zW8YBKJELDsnI3zp
yX+s9pJDw/PhC6i12Jh62FYGPDBRPe1AmQoBkDKPAaIgYTqj7BLSZA8gEjOzn3kU7KVpqmkyQ5Ol
ihb5Mgi9qx7Mr7tXy353YaooL3kR6m53kG3yT/8ELiUm0YeihRysOZV+uXGVPqINhUbOhl9eNK48
wcd+YfiSDcSTNok8ENsUqAf++MfZRDBKPbhGaKUKrQniaaju7SCdlacYtU89uj5mztKXbJcXKgO4
2VfegSIK2cZGOpgk+sqo4Kjvv0Wu/TmivryIZ/aUesGtpCx6b93A3lpfPBsoNOn2dFGcyPgE1pgD
tGQAXISZvWq8joJAg18DFf17tw7HSE7MaX16GQSWvv6+/uZ4GUq245KNjx2ixFtkyIaJHbjEsD8d
yuIOYBw4iDwB0lvcjUAyg852QDUhVWu3apvpo7Vo3t+pTqIzTCwtXENCnFTQPntU0Os68bBvnQtL
k6NA2x64q10dvkEgJBPTIkwAOU3JC9X9u/wqa4dgAkD8+OjBntFG2RJNnd0prqQ4ieUwS/5Ut/b6
LH6J4A+Cs6UGgubJ3IlUfH4XTA+8KDk/ljZPblOSnBtWS4sTBr6w8x7zU218qWMeyZwM32Iq2q/c
rNSJ+fqBD8CFJ0jE+p31Iw9HIaQcb7DCph2crmCzz/BknkjTxKLdm59B610LPUnHIftFA1jcdO5L
WPy9kI5gKzoguPg3ciEWgiBP7EATHAUo9aXIAlPrA4Z/Cycjut8NniZ1Pj3KJ66u5LkHmkLzw+2D
dHLrKJIyjz7DEap99vWnHt2/3lj1MWHbcrIITNUup8/YGLj2HP3CuIAIDgguYP37sdMONiTwWZUF
PBWdH6AOycvvf7iPnsKQH0sbb2gwnwAxQGkWba749M+nGn8ei34AZdYNFLTxGI03/W3AAstcb9pc
+AxyCrMteeTaq2IYsPLDLPN+8vXhb4sPIYZfwydJXHkdFCEcJWQ9J+ONoc3DB21lk7M/l4kU7ZBO
0PjpirPu4AAeKLC4QZPzqT28OzcFd3HbAZ/BfGezCoOmIq7WzBnumZNR3MyRKPZu1J9GO/WawQ4l
ggDF+a+JvcTsjlGmzR/elNgc1UB2G1HX3YYRKqFvgVynRkYCsTu0Nn7qY3R6VnLZ6Rnt4H3vnWvG
YCH5nXXwIE7M3N6PeZuX21M8A01+lkC/rkaUfPOMPAL/5jsltaHYt5SpP99k1yusZRww6uCvlv9/
Z0hmu9VHqWX3MV9gLX+rpLVHyOUm2NawsssFoJed1hdK1VQU9Yr5Y/qBZyu6YHA8na+PMRNo2bMc
M8G6+4+Gm6UPjWSSCUwmRDudqDw8lYj+RUnspJQxBy5zrn0psVwQJ7iysH/KYnD1TOPgJd2lzjSU
DmeHWOQ8e4VEcuuVAsVNg2LK6/lOlocl2sy0jB+v+i+GMSehzxeRxgxaGSJrqPS34RhvLhInIoul
2PsTRZFswVIqpDbysJrwp1LiaTHHHjrl2TvjDCZlhGtDrV+qZH2LXw7Len0mMwnpwt//2P9LNsys
ykK6WkYInPGWKDMeASe5k/ASiSJGMzO9PJWMj04cEdHP22UXwb5hZK6QsYgFs8AMD/kQJAu3iURM
h/q4o/TUGHwX096jKtNdGmiMjTUDXQ9GrfQNLYspAnEF6Vj/UlVLoJYITa577i40U7XdCWj9ZI5o
wXG33RWllnLy8+uEDs96xNZGUgV9StBGEkka0gp3XhQaaKCx+QIDigYmUQzIqST0nlBCJfyxJgPD
sNo8lwLPgFcRuNfnxNCu7vpa2/D51rKhMCCcEpGnHoDz82hIU8x+nqQmslpIJ8XZTxC0IXf9IP0r
0Zr+V3zDoJacDLguKuT8rafYYW5ERjSbeKAEUsj8kvuVKHy720I1NuCi9qt26UR4CUEfR/AVgn9V
jUOIP7lEaVlB8f5bcwnFTZpaACkAvbm+WZ0jlBW9Lv7B93H1gvd6NCevBnyCKh9RWwDBJjp7lMnk
+d6oQpdCVWOU3WaffrLxsTQATPNO2QOch71Ma1+d0wncHrL0fxKi+MgeM43fT/bVOYQnUArY9Jvb
kztq7DnYJOY5DB+dgkNDpGYqNLGig1bm/4o7LPmDFvaRFwkLo7hHqVLfAUAR5ITkmvP6FcqxL4bf
uT49AfgTmtXj2DyLnefoblokiHGwHi/EAkjrJ5ztLluqyp1/SosFhLmgAdr5naAaJzwc0FhF5gUJ
u9nR+0mYM76Cya4Vkv56Cy4GTX97ZJ/Ae1farPDSmzQ7p6qhWI+7QKOn4Gx0+tupW3IZsfKilBKa
+VMOHdkkebSF2sDnG+G8ilqt334Kbn0sjFdBR7JMxWgi7kT9ShMpu49RWF3/RgjQeJdSo2fLDBia
c8WabXrVPypTXBOH7HDLU28SH57XnlDhjvJy9GIVpPA30n3kgpqyPRG//gGlqfO78sklxpt3m42P
sPaf9I391N5+rKN+PM9o4YdiotUYEO7eo4d4THtDoy/C0Q5hmr7qqXCAMh6da8j8I5EkBR7ayJEi
PqtTvkTd/bSLqCILqijktHeb8gWo9COpzXUBAoLT7aWV2FtxyTe/RJbWjqWHIG46wJbx3UnN5THk
uauTsmYsJjs072WmwMwoBdZdCmxn6eNzcx/VLKzfrywbl7CCTkS4mfQ1B/jucLJGM4bgKbjPFeI8
+vWHFVeQrdroPcwkOwN1ZCQTNmvkLbOjt9QweCwbCuxf7YXPAqcJLjfKHt/qzx9P5a5iInmBHTvw
l0jwDrqJDUwIvRiPgMPjj7mM4kxZMcRA80t4RbgHXJ8Va+oLuSYYJ2YJ7GdFK34vbnAAQ/vmEc3M
SEShU/Vt8V3ZabAWQ0dNsEy96Zss5q5FaQfHo5moMUcoo6i1pxQquyou1mmSoebTGO4VzH1xvyOk
lUFaQKpv/K0hBOsImrJqcSZB6JZDpJvuf1SlyH9WR7VSgDRCpIE8gkPmMfXhDqvDixLjoYasUF4b
M6fzWIJZkujcoB7aTT+O/My3FPIk6kqz90WUrdqbeix3PrvXE1jqSHjHGJ0nmhgfvLuezMuJaCbm
lWCDTySQOKwps3C6wmK+wBAOWRg++MAJcsERLBGXoBIMx+O1Mr9h8dOaYHjJ5EgPmUggok+/ULyc
JOpAt5x13SsTuZELuqQ9L//rlka7oShYskyibf72VUhZrT/w2EygfFduMsplBF0EzfEs3XLm96sO
3ssyseuphiHf26Yq2qvG8j2phbf6bz5evnb9X1SknyaFjI3Gw98H3OQG6Qa20F+7zD0/yCA/SGWN
/gG8e11F9ppGaOZVOblV7/Bt2x64s+yPeTDZtQGs+4StULJ45ZwUuN80ARAKgSKgrvUlNrfZvEbF
wUTe7t/x9cYoQ4Y3Nhogiz5vLV+tZ73Y/XCdz+lwhe2i05xwJLI/jxKM38keRRc6PfrzdVxf1k3/
TlcqHBTTmLLS+Fd16mFDcJ/5AS/gEzY6y1GeF0jNjCjewfnzO+3ZNUpoIBkgR2uarNBSIJLnnrPU
TZ0v9JYM8A64/M2modXJVBEogRVEi+N6yA2Dio2pnulVb594dFLgfxK5p7ZKOM7HnXE9AiL1AFUO
jeQS51ifBx0YmvhlUEE4SY4kM1KrRXb8ii07zf1HkPx8vq0zT6/5D6D6djR4gP1KZHfkAp4/1SpO
es+3TYAImX3TjEsEQkfXn1eXEHiZvM6kgjJ0T/j5G4Y4tk5qes4Itj+0SxYcaBRrD6KLbgL1gk8R
wdaiVgoplduQGjpS9MymdzkV2ZWHm/G2B5xTkBKbfhENH6ZVkKZ7fQzwlwlP65ChrxzppapjhNpb
dbw/fr+S0lu6gU+raxUypLN/4ZTojg7XzubGmBBXt9uMrszL/f6Wzh1CAOcbw9xrJXh5fvDcRono
W06rkKQxrcF24/rX5OZbA0qf1nW1agUVa0vuKjGaOpsOs7/1drHKb5JkeAn747A7ztCYUFTCsTQi
oeM9eiStC5C3vazUyTKWH2Nxx1vg1X17JcM81fO/CewvKYUKrq8/3v+NIGdcXsEKqzmW+fOCEA5M
PeZLP1nkUG3hJwaZiN87zHjbHpDckyN7ccEXQaoGFGjSMBwjC7+rYeu8TBBmK/6e8ij0h+A8X0Ft
G97ZbQE35j/Z8LLSpM6HZoOiThZ5Pm9M/JYuRMaU0ts6PGTXApQhkNee9gMIwOYyhFasND3Pu3o7
X9Ub2StLWe26858+k7Sq2Nz2iUf4IaBHRo8/+DF3Zu1xI34XfpQXbcp3FJ3iM1eR0zldGOAjvRaJ
YMKSU3vOMwLJKYLyx3n5baffSjKLs98LSDeGQGvSVSruFqBck0lkk+l5W5l1Wl3Z1lWRUKUUACUY
SWKXs84ZnM4VE9WamgFoCQYTOf/bit66fgDVB1EFOxRNqG04SRnbWXc4cPYsKoQvSVrHjTu/kiBx
+Vm/WwDS02ISQAp4wuFI7puAUIaLVqKNmpZsT81yZqLEWluFJ0HJDC94iWQmwZY5Tsm/9Go5zdgx
KPIZdZPcYeDwC+hVDB40KNVKK3YjlK76Ew3P5Wg6TPZF5ayYdNvSeL5nYD5yma6swO5U7t3mEdBm
1Fk0ksW/v1rHnx4C+7aRrn3Qsenb8X1NoRDhqsrWlcFRvfDvePer9t6JOPQk54G5d5ys4vuBYMHO
oq9yF+qtODLOlW2uPcGiIlXSsQCT1p/efANTR0J+pkMwKs5MTsfEKbZWaSOZ7YjDL1ja4udpO1kJ
vzyGhgV8XnXOMtpISZ6NuYYs7WZvbXfH8zjF5PMdoFHJbA9VfsSzoeSfA7H49PQDH1BMV5PUHJnv
NAXbWW0foXuI43+zYs/1NNSNGgqYTELBxlgKHTllr6TCRMq3NsuEqrsuRPHGVR3RVxvHSlYcoe/7
2ZUTiIuLH3nDS55v5To+LgBo11lw7OkHYA+7y62jnEEkiDqYO+YeT9ec7Y3KphJaJ3MEJz8SQMkj
UDKQsULOmoxtzhIFs6OIPbNeSDfLshrkzMzqdqXF1qP91nt8SroeTcqyDEzgbnKWh0uv6Xwh8hzV
OBav+H0IGwyCOCxDCI8m0Luj/HDXqiEMhCem6nFP6pxkUjY1mYdnDUqqTUemxih0LOiqMarSWklv
t3+SlvaBjxazKTwcKASHVLedBGWiQbXIgzXK6XSv+muu9zbY6OT6sBgtj5cJUw8UQoWBlryUGg6u
BJ4uPWqegm/rtXmIHcKsr5dxDqU5z2qxnT+bNLPn6K7geRLvu9d2725k+JECxtjm/Jo/H1n/RNFl
1b1hQf2NIFvKIdkXqIDhRd3EViD90Y1C3GC2jkR8zKavtZm0fcPZNyhhNiUvZnNXuqTxwXEEvqhH
s0a58N9Ow4SBaIUfDThJtPmdfK01lBcVDZ9o5VMfNoZrFSfOknJZtpyZP1r5cswH0LyoczQR6hWW
p7JTohZRwquwPWi6TPVdpQbc/+8w7BKTaNZlR5d1vh0dfh8DHKLnggFlMxBOcvsm7e3ivymZ4oBZ
81MRiQZFcDlENTLwyIznIn9HD/LiOi9VemHwGcE32w3//XeAG9CvkgzDCGXbYSeuIImOvjl7vuxZ
4WwkgaRO2FuupMj+FNMqH95QbJEeNYFE3jt6EuspzhjSaOuxDuUot81j9OixqN/i/vD7RiO2OMB0
l3JVLoOUW4dHHn2VCXKqrMNQNv90BwUSoltZ2vj2+lKgF8jJ3elYrTpMJjO3Hxs4KhEeitO7TpC2
9bdW6b7Z48xq95LsYhEKxGegfGsfqAFmhT36tlt5bZYxLs+PiAKbgt92wq3cLPWNmlfvDQlwf8yT
3k0FTWLFgb9PET/aoaYOWtIcRH8QzYvCjUi1ITcrxTlk++i42ZjeRaP/NKuCo+n8s9+gvmCpQatC
Bg/C8J49WwI8dk6n77FZzgbFDGkAqocHo+uMGw2EiZcZnaBMw51+5oMHcUUL7NTtkAbWxSbdWOVO
ipnKLg6VCZV2jJd8F0JE2OVKNVRinkky03xNZz6m3Jrf130LPvbXJrk4JxTEfDAep52S7fgIBQGD
FO0jSh3CWpDeZS6n5xMF+5ixTEaRsyR1qi4gME6OFwuJiT/AdmCpmLwLgUW//LP4euVFC35WWL6s
E2aQvW3HPN2e5iYkKx4maic8LRVw0uub16cF/SomWMSJk5i5gVEgZNUZRwB6M+aClJPOOY/uIEP9
Y1k1tfg3zkwITuQeoU5HUc3s+bW1n+DUX2ZlPC/Q2DjctwRTWn+v07LWd9XN+2wUQF+BHUG4RMl4
FTuj0oNuyNN8vb4ZXgtVNsMaY5cMFVBfA1MPYc8QJVfYOmAroV6T0k0UDwe9yvIqPxXuTci/+FHo
v8t4UFvB82cpgN4wHH3l4HLs3IJJkAm0d4JY7f8MzNPZW3CbXcCDWpgykiESioygTZN/idwizOrI
WR4Aiq7pBeRDjwRiU97TOG/yORAGJiDPbeaUKYBuFYPmNqWGA/8HgjEH4PFWIBFqNhOAryZZRhnB
2Zr10M6WsRcv1RIm76VmFRFXJGhENtuR9iVyt0vQg+AOCVYTarOo3zMAM/0r8NduvdLL/Yyiufq2
gomALbsYk+AdVLRjRmE6jd7+mGWKCJcDAnfLJtYl4a3Akxkj2rBb6SD+iGTbskaJy/gpAVM85dRh
f62XTFd8QeqqA4yhHuqHpl0q1KDbBJPrXxuGxqz6sgTPVFKhtOScg95qhs+fxCA2Tgn+mt8fS0BJ
mYWwB9dBXOVzGqhEDBq1LVgo62jq3Up0JKB87TQEPoPQw8trumlGEaAbckSvS6AzgjJu5u+ZaTTA
Vpvp9gGZEriSxrQo2v4/qJTkRppUtwc/V+jHkrokKmXK28dIgsfHe9smMPo5nk5oqEh+XIHzmqS7
PQabEh9evc2R0Ars1QqS71XIvHu3vjqg2UkoClB0FoRxB2xF7dGMFbaTzKt/BY/I/rnYxBH3riIS
OG4Lm2FvgxrJ+2BEQjSEnXkSnJb9ZFQr+hodWtFr9qCjBqrwHOnicyjzJ++YZjoaQQb8ea2UYVjw
IkKTLP+3mo7QcbfmNKugzlUMeHmGQtkPyouVq1Z9NBnUimcTvgHFbszZQnB5kOk17Lp5APTxQcDG
jnB8h/dgM+38gFvqpRLKo6wD9QxFKwILZ0ZrnhxtfPWIrBraE1K6LgGwvAbEdqFpCajDAj31CslE
H6Hr7TNhzK2JK9+KJqCryQ/59qzv3mdI5V3P1Uuqq4L0qHUPSWzBfZGi1R/6uiQ3Z+0pwockO7Kh
tAzLuxiQIQhI56kyAb85i8KruzXTjlSm+lZkm4CE4YAhh0VgkO7GPeZJUtDWO5UMkivzN9PuUgck
je2pqbahVRtEZuZePiWLbzxVcUif0u1iQ7KoAAzstr9LB6YE126IRncL9gqJAWrVkPEGXcq8TEWw
NKuXKCWkYXXH1NN0VY2Ru8tl3D42jeTsF+/1gRZgsOJqn1pUlCV85Mgrb/by5DpMeDh63NQKwbOF
D5dIjuGPQ99Mfrv0OY3SuAjX383vpFHvudPVkprI+06uvbTHIu6D5OC4Iy3s5PY8pvh+ZMlGw6yo
sVFCMUGOJBXO9lLYf6qkA/w4x0DhVVVEXlQ12ccOjEF4AfNC2mQqAZbnnsgSeHCqf3Wlkvb21pl6
meBr5RJdN6+jDhikFk+WSDZK+KChO+tnR1v2vXsBa9zdlexStx4ySyqLP3xc2E8askmgNZyjdC44
DEUMOoWZQkJNeeCDTPk7fYK/9t6FJkOZhnxEc333t8EBvuvtjV2dhakgVL2phvqboEAS0V0OwVtS
xMLgZqksjW1MgFIXPlh4S3g1vmBIBnX2jOSnAeQvcYWGWYVFq37mrSuzNB03hFnJcGuwLCiNG6yV
R0vlJWtvn4eClIhYJ37rTYqzLRMFmDi2Bp15QUBn3F91xbphEhFmPPZdLBbnEI5wN8B+Hosxfz/f
FkIm4JoCB0AGGNOl4PB1SjJl5BoqPqZ8ugpZ61enijydKuJA67/vzXaldnukfKZwjS+impSgTNaX
hNz9WH3yJgu+6DHi3ayH+U+cNCVhjuRKcxexIcl46C/GuUc4rL01bF2mqVBSRsfWpzadlFy7OMdz
rRd09e7CyOG378SRCj1HhXUA/CT3fGmwX52UPxpayX9wn4wFRRED8y1pUpM3sN+l1RoDuNvZNzNm
znJMXzOpECXgKdyf9FXksETIH79UxcPJpWILCT09CQdiqlML4KWdxtW+NBvRKXrIxxSwB72OuBO5
IR3o+Q0Co0DFh3ieUwWNuC/rR604GZtVldAy0A8UI6rqXN4JotiC5Zj/pAY6dmO9HKxnfn2Z4wkP
GcBR3l4V8yAHjcNfbEAL9ornOF6nnOTVBpCb1nFZPqJITDolF+AV9NJk0+tI9qVU+/PBi/wwUGhX
Lve7hP3yozt5o4F+reuIy36BAPsQpJSh2amXbgwhS2gnOpfuuNNL9SRAija+KrFKJQz87mFn4KRn
o3f8l144asD1bkqzKuejMizAHlgdV/vS52y7CAvetcrIf0oWI82dpngZxpX7UGBy/jWvXuIZ/1Fn
yfkgqhIvBarBi1Uh4nUdtESabAGWEb9WTnHciyLSWqdgGfwBMsn45zT0kxy3fX1YRmGM0BxjCI0n
/P1X6i29UPqIFga1ZryvODfUO9ofUUB+oXWqTKkcr6j1xhdKQqMFhJec3yT4wApz/NQIRaF3PtFy
VaYGoyy83OnDBp0cB6f1jh9vOSx65UrAFCZAojCk9HOWGfQhq01ZUD4zlciOQiIqL+2UiPNrEd+K
T14qQAqwcZI2PaeEm3p45t6S6Qu0zRKgOoaP3yjkxSbb/VaD/OFhlgqSsLwC6t2XG0IdjwKpVedu
TuRs69RvRTGiw8hAP62OWjqU77amzA/skujHEfEzLijeucMpRVoaZ0J6OexrrTcF1puBmxuC+uaP
zzsCW/upv/yD/C6lu1gJ5cJZ6fsUuN6W5HcM0W2L6TmV64V906oo+ak/KdahGrOy6FXaLdN00eeA
lGWHhKbB5zNY4BwWBsnpRKkmjKBmlo3xmIU0CbaHVNydfgO/ZAZqo5V2BMZICZcDgN80sLoVCcVP
/SCGHSGGUToX2gEaGsSgvElDXKYbzlWeuCha0AoJ+BXWDmRE/YcJeLm1fBmaKlMYiiLGQdUpdMPC
ZQghOBjxcb87YN8C/kHq8/0KANUvuOurDUBQVwLULmNEzcoP4nYZZFzCaAsf1Oi0uGTt/1DY0k5/
e3N+L6g2upjvcGkUZ+P1olIYWETuFPlqybTkS9vPhU+vImz6Vnyi/CsJFmaXgJItsgiXcfvXvD+m
j48icrd5XSAdELgfN2/g0FXR5DJMTCzud5qiqSSVL2wS54rOdz+FRYqA8WKX5cSiu6DEBAxpR5U2
lgQcjaPpDH3XTyc+QyYcQCIxyW5Ec44xFPJgyAeZRqjH3QoueuIxZGcAzIcu2U0kdVP9TGLa4NoA
rMG+hvwihn+v1mFLzeI9sX9eqg6ysnX2xzY3mmG6IQL1MLpvPu91J3BJyt2C5sDRfNq3C9s9qorX
6fhANUzh/naTPLZGMPgwMqk5HC4ZqBX8qV+ggVGGcEB9dQTmwwVuMW3cGoEnWphopdOnGhazKTB5
oDfM8F2AjhM6R5tVpaWbi0RVQ+s8NSuYcthoml+hdVd9JvX/doFhSIewNQ0wTYcVIuTS5Pe8PJyl
vuxjEQo1nPjVlojRPqQHkebzAk/wxWDq99VP/APeiTm8j1pb7XFsGZq9pFsd/fjG6xnOrCknG6Rn
4ay6C3ZNts+nLkh2op67QgMCpVlwyfJzONeFxhnNr+D4smAQuGRw26RS6RIn/mgpPAIMRL33NzR9
wIY4gb1bTLWh4p5ZVss7XLEcpQaBMJr9FnnCxY2BMeHN4uLfOiQkpPvn4FkOQxLVYXc7HCAmoRIs
cczT1ycICR/8VgbgaDve4T8XlCAaV2kSGKH8KeaAs6RpRgrkl0V4PeUyDOSLA2mgthG47JIVyyVl
1Flywuvsz9LKoWzXIO06B/F7gAp3IGwLM8tNn/GPNbq81wvbcZhoexlnOkoxYBcI1/oL9FqG/PEz
0CP0GFw7xDIXOrkJNzrjo1STvjiKoaR+pgW3jHvUaAEGLBxtPUuRTIrdt1AS4Work0R7OoEGuLn0
Wfu+SfSqf6WPhZQ+J0CO4123m10DjYo5QfbaT/f/N0ONY4rn/QtD9HTKz2iaOyggtLkqGEh1MAZV
ew/Wz1bAgKGDO/3Lqn8/euaWeD7cP6hqZ4GMBQfxSVJNSxvadIp96zyQpjrub1eyHx5+5dCetaoy
3sZic4UsdwBCATaO2NViRA8FqM60EnxMR8M/336E2nXI+ypQq1RhDIa+1G8uoh3EuXpRKdBxKs8C
MuHvX1+Z2nf4rvYnaOWo9QY0HH8RiFYLKGY9jD52C3DNjX8Mqyqc5EFB4fXcRPwr5eM2+zBGxyjq
hD6PVElCLrSHViLZMGYsL5fqlR5FSgGngnF40wBfLG+ys9PyDLboskHD9z1tHTgPI87r2BhIaZZS
Jv3hYEe81j+ttwlZJu6ekut4o+oPeOW/20n0oO72n4tsYU8yr6kWI5yt+5XlmwQ8dQpEykg+ku8d
4tMRcnGfZ3i4UvlM83CoPg8G7lz45zkHFahia/KpgqqHJQ5qEze6ZMK5kwe55iq2nkCUiXG9e+Vg
ICPrPdy8M292I6fgUsCMl90Ufp2WVAAoz8R1/QVJuJISkIOqTZEqu/xtEaAyoHXtMKM4mcNTRBQE
OLr7s/AA63F+gVXNTZwxMb2S7YTiCdTWHY4Xjdd4pIwEOXjhy8lwEOF+mdQFxkwAe01TeA/DRvB5
6+53aNcd073ePHaOyuL2XHmQn0TvjDf9GSFoNnjO8BRCbkNR5TZNgTa1VhMh+D9X1DmncV6jkvPU
6uA2N3AxOTodNQ5CyctbpKlFCp99olxLaPZ7O11cVACmHBKkQ4sv2CvPdY3LQ5xnBtxpvqRACKyv
ljRKAMnQWzOqUZyh40vf5FZF5W7Jwjq8Q/IJkYcreLAoo97bUNn/eWc/lA9u/viyVxeQV/XxK+Cc
MiIxpFnGb04TAsQ8fOrC2bzd1JDy5/AFltzchYL3nAlxodQ6iR8sxBO+SXto71yAHPq7uWhVkimX
ggDtliYT+v3edMk3X3Ztb3oPQUVxHVpJypH3Ypa54ILcTum0xdcM9a9nbH+bRVM49x+N0ybS736a
hs7oM6fabZRIJi20Ifp5LgHpQ9F9+zeH8NfBvDl/3YjoP1+w7uTGf/JxDO721619mumuXr+LlfCw
0ICtjK721EpbpyieEQKJ6idPF5LYD6jsc3etd6kcMrZ0XIVToh7zVItvW1l90HpyAfvznEAsnyFd
oabeIIzWf3SM6xUDZjQKZ/iJuIkNtxHb/ZNsp+WIkBlaPa5HSWVYdkf2WbNPqurSp3aw73RJ4294
sy3wA+SdJgTIvU/ie4c/UvQk102P2qN+RkJPOFSiiLYx8Hqcz/HnETT6vI/ZIYddvYWAnBG1m6+8
omD6MRP18cu9XKm1eB6MkIavcDgDcukkR+PAT4KNw09lBh3jM6uod9Evq71pWwHzRrWz8RCrhxfi
MpJpLyQZbvWSyXHIr6jTDDYgQBhLAjv6nIDku9yoissNs3DXVVNebSwdyJevxkSQ463Ferda43dG
/AoLw+MssOJ2CMPaZryiaMNRt4fuN4JfgPfkGNR/5qILzOke4/fp0zT6qu0RrPzLXvWH4GZZhfTa
2VEa/GAuDqSXOS8NE7VD0H3BsF4Qkm/dJtpa6xNm+vBFj6sUADAyM90T/LUgSLVR2a54jO7yjRyU
To98/r9TrcJaDR1brPeSwPKjWm7T5uFElrNJUqGwu4OdIf/o7qSVVERbg0nfeRfL60f+ldFlOppX
N7ebynObmOx2dWt7f8rmO/fXXrt7CBePUITEMvif4rmV+s9zQO4rY4pKPtng128HGOrv/84VQq87
7j+TADamexlPdWxcNTCZuvc+LJpugk3I4EJNGGsAyOfJAWrZu0zwt0otns+/JU1kvgSsJOO/k42l
G24GFYqN7qJS9aPSbELMJ1n8FyDIekbQE7WONG8xmVTdlVqtiLgBZKqFxK486WAX7iK3ol5ll1uy
kjEnixC4mhop6KhI4mAQvYQDGWseCKpswc8gQ/Cnj+9MCEh07SnMTCfV5ntN8KfZ8oTFPszyG9RB
tzB0XyNhpPD62IwMfKN0CJgg6kEica77YeIO0595kUp+V1J4Q8CqfauNPT6nLmACEDZWMrCLbhd/
TT0uGqTVtcNaVtLsgHqWAQY3kTKCHQQ5cxn3crcKJP+yI5LRYXJmyXWP8rxhEzFSydUXQHV835by
hHot1UKiPlUIIjX9kEEA0rKglbFkf6vbZ5Efnyma491FpM7D4q/WcHZYjfQZW9d0HUtoyWG+E72Z
ZKeBTKOmxw1kAmE2RtOQooDvIaCccddfus3UEQSqenEPsfwgQFzbsreR3BRTPWTgzTSP3S5AexC8
jLzbWvTPDoB7S2HTdKQQH6mHdJbFxqM8j9ue29n/dh2RGsJuSyJWiybW/ybeF1enLxonWKlo0zRB
gtl63uBrmiYEGqsiZZKWYrue5jSMam85V+SOXMlz1i7Ozqkma4Ck457rOPcWKAb7Yr4o2brx8WZI
6S8KVtQavvmCTn3IOaNY3uo3mGiSZSNJUqFeIdqiKXwTC9DO/7jJf/Sn54J0Dk4HZyJ4IvXbJEVL
l4UKyE9Q1HTzbgT/JLx2H/gBDIU36lCshW/CahNxXCpWrmJ3M68DZfk7afMQ/+uHq5wkSMbj6RlA
cqPkhmObYnbdNSpvGnj80+T91LucrvGb2WNXe1zUIxq0HLgFVoOmLOHrJzCQSgGFT+L+njGGFkWE
r6a72ATKtBuH8kii2Vh/uI4ZHJa8ewqtoCS1ZpuQh+IvGJbtjUFwMIf4zxH47ynfSDtbYQ7GnsAG
kcqkPPlFsM4fDf5QTgGTgXvLoVgCkJkw3UlPZfoR21hy35dJNRr6d4Jl6qhHzYNyQZvnjjSl1ovZ
2eWalrJ818hT0XK9PL70BPv6Z4PFTJ5aE2bhMRBiazZE1qDBtgoLtMiXPSl2O5n/YeCYwPYhrNf3
aO5gX48gbQFePkKcHpSSDDIyN1ThbqdJQw9sdkkG5SqrxTDjZqWdz3Ge4bIVXXsKOukkMPitAHtd
ReRnhX5OrdtBM4gei0bu4AEDgOA+SzFkNkgSuA+f3r69M+W3x1bmwVzPf6nX0itfrBmq4hitsysF
iMTn8NTWud1Snd10NbtOyNg4yWdDbmTmJyMZAzL0MHevm9qI5cKyLX78+tTZfnWIP6KrjMupaxlk
i8HbyMmjVEVfwdwpfGWR6Kgz0eoCrKblP1fmx0+IT+lK+miISl9Qwxn8/rTeDwDj9Gcq62ZjisM6
YudpGL0D0E++5njY9446QKF61zRHjxvVmfile5iWEJmbx4mLzq1OpUG5yKQYjQ2pxnXus3mOd4zy
z+Yfa4MJk5onDsMRLlaGHYoRnqX6iouKB05dd3UiRIyYl62Jlut4U+320DJLQXbLR3IxPRNlcu9l
LTxmR4BzW3LIJkiprWpdXskuyI1XNn2oeA4nHG1dZ/w4mW0vIVLIylalQ7VT4iUC7CIzCothdWRh
Dds+mNXuQzdGpDyYxJYzbfj5k9siPTVxsEp7BImXUCjsNvrh6Da9pNEZuNkqpp6kWFCkOhxONHP6
areC6N2wNc0Dmp+nlnmA2fSUnspY6TJge/Mdte9qhzEQ2QzTL5t7NygxyNILVer50OulU4Mlv2XO
L7K4A6fE6GuPRUwXgNc3UcBaqg5Q+bnqVeexbvRUgry//SkWOCAX6q7hDHAt10/lwRkft3IGj5jy
+ZCV3v5M42OfqyBMZnIhd4SELEYCNigbS6M6Swg8Ts7Gr66fp300O9NzAMFmsb4XqXSjq4U/4893
f5VMiLzgUjcTA+8Jj2snb2iy8vqs78DFniJcwiXyU02myfRLXqdwGdOzsyrhDl4Sem9iSK+mifbs
KQB9y4hlXWddnSL8OqU4DOFy2vtH78VOixdYpxQcir6p0l9JkZXFLFEDfLl4/AwET20x297m1nmx
ms6xbZiJEsjPIIj1Y6OVXGl9R21YQal76Kw85Q0T/P9PbI/ozVaNvpQvJBb6xngcBwwNKK+t8CPH
fHWdPdR3NERkcQRaorWZS7fUCkXD2VtSUv2lJ/dDdGr4Jm5HUVETSfEMYD2uJ4vTopxv7WO2jGJr
wuvZP6EraBECQVCgSwoFTbmF4JKpE8aoY5wTlU7Mv8a2HcduMoHhY2jhLY54/i6P5hEWVC47LpuK
JHLG6RQjt1F5K87A7JhqzVtFlq7cpP9IvcwsJJU6/utUy3jPeTQrvLM35zAdLyDZ5wl+i5siYbyk
UrJU8BhN3BaGS83CZS/W5PiO0RUYPSAPNXihBR4F2mHwAk+b/alFqX7ade9Ri5kxGCZeYD0a6zzc
GqgvQ9VpfgIpBLPwyhvPoGzXCbFaFSJyWCVTsuaosSDn7Tpu4iSBNIQDx96IImlOx0BGUhnhjD0c
wwnnJwuXd9tov/8vjaFW/eEnvUwN6ddPnoTQLLa/iurIXSDOEirT5HuphXF+tg03Pi54KllfQ0PY
RX04tD/eSKm5euQ1HM/CF0V5ub4gezvndiuRyxbpHZTHUjOytsymZO3oSvzkigGrv+d0w0c7J3Pn
AccE2OAyBNz3pwTOWu2W0xElKJenU9zmF44A5xWmQrc3trYVnMLXsmg1GV7MCP+aWXw2Q7midg+a
/vY0LwqavIOMyETa0cs+YjGrz9cc/sYgMPdgQriCPr1XPq5dFSThYu6VK1lk4rYNN01REn40enio
hGXXis1NLXeCNB7OUucbQwVxG8NALKPlTyBzB+baX4fmhNjQjm/3uvBfXiqqxvfYfQJOKQ3FK7IK
Brd2qnr6s1wz9q+WkfPQPVkHMo9Q+zeeY65nCCNMBRQC+0qRuhnEV1c3+bk+1f4R5VFOKmAd0GuQ
+V1z5KeoOpwDLZmeLBDLtkO3dXLmANy5n//oZZniLqFee1QSbGwQHdA9h1r7AqFZW+Zmk+QV9np2
51J9v5dW2Yo9Ckl4YXhYwAX2kOQRjv7wnAraDw/fHO660adST9Hhxp6JHptvg2M/0gwdnkDFwgb0
g17eUrBegfid8bpJ1iPBf5O9Jklxl9LT1GYDh5Ir/R6p3GqU0x3cL1DwqT77j2fQCg9Htdix19B/
MMdCC1bfF6K2ngQyLGqiTBdLHtk31Pl3yCkLoWEqr9fivVGAuhg5Ffn4RmqztCPSCoZvm0p0psbJ
ryqctLGCsP1js+vQrAOKSKsqkUG96zL+hXwvFTMjgQRFpTXs9Q6zjKmdb8HniouT5c2Y9jtrMUOt
ZFdiDThobk0fHXnBuQ9E0wJzQDgzzpGaT3VauUif2aLMgB+0r20xT11k6BuM+XpCJVqA+D6tPcqJ
E8+DTcOkOXrUXvpLBO4o8dcRWpv40nI2DW7a1GR4Xf4QitMPxrnecjkl2FKWaeXLaDMT5z//gtck
nVygxJ6f5uoKSfqVvtQzzZb2L5hSP0J4wLAHButNgyb988995QS7dFtvlaSy/Rm+DrcJmsJX6SSC
uAOgoTWbOZ7ax5khZEoEneLk0jBX+1CI/qgWoikevsL0JpWSUMOPXpXiZwoor+sggAWQ+wlsuoxX
/R3L92na7br1HPzs1FgNdGrgSGGQgx5GLPVdR9e1GPOecbcKZ+JX+yVa7eyjxy+mU2UINUf2Rq1F
8q5CXeAFhmKynm1pX1f2gf+KqtfTaoMl2ThqSuQH+0XKe79dHIlQRCaNdROyC6PcqvvI/K1RRVAj
LjLjSSmlR7kE5MbxO7jknBpK3+thSijHElArB/+L1LGgBufTqtKi8q4yUzQGXky3wKwTXVWfpa2c
ukH4nmjRtHCaWdAUGeoVYvvfomNLKYuf+A+i22sy1kMbS54y4wJyfpQnKFFPgQBvuKyDVI8KDo4/
dAiCcODbKtRN0M5wvlnurb+ouAmvabIUVkfkOlJflLPq83BySDJEXh7h60KMEyJlaYCaGhvMzhim
Rh20R4NcXki4SkiyleyX74eVZY8TrtmAs7Z1M2eqr5qB0rLlfYYUY0J6z/BumqJqE8Fhtt/bm22m
qL/Y/y+3WmTOL3vh4s++aM17VUIqy4SzmGMaQmyC6lKajEZhDFTjHZo8AEdxjIM+M5ccJJyRE8+/
RErw+Jub4f0HPjk2DIkC+G4rXmhhxbY+6+KDw11EMxc5PoYcfP4mFYE0JwAn8LL/kPZu/MMTXS9X
WkUIQ1GQJYi+Xap/QWqxDtQnNC6ux5M7YcU8vjnYCGbxsrdeOq8qC3kxBKk1LZBizxz/EZIZz8un
v2XjVhzZDO4aqJ7/M4ZihnwO+vsO8wpz+/FyClLu5I9SdC3N3wwgLxkwj6tNc70QaPC2w5G3u9FT
xwJE3MncM+T3D7/SkqN3z2YeHEL/XNOseeQo7PP90tYgbWUvR/hlI0VJd2bGY6L3JflTLHT5KqEl
6cA+5m+hMUe1j2pmG5jBAGd1+I/zCF4NtnCy8K1aaP2OVnppywu8jALa6wH+U4EllQXd58UeJhm5
eQ/yKFc40MRsmRdbRVP0g8C+oiko5cx1dtGX7NbVFkZjNdkQdhIcXIuATNebU2eHp5o8QNbglY+f
AyCSm1GdogT7DoGtxZyqlL9e/hGGWHkucMJ7mRceKHRrc+7woh2IJYUOFpN8/pzi4bTunnIJTtlo
WJe6Zkrlm1eTT3HT4swCIl4gtsepCC4O9kNF3leL5NwLJrnYuHegtG/gDoQcwWbzIkLZdo2ZEOJg
ZIJ/flzMBpzfVOf44mxd9woJZ9OKdrlAHtabIY+dE8eKV1dv5yM1X7fzfv0bb7rj6alcyNDRcswu
h3cUQiPiaqRefHNAhRI97eqbhNnKnEoZAoVCyXeqsW4290jNRRWGUX08UQysM08OzqiY1kKaHS9P
AVUGGbF4DH8SLG94pqX9FOKA+RJ9/Zhuz3tFBNCb+Qzh+ow451M3JLN3pK4zmwXgowKzZ+gaGe3g
N37bTgC/iZCsPjbU3SzfgDvT5sXSBdcTFPq2GT2pgiLfq24raqFSWzs6IhGbYKbdE4yaQiVIb3bn
p2aN/cFdey7hKBvSVJLoBkid9T1WTtCLXPlZvd9UDnqJnTPG7c89BgzZCHfBSE6d4JMN3jbaPzDS
hiBPPu9iPeXInOhXjamQHPR2wY0pu5ofi7LOd4GXj1ZiapARiwx64XWJIRCMl/pNygwPMxyT8Sej
95C46BgRs2SNOU7bvh3E4a5SFJwKV/L3moo8dcW9DCbBMySpiRPhXjNX20gY1EbtrSERRiP4Rl2x
wHR8IwJHdg598mMX6vp6IQU8OMW+waR7bpZvrdnVtRe6jQ3n+QszKQc4W5uxKtmm6Hs27pvKuwQp
bN4LZT1zV7Z42WjnhSwusYbN6HOqVaTiUgV4ZW+UgHdAjxH0J08YD8BKl5Wqz5HJUr5P36gT/ryC
g1tEmayTBUIA+VCy8EfGTXHTl938WIHIk4d039vsaMmohLWmSwcdr+5p+RID9rFfKVfKnQVPn4/q
0FYqQqDGZPz6QOeipONdFwqw9z6nhkaT25fTao1hI4fYPjrbJ1Rh2+CLObr1Orxp/Vcsi3BWx0my
0aQ34Gx4+5MDuA3IoqiQKZGAW95EBNe3i4p7dqeZvoOcondNKXnVkuMJkxPJDfUbyZBQSC1MtvZf
rbth6DP82VH0nLd4CrHUW0svgfQ72Rw6oNylkDd3bDOBPIgB1+8yBxu9Mc7pMRk9t2c0k0wyCM3O
iJmqK3Wyt5MctH45N0sBoClqZrTh+FS3wvXIfckOIDQbqAiQEyePEYaKnv0gNipS9RLmFVeUydg8
deshAK7oGodIoHjRdV1sPsARqappZPxjO8nFGNatJ7uLUDbb5HNH6nEWSn60+9B+IAQ3n4+ILm66
3INjGZ36szdUCKY2t1zvE/HUBzYrDQZ/HJ3d/cNSKbNSMKeRDPd11Od3QK3Bk7jlo1b/1Lfi4892
xCddugWAn9QxtxO/80GcBzfqyJyJZwU2t4z70l/6/6Oaacu/F562goE22jeJoVFcF12A0KMZKecD
LeAFzoQFwnLPaMLim2dtxrEoJeLX+cQy9fSnVbVM/nwUKSYJU77Ht8eyrSON+KifvD3attWFbCeZ
0LBWBWaa9E8mP+erINJH1z9bZsaaw6ji9EVPECOBUOsXO6v7yx6u6AebeDRsBVKb8s4yPhaaZHI6
sWN2EtYa61zqZboyK7IwaIgpgGg3JEnhQe66O3ZB5tmmGkh4MQIp32fllTMX1qhCQgzLmhyVzpU7
Yl6qo8BjwYxPfCTLE/4aFB/at4F4gw4kbbl57kyVOU3pdhJTCtyuYYhEtCObUUCAt40P/g0kND5s
3I5qtRRSc97+z/jKmByEmxec/UglJEn47ej2vRcoQTbDruO7CVbSVWvepZs7ImMlZxF6QgJFL4Zu
gXEhL2kQ4di/WxB5kGLhEhfY+ne4JsagTMEk9ahW5QYHcAx7bbOWwx5MBr56ERln0LAtY75uUd8S
ah1EnPwBZCfigact9RKht1NUbKa3xFGvg6qY8D3Q2b8nYY1AJJnP8kp9lVP9vlzgEcxkI+1oaEd4
lLyjujBLf9dXpzeyO1vrawhxj/fSaps1RbWmNp/ch+EGyHTZEU1hd6Ik62c165CzHPTUjvdckpNE
N131t+saIwdMGA5U8Js/cXMS6k5vbMpTlsfku5OCdUPb7cY5mTxPGm7oQTfBqIOjY7hxEyhDxNxN
iSBCphSVhktFNlHSdhG1Zr5dY8zdJ5vKNAOcsclLadyRpfeD5FiBkv4SYirewygmEQYCU5t2NSaX
5aclfcCWk0RUEl4Q7Ecu78cqY2Z3fx8fHJ55idmY6Wx7U48Kwq4y7hSVXglMyKkMIzhQmWA4o83Z
J6OOtk7PthGaX95/khGyGa5LLS/lTuEky52N1WynDUgOdx21vL35A+pzKqvB+UN7nZ2FVvi7v00o
7FYaYfzhRnuvsISOOcVA/6bcvtDB3I9R4YueqJh+ZPrSY459L7kh3LWoe7feFyMGOVzhtvFe+4I2
5wMdyqgkZoGIFKpqmnsLMhstNj9HfrNZ+hwGj4q6tN36lQHzXBffJNRUfZUjTKpNwtyWa2fzA1m3
w1KTo0vi7JYTc41HGHKCPzJ41ozhCXUiKn7jGD4b/0Wb8cDYtmKivNu4tOCja1EhXkG++xURobp2
lFLFFMbu+OwH9+UbKdqg8K/adTV9H5dE8WJAB34zKvp9JDJ/4+j+iHAnBqYrC0hmZBru9nPTbcZU
ib4wOoTxw/+Exs1JfjI2Y0XGTmoXBSBTc7KnwQFHMKq9vXJcAdPDGFnICKN8wrG5ZsnofFYkXy17
wTPhaSZly+zkpXrn5KvvKG61M+IRE0SGooVq86kwJoEQuirsl4/v2YM+YVnRbwLzieWd/FgkJnhg
LzXTjB0NkDAIr3RMaZjgk7wboRefTrHaBbkgDaFykTQOhzLQcLgLyjt1m+7KE6Lh5RffRh0OdeWF
sDHDFvarFUo0J5oJeYc4ebbe9dawKOXhsYd+QQ1mKc7J67lHFY6EtSedcySWud0hf4t96+YV0M37
BRTPz0ma22mIneE1/jFGUdReRoVFGk0cBh92jEfU1/MVut79rVp0YowUgrApiHRkPQYCwJtvqsbt
s/SW8p0G1fE5tB6KT5pjJjD0B3ze+BXxl84Cvvo6SXTogye7P8nEjNPz/DLD0fMzecxrST8IyrvG
XaRZvAt/Nw2/4kAaltixjoWVkzV5ARgehfYEXxBahVEckx8bAO/Dc8jpvUB3OhuEiAyGbPu3S0mu
FOeLWeTFoKxHL2/SMwyim84mBbL415V4hBSEoKiy4EHV8o1nI2cJL+m+1yg1SqGgV7jkBsESyQPt
p0g2JYEVtVViDpKbqZxFO+E8uj04YPiCPuy18sdjWBYBZ1LSZ6xKyxWJVepznFw4U0mc72ZFypdC
D7f7n2U/9J5fdyDsrCUJWZo6cd7+2koQLZ5Ht1nX+gBXuZUmBcBVMVFIrS4WtkGkpyXY/u1/9ifi
61vZONcuP/GYBsvIB8npaZXmUCiHveqdFuvgpmBNVCHZ4080qRWqHo8oz9Gf3mxlonVbvg3riUO/
h7IJwNwso3oskeo1wUZFagqZBQlO+9oZbqDhtzTd02M+/W9V5NSLRCVlAwak8s3zlOxFiZ5R1r0K
zplou4QKEQb0yk49XNA7u8N20lvJXwaaKKL5WvjqfUjxZVKFvsGjz6V4WqAvc/YNCVjji+K+9mVC
vPHDxv3l9MS+bYKM2EovhPAuXT3IutpLc4oM6ntOKBAK6z7vfQf8WL3HUuiCJoDDxakQ6oWo3MiN
zkmhyHqLO/K7oKE3SFlP4wsVuBzsSCHnOLh7BQw9UPwthGWAxY2CPyXnV4qUSnw67T5mjx6hSJCn
/rM3dkZtHhb4DB+lYrtcQsgoGuyj36Y4HR2XyNHx+d3BUnLBGpcNJigyS0PRNDlnM8zmofIOs8fc
oFjhn2sMW6KQec4ADJNxIcoeGbaLj21F6IV3kG/sj60VdJNyb8joBBnYob6KMRMwcjaiHfn2w4yM
aRy55tmsxhnbxzLg5vmpa6Sf5u++KDi8pHaqrr77yBbO51k8LK6WuaXDsh0mbYRMforbqGpVHZ7j
yWUQ+EdnuLFwe+wc/eDWsAZhFVRhMHB91YRo6ZwnBnhpitGM+uAgdXmXZ0zfTOCt6DyKmHP0Xmwp
gi2qyMceo56zGn9NkzHFjuq4WHLqF+ZBC2hV6AESVf9P4qUF4im4ykqyqZFs9guk/T1y8W2DBspI
ZwwnRm6cnl8rVcWW7jCJxDalqfAjnJA2ggKDLC7Qdu650RAUo98giUjAIEsV2h3HvVh27FSCKp18
vkU2Kgs355JsWB2KBzjNg93v8nwGSdfvo3VaF7NaZB94rtK1xO0ijUByFf6F1cJQ9FDlFljD5Hrm
9Me+sbwFb+GGPL9yTKB10p/m5f3mTerPAVQsv5wSWnnr4pCI0SRl6bg469srbrVDGDYFWq+QhZQ6
XKQfrEaKR6Nz05nQksHrXnTsmeYTUr2SifFPaMCsUvx+OAV5iGvGH6Q0zx3JnR3AI3h+JQ04t0Ta
Qwmhgq1TjvhtCq29Uh++Jsbn17ICBwAma0XvOJ3iEux/6y8yAxmx6syls7ahOVOIQB51//EWgW2j
PocxPmNBsYUZ7sg3XU/I8UfbnE93XO096V32no2hL5PzG9pdoI4j8beslc/qsvXN9VqeH+M3Uv9R
v64bvbmji5e6PW6vmoWbY1DdyKpSQoWgR2CjEHcf6mcmkq9zYnfbJgxsRXw5dWzkWbcgA9awTjl5
OgtVPKlx5oOsp5YBJxfOa/LQxcQot5UOqSguP1S2po+F49ECHo9IMvBfy4Is3btkzL7DPCX69qJx
Nk43oRAa0rd7lN1ob02rbYq1GHs9HxgU27nTaWFme9Onl4Dck0ERgWIGbW0OW1s0qPXBoe8U6kNx
8pgsrveb0eA30Pjl8VUnjl9+fSZRzoon/t+KCf1tqjBujxum7H2Tjs1eicNjdkq7FMo6z8pXuc6c
o5yODGwyw6HFs/A6KiPCSp7rhHwSkY01NDBCtK1CBQvGj26+GhGjc0wniqY1eNPREgBItXa6gUuz
VeM7XcySv3+u62j8ZtNAdAkPH1x0Z4kJtzDRvWn2CFm+2IEgj5v/wSjJVqpKvOftWx/A6Cg1DQow
BQvaRk0A8w5GYdpgMnAx4kA3Br7zwTh7NX8cS1Z7v2yijVXvixXBSCGEDdP87hupXUflCwlRGkfk
oGNA6XqeC9vEIQOIbrjwHlFF/1uk3vQQ1Qn1v2lnXzx6qLhBh6mUFtEmr1ewHrOKyZ3lZaE/gzvs
o7/flHw2Rlj8ukaiIO99Ff9sm2ISnMUJUvXLxkU2azIJUPOCLvSUhlUFp3nJ9qGNEcEGEoVNMnUt
0U8lXPaIkqwuAFaWf5JH65LfKTj+UyPUOZaWfTL5vvVsjf6xvzzF+w6MRic7SAwIpOuhPBH/Vs/B
uMJ0XSDAF70hJm3DUBKr1yt7y9+LupuNwxaP7iSNwWQlCalEoKk4VtkAp56BlnsQOQBbRsyMS+yW
wj4HAMJg8kPw3qccNRcy6NKVb2NO3mBXO5fkORDazJlFeyS/x/sw+0bcBGMu+PFQmVhPhHFptmzD
kiXocf3PVTVQ35OJUv2tG5sG2FOk9wp7elTP7RT9kIKLCoKFqU7a1GJuQ/bmRboj4Ew8xgtNV7ao
C4MK6OfTok1p6nXRgaGUke/JANH3w2doHi+MGdk7bYR1rd9rDfqynNXiuB14gFUvMQmWuX/a2X3+
ikfPIhKM8pnr5yD4UyvFqK7boJVPT7TkIyjfN+Sk0tmVQlvVAK+4IrPAom7Q8GZJk4CFeHCMGXpa
9hrWiirv3ElWfxroG10Za/8u34cTpuTK9wihd82g7+N9e10UKLcjm+nU39hQDFG19SUcD8uFWIN1
dQANNPjbY9o/CJXuRnC/zCTOW6JSN4uSc5qu3MkTxw/+fGgPp3XtSjJYAtQJ2VO+z/i3Stjp05Rh
xnariGHI2D+4EGaWCenPQsgsqKrnt9SBDVCmL9JJaS8cOPt5A9qKaZ1NMHQZ9g5ozo3bUBM14+69
2Xv99Ipdgo1szfwmjeb5PMcOkThbGFHcCfXT4b57GoVNTbpzlsGdxTmQUWXCQH7GwTECEq/WOTBO
1V0oXZqFYqBw6E/bYODMAzMb/Udf/Ye/GbtYCiwVuJq9bx0JLMKt00oLCV5kl77PkgDC1jt4iJMX
msTaTOqDA/nmButhysYI2SQl2KHM7q2bkWlwvF6BgHoCiy1FRa+2HZQleY3XGzyjxiSxCDwr/9kP
jjfq3GiN42uXdMt3G/OEJ+ByXrL2Wxn5fMUIgbATbRETYBLlh7vybVdDIk2QqY0MePfSY2AX3YRL
rsu940/Mzemeya7FuyvLUxyfOV4Y39FuwS5g2TILbhDnDIeN3g2sdrV+f1y2l3pt7icVP/3VS7te
JH0eT2cVny4JH9X8/JHdhSQgD858c4P9o0sB6nLCA/pGSaSAeWvywj7BM0PQT6mPAosJexTuHhnK
3vQmDJ1TwKXuNF2fTg2VsR7XbB26BClzHxSeKj4xEqUwQct/eQS3N3WA17n/p2tnbMUWLLxGjy7G
YtgEEX0+HvKWodTksraZXEk0ux+C+99oM7s2nnZQxz2j8M/KIEiMBaUVLiGkUW5za+i2ru42WUdE
ZQ2a72c3qUAi4DmZeuS1LAchFKVV1QViQ0aOamThOJhQFbvgzs9mr+R4LeK5i4cTD5qSiLu7ZLfC
eMgMLNO8rpfQ0/q8RkBiBhvzCDD1OKWyaF20mo/jxk0O+onSTs02c49yrrCiqSYxX5GrNsSbv6TG
7IgzqfRWhthTkKO2bx353uGs2edeuB7+1MbJs851TASKeJG/jQDuUUZLVMYMmJc9ZzhskV9LjQHu
FnhAwOmOXMwcEI8SuCoy7nxhFUSKOO3ZqygJKQXGN6SatZTkHw5XlJnsqv9sZ8XzYZn3G7ZosWDL
ovGVBQwPWBUunw/LIZUHWXFQx6Ir+/tOxYM9JO2C7MNVoOocMjkNsOdCQU1Yb8U74wWftjs5c4hC
EWNs/WiGyxDGCC5SrkQAyn6XAOnsiscq/WuO8b2r5QFw1LtqRmUHx3ExLMURfVAwlanbLl865pum
KUE7PhWz3OVC8k6BkGvhKXcLQrmPfNgDChV1BvOqd0R3SJmq7GrH+OoWebWJx2Z91jEHw/dKFiB9
TKUJy8Zuo20F8b638kZ/jzBgO1pX6tmu2hmtwiduI82M8KC5E9BynejcZonKT9RPppET/SJOdo+v
KVziyYygDSJz2TwY88px8zUmsQJsMcU9+Cxr0SrLejT4JyMsj8ySbCMs4aP560MNeWJuB0RxD9n8
JzkLC8OxtXM8r4Zje/2oz1lJyVp1/7XzM4H/7bbG591jbL10cupmOFrX97Rdc0j+GuWHAx/AcWwb
P6uz2wvYfsCNAaNSnovUk7TzkiX7M4d5Qr3J2KeiOBfVaqWu0LHo5rYrQMrB9Vw4sd89PCIvcnpH
Ui8aP5OR/owKtcwLTaJ92yLMXogbexKnzyGvRezHF9tZbpQPvgRwtfUEiyvAJuXx4DmTz8P2wPnS
vLL/joGY/v2MP9bW4OiabiEJCXafgH9ozSfvRYFA0B+Z/iAOodG1orav75k2zrvxZsVbYKDSXm3b
/AoJAJ/J8Q3xL9yYHAMOlWQ/m399m9D0tX8onPqW9WxmJwZTpMAvI3D3pBPuHJZH/UjZ0hYloaoZ
epnjLGEWMeY5Vx0r4ed+LXvVGyEv62Krs6HzgKygze9nio6QO4k3zUx/gKrprJN7p2qrOpYl6xPA
w4GIddvhETMg/Vvrlo+HAnuwaCOuseoOUVJdjAzsoBN/5uWuPAiQhj3SjnlrpJuaiCQ63Y15wwfM
e+pHpsb/xAYATnbG+AYfVAjuz4ZanEkQjGDm67gDO8LdgVRsmsD3fgGC/vb3IYKgUMq9Sa1HZEe1
aOyuf2HbqHW0sFVtDXu8sV4k4MiegeKU+ESKY+CEKcDTReOeyvDRVzImjVE7ctBuvqJ0kdvtj0Fp
BG3keAk241jogORTW3KQuYoC8BGschTSW++JOxSBjk58oPQ6y6k+4CvjrBp+mftQSXIVQqi9VlJY
DtrFOeBn5uPczr9btaMpvDV/xNzrzDZigk0KS4/RtoTN2RkVCcyx/wjlBHFSjefFJGg8dtL8OBG1
/Xtu60Atm707Aq5QNfM4ZOx8vpNB1ogR2Y8aRKIzu3npt2kcyvBpsnhS6gS8B4wco/nfFy5PmWB2
tEInY08M/TGU6QXnaEMgTgOgUypv6vddFRRQbHGe3Te+BPKuqRwh6uiqVa7Z7SIaexbLshI+XzbZ
9ZqAhVogsMefCPZstzcjYpcS2FpOLyue2+A3wsbkvYe1VezO8IUuXLPHvqyEywXOxSH3fcpro2Xd
z5jO3eO97oL6VRsJmnO5+O2AqZlBlOEzYMtyzAy9ZkUANgD5PKE4878hsYgeSaqxVPXXuqrFCIOF
mzqPL7HzS3Ypzhae4jnJkkyGvMcHxLhnVsZ/zVaoY+WLObuWuPiRPLRT6er8b3Gt9Uf8sfckoDKW
KCMgOUfBu5ox5K+l2A6q8dtCFIARZruphv1TPaUu2wMMj9LPR8V9o14OQAi10pa7PEiMD1S9gM0c
TmNyFe+GJZiM5X11aG8kXIb60AxN198ef3vXKE+ABapuMfRWEf31IqxdyuiaTda8iDik6lH63g7U
cx/KLd7/46IkU8n9nOPT5h54l0NX34PTlBKMAQXegrc5XKfcjqWg9jIqrZ/Qxv8zuVFHpKoUaqXV
9ZM0VNpyCUnkk14c/0aZALKvhJ/o/EcxCPDDubw2A7sXiZ8UyBJKle3MeI21+cRyq4zkGbotpb+8
U45FR6/YNrbzzt+gsnkfGJrpygSCDwRGJ5BxAfUywCmjhmHsJ3c8kIQa4lidsCAkUeNvVx+t6y15
POVn1enQf8iFW4Yc+nBvQuL/3e4IGOBNfWTHE7FGT7Pw5OJPeU2f22mB86MMsNmNBqIg2NehSXYD
qB6gCB6JielRtm+7h7it+WMKT/g6fDvWm9ZpNvm4/0i+mp7VVjKmvFm+AHYJHyWLrQ5Jh/BXFGdS
9oTti/ErDh6ELMWmv/iaZE5xYgAnOFbs6vwUu1FH5xVqSVW0G+PfA0UeoFkdak7sDudPc9/sAur8
34X15PrFjUYFPLN8J/VoTdEtw6mgvdse0KU+2nreZ7AHU+jAmaK0iYl8Z+xnjq4PkEuuB0yZ01DM
5ApA15AmaU7nPe1Xe294Lqnyil/ZuSeuVmGjewIREtqmDxOSqVXmvCQh41Js4nNK/5vteOjTsS3y
CTbshOIKet+GVvYUrVE3MCNQFFXDM0mR7IUp9Ttac79ovX5UrVMbi0hS+jioaC1GQ9q7lXvH0fO6
cJ+mKKjNR4Sp6Yd/NyGN0ijvsSWLRTVNpg0V0DBR7bWvCJu4CGg84RtoDJOehS0iXe/u/C5t8Rbw
zCYNu7o/aEm9yW60ZQy4/GnuU9dVd6JioeW8nEPAx9vukesedOwB67BOQ1gbD8OLcPVvuAMltOhd
CBro2JLLj2CDKvLoQaSK6fYj6nrm+v1fUv2NuX6blzoqv1otUMciQZjQJxfpAXQqalnR/ZLebxCH
3y6s5ODrpzdh5biUSQlBQqqO1XiLEiqJhcjjiaxf/Ofsz7wdgRItR+MrRBDSe1kq2BicCPLXdx9X
SInHTItobbR/IUSIsAQlbEaYe8JYFvWUEPsl7WXHL+wYMDSfvt1qOaqP16NXdEmXW2XuvGIrnof1
DXGcU+A4of5JXA0WePaGMzvTCVARX5DBjtYG6cjM91+WfDgd31a47RJ+6J2DTO49hf4Df4MuPoLA
ngM1Vqp7PMrWq04zGjsfOvi7f5JPwspXYZr9hsERdpBO35//72JUGya2312uPAzInNWcWO1+35IE
Px4Oa+1+hC9vBEVp/a/gpNVhfwtPvaniV1qETOqLNgrt+5Vtlq91XUjiFsUvdAUC0d/FsSnjn0Ms
tmuuANo6Go+E0/gnki1wqcA/pXuPaBhMCEf5zhNBw2LNK5hgmBVokJLhr78xsVBZ+HsS2QLdRrJT
GHo1/oXHjwtQAYTDMCshL+9AVMS1eMGkxDrXct0/m1INpg1+IXLlwkTzfQDbbwgfpmB0CV6Q6GYw
7wb0wLZobiDdHXTWO94Dx1s/Jd7fect09N8j9mN4d02mcZiydye+IduvHRJZAdwfxE0+4/3S/4Yz
UkPi9yU0vYC9wWIQZfoFzaDLEUQ7JgKyzobbA4LKnh7PjEdK3Qbb9hi510xMKXc/HsPxLo1VSd5q
Yodk8Bpa7Zs5KZ9OpPUm3ecvez5v+af/EP9sXa90vdxsWh9gPVITNQofUd31jymJ61dj0eaGjf5f
g41tvzZziZYyVzeRCzli2B4VqVaTUyKFZUl6x+oqA2OQwUQZ5+9a++qEu2bPVj1rSURJ3Zzr71Ej
SV3JQMFNzvEIAnFnntVIS3KcWmrSj/dy8ls4I9u55K5PUL5rEfOPjfYRsDbKG99NxxW78J/h/MfS
bHiFz81OADpcnI0+QHtuoceiOcj08WO99FAwnZdT24frxmacfEtOg4orfRGU2L8ab2bHucPDTQNE
xnuutewyPpXCyahv1XHiptv3PwnAImczBB/t4ozFT5wNMfbvFiIm3xVroq5dwkHYUnTyx/W9grj0
FblOlEItwC5hm2HTQGwAz1Y/vKIHFTVzEgahE9SwT8ge6lmmtN6ZyRfzxK19I/ULO06Cmd0siyri
Y6AFL+dBDmml/4Mc2PF0r+6hm1ja3X8SDVQTvPsNnRe5440ncPTmd6L4Xhaa3evonO5jsIJay/zk
OCuz37U07Z6ha+dsq5XYSfwx64bNeIzMHkccqd8cW5lgzmJMs6u0LZiS2u0ONcUMSaOFoMTc6nGA
j9BRnDn69TnTgKawkjCf9U7jJR6B6pjEGzDnbVRa8xj43gMTiN8jxmBl95ZULfhRdfs6GiIn5NVv
t4dpvNgz2pRwo++Zyz/dRawsl2c/OVXt06dOQaShNBvWzqijiCgBRcC2FDqd6cZCZBKJc3yaPWp5
hhoTBuKgaOl/AY2dKxXSxOHTaoZk6Ovf3ao8Z9PICT0yw2ljKRC9vd+qgWcSD961s7v8fRW+8gxB
qfgLXCk7Zg+exqRSCjovvnM21W1FfX1X6BTi7s1lP9MPKq+crWsh8a960Rgxf6JI9/rwKB+OCRtd
WpGrsCHPRxdHWXDMnMbGYgiNQKpPjwgubXJvFrkKONmiEH+OKnbI3PffgcuPeAjsA+m4KL70RcGj
bg14wSqCafg/NY/97/u9mMJvN2diLwmG23d+TZrmjx4Yuq3ouVPy0dUXp2oa+F1XBkIeL5qzLgb+
RU2wz+MrZKwTLaSBe5X+l2k/1BZK0TFj8PlIrzisQcGpXA7R4JZNmoiuh9MnH5TDaI1FSuBRK10i
tSOqbapiuvCnzwcv/9+w2WhhZc4CMwCZIMx7w62oFTFvDOyEUA1oy5b7VDgCThRGHmGxsVrUPaXi
5XvHZyScq4/eNBBjNdlCf478WEw1qyk5tYDZ9Kwl/KnDDF8Ynz1kGIZlDXju6QOnEa5yaUhKAoB2
tEI8/SAIeyQJbfBV9/zYRfbb591RmD4zUR/MAsDr6Uhuv1XTc3bOoOevCTxiDLuEtvJUt2dlzjcc
2FIipXpEHAC+KhIzpXOruVuWnTUVOs8fwcJp+6Ar5DfQYoot+TBJn17QDuV8s1jHYnqKK3G4QlWT
G+BJHRYZBa+scpkx6wc8qtnUPJWQa+vv6I/vpDhob/k1oUMJr753otTe/GsCHXY+JyVX41YRtj6G
Y70vFf8BuHZd6TXaf7NXN7cTITmljhByAcKwalbOL9SiUN8lBSV+cKW71oDCmwyNBQrVG4GUCAHM
bvfQZWb3V5OH38+34LUQi4QW9cL0ERRyqPOadr7J8wTXdfhFVheo1NmG2/sEU/kL4jyVXRNp9TJ8
b2P6BIcoH0Oc0mWNi0YAsWLIql1vxCn0gDpLXDw0ubB0elnEVlXB63P+/m74eLaGIf8Nd7Ib5+lx
7UCDyK/kZ1JC+F2uIpOIRGHWAC5J8EWUFyBjZhW+9kCbaPYrToxOjTY01CSoT//VLmsyvQbIsqIi
bLWwD/tIuMg6jrI5hrrDOpx2COyOT1koh+Amtwh3St0Sbon3ztFhhSBWXAlbDURey8wnJ/1CMO9V
XDpaYThU3hII9m8N6ej6dRacySAmlDRrrJFqM5vLGjsfJ85tVekghy57bMYTKxwweo7/9b44ntl5
YIkuOTsuGC5uvVc/wW7lyZVl2r1+gacB7RMYy62O/4uqxN5xS9jr+6O16idZ7l7j9iybhdjxuVjk
b+XgicujLjm1EOw6u2t9hAGPz9wgRTaiY0e/MvTn45ti1K/2j/J2GZex4nx/HzPwKn3p7YJhmwSX
4fmmIG9tbTQhpXbpLzDCp4fEuCbV23PzYw8QvilrOot9UJw9h0RhvHas/MYafWL3UWxrR5vQWYzs
UMZtaKNyVqdAwE5mgy3izjdrEuKUFeAtWZw0JejSaOUAR27Ufq2V5JLquILGALmkjj2AFORS713L
5wHET+ebGnTuPd+GPLEor61ZMCg9wk43qMrWQwsZWLX/hX0qRWQgLAxsYlvzDN/BZtJs0qdPbGyR
/jWQwyVjsaP4dvXszwWst7xSDdGZzsuWXpy85ulnRdW9xzlD5oJPl/HQgcx1IsC/W9J3ScxLeHGu
Xv7IydFRKY8Z9a1I1BrfwGbCQHq350v5Ifmb3MgquQfexFuezayxC/6MoYFAznDwWRSvNx+te2US
9L8ipE88CJ1r0vq4bcGBy0nm1ZfQ3k4Cw6b6l5Lj0p6C6SfuBPxjjRxTjVsWdJRnBpAQGdqgPD3C
ATWNnAl10hE4yhVe3A/J2RGwlWySGmCnvhLFEC5ytcUrLpwsIxJ9IzzrGO9alqODcNypAVipgySy
rJ1xL7ipwLUGDcgHrl13YFTgaaDlcyW5PpfCs+oV1uLyMiuUNwOPePKcEUGWaFQh2OM/8eSYs+At
iAWjI1bWH6p+JdkgRB2vNuWXcLbDqphD9GLteW062lFI1Au/+BnukZPKfLFEOgz5dvu6E6aaeYLi
WT1hhk4AY0RoQSXmzi0sSpj06HepF9H67hRvqdNLuSvixfM/p2Kx7htWASO8wUWDtTf8Oxlx7x9c
tUulxZj4OgQNtl33w3P7DZ8k533d05BewQbv8AeLRHvvD3BZb+huXPLHUEu+TD8RdhjZQBnXJIfU
a+BXiXLCfGPWr+QcYLIdXWqoa3T8vVvBgN9ECRyQEW9PCRP68mjy+V2Y7VQs2vO4NtL92CgH91Wf
EHFxCvb0Bcjols+75t30gWx7kGn4/cSQXU5XrL/1nEt/aGRdcFz1niIv3gXQaFL6pG3DC9bQhUoK
A5x1IhnWwTd4+rSpukzlgKF9yX/gDZPVqPKVZkZHUefp/lI/grGkkEzjB1TZ1XNeWnXYjZNzlVa3
gvGlodqlUG/zTlrqnDTIdtP9cK35aC5mTENVSQRn44wkOyTlEPEXTzE6uFWzUECWpdDl/2h0tncx
yR+wmGcBP21FnsJf114DLitn02Y5aqmWq50uRqu07U7BU3/7l9ysGLkjdqvpG2FTZnp7An1mVKh1
A5IwuSZkPxHbctJzIXei1wQ+lXirDDmd8kee+41oxUaRrRFGWk1+sC8uRHP0EFXP4QlTRW2NzWGb
PPXK+EXZO/x7c0GfoJ7OyzPH/5jNZXz1bZRh69YX+Xt/X0lRjSresUHt41wQEvKDag1gL673kL9B
Sj/xnkVoa20DD607E8GLNtAB8lpjkJOWqP9jsxJtZG9BVOwo0IN9wBdoKFmtaOKjlJtNaBesPq+j
wjJDUeyh8kSyRcRY/si25TYR61P/+jBUtEPysIIVQvq8c0vJ67UYL/L4xoMcidpKTwdBjU6diS5j
UPiSJ1SpnBHQyiODzgjOwuObktcXJuB3aTHf/k4GSPaernRvSxcTQb+sCxON0y7CQ+IyE9+BmBzH
4ZvCc9+yI0xfd8IgfHsofZWzW2SrdmKHOUsJZp9VU8DJuLCcJ4sz0CElGgO4f9Pt5qLc02UJVAR0
7wPmMSrHnVgXUFG5Aro1MeW8rCfMSpG0EQiZ3NH6P/Zt7Tp98bHKSF7tNZeazkJq3kJpCoEHzS8t
E5qW5zPxIiy/fybYgcj3vLTxYsWfHDGwK9lNPU9n6/HAK1EZomwccd4x4+jZIed+DmImKgzQbAIo
mvRUCmkgFTa+0AbB+35dlokvIMpMA1qqCe6XBY3h0FnVQ5OOEs8mkuWwEtaAn5HdskWIEikBQ39f
TnHSFd/z0RMS3Wzw4Le36hXnqoam8Cxi58YTMm/EOwLBiXiqwkammkxNup9bLfccWKLagBde2OV8
1QEU0IINRAuCOiS/3Pfabevq9Jc2l6VBlYYMFlduBb9RMJbuglRko8M98xQ4Cz0toHBzeAqKDQf3
PrFRzlYUI6LuCUq2r72prYGA02AuKUPsrg555i2dscqZ72ugwlJdjceTIk7Fc+kGMomy0CoPI04e
3hJVkjdAFcFpIGVbM7IuvXWN+rtLcZ1GoBjhZA1xq7X0JeirkVhBDebFkOWr7uog5xk3wMWCKci+
zs1fzybLqMaISlwA0cBK4OZVPJcZj1i31sZ6J6aIN7wRDi3VwXaJRLpWjusdmOQYaLCtSga2JbET
A07YmWOxOCtXobH7aJj1bB8BlA5u3bJu30RnuVBxuAQ1prmJy9x72g7EpzU7+5SAkpPLiUg6buHx
QrnOHy8er5+LNGbveuoAPRG1wMHkgkxmr490tEsMPG20Tkpf2RFJ61ZOhxOFWbe8bU+wgC3TSUVN
nLtttRRRekJ8m9ceZEIIOD5nYORxkPnyU++A3VwUfQdxYjbAmUxG3bN4wJfP96sd0ODzXHiBxMsH
YEkCWEkId7pgd0wmmV7uMMa8WS25fJsZLz6Nr7dEOGg4/it6jjc6XSUiov2HsBqsrsffWPkuow4e
yvaHgmDuywIH9j6dsIIA2Fpt/N54VVIVb/cDW4p6A3Pm+iHXz8PuVHkXdCQuItl6a0Od3Z6zAEGZ
/b+I/tOXAqQQNutyQrYC9qC96zRCepQ9HJ/CuB9Y7zpfbm127kRRLXqzF/GpfkLqYPMTK4Ig0W34
7QjJnJ6lNJHmt+8aquEsXPqb3izjqvqIzHCctj3t0IsWIM5pi7RvQtUscSxPBLcVxpRUrsdSxfpi
BwOuNxYajkK56gqsDWeFY6HPqVyJjXmREQZ/mhnE1K3h1SCD5vSIUVml3Wkf0nk6rEBJgIpH0mQj
WgDogBGTPHklarCxO476ZLJukcOF3k3liiB3Hctv69yiQBPG/Tu0MFMxjd9gMgkGry99Bj0erKR4
H5QVtWhYqwqbFM+cLe8x7cLc53TMPXK228HSqAuoU9fCu+dvPANdirXqSnmQjE/OTACL7ynLtq+U
FZhZ+qKIPIYBstniwWiLt878wO1JJNFGNtmpXpi0iy7kAAQcnFaFmP7NFOd4gOulGpq1Iuw/nuxd
rYUaX0z2sQs2ZN9d8Ltfhd00VqUSyZaH284hL8XnatBS3XOW3MOMRhdXt98f7u3E4ID/llM0C4G4
kH9jDa3sIE+zSZFZ7bV6l8z+AhUcHXNX6edVMEq0nUkYdh6RX8YHIRnPY6xYuDeigJ5XHO4F1HRs
0G+qIgYPGuwrSx1phTLt67CBr9ZYxWNhAJMBwLf4uYNrCbklME218CN8KE9HiqOqwcP/8evFtDPM
VbCvwbUzoG+zX+Zslh0SMPFtl/poh6uOjDKwFUhOGW/jFKWRNh6dj60lZEaFJ5e9GsNR4uwafAsd
49Mf4fweeo5Vmh2OHm6kIQIq1o+zUTp5OXxCVi7PHlZkfNBi3+aiyU2Gt9AZPDyL9Pp3MtCWsRqB
Pi8SaZXL/NlmTv0sEEnCjMDwAHp8mub3/vMmarjlZTbVPQbgV0vEOLiCX124OfGJJbI1jKPgjj8b
mxE9PGqgqfUhC5YMjmiXiAec9Am+CIcF83h5HCqgYXRHfmc8ZuugRGQZuyODU6qQue0jDbXkq3X9
007BXwT+EkbVtjATQddmRQ/CFf2fFc/JehCezWpFzL7kL35qCX0yI/QVfe1BOvTZEZtxmraJqEcT
YUD86J/R/u58LbrHslyjEO0NwUs1UQZ9hAufpHkiJTfqNrf3Ur6cJ/FZcaiAA2ram1LmFFdgAv0P
zRPjAIy8O5wg0WoGdST1+nWi+lEIY+fKV8Ymqi7YPFm0Ndy/hyPxwT0AvkQePhy6XBpTHFPfM53D
M54/rZOruGl2/GkdrU59VLhzTYIvJr2TQby9Vk/F7uFIJr0UPLHbe1fcjVXfJ1kwjxZ36XyiYG5O
wvIVt/9e9zqvwBZz5l6fW3vb09zBVOVqrvjqvVJ5Q+6NNn+EWQuLc/EbIH50fKkGrTqakdl9uPWS
QPqEm707JsNeCuawEzhhDcVjXb2oqlBKpjoecXbUIiYXjneogDUSvwQ0qOgl1BgfAz3f9PfUZkTm
UafG+V2VinkBiGvPLB7jLcDwWiOeepTTUdgkKGpH7FiCIn1dzqyKRuVYo5JIkhDsop/NjO6W/ddA
pza1Lw/XlszdNHa18631DBa2qAnrRgCqVD6x/wnbNTDODjtHhvY33bO/cvxVNT857uy8Of60pcjP
bSNUK0j8TWO4WOAKi4iFVgJ8wPcvvUwLd3jg9e4J+jLVhrXbf64KT48YkWCJzc13Fg66AerS3gt6
jfmFGAsT3Dh8Gu/gYy+r6h1toFsehRE1OvlWLGv5PDP+hJhBDkEJLNYVt6r8zQGWX36IRNtmV9Zq
Su5bN770x9uv0MuYi1JO3gae9fMMj7XxnVy2fap5qYg6tRjrZAqlAOcXTeufoFhti8Wx7zK791XO
xWHl5KcXJvFHQ5EGc6AWXs6mZ0gYPJIBo+C865CUx867pD1ZqYL2tr9YAxEzoFozEe0Hgx8Ogg9r
aSHcQS98HPgEMxOPWddQF8py8BL3MLhSCWkV3j6072AGHuEhaB6e66i+OHO6a0Q4nbfLMcLZzntQ
/nZlFecV4rlsk42L9kQBYaVbxWBhB8YH7+ak1JqQmPlaLIBG6i30K75DNsj2FkMRA9UaOnXPdys2
L9Hb1DT6P4BY23HyBzSVxU4gztB7Bc10DetBqlL/LG0xei/etoJZnzyXtjOepYSou8x7lpbGL/Cg
E12nnE4fJ2BgBuafxeqN0ghWgjsy4osJbMzXMxaJj2+kUU+2+BrmgtG6Gv7NBsY5q3EYy6h4C2UM
2sK3gKqLVC0DA5gW8vZtWbg+rg2YAiOoG7AZgXxD+4g0dgRbBf8Oo7Lp9TUu9XRl3HPPHQXBiqQh
wrJAqY3zamjm082pAzXVaH7AUhIW9UMcnbs2s3bk4VcfaQE9to8ymTDvwNsl7nBiPBhExJo+j1/G
l+FfI85Y4tTOxHeYxXqs9T0w1fjEIE+MdZN7xYgX4MSEgPcMvvbm7G06aI1WefBoxcDjAKJUN644
ZGMH9FlPxt3jfBmdmNKJn5XiBQ35d/LTFz72KXpQuqzFjNQZ3irgM47SXBspbzrYk1/OFB87aIdF
oAFU3Bkx7E4QKq1An0KF164or2te10gorXonzRjp9ZiWyBiWWO6SMbK1Nrd4UwadrBdFUoFi/RfE
YMguXyKxhmFmdlVOBrOlQSLi4LmrUAhGYvBIsOB4GZkqOFaIjT5RkiR1pj3O3qVBO730GYodD9Tl
Hys3b9cIL1NFmjccJSOAvV34nN+pO0kzmn2kuvWvGeGRlJzU8nYcxzq+j6g+6PIAxA+cjCK7bpXO
gBV+Ort7TUaxr1g+w6rHDRU3PC9Lk1x9YZzFZEvNgrFxpxiP/pwHNiBQBtiiKl0U+17TAvJqTU60
6RTXuTB7rZ702nm5Z0+PVuUMnX9r/5UdZv4buYGHN+k690/7LDoYYR/TL3q/76K6ppdMQWfchg6t
62lWz/PtFrn7uwEtQ8nafGLtcaZbO5UHwbZmfqQh60VEIfO/ZXNmwJmA35vBXvMwAgarYRGcuc3d
Ry4dMcpTuuLvmdn0lRpirh46c8aSGkB7PCysRzRtD2zalw7vYHaLVgK2Ag/qPCl5jvvU+tvbzGz9
3kze+852/3cob8iBgjB47gtPBc+gyGjoXwKUj1xMoTBiq/7fHbrpCos9SEueWoojtguSQhDSfej/
UzFhT8r7Gbpjbg7IFytgpAOmTnpV+cfHunVfyQUehwSbumV953nLpeSR3bTAjUNEUCMQFAq9QwCO
bQElTgoKCO94HXi3TNNXSNd1DQpH1eaVry00PIvREnYTWQqgKvp0pIxvACkEZW9oYm7Ee5XyZW4o
efWj4TvdCZO60zdJCf0/eOs9xQB3eEO8aVVej4QtL4tkiGKTfOvPOLURfKGIAnOEntufbTmxlujD
WQA9mCWhZgihda92B57EEdpveu28g4FdQhwucX45JM4JdFIIDCbCome6ZvwDwhXb7X97DMBb17SI
qUe9HcnKrSdeQ1vH67jEZ4ho09ekQ7jw9lxTFxHJ+eqoJk903rAuqSbdbzW5O/+5u0mIA50GY6W2
UN8l6T3xA5QB+rVzNYHGRBdG1WFsLtS0JlUvfecA6534LkwOvzfMz1FAYbkc/RiRxqp77oBJ6OAO
uI2RhgEOOplFLeFT17w9e9iGqe8T4e7tRdo21677S9xK6yC/ohqCs+V6r4mklSwxzeB2VEOuwadT
zBY/ErGWngJ6K0PcIFaDBTmFkn5aGIlv63m0bmBBsdnfgm+1XcjM4Ss0wIyYkwHXCHynwb6uKkWd
wAnn+VmXTL8SGASD92aPTYHH7Pyz+ysS3+ICf25+EjsHIR2bnLo4qR5vfog573vkofOC/yX5IwEw
yvOZhAJzY2my24d4zp9Vyv7RHglzyCIigY9MG6AnZZjYHJjOkme+ITJgPLM+8SfiQC3IWY3EsyYz
z/D85z1U40Z6e5NtiwsH2G95iE2qHCifgDegUmDz0Gg6tDvKTAj4ga+VlvjmsIf/PGJzdtkoFN63
BVP5bZ/uQQhIGZ/HEnDXqlTgPNQJfIDyuWrGSEDu+lMXAkZYEwOArIXN6HSBS9CCwxUyJl9AWyDY
jLvSJ4oLW1KdrEuuyXU9SG7efj/NuHnkb/Ofz+ISmONW/F1kXudlAVqBSq3QcUsYjHQxSeXtkYir
E3alrGTHi9wJSWE7GKuWuekD+FoZq/ZndUQxDVvrzQMMwiukoE2Gk34TrsowYUVh6f7J0iXuFoYK
vm1dqnMjp4+pSKE0iSbvOo/C5lmXKFIDssmbVDEJtFhS/i/uCfrYj98ZotFiWLbxs1XLnsbbdB5e
aTZJaVy/24gj1I0cOm0LyS5my4cYMV+JQa+kDe89ctb0+8HWylefF7FiLobPqtnGMTv7vIGlCY0i
nhUfrLAuJCQph0C4YuKXd9W3Y5jIRhR4SffLgXQoIZZegbgWWJZ5CP5LbXwujAK+mLbQ3/K+tYGE
bZSOGQySTQ4OO5MstwxKo6WMxCZnFD4jHBxX8OjMRDEZKMw4VqfgvAIyG1AXFP4PfalvMbobIprC
82OYpQZWOBVj2JcP17v81N0NRJLnEQzdkXNtpiwFcmqAAtSlkhlTttCiPJmNCuv0/3FOSEP9yYFC
OscpVTyDXKUGjzLOXF3pOf5SYDr0fB2PcTnyidvTMR2Z3U5jk9oSawMf7jx54k4TQ7RrDTzSdR+X
g97chKSzXPpo7qnm+YjJ2DOt+3qHKR2gMmA0Vyv55I6oOxERTpDZGhX4IEaJum+Mzh72KhASM+PD
nNvPnwe2257GuEXgiFO1L/Nqs1nLQ4NMW8ITKK4MHDRQcyJqjfRlCEuHr8ut+HVMuAAxIFvtct59
ScdquSddUqGztCDeAFIlzvO7uYuUWG+c2rUdwMOa9l21lLtTCuyUHYkvCS8jrlPJhGTfZTcRimXu
AwRv3FRu3O79XFVqBPHPaySE5vTtdIHGZY22GAzBMvPqGy4xY1Jel2xx4tLa6EVgWUfQ0Cig6Djq
z6ihYBujtEgekPjQiGULS72iWGbrli913QwVkIkC1IYDLHPze2kW38Gduldep11zraFQ+/D5UpJ0
yhou4SZz6Ic9rSVCuyAd2aVupQ52CSz+vY/M+towYo1Gu0dDDcDxWXFDbmDyKg2NogoPJZoCm4jx
0ew+VOCFIcTWojVv4KVH7jmaQJ4QHrhwIXCIs6W7hDu48IcpKJhrufN2kHdpYSqDvtL2XJg087nJ
1L8uqjC/AmFlyJ98cQRhceBdoVnz0Kf7Bqwwxd1wa/Ax2px63fOxjqQwqmw+LmxXc4WJX0G6rz4g
1QTQCy6m1fDnRidHov3oQdnH9KL7Py/Q/fU6e+c9wZwiJuBGH3QemnI7GXhA2tx8SG3l5YYq/TTM
EH1f1ar//oGr/QA02XXnR3WWSVEi6FXq/PGHMKwtK7Welv0//cf0wVJxmw2MH4NNFdvxoErvY/Vw
AxmLkXWCUH91ZmtpJlya9Q28NebubuCok769dvIXAn3LVKOByoS5ZRnu9S0tddE6kO2CnLqmV5x+
afJC56T9zM5bsDyUVwC+qe0q/2DinyILXgxFQv1/g6tmj59k2RRgPshx6DQl/yYERILCnY+GZDaf
ST+nuYjpCH76OmjQr1AlanNzcEE5WQ31pukzgs+/Yzv1L5+IUR2u3xK5lJAEazwyJQAS4+ADS24s
+6abs24EKenQh8vye3Wm06Ewg/3aoVlggnMBvZTIvuq6xLkM7icXeVz+j4P3gIb/7VQpXdah163Z
5akL04kEFrwywhrmzTfyHcQLWWa2kgo2pJ5JR7mNVzmQSSpm2Buq4SHcTPPUx3ZbukDs+fSa+hh2
6ND7sw854PTzwQ4IBj7iTWOjdy4waxGgu5fFGBufMsNZsHxtw5vSRUhfp4vjXpi51pvEHIBkUaGz
QQDHh0UqaRrp0TDH/3N/N2zZe45to1Q3odwdVqlAyzs378ucHeBQ005hBqKgrDBhSIQJWkKw9gTy
boIpGbOb8aVg/ilrFkzbAc3nWefmeNegDQPjt7Rru0NuaWJRL49YKPsOULsB/cd59TavSUdaNNmn
F2wCNAog2w1CKvZ/YE24ir3FnwatMCIcJjr1YkzFzu5piZxKT9LFSMC3rripL6jFaZsmWhaR4VRQ
+rCySNcjGKW087SPtNd3fpEt41AokUErasKioj7ZYiNGdMkfXc5aLyTexbHhe/h+puJDtuEAVwX2
jh3+rFPv+GJwXrrIsgxI+8obIlGlr9ZQV0EqcVEFZ38edLOJg0g7pzuV2IhRs5ocaWrzBz0p4ysr
Ufcw0SWps+dG8FI6zYg2vTEkp26gV00iR6+hMsSMQ3Ce6oae41g++PNZJfm9oGrATH60B4bsfOv+
mOqHVLPyq/Pd7+vVflE203R5Ln89smFDKQ9/BXC9wyZhdMDp+HokXGnZoe29OxhoXzT8I523GV8Z
U6pIAYeoJpp6FHRZCR0t1Z85/hPRJs3kNk3Dd62um5eEJQ1Y7lAnkRXTBTwvBTkZ9JEzr93q/TDJ
SoFq2oBwsMt/gSTQf+o5WForqWY/DDok1nCzr3cm6ZsjmDFqWBA/ecG67WsVBlQMSSKPoJjrS8/b
//esggsaCYOHbfOf04vpJeAflL5xMNrMvCaKE4fTgZ6xv7eCOSceg2/YpcEAjNPDgJYREYkxDUFg
UgPZfidcLBVxrzJMXHd4J0M473QpVuxts5AcWgpctvZNKTmPOSXNrzr0Nmc5yeUYNWCaFg6DNkWL
5RbPEK5fFUmr2PWiL7tl5gkn6UnT1/CTFvpDCegF/0JFcQ1HBYsvOeS61aED9nq4Ege1sRoPt3HR
1GGJHmq9em0RgmWoyzDzGFZh4b+XMPpdXT5QuqWEizDQeBNS5WzpvwujaUoSUKn7Y0H+SHlHtW/A
eFrjgpolqV1oum6W3p/7+mLusDi32y5Ksr9jj0Q5hNqmyvDu/BqCBokVi/yfuSOs6VjMNew1p14a
io4WnDdCIYjdjNbtHrs+lYHtwJu2rLM0aLmNrh3OszYr/MyLl7igTq0om5EVJOSOEbGnRKQEaPQd
mAdVaBy8NEEqEbwZ4O01zlLM6KXa9nrWcCPGwmDDJhTHAB6Qzu4R389WP1/jXB6HF0snLukRnC0J
ij6IF5bjhWW1ZhdFEdarNVfjvF2kzSniZhyI7keoXeeNbWBNwZ+OX4n5/saViOFG/WIXAZeh4Xp1
N/O2ntXlA8AbFEWDMj+SZsZJHV67zOLm3KPpWdTL7+2zRdNjrGIWdt/r+xtskwKV+eQSOEz8Ncsr
8iwYlS/S4uthYsIon8+iPvDBsmCRGpev/rAP00NWCx/h+tVthriA4zgQ92axdTlSx+Sc9DLupxgO
5OqFWHGFBjTDkjtvaYJSmVlcT65b6iBOyDoP8YMGU4dzzHPxxFMGdEJzyD8KJrrhGfvyMETt6FoQ
RY8zWhFFF7fDCz35Oq5dm/pUsFb+oPWtrXDHw7skVYgh3irw9TlULUTpKzdIefd0nNsX2/tzJD49
v2LaTK+cs8H104K3TCJcC1txXoQXDJf8j0A0UqBBUKcU5VKqoJKW7q6popik7S2PLo+Ghgozv5hS
DtW2Bc9yqFtdc7AgqcbBHHYh3WPSEMeZcpK4ZBF56niZ/xa8amhz00b3XoOsUT5WlwTlj3AM0gBQ
S5rCVduxIHfbNhBY7aggEEhjQYAMcWEYolQN63TVWs9j9f4b/oyAiHDgMaYNIZNsV0SCXNpGjWnh
jNdsQ3mo6W8XiqCQM4CEhLBFWrLiuhjghjZFIhjUNlaQa6ZLTqsHcGjS6R2dBy1rqWLRfkSc9Hut
NSKwVELbyGr6agoAqT9OWbK5tP83aRUDkxQH+EK3StPo2WP2RLREQMr7guBi0//cFe6N//+Yq14o
Lbo+BsYgynfQXZfj/pKr+HpOBUrDZ6q8uUirxEnmAOkkz/NCRjiFxNLNmMC4iqIVgH+CbgO9rwd3
eTMG0Qy5X4PS5k5CDStlipAHrf5mf9TqgBR9Vxzi3lz/H/C4L3OWofxOQcQCikrn47ltoSRf1kVw
8H0Q91qaywBvrGi0pl0MKZYSuWwMFCyjAvS7ShxhUmpuzCtkiTngXP/vG8eT6EXx66uQw6oLZ+5D
jpiab9P4MYUxPHYe0M8Le7IKykC0eDp1x6BH4h+i7cXMXjJXlBfyN3dcAHjH/bCgW8AEL2GriN1S
PG6ND3D/h+s1wKeP57AfFBfUxbeCHH7uPgftqg+G+kskSfeOGgkNCnq04yK9gyWti4z5NY889fzk
J/vvyuIay4rF1efgS+7ACkMLr38KYNE3+ukw9oFezUqzJ1VbVhtASVtaHGhVQKrfEsFUPp4zMFeU
+NcDrTKOm8di7bsCgtFfgzOK1InyF62RW3isTA6bDfGECPC07A9X1327TEDM8rPK8Bs6Os/pw1cL
GZN6XqcLdtGEQOFW17LCqbjzY35q8jZppwjD75NovlqTkiwc2UxrYKeFdgwQYE7cFPFwLze0zilD
SQq62S73XQ8BFzHJXZwjVpLRMj7OqZIi8DhT8SvMGe/MEIA20aH4grVsUknCre9igl4fZ38Fmlvd
H6SItfnBFfRYzfvJCj+mp9fztxWn8qn4XUgW0/80X3y7/WwHkQOSq4HYkZfbxe363p8sH0xG0Vac
MkxuEo14HdFZZDXAmn51CWLfgKufjnC9Vd6botteChQ+dlbc+x+eRTxEJudvEgzCjp4X1TRvQaZ9
pJaFCZziO3oiy9lQ9fsh9MRocqt3Si27EzeXGQXKaUZ7x3i6J1vnYPiyv1Xt5MZ+tQVqxWVKT2PS
04HtaOUCkE7SfaQjslxVxtVHyGS3YxWrO7LeYC6uJEi+yT7AuFGqsANh6kbF8FH7l4Q9ypvmM+ui
EEEtHe3O3MVINe/WkBfDs2JzdkQyB8F1Tnl0DhPvQgd4dwF7hICTzin6nkcKWAceNhOA4LBJHtAZ
uJg9qU3mnHsf1DurqtgQiLQt/htrA9iYUtiCorCjHLm0EoVr6uyORb5bRrt32PJ7uyG7tbgyXTEq
Uq/V1zeMZCPEeui13mPbm21zzIRTR8/0FehVyUDS+po4y7ZGgZGW8tSDpnJ0NYjo1P2pt4MQXomK
UsZBJed8geld5RlWeSNKGw0SORJ5nIMYTbdvUZ5rBPROFHYAkQyEoVcq9AVWoJ9c8wy3tzCthdUX
PYJtnOSsVGDYSm5syJufV5qeI++2UspVXEmGtFD4isNn4ktZdaiudlAEmT4t6J1lw7geSxpF7ydi
9c1fpVxGMMC/wso0SmqLKOo6p6RrdS09TUx0e9Mw5dmH8k3rH/qmsF8/Ds5X3K1pnx+AH0d9iTTS
qaKjWQ6ueIK3vg0sjmZK8lFs8Bw2rsi1F6bCqxkDfEJ89kwMFkg+9BG4oVl152u60ufT0eJxSlM1
WG/Wwr8sGB3HWS8llzQCHbwKbpM8U5g6wCSbAp+kUy8FP5JAFMtH0fGNc9PW79IcnLs99YzUFCex
3UjyG96U8QatCw+kbJwH2O7KXyYGCFGFlfPND7W5PGlQffV2jaSRd76N1Q/FsgREv4tERVYzfSX8
GpLXr5JoPpDKoIYoCI8uNhCjGvmWG3iId2lwS5Geac6omgzPZ2G7t4DvUFqhhCdw9elOHT85haBJ
c+RyhWQBPoOIMUnaAoZ4vmTxLfbKFfCcPpgVVGK4msSHIJlynH49UjfZcABkUnWYsXclqjj+x8Fx
z12MHz1wLHwI3dKUSVDTHXur6hz920HL+J2f9m/83laMCJs7hR4iMHB6lbZVg+DL6+IhZCGo9hNe
GAUH0pZHj0KOk6qWyXYEVKjWxVOULcIpAFY8jc/MVePCR9P7pPCU+zorkGI/JVzlb5K8e93vEYWE
Dokmum4yLqnGuSPulW55gUCAFNEbY1NzaihFsyBPn8m4i/qA+TjNGFTxVOCFQFn8spt/xjKwLaG1
phWQQIyq61oFz8SWuXMwjKrPJBzgeG4It0dMpy/RMPHLWPiZD9ybutRTwWpVUKF9quBIGh5juhlo
Mbl1q/766fbOpiAoIq8eZfSoeuoTQn8YsRk6aUiaLaZIqrt6Hvssj/bJxKqh3pqYl/sFGawo83tv
jLMBNKzRBZR8MbU+W50aE0T3EB/qX3dP7WEfu6HwkndqPnephT841Jx5DfcQbZn15xuf8SW5ObRU
efoCEoDuHk3PHyOk+1acZfjvvCr6ciARMpcxJpxAWJiA0+r1V/dHxNT4jpAXLwLlVSEHRL2kdfIE
WR4YQirS6Xl984XTSs6kI1aj6q38/ejFcd2gwzODiNQu32erjqCgyK8yt5K0VMKhJympqYmY+Ijs
aT/A3smqWEM6zEqbdheea7Q7uxXvfLKi9REKawDu6rPkYtUXGveREXmXqcgCLQojLA/ggAwLeJxT
JLCoA+CF8l5v+9y7ReKlPyKRDf8MqFXEPmF6MypZKV+U02AD+GQAoxs5M/KlwXpR9Av77Jp4lLAk
KWe0/R4Ww3KccZ3/5b/LvqfEfef9toiH1RwC8X0xL1twIaGBZiMoweF3jSuf7qQu8vjpAIt1clDh
w7ub6fo61zlxVqD+66KOrFbTsxYm8050Ldc/S2UmuFYx+MF4Jt8RslL/7xYwvzQpWkPQgpwxV2Jm
5vPMPragB1N+YB0FguJZbKjgmD8IpNWuO6WuzU7PKuaQ8hvMZ808xcY9REaVUwX2uFJ8HyL2tnDT
3/sIIWjUYiXnAXT33kRdG0+qOiJgBTExr0VcrJ5Ehm4VrWJ4eXw8w8JyrpR08EVzOOu5xPMWXlzM
zAyC0vLBa2+r/K9Do2pwIBEwAe57J2QYGM243UaH6jYiC7hacTufbltI3dh5A+3Nun53ujmMTQ6v
sOcSayMwG0CH5RPLZWhH9l0VTMnIAMFCjvyiBKRH6q1zIylJ7Zr0dSmENmiLTC67BxRCprpnvmcF
5MRuL1SL5Tt+2onRRcQfYvVcrKGlXT7LCORbaDr+eey/tuvK2zFZlccvSpWqNyX73GDCMQjGQOzR
eM0EP7hGvaCYnW4GNSHSvscDmolyWfe3oMqqKzGcOB5rePoFSlODAMerNUKhsaoiptJq/CHFLPyf
KWlmojG/PMOhDuIPlrruMPKNLOB3klY95jbiUTLLJYp4u7aviY8q67sCkfB77yddHWn1VYDjTvB3
I3/Bl0rfe86EsxT+yNLcqrR8Hh3PIYQ+a9BsPIYkyGkbqzxzpXRBzc3ib5X9NM4NjvJ+AJUM7nbw
pUvEwdV0lzE4MYPI93m+Jip4lReeix+sRI6nHybFtwKz4A5tM8TReTIHcIs6byzA0t0pEqFJuZI+
ahBuoZlsJNlY9UfFxjwjw0OAcz9IbBtHed9Sq2lO+hrj+tsuW+JBRpbUIkW2+wJNae9b+wfR0CPN
ECudjEni+bMHZLZP9LRCj9PYQxTcwabm/CDVQyxrxTOCkLfif0c/iTAdSoGBBgfcl4lPTij6IC/z
9gp4GaIu9bq+fHeDifN9GbKi9nd+RZ1VxD5f0d0td6noJrX24ssMkspryNGu+yDeYu26bKWALJh/
vO4EuYARlqMAlY2EDU+/Gkt7J0sMNh48tufE+2zAynWbHPGXgMSIzxI/ENUJu6C2t4+81lkJYwG2
Y9i+INwH5bTxWZi1D6gAUNOJtAe3TsND/7WnPsyp/OyWYC/QmNPK5j+G6WhkWZDrQ0HUFAM1RLsc
hhRWOr/RanUpifQ2oH+xwif1XGRkIYEdePGOHeuIRjAfdqp/3vP+WWM8qGFsFkPUU6NkVyLPj1oA
Q6zcImEXHsr+OUDO1/fEMh46v3mgbMcLRsaFu07RKVQDYieUW/PPkpqheHKzcfjLWfDX/ZiK5zlc
9a9Ga6Ecu2iUxcXjtoMb3HrntzPvXnTs/7KR+6pgb4vQtYUILOnnNxnJvLy7MyMrRjN2VENk9uT/
Yls+8CFxlrhqHFiy7y6GuGcaxcfGrQ/Ws7OImhdGN6iwdF8brAlxOoGqXeZsFHz0NGbc1170IDRs
5t94DI4fP597W8yGp6+mLZw01ASbGV22JDsfPuHhUTu4iJu3uSvhVr3ySsERQBQGP07dCKS93qEv
KGxpX9vQB5uNbN15iARDFn91G5zv9RQQcIkd7gBCX8vury7vOyB+SMTu2aSKULp7Otrmkt7MiaoH
YnGNi98RhJ4caIR1o2iGptRdaLGuWmHryewDVFxHpDycOwWmqjZmlBvcEjrVXTQ1J5xU3DaLgVZa
QVna3kYZqlApojTAYhsIradGrAgePIH8h9AMnImnAeTsz5u0qHiAgX6xiSwc3MgEgyR8EDIMze2q
9lNf1afIHAemoKpzu6Fs4BNJidavgYHQ1sAIiRTWWMnD4rbIHwDkqOdTi8XfSifqNnW83tFDgY8y
KiqA6hQF/05T7rvlknX6P3Va0+cNI5tNS+LGtMypCGUUMakoknv8kc/dJtXs2fzZ1Gy/NWZgJTJ4
8VUhGsSn0C+UG199tKIJ/5u9C17aiHuc0s+/3A87UKeudHp1XjKeVvNNMNJiqla6Yzv+27LUsxdd
SxXhksDo/DB3HxeVCULjZldWhcNqxGZq00LYcDnXjsf9MnUzY7IWftYTnf+BV5fGrwVf5snBauIF
H6GmXjwqBqCbYeMKxkO7wCRVT1+USvTd+LkjjM1EF8ERuFDE8fIQRbGtjDK04XfpPJIax4UOe2pX
c1wo7CRdBDvXK0wvioL6AfpLLx0NCVebdO8sE7xO/xBKtLbUNoaiWsHz/RjHBOaRdn8KiPXzJUBX
G6mN6mas6Ojwj7II3YrxxRufDTZ1LIhXFO05R1Q8uPbXtTjv3ko+yfxVjKlTOr5nubYeVWy3te/X
UkPBAQR3GZgK2YHHVVF9byNZVyJJGDSohKtieeJLRMy0dtUsnaemuc7es2XqyIpeEDIGBZix1oFw
B6n8JPoXDiESoHXbAgYoZCwwp8SKrEAijY//IvLp4Nlg8esXuMTBlK1F1CIqilxrKNDj1zSwPJ4c
lyONxWwnI8sVf3Yj8nYUzjni7WYjmZL+NcDqfEE3wfprkS50eRRhc9dZ+KrJs2TerX8xszRvSuQC
WHcznT/ybRRjUuBV79WUfzpbLEO6MgpIivIUlbI/Z4RafFnKdFQ/GNWNxTJ5wO32zslvo8gEb4TF
BV5c/GreO6rt8JKgdADxPZ9hgnppNRlJ4FGWn3m+1/Br5Lter6f4Rq4Lu+jxpOKgwwTpEgaTrZ5G
riKT/7ZI07NqVz0xtAkmVW4sdiD/XAP0NuBNiBIV+/JAvz+XE9dhhFTg8A+wEiVx2WdPgqKn96e9
IwGLyY2UrB9lVSiJ7wuk7sdiLpGVYlsv/zP/kayPKegjDopbWiH8zIyihkg2iZgygPXmuogvGxW4
qHrhDimFv9eYElgwC1NW0P8tNG62kXYTNwCkrwSijk6mueYorXg/nADOnYE5wZ/2BDHY+JYvX2nw
jDB/3+dNExv+jqjwSw4tIgB3wjUxtWmsfJwCgdZOVsq8uNz6ZIOW8VASsBu1Dohjm1m+yo8cUfae
9BfL9SjGwKK+xXxplwPXbYpU2x0UdYKtV6q2kURGcZBCuWm8ugraKl2P2cjNQt3zhASCpBq6zP9m
pStrU/6QJ6m0lB6cm9k2sPHCko5HWgFuqRp7FGyAQmPT5Rf14jwCylRBF+6mgEL1Va6H01VMdkKC
VE+qCioE8XuWFeW2htGSU7aTSjqzLPJ0tPl7YqhpUd2oDtxjG3tJ5TNWV3wmgmzpnKzu9FyYJfeU
mk6irPXYLpEraf1T8q/nMD7TGSykyl2RBXsHosw3QKEW3YIq09njPTypHehZqzptP+bvjkqf/O8i
qAeJg8ij3KHabycob4XtwUwmj8sl+3iqNhJFV87MWUA8QPbZYpVUMdez1hRzGw+X2OtZafewtCc6
GesN/Q9TICB/rBrCO4GS3SpChilffUWBNxHrsZ8I6CT8GzI/XVKaUHRfzcdFORyVqhbaW3m6wBG3
pRVjojaf4NtuJ+3lm/Zw4LnkqudIeP7H/CGerHWjF0y7rg2toNfatIZkS2sG4o0SFe1jlB7sGTb/
W56X+GwWTtk/BMfw11roE4BXgNAXPHClebzmBliWDDJrda614BDJC9BMfMnbHWK2OX+hYWCSp2Tq
g9LMY6GR1FnVD00++fgKjvNQCuJkU3VUY6ArpR0/xtlMiWZq83nYtH2ODty9k37t52h6l/0bYo8w
mxgigDUGwtFgs3k1P0v2tOoxKOlXfFaTgAyEYAnfw8+HL83fnBctG4busdpq3RldxDlm4r1W3uYZ
eHhvmVTwv6yR0Ev0dKkhKSl1tAngOIR8z3LcXGtVCmlOb8x5S9lGX+ofMx/kbzwbZjPp0yiaFLvX
NaLpd2qjUA6bC6RkhToojwLUkHPEQpX9nhtsCWt/KCRvsf1aeawkJxN0k/aIW9UQ3gQU5W5w9JAi
9BB4ebXgQCiJTgSfNgL7Mg08mOTHrChkx5xu9W08NI7GEr1CuMJokZvQuo4wy1V+3R7Iv0fmBoga
I6+hwKQ1gyEUdyo2oE3lvmTLzvEINYL3RgHUbnpFVk1zyk5AxVCxJu6kAD2m7MVmAQbumEy0XcjI
ILoezyCTo6LeAWsf0TeeLKlQw4+BvQ+ue1epadYw587wB7fMWQEu414ZVb68Y0IlG2i/BH+cpjv4
2tlh1RXtJMUVLhFUWbSl0LIrYSuR14XofrGj/d4/AaQ36aEoQtApSSjATdrX+j78yTe6LX9jPwTw
xZp31jbrVVM2oBMtd8GCf9+HhdERcSEk9REPMAEcsLOdCPiMywtRh0fHBg7ctsTrcFL782l9us6f
dh4DeKXZNMAVwNY5WO9utqvQTddsT3lslYoIbdESCAU8mXINQgni/ujoe2C0OPD+Q+X7mN2ysw6m
B53/tegnnedx75OU9ZS8019i6RoDdzCtogvn2KCOsdq7ijL6xCDwKYd5uX8CtN7J6vt+Y41rUU1p
Bt1zisR88SBxVcy1/BT3f9Ix2bC3Jcm5qI3U6H6AR9rBIK1O/3RolNKKv/iR8ZDsTH1IJYJCeDUQ
0rmuDDJVvZX4BrjSDp1RvwuKT6ogBMwoSRQdeSfKGwS7yL+E8E6VFdpdtxGIu3WVAR/hThvrvpO4
DpFFVjg0AbM/xo7RATRcvHuhENYQNBQTIiyqMEHdq5RlOuzWcwCXnbdwU6tRrWU1j8v/DSqyuNVh
qkncd24/rouBW3ltEP78I8d1kKLpNJ5W1FhapjLrGAbRG5tj6lUJjZEAN6i3ZXavZgvhuXd+dflm
Z3hB1bfiNPToZDr7dcrySDEeK65bxJ5EFCGvPFPHwxLxDtTj4F6Hqr1/g1g6QDpcYeCAABo6f6tb
qMvSoLCrtoYusYSZwp/6hMpgwdBbrVC4f4XQ/UKoMFCzRUDkHeRvcMZUx5gD1EDb34oluc8Gm6zi
CG58lgOIdSyaBb1KD2FygJBPGyIT5C2nHVtUOfma04+kVJJ8igmYIY0PMwbJL6IDDBhrkqJMdN0D
naXRvTVbjibjnK4AYd9RoK01acgc2/CU0G601Tz6WNAWq4p9XXjlroPcl29vDTd9cxM4NBuv0uz0
g0SjqFdRA+VPrwgnAxQu6lFfeF3/j7vTJqPEruwXPPmFRXS93P3QGIuAVhcmskdaW7O+2sVfgGSj
DxJIEUSPA1B4cd67FJIY1IiqCXOMShubVxJtqXbDmVYyphD0oAMAZvV7mFoGZry2wWLNYCgsVqHt
/5DbzxQG5Alu0DrbiJb8OSkw6bNujqZK8+ldQrgRnZQyDFS6l7HzDvElbr/u/JvSZ9OxwBNfrI+3
5GATNj8OjXdL/bVJAi+g+xmX+8BZhtvP03x2gsio+dXcvgLojRclU+UTTt/8HnHXYXC0b6BDY0Eh
V7JGr3HrAdK0cnRAjGquz2QscAg5+gqc0oBjDJNUu9VgKc1IvFKNvgotHWrH48OULPf09TRyHzp0
oRmkEK6UQc+scb41hbAoD7MYYMDZ+UOxmOp84Jxqc8aPn4unUjzhf9cgSH8NBegdWFZ9nZFfkmuq
/BwxuzoHOUH58fh/rlLYv2UG316Pjxfp3tK7Ww+MpRhupA4WBUs2PTqbQYYh77pR0Zo87GVmjQBu
sbT2OQxlIntcZ3joexbFu+SUDK8L9+KcRPXMyBHn3tSTYcAAGYRvyUi9pypDFO9YaYm7zE5XLoeD
d5SvT9MJP+UvThyG665yFlTlR9Vq+Eo/juBXr6SPxn6RnABafiquWI7xzvRbQwhrUFGHYygI3K7T
wTOeDXLGScJ6ir13rox6Ne1D1NmnQ/GiLJ3PI7cHYZ8YQ+tqlIAlnpIuZ1X7jB3uLm1GvcmjUFPr
XLyc+W1eWeHbdBiwnyQ5LQxB9KJa9ykIPj5qjr+bKqPt+eKvXpeJJn4oJ9OrjDopB2l1ip+zEUms
jRvu0859PcyJ19x+e6dCvUmdJpP/W82sRUGipqVCLMho/bPmoyZOxBD1ngdJQislEP38srfbA39f
9M/cOMxuPzDb6FZCD8J51oA8R1g3qyk9ZcalKTq2p9962nd6Yq3jpP/GvI8CQm0YAMbo7Lnoa/Yu
MGohYWLLEwnBLFDcwAhvREuqzLDSO1DYkEtcxXuItKhYER2onHc1O15BXMIEbIyzTB7puOrW6jrp
4yCvQOvnrBz9mWYX6mmz4ZHbRiqxO8Z1+DPJ0bCZvc3NjUVOdC+G9MI4OQw1k7puTLHZXpuPDEUx
TC9tDS2ilH6PZZFZaFNcmdYsHGlEUN9kb1X397mSoOsPev/pYusJYzaPHlwAJMHld1YPbp3fhVWf
W2D2weAD/sP+zxHNPhtgUCv46H6RYsFBSvXPsJ6OQRlEbebGS0rozkLCT9rm1CgaC3CuV0jgYp0P
SJq9GXotCONqADl4eznD7E3hveQoQruq/Gj1Ewp6yYpvibQc/lvtS9mpM6sI+HtbidNQS9OSuaJe
cVG9kT3kJAQ2D3+E/gf7Ry1nzTJqBFC1lUxD0Ro854J/hIEFt6PUutCCpNtl6ahNfjTFRDx4pQ0l
DNjs0K8zKrSrbCKGhEOBpQRMIjVw+ijzFO21zlJzEg5f7QvO0YrIRxvqGmVt3+1ENi+12/Ew4cDU
+dPCacmAyg3Qiwqtg42h0K79YQ8x0YwnsJCWHkWCPnOlDsmw7QqEax/wWVu0eqGbbtmMQLjkHmA3
43SUltdeOKP6x2CXyOS4Z5+2h1XyL86lKrG7AqqYV3WpuUgtCcljmjhZqjSLPSKjAyi0RJTUgSZa
tJA7E6UUMt9xaeRT1eh0AiRFyikXJYfdXGS/Ot2ReRF5ICbdQF9sDYio+phU75z4C4yfaPMhdXNe
s4ArCXBY7mdPGkfVDDy5h50+w5EEjzJ/sLJ6aGa1/wunc5QT7G45RYjg+u1tT7SralOouJRET/KR
uTfqrORVFfnhPouUatNWytQgaiTK23DnuneY4wY50Jg97dKcRRuwvYwPB4ETKDWHnvIKAnNUcAQs
GSWZ2EH++s6HqpsS4B6dGOBym4x/S7mW41vERbYF7PpcPKFEyVRkRjkbvK4tud/CYNOn/PKHhCY8
9lkzMLmvdQt4feo/WZZKoj4eDGYlZoa+skqNJuhghHhUNmGY6+qsaJ8aS+O5Alf+fzAHY3ZkYIOO
oUriENInu7cTLq5PEzCE4GOqR2uP99Pwl1X5y2JZeAv8XBntME1WGaciS6SUlYe275as5t+WprY9
SACrDSdMfIeIlofpo83IqWLn9/bzjuxOkGdVpgHZnW7KlzclezF8+Vk9e+gF8kMHdBveCby9XFTq
5fAe0VlBGi72xqFBj3ZjBUsyzZRIvO43MeKNqXpYdsoMeL880ziBY4eox2TVTAJoy77vrfyBAKzV
1NWr2mm52YT2VwwXm11MnopHjt6aKECEMdpoEJ/XtlX/MAmP9cLRj6MkzwJlV98Asb34/TtCHZ1n
3FsTXD7UqzGQ+HWSgbmiyU+ErY79ZleeCANZCcR/xfgSX97HuPvGMeLxUBb1NKIbSCF/tslEIh9Q
9OVvEbxPA2Cl0VAaj2cuPHBPRBuVz7qxJYe5Kq3pDZaDmBkLu+B+7NX+pxqtnfoqSc0KK841WZ54
Qg4gAe6nYlz84NA+d9TDVSpbnmMwQf3e23U/lucsAyhKMz0AbQfwkla6DfdmDVoPU4G5RUZrVAqK
mh09ptFt7e2jPd+rjq0ZkSWLydTo8qDiC/t/RtKIUOxn/gRFEi9Bpjvh4F66qQVdacOoe2BHEn2Y
5SuSPU4sKSsu3tYHCCtC7XGUYnNEjnruQhPefKlIuc7fpXd0Nd/XrJgiVoZTKs92b/mIpGhNV/Q1
Mlgb715K4+im06Cp0VabmPBX8Gq264SekO+nlpOBcjs6XGYRFj/PgnWb1m3VhOxgCfuzkpK5hUdV
oBkcq7D0iPy+lbadrLo17RvUXhStC+2JOCJQxzDXEFQyEuc7+lb72kVgUbeOXOQFgbNue64uz8gB
+D+WBqWmy98lPLwuQqBAdkk095IOr7KAXctNh1F7KlVxWZWknl3vLlhumHuQObITNdDoB7xtyT7i
OouhVsMLgN6jPFbn5js0AS4PmAO5zBCdcdcyICZZy8x1pnOvPhvOtbCneHRmcv+BVZKKhUq0vbyN
dRm3YIqDeF+bMBJ9val96wL0leqJ9240qgJenPAMtiKCQeFV4BfozikvFo1jjKP/nqe0JRQzUDf6
qItE0q5D91i+Lj2hh4mjWlDcX7Gfyb6vl8ze7xpBiZLjzqliZicPCMIN+okUVFPoXVyKDIYdMuPs
92BPdGL5qUrSDa2CFVyHjPW33AzePRu5SYJlgAc4WlQH1pzFbtxqOeIRMcrs8q/jXMn1i4d3pUrP
fEVz4kzVp2eMzDKncVoi1EAmwyrWk1MrnKm3ZkMlTB9xkjrKULeIH+vcymOgNb49YQiyy/bAUpvY
md/nDCT41sOLrAhbITGemSCskiDo34F2nhVJQlzRJBrNya4RwwjAP84p5xYF9V558l9aOYk35pkT
8/KggN7jonqZ/Lwz51kBCtGlyfdl8N+FlWJP536eUF/ZLpiLv8BwCJ+jk32fjYoQ61qyzljyNEZ+
CFENs4N9uqrTM3eoO++XWTH+WVuPH7WKvFoIX2tU9qa2dUMYSLgYGE+WOEFicbWmhsuGv3MkT2oI
WN+kgtz82M2tJQYT93lAnLmY/rGMJulPYHX6iJtz6kNNb5fA2mh1VP6TGqs/AvwLemkprNMeDLxP
zel6BFZqrYAXS4c+RL9x5RBcW0WwzuDtHlLjRMV1uGCtIHCScTFx0uyVvazGWAIwptYvjxy8+jsV
HEnrQOm5GRcileClE1ye4R0+qahmmrrvreTq3c3UG7VnRQXPYUmEvVrtlXjszgMT6v1TD5j3G7Cw
n15v47pm5HzmgtPbdShsl5Oev/1Z0RzoJOCqDXhIg4R4LEFUlnx7PlRFIuHBg9Bj5OX4cOB7wfB8
kBzxQCtyu1ZiXF4KZGqz2cSkQcBNC8dSN0fxGlEL/D73Xj75R4PLrmH5522LDmhAvez7c3pSaQqK
0bEPx6+lk8NLbOGRa/aPYCJeYQhDZfjolQpNC2oSaacIRKQbdwgfViutYDKnCOAppmSzvcfEtiPU
1okutUNQkHKCR2u9jXhTdrIB78mZ+aPkh5Bx53wMruo4ZoAEd5XWglov+KGw/HoGiRvHP/r49SdU
sk6wTikMZ87fYqLnA4G0fQSDmLe7M114ya32mE5li7ltN+oJ5Eoq8v7OFEsz8j3xj92CAlZGTt0Y
3tD2RipDJUPTOqCcnUtkHLcFSI/SKyWWx5cPOhN3j16+Q6Hm053zPMSCw6SdowKFWEySRCd+bUBv
NyKMGrrCvUNJwuz0s42jR+8Rq+L13eOhFKUm7LF3l00WJtiMLA/dObWmaGx8eyPfAdRpKykNW1bd
7EpHbEMn2ULXsX56e8vqCapS5hVdb6hOjT5bz0qSAA1fYNEUOkYPdMiQw3yxS9WoFXhE/cfw6tEr
kUjn4db9Ik8IbywF961m6U2Hv4jHgMSaFUe12ayR6FP9npmqcWu+H95MQfL+00en27tQM+k4MBtk
T6l3P5LIyQOp15uVKANnCWAi4PHms/Ml1yxoWGkh9OVDhfjpdTWqfYnvO68myLbbs3JBVrf/dhke
E7Z9E1ePbz1EKB194invw2Y/t8bSCLfZWkpxndplc9x9MxbGOSaE+LN6izkLbJ+VG1mOH3gzRSXn
3mAmymQMVD49qF/qdKIc7tsE50mtosfWKrPbNVcfQGd/XnK63sPJeneNJd1jg5sbQ5hgIkNTfyhl
m5ITdd0kVrnfYHt76TTsbel9WPQWCkF7ZBlWtK3QBOmp8ETbYcpjVJbwDdM2+h4IrqrIIunc5gVQ
s62fXlgydFtop/kLYRnvONm60A050/YPXhV8VcpxM1KRmyMxMpXWqWn3lorNWwzBo/FWYNLaIJ0E
hAjEA5EzB3U0BCv42u9rf2VLHOfqglQq0pr3HZP882ypv1cuysHXSI3lSXDpG8Bx9GP0tZZd6WtL
UdqWQ7ASA/tCFw/9bT38HlRsGgOI4lCZG+2H6si2HlSdlRbF5nbHlCgeA0QQvieHdRpcWdmqFMa8
v59mWIXyUOZ2ZiHOjAwClOXgx0+PyZXlSsxtXBTWh9ExvYLWyPPtQNZu8FIxAGkimL45SPSLYKVe
BJi7+SmYr+RwRjzB6AXou/+z7qgedHY3Aq6J2SONZtAWrsZB07fg/lB80SJFlSdbvbEmR9/qGbuX
SLdh25SviZlyJlj3q18aVMl3YuSwk/AMiH34QgLV6UDYZ3Q5hUJ9d+OuGw8s621qaUw3zWVXJSIM
U8we7Dz0OC9d8m28DwK36nFYymL+ipEPbFAOHlYzlEtrURd+f51H0rAuGZ0COXmwnUCYeT6N51ce
l8+/PRbP1zIT/mF6f4XDCBUjLDP7l/Q9tTJQLn9iA6cDqdIr0wAfxnEgb8csyYvq1tHi1DCpRlwb
e7Ok+ZkWXQ/d0jMn4wyQQsJN9SDgpW5yXoGz63b6PtTa3W/to7+LhXkV3dAmycJTZGDyGrI754MW
LZosAv+JkRkvEd4h+PYPpGIMyn6ByhtN5W/pS2AWEjzNeYGfYf1eOoqjMDLQ7cfZr7TSAbf7Gnu+
zlr0+NGVzdc0ynhJcl8pv8vCvG25B0kdYoAAsZbMTTx0GKsW35A73xXrqKph4zdjNT6BTTmP7hue
Rc+q9H4/V/mYirTesAvXO1JtmeQI5AzlxOPMRfNzVh7jET5n/1p35j8d7twVn5v6QgUH14ifP+Y0
CM8gGbNM27w6Ew9KgYav4uQeDBr1T65Uog/M/Bwu/fP3tSJGpijZuRenO8RYXrKP0e5cFELke5Bn
8sf2gevoxHvxL2XZezFgG6kL40+XVjRaWKsJ4uIlEydg4s5rqkYFAxqgPNUl5yZhySMhF04VgJW5
5TrVW7Q6/lr585JGTDa1wMw0nWQlUf0OoqWBIUNkVrPKG42pLrLPmLzgCjWKV1fB8Vc7dl8Z4Qa1
+1Z46e1ssl/Mz/cuHt0/mWnGnl2ordlK28ysN/aA+TDmDL5F1r7A5DCLvUa9pOkiDMwkt9qENQWH
Z3FNqXgc2p5CknSnI8I0SQvhWhs0lARaBarju26mKxTsx+1+/TDiJGUUQqXHMRakMYvJR3dcatGp
U7nX2Tt+w644hTJaJQKxVCmj4S6F8BCwaJD4eABIurA1WXn20suRkQHumnmKnjVYifec1taj7XyE
+7sWmBUYwB3pgRzExDI6v/pV8YlhU2icu3zh/MkCUPqsAKR1LWS7vvS94dRyG0S7bSsWhvyGzI/G
8Y3B5HwaCva1Ep90yrDUz+LhJ3PNQkfg7OHipxxumeEomPoBTzOtzQm14S0GPHhbY+bly/w3WQhW
4Mgx89gzWAAsOSGjyJ6LGNsiKuakGybGjhr3cPEUxGGjj6SyHk98sp61LM0JJMf75qGJcSz2q2Tn
+48jpvqp3LlZwshMRxp6fZYXbAQKWABqnXKVRqQpYAoU4Do6SWjBtXg4jqcWp+Vfg0+dfrsO4fXU
0gIJQVZlnoFQRmCFg9lVdXKmLyyO9J2dR8Prp/GOqlemnj3Of9LbJzr8e0ngd4Qm0smxiTZjfTjC
IGm6jy2AFs8RDunR6ZyueoDDFumMC22IvL4FknPi1qPG6NdJCC82/3u5uNAT05VMHyz7libSDx0D
IcVFOAeoFDzOmooo+kNUc/p+f8Bp5vCC0MfaWVFIC1xgrQr2Es/sWKThfNrnoIkQy1p51nhrHORj
1eB3+Pgk9A58nmlt5rddaiTLenlo5usw5eH7InN/7ncDgaADnB9z+9VIJtU/4BF90SSlVJOgrZTN
NYSJMQhJNHe8FQlsJgRXg7wVoEHU4g0Fj9ghsKGK1xbKYGDGjO2ldiCV7B1C5Qvjm/8Ty+VqbDQc
lxvWpZ9WRUftk5fcvvpajLZDaVGEq8321KpKVEt/Ua5IiIYMnHd9T0ny+Pi5M3b+PkgNr01FaX6F
8HBXCVo8aVk6K+j5xT9hl/UtNrodRqMQJs6sHzb8meP97VNqouTPqoyqsLHq2UGdmC22zjDWihuv
qtc31AM15zVurIkEUIPeoxLMmGyCetrLbZ5dxTz0DYUACiXl/z2aEOKU/NdmKGCd6k78U76HwnRa
6g6JZxiQVluv+aoDPflnC5guRAiMEBLTG20Mj9aqiONOnWMjgMTijDnfoWUVvrJWWK6q72u4HPV4
fG0WTJGpiLdUoaGT3wSZC5ISAr8OJZfQMG71mM5ZFsdqCP7UCKE5YkCQrHknsmO2+AQClKI8Oprv
Cfz58XuFnxYLPqRO+6fHXVjN2eTYEwQscXfUj+APcU8CWVo7GSO+gtNZ89CY29yYt6TdiWsXUcFB
UR5KdgmHS17dwACsKtA83tdoxlZcIWHUFQBHyPKyOlvuTaCDeLa1LEbOX3EGe3dfknfIczX63vVj
dDYk4PAzXRc18AbseS1X3RVcyiW5JlDICiOL91KbmLoV8iYEW1gBDOxQCnrqQnEhQRFMAk6a+Mk1
vGJYw+1ukrkucc/U0O3S9Bi+oZDepHBhO8Kysi8ioXVs2GmCfULcMmKwKxIjcXlxCjDWMpp7/ebp
RPY+zDob4w+7WPLTvr5qM08sCP34BSCwVRIJ1ph0fB8s8/UP42Le1xgP5RcbmvTSUBFKTXum1FOI
6iCA2md8mJPt9Q2zpFwq6wNYfHZtP4RN1r56arpsR7HpSFRfMvL8oAnsBcxjuAZpIiT11/oV3+UW
sISiFHV6Zm0xwCWOS37pFQHl3Yqc+zNoKwQNJx7Y8qoBFow7AwM2KWMKWbcPTJDN9iBSBXh3fWLN
YCJ7rxISRcf9T/Z8/Z9uSaUqXIiInagpNzdtbsYGe71mqJfgL8aCIs3BDyJf9+zMypTy7hOduKo8
b6dWS9OlnBKdhpDbkVwcIKLTASfmR3q+FHfeC1tdpUql9BuGEH8nrozgseW1g/M6fqV1bxHBXwWd
cFFSO72NZD2V4jqd00UOAQsgjYP12f/ICLBjgCFm3fv5kE02dVzvRP5xcwqWnwmlJ3Df8UPKBAil
WX8iWRYE/enI3vUDwVgGwcVTnFujV04WbUHbJOCrO9DfEl9KTmLILMvFDhjtJWEa4Y27RKKipK9D
V8qD93ap671VEv9iagnp3ql5QMFy5S8ESd1es/MKNf53sImSgHRzFEr4QG97WymnF1Whj/pRFy9m
2vsQAAxTAXLSInnRJNH6jQbTDPYjemPS4dprzwkTQmnJb/qrIRU/Uw0XdoNcAXioZv6Of/P1rSBn
62yw3evNhXvZwi+spi1bKzB2ngD9gBzip2HrSV4Ed4Y6MBnURHysElH9TAxPUWMiKe//7LF8nWol
62o8s9Q5/rp8BtTm2o63PEjloINUpk3uR4IPp7U5M227jVGcEwcHRa/CWLpahVxKRqPQrentbgWn
vjfFWJz7V3OYScs16/bXTDivqG+vMySk1msRoC3pKQaY71uTH0VTM9SNyvJphhlpJTYrqx1xNXuk
9kR1mGXB42CM+lpcQjjxghTbxRfEvvlFYQDE5wzxv4CumFRa791oITMUF5k6aLgdqAKZxaunkQ4n
8TPO0z6zq8UMOY2t0VvbYRD3DfM98/4qPuqvcYIAI7xx1GSNpMcnGZDVtSBWMDQEzgUunBKdm5v6
RVM4Tx3HdWfJQEITTq5zGck9DWEt4jQEwQZpRhUU56chfB34BzHICHBniJGNQQFuxfQo+l7ChfpL
Ux860EhKE8EdGCCZbP57GpdjpOAH3gQgkn2KOUbYEmGz5XSxEj9nXF7OJyOvBzSuYZByZS0PKrzu
IF58gRE9+H1Rz9tgOXQl3KQrM/PUYZ5gs6MYYvtUJyVPu4PoLYh1eNnlBhbIvGcObZXaKXUUtHgX
pjJkX5rtDep6vgAN7k2+iO7edILl7e2z9L4X/0XWBZOyCC3kCYbKLOfykPa+kPJCZRsioL57O4KO
wrJcolR3UmBd6O0mYNMPKT3YsRB1rD+8AXC6WFh6loG+8Wx4fP97CweQJbHJo/sExwq1fjpi0CgG
BoOkdmklUiO+8PlFtQl18TKeEfgyD6zg48TVA3WFLebnBsyJNZKS+PP/aHnb6vaFGbGYOtDibn6O
J8eTxmk2MImWyamV78fZ70DR+35ZA8Yo4P+pHgNKny7q5avCv5juNfUhCS2jnD7m3dns2RXbra94
y2pbFdF4CWn54KNgJsAsoX2sTL7kB6f3ljYF+z+Ozq5kGXFbI5YQ0eXyOv4xvSguOK18aNGmBVz0
H73G/rgRbj5JrODmYlul5Y3i8kCvVOfPkG4JhrnlYGasoWF0VITELUkItjykddO6NbOY/RxY7RMu
QbBh0F8X/O8gb4dJedddrWDPYjc8HkqF2efL9toRwblp5yCcAlSTPM+q0swL0tGFNEBX6HwBXLsa
He9SkmRQeulAPQWHUJXN3sjCK2TLMNVgkUk3HsLl7V7yd5K5y3VkmaLqZUSp1FjfMjjUVvs2zJRf
4H4yOl2c84roLgPrfsWgKZL7AHCfvuwRkVSzYk1/jdSIgP+TDRxtRVU+zYIFTUHpDGyCoI4lZ0PL
pQ6kBsciq9jozPUL2L3Wt/WguMmSbLqr1YPt2cNaCU5p024UXR5Io6Rlitk1GeBO8U6PHItW9cYc
Gjx/XT7xwdrfWA+Dnuhb/htzjlVba1MrdwdmsqWGZLxx2bsiEnr9zjjd3gCz5zZGA60oOWBGJp4x
R7Fviz/BZwOh7Ojw2/G87U2enQU/S7YjOyDnSLkY7psB63E9WCkyIOigvI6Gfb0oYTanEtmdX1LQ
K2eHSbUi7n3trENYhLfE4bjcf1NWL3bnasKnnp2Pb0JxcHL3kTFQl+TN4hFYn2ZSyj8r64Ogfs8+
Y8KW9nyi2FD1bKa6HFuDB5a3Pn0cJNj88Hk4ZTSi6fVqxE3B84ejohVrVE6s0bZu+srZXNSXCHBi
k0R7AsZdeLfbIDokWxqtRcgBsBUw2J5lO9reEauHCWIH4Of5OiHDiF0nudyba1Edztto01LGqofR
Ocgt6Ozu5bZVjAusqwz/7XIHpkR7LgksFdmsXa1sIKh1poXBFJvuRGaytLLgfvsdjQ692wyFOIZu
1WbAPAB/QlueAVSFGaoySfj3qQ/NXKY0mWnK1k3UmlCnmcL1K22aQcOjWa58tPdHPTvFjpEHaT98
uFGpIwlsNve/95llUKcqT5VjNtuWJhZa7ssx+DZm9WsVh9YP3j8W/mlN5gRJr3UXOtgA9rhrKJ3J
PZSqvGST0BzRu7k9wN+w9n/xaeUKDAGB66aWfQZJHLKXPKAT4PfukK8AeW5p+CNwDHOgP0QzFOsW
20zweTwKUtwHEfQjrFQSojtlcIQC+7Uk7L8rjKVgOuE4gRuu2fTKOCllGOifCZHsTJUpqlouOART
k/8bEOA5tVT/pGWmp2TjJOVUhCoWZZSEScXumc0FuMUhjAW0lK++3Yv1Cr5f3sL+UYVxtMT7M7s5
a2VMkBHAaCnzgO5fvvj0nKw6gTLCs2mLSKHYGJIoc+gcbIgpFr+SiMDOC1ygMLIMU8sO8xDuHfYi
mV+VIYeQHR0yU13Bp8zUvVh66vlpQKJPxzL3ROxQU5hcaTXxzzGEVPDH03zk2BhjCBFupVKC3Oll
rl3ZvyF4/s0FEctSJLgh16BycwsBQ3WEoEorbhWoiULZFyhDpY8a83n348mUEsYSr94TIGKBWR0S
WzXSvVFNg3XVQSVApQkUnMpn06FhQUyv23apDUHAU/R0UTztKhz9f9uMKstTgEB02bIRSCZHYXxZ
Re1hqFcsaBF2q0eYMDYSEBShI1BuBRAV7cwlPHWi21IN3MpsVPiVEf32sLjCnaESNbBEQ+oeOdDE
qpMl7KXI23hNTXbTMtGsIAkMHyY+buN/3xrjeeAk4BgWO15DfeIbKbK1e5B98SkZNrn7jHiXab1u
63OP3p2wO0pkHkRfXvq5ZN5YoLTcgDbFGVAz1PpyuAPxkJlVAducqoH77TupCVHA7dnFjrgdxQPu
vNM13oeuiDHuxv880mA8ibMBkwE0jlTgkM24A8f8QSNW8LnHwegmX5hujmnf7gEgMWpft530FubW
Xt5fxev8xKyLIAiwc1ghUtdHVeUfbb+FB7Liq3PvNhVakEXlJsxcXlCqcd9/JTY4V+2hevmVhBJr
/aVIg+QJMbv5astyVr0EH7lgjdQuih7uwwqN6HBvncXMb8BMhvPNQLH9qDthdwYQbkn6+YUBY/GS
yioHqg/NMBFsy8P0oW8zQ3W9yg5MV0TWcEgFgpbLLbcRZbu4afkql/uUGgALvz/+NoqyZ+SimhrJ
H+xUtlldPbgHXzPnsohEyWyRDLKCj6Ia4r+V7tWXsOo5lW0qnj764KmF3U3s37k9+Kd9hHftc46E
O6i8qx5bu2KIf8rLVhp9QNFYzCG6IV2kj6EmPK+J2fLvvDTst03ck8mQptRuxUcrsCTVJ/I8F21Q
DO0mHXSu1O6I60yP8/uoULImKsFAVIWyEtk1bZfd/zAhml59zcquLK8DL+IBIxbj18ApvLJLj1mK
bxtAr88YFqtPvXOtxYe4fJdwUmbxtSBUXNjmgASvIS3hNyh4tG8BXEGPOTfFu7kcLkRfIWYB8bbw
jZR/OnilmabN4PUHhYSnvrGnOXrsXi7GWo+XK6G/HgO4uqxYh+/ULvksTMZCBzNDOoix/Kl6hsmQ
XI0Chi06F/2v4+K6zS/O0mB4AI9Iall5f36KQba9mO/1vpKTkPpzMMSNb5Y/9Uhcx0nUhXvt367e
cGaQyYVhrkHR3VoqRcWG1n+j/7cPNIqRlJt9P/GOHfS0IYdVyZ//oxJmCil+rc+wnBoG0Vb3dpS8
1zGbREEtq2vMMKBelvsEJdKmuRTZWGON7SqhEmFJNezciZkvnx78dXfXOLy+Z8J6vi12BQ8E0yNZ
yk66sbR7JqaiVw7jzjqYWh6ewH3GlfYIe2J5Cm76R5JFBBRk8IbPZXKYej2C9qa3Jp+R5mVjc5T5
dveuYVJXsFIh3QlxKAQtGfV5SLFWFOeMc5OYIl77AWxR9AmV1WCj4nGWOwnDDUDLEOLnlrzrPjiQ
6atweez14C7jg86jDt2x117MsJ3k0LmXbTAMAR41dbhTZQ5F0ileKuK5uync0SblJFJlLWyEXUoo
3/31vrGNJ2Gst2uThXPW4Ukp87TvbtyeV8MaLrfdFIhYASJg3PaYIf9jyEzjWLVXkwfkpGOik0XC
8VjOYloyuTao/GhWSqaj9NOtsvltjPD+eoCMVP/7UnZiCoauzOmbJrDz/SWUv2mCSw/Y26FX9fNN
LeItQaYi3c2vnHJNL3fC2WSVfL1w9NlvIStVs7MnnbZzfh9TLJMgUwAUVXq1l/G722tSbHkw57tl
KuDIFnRIBWxwdzWJOu2LSuwi8r6so/kMs1RwjWixZyeVhDsiWC7MRNGNHcaFhlsivHzbKGNqp5ZG
1ljGTlxAb358wmQAAGES7u3TO3KgBFFKPa/HGtVBTL35MQWLqkPNR4LElcVb6fuoRTtlTs8Vo3XJ
hw0ZFPcxo9zdmgd184XEM9rAZ6ztZS59WQFajYz3kNgOGxTNCWhSNtraENTEIOf8xbdZ4sdGYy82
9VWrn+TjWA284peB37PZrXLjKg2UiNOEJHC/23iTTu8c5vZ8ZksZSHXGAdhJbHf3D9FBrxqtj4Pd
z5KZa180Dl7N8NomwvL5CTD3iN5R1yBDyvZ6W36rDYjdPWw9Ky4XZxxT3sBuekb8ItJal+zm5Q9v
08f7ZXExGXnhki3iY3DofRL7qQO5r9cjM9QUKxQtp0PFa5oLLPR3zMn4L5zNeN59/MSnYi8eb+QY
ciDYOsdEDx5xDzWvIrHQ9ZnwkeokQT7kNKZ19p/Qmw1qpCctVZnQ5VIcLImDlmOW340SvlytMXuV
9GP3cmKktQ7H7zEJTOXJvoVC1TC05CUQRV0j6tatLK2xuaavUv1A66yILCQdVqMIFCmEDVfAJn9f
TRdHXMerRRpAVIQATTseuxy4n/IrH3UaAPtE+wToSynmAS3qamFXVl3g4BBrZ0uxmfMcq8t0JEge
DJz3j72/bS1Dq5eGqjOdGbT7cyasDyHsgapsbXemEDatIwiwj11UWDTu/kWGeJQb7oJpTBUW3wtA
ruc9T8PLtkUb9pqGsI7WiAUOHso3YOudn507LYvQoGsHb+hbGjD4/uxUGx/ihQSS2x53p4P12uj+
Q0UUcccYU4782YJJa13jMf3ZBrsQKav1Ym32+GLrhZMTA23gn4J7JkhwAueRM+8XOeLS9VnIDpN/
MYzeZqJAM0CKt5jm0d3oi6ncHmtFra5qFaHYcjzuUiWGhyoI+lJWiGa0fji2vY9McPZSAWAtcrd8
BjNGS/Fl37KPNuQDMPsSaHAPBV6zfyNNtrMnDnXcPFKGC8SoMzomna5rqFLJAT5ybZziJ4EkJX7B
VZEzmD0XJh6q33bMmYX7dIlZj5PvPpKNh2Bq0Z0QGY2zjg372bm3PFFKKpdYsSYQty24bd0nuUXG
OzAUZzw8cjZ3JKVd/VGnsakhOnHqeySSWNn2IJ3W0MLv0xgz59YOzpNCmxHo4kRnCCqcf37tgxzs
ntISvg6e0qeSlSuuIBIag2QXLFdN/0+HnNVQf+ahVd3vIuLVa6dibyWZz2IAwfIICCwuE89cUD1G
PPJOyorP4OXuZy8frYmpf+VUmZFylGTUqwJLxOyD1G8iSspNGV4nWhelMzWCuR/jodQuOPGqdp6w
Qtkm2t5bTdXUu1YeTBmXVDf/TVV1O+T7QYqJG4suLaYgaJOBB1P37lYPmTAQtsaum4q96jrszH32
keXOSwJmrJOMhRCMAyf+ikc0GKNySNAuIestzHBJq3hfnSLgFFi1zbXcV1y3eJyUjjx6XqJ2dk+P
iqhzvia2KdO4w9wJLNDDncSKYPcyXudB+evFOwTu4N33xltkF9YUWv4bNElIlEdTBNYeTNFTa5bG
NOwWB7M0hnYlhoJTTZMD/IR+BFHQF3e4rl74BkMU0OvIfqo5zOP4S5pB395N9PhFdMcarVDEC5zx
9VKHNWW1PJ7y+SS3mAO8847b2uKeLYa8VsRUASX8gimZ/7BeJlxiF8uM6UxAghjnYhjeZu6EiIFp
SS4HDO8+iOCLU0co8IvAhtjdk6C+7sWgOeI9lTRUUS9fypBKrWvbwyh0R3tpT58CjHEViYA60dfJ
Gr0PjVHqRIhAj3y2L6aWwkFXaFA+Qc99+XlyRCIiJnfBno3c9yNlsoYEw5jn5R4S0yBuZf9IlqpD
om2ERPcKAo2iyj2vaZWJ0rF0ApIck7VqD71KKHa01O+AL6tidJCJEecHAEXfei9c5fk4tkzfa59M
WCLKDFIDU2y6pmpqw7lQOwgV/8rfPgw/YQ2sk645ESaM42TFoljZDEx0reuQYpog5dv3TS0FtgQF
GxwjYLQZd/KHbrjMnNSKObrx59HkPRIMGAqyY0e231k0CpVxtqFK6kVa/q4+nX/Cb7JAsy/AzbXR
Im2xzrAQI9c1UJ94Z87QqSJs9zc5cpxn0ISEbsmF/hh2QA+B/LTKba9WbUso/gCXhHiD5W7g9dYz
VqYYS31Luk8P/zt+Vc+7EjT1DZjqo5xO2zAcPfNwN4nrgbiCfxhR3+a3AQOSfbKxKcoESMvTilRJ
ShibBWD8RNPAuaghyI4lps0rzW62JkrLMkGS8LCYoWZbss8+ZyZy3DEYVs7s1ZDol5keoNbeLiwu
uaUnP/kcmjxlVUh+i1FB4hiNEKRsbh7XxuG3+7eUqst93jcWNg4bL9Ze0YMAFzEGwcY4osHX2Cwq
EBonyNuFr2szy2IFfLYNjZ68WYlFPSDpQ5fKpSVVZES7ESKK+JumD5ezwhcIiES6pS+5zhjgy6Bk
+2tADxQ7lnFM3h+JO7RMGGtQHTMc12piAu5Bevk1t4SLqZpQOZC3L3cjkNlgCcJAhrSLbWd6G82z
3yLaHMafMF2wtOTpmIzxyIa0qFvYGztaUT/7RDDZb9JgErWNTZ2Kb5a2xUnnmC6g3fiCHI6QS02D
uoDZTL3dmYZNq4VyWAnDq5/XnoBLC63Qp7khZU45GpgRnOYMNRqzgT++yIZq6VRNyFl/L7VM2X96
gDWchTOw+/S/CIkGPuUo/UKdvmmyzEl9poSDDx21tItWbaRKqqOMbIpVzZAc7uTRs0Z7dIjBzVWR
4tDIu5pGjcO/MfZihnVuFwpYOTGL81MxpE4wk7UZiIfSDNAXNgSNafor9XBpNGmY0jvNLfVqe+dp
+gm+35CIRaemKKR4ekAVggjc9YlbOEzoYZAU9eO7aHNN+ey6kFRfxd1GgINmb6yjeT4vnH1AjnG6
iAiToy17OZKrA5sVNBJ306kZp72E8XyQttk4NaKmPdwFBpwi7KSVkXBkTivL5B6M61xa7Nx7Xz5z
TEzWEEU62OAzb9zwQ9zgH2qnIClNKtbo7IGcjjilLsCqFbfIe4GXINYsN+PmzCTnTkfdLpSPnptl
ZIwwm+JyPDv8F1GXATUFzj/xsQODeuu0mfBPQHrPasRm2odaAb0EtPQ987b94MTWewaVWdpn8ssl
n9tCRBHDeZfSXyRcpbw6Q7FgVoytFxFIHdpctLR1G+7V7zNO9v72CQDDAU7KF7XiXLfq8i110W7z
IhjwSjECcae0DPBnawk/bsFp3U/UMlgLpBrbRE0G7wCx8hrj4nUtlUK7iJX4tAY/HVNUf9QlB3I1
cgiLwg78L0O3K9hP6y+g0eHcffqN6TPPzAyGQqveZI9GAuarLrbYa3cpJ3ubcCca/oPVPqpJs6yJ
fbsTGWDOvXVis6hVtKW4zmDfTyKHt3ID5O/agXG+Lv0iZSsbiQSjHNNkVlvTE6EBepTaeCTVJwB1
NewOQeGXVFjscn4IfPPDsQGD3yStXfT5qof15HCy1Glac1uws9VhDncu58FNLUdRk12QotCQyIXK
pvuejj9LRBsxWe7S0Exq0W+0CnKvqIIootxTf/VqjZWnUdHVJxdBc23fRUsOBVp7NyJKH/Zu8f4s
gSybn3lcRGQbgPPlIwEoO1iim1E7F0cnqvnHRGBvWpp0BN7v8aHyUW3vLYm8NU9Q2ylMxpUZ5LJ4
flGOjDR/jUZ47Wf3C5U8bZM+YFdImzJ5wMXwELd/8UcuS6Aqt7XPcsZPJ7irQt8V30xHNnWktMzl
/cQJh09K6Jvk4xbN9iZ6JvWyC4GDzXKg0xg2Br8qa6Hcal9GreC2DB1BCEF9FW3ew72/+ZYo03AH
X2DAStwdm7R0naoUO622iMK/6tLFZ9JUIv6SW76r4qvSFeo1y8Ji0PaHTv0Bw8HHX81Vz1RMQJVr
EoLRMwFagiaWQPaQtXql4r8MYkTZ0j24OhbV+UGhE9FodF71lvOHECTr+qRPC6smUgN0Xvagkhkh
pDwvDPr6yk/u3oI1uhUrl4RdxxsEda0qa3sCabtTutA5yQxaOtgicaM8klWdWU2lpCNKQGeQP7JY
cnGIHpk3HIimayyB61q4Zy8TXQFT5RUYdFNVXRdvCsfaqwIMCRSqcYZe4hasYAQ46RkbMHEfmuk6
OWa+qWt0VHGAkqpOkBkfvDQW3reUiUpqTU8aR7h77Th2ue7R4Kzl+jI69yWezsqrytTtec2W7XrX
kAbAZa97CRa6vZ2g13sgyaqN6AXXorh8k5UYAek8gwopoe94w0/UV2IvTGUQfOTG0eNGBilUtWPY
pAx27GhtahA7vFFxN8jC9sqzs3xusmmO295+PqOzkljwmbXd776IzGys8VV2Rykm2ZzB3WZv+tZd
jL97Uv3Van4f7Oud8q3k4bW3UMHiT2TvtBhymSao1LIhfsM9VtvJqPdo1CfZNldWH2I8zfoWNbgY
TqdqgcCoSq1brG8wwzbm5pJFQLVmhFvHLPxtdqBYIhay6/XswCyknNVvGEcFNgfvaN9r+Git/nah
YcMv0pJTdhMkykTKKvI/kevh8U1ED3KR296tgUEn8Bn3aVJzWHQ3oQPUZWvCq9x2ohG+Esurv2vA
iGqg8YhPb7AAKmLNa+qltEaA2jxMHeWJhox8RItjhDtxYX2SDnwOKF4MNZVS3GDLrVWscgIfmmYP
0Qis9gcO8YmJxVyuE2CzvFfIwUG+7jPksANmrRcyRpMfYzMmt2hRdUuodi8sAsyUf3ix8GuW5p7y
1qKavoalizbiRyKjBjWHKY+9xpXGxfwOc01ka633SbYzz6U/d3mhjtPZV0gD/H/IpTlW4TOzj34S
afAeGizu29Ku+8ucodOypbpIZUEUQHpLSnrjuE2O8+mifrp+xyXUSCd5NWEy5oD6RIbT32QsyJ5K
kzNbHoesgqt4prVdaky01ZyqSOhRH970ert60BtVs1X5vRWv72T75yq53Q0VHIoVO2foKpqplTkD
jqlM6N3pK1aBkSMIMV+riAzc+Q4+5bjDuL9Nrm/OQr2OGCCEyxjjcVFEakHTBoXWv2dfBg5SwYEh
9oGNaf4DV/i4Sjn1rmwLdBcSNooOF194khqqt8e0kwFAABVJwcNya+0a4bFsH4Zej5UdW7yW55BO
w7om68F94/LJqgjDHhRbm8pFov1CcmkgamvU7Y5Z06nCKxQ2rUhmomqyVTrM7nBHgEjfEPFRqpj/
mkLNmm1BDwqNcEU41MgIOIuLLGlza1eYpEUedRsasRP5esnfSf+uvnEAfpdUY+5ZkfVbF6b4Mt79
s49maPjRt2VTNnVyvQkxF80sYlCXf69uN7tQLhCXx+/BVQvm/7qnBGMr2dEcqS5D3DtOQjp4scHK
y2OPvdsTLUCdNeWfma63SSuDCqh7xVsvOIu6BEvv7M6dp8P7gueRw1LaDqTy5+/moyMdzHVATCq3
+va/7oviWN6htfSxyyuZLyP7BADFw9DS/sfahHUZvMtLCUca0NcO9dILw9Ol3RyhF66qtjfB8cDA
F6T+KVeNl/+iKxuoi3hl3s/dfa2mEYGzc3VeJ02Xrz2sObbwxk6wIjc3fOdQr3coELDIRhfYDm55
RQIAjaK0OXts2iV0W7qYoGKimwvGFFxeqLdKuWeawVng1Y73+MEyQ5ODdnFoSIEFaD1IhlPoBL8/
PnFaA/Trr65VobMFC8pD+e3nDI9EjQpbG5DR+m6urfHNJwKhispvHToYGvEKtH8ga519+Vm2tEO8
OXyXM6OwFUWkCxWAW6GsVRr3IzbRy58axnck3vDmEwij01OyM45fiMsWaQaCY6KHaZi7K/bviF28
1nLIwaWazlx/+n5D6cDDOBTW6YqPosJWLYvV6QN2J5BIrHMc9hTiyFwheqnWv/T1u86BRwjqvZtk
D3pxcOfZqPCKiTlrW2F5gFYFTJebiiKleRN7KAPiFvC24gWnEjKqlebC2AkgWuPevLOE7Rdzr/yN
XlMu7kyTokfnOK/qfPOCjxY39xYV3AHz28pCkELQXcSu4iFLoEmMBZaO1M5cfmNojRWsWtDDO3Jv
VKPioBZuxzjpG4pdRy5f10Y8tkJ1yYsHmtI3zrCaOqq7pkn/vq7PK142jrZ0qtNUh45FdQndsV+B
7mRgdJ7Sf08wGsd+Ip7gksiYJ1Dv3mKxQIBZZxiygxoBltcG83kyZeLuNHTQ54czUxE7tyrLO3f6
1i1w3ELCMxXxiethMUvCUKkE7nmwFlk0pAUXd4xN1p+v9q1z1i2K0+S5500a9+vFxE77NhT5VSpe
YWeCHbu4C1suJjX5ZP+FgjpjX7ln05bKTCmNygaEYuxoxF9dGxiPQOUnjkDcJuM6q0P+ZMEAAz6+
5prTlCJVrP08acErHVCQ6OhQPrL5JEisRt4OusuRWThdJvrTl8J03YBhPAjEKHxSAjI9PsWU5q+V
OEXxjfzJ78wtpB6EIg3jF6CebV+4CSSyRIIil/QJZQuCeGzGQVNiLV9pZ7c2Gr30vK7aPLynaEOt
cQIswy+VUFhX5VulM07lau5ESyDCAo9eY7Gv8Lk37lGyrZ17Kigv47344kiM3XQspDrPTyWKBWCl
xkGofRO5oYFdnytKwsCbDPlpm8IXXTUUufGGbPjOunPxvmIeSKkHTRI1gDqZK0PHjZYyqz2Ikcaq
Udue2MGaNg0YmuEUwITvveRWCso3yRpqO4IcxaHcPCGHuPglT1J4DwKI+srjBi+atcQj+VdzPnKZ
xJhk05Tafmf+Nfvstqt9tUlxXz+hdSBoi/DA5pWAQEDSRi+6PnAVAsBtkw4Z/7f834mB63mJoa2q
2QAZJ+t9BmNXoopuSxmy0+g5JjEVLoCkA4qE3f/s5P5OKD6tBgf8kM932CoN4bw5Go2zXrnLv1Hk
uJ0iQ8JMhctXY80GSmgvU0SuUQDEQpiDW1UCNCzxS0eIPw9DIhpm4l8i+lwvZahTOdY5wBy6spJV
clLM/4uGuOr0BLOVaU+w68YtOOKXiuDK4XzqYL8N3UjM2zcwx96ftipYmdcJx+RtUCHHd/1/VyYx
HyqsC/8pHv8jH2jmjSKW8EiNoe+UsqGDSn9S09Ooc9LZM7i7UvDPXiNwO2PCXGoxYb620jV7HTsj
1jDbsYhh8HwtjJdC82XOPLsOgWDVwdpKI/5IY9sW1UcfJVocr3uGBIhc1pvEr5EiXpw9Bkehrrnp
TBy+V01EF5tyBMGIKBMqiVg4gF7mLC6MD708VAH0C5tP2OjtLYzKF+BJMBXXbG4jd4TkuJ/8WqCe
342QZ+04OE0t8XBQRgT2M1h3qpJChrK1Nl91Ze/O2a5ml3LEfDCC9fFbCGwK9qq7t99RiwrZ0GEh
dtlIQMLm7UXxS+qBSpSyulUlhAoSBpWx9KLmRHn3Zx6fH8EU9I/E+cRu4fsyr6r70tmuiDUFrq8N
sL2l0bO89b9In6XoLvTGSw2R8tgzm4/5hn1X1CItyXC/zVAleETVM8HatVK4lxzIOJO96GFkk1WI
/JbaBMLrxsfAimGp2Bwmr6izZ9S4VZYyYqW9Wg62e/Qz3CeeDktsvZsF/moRr8JohwCqB9vCza/A
dc8D4rN2SByTsWpjDKLnTBl+0v+WQ8pQonm3cjUuDhadroQki2a2y9eKhjopRU9afC4ob3wln4Ha
+vuQ0c9twIOEzCM+sa2BqRjxjGhsP4B012qmpGVJ51JZysgACfMGmc+L3Z0NJeT22NNiF5iVbjnU
hbrzuTFURtT58qYYZCdMooKao3pe/QeYeGvP/pYl7zBWvZ92AoxbYIC9Zrg5q1Us+XV5banNVfjX
NjTfqFiecfmIty32vbGJRBL9ZT4xu3ZWsi4dbzHSsF1cmsrvmfSizVmBLjqoE3qhx5g9iSP8r1kI
uJFg0GkW5UcuirVCZYoMJyE5tPZSEuY9MoqfWVCNV0+mgBolL3wNmTSspZyJbjGMDZgVJDzSSxwF
mdljzYAdF+zrrB9453z2CeP6U+EU0/rVuq0bf9sUJ3O4sFIglKX1d4oMgFZK65Klp0JhKHwVDoth
nxK4+JQ+e+zNdAFV5Teie1tEt7bYa99ezJcgHmx+NO9TCTxP6I91utHXen5EVVEYV1v1v2Rc/6ZX
k0dVz0V/4bfeaRrXb0MjV2fWODUWbDL2KDPeb3vYRAxuWHD1A6mpE0Jy0DgZ58/V43QzkLRxYYBc
N7QVPxoNgaVK/vLLd+53MTImjJQoRIDh0agUFQYYUEr8BWNXW1e0R0QeHGxEitKZQASRhaHFhye+
UC5Dm7SmExVnH3+EuC5g/+8WkKmLwPUQj29d2VfRYXgDt/dgRhngI5I7w36v+IDVENVetxyoHMjf
OsY3Dj24UvIbK8qZSbtdZL4wUJ4VZ86OncoaoLYn1uHYN5B7xL/fkReHMaqm6cWc1NP7c7CerMGA
QXZzX7UogmjB6GCbzlyQNrg+ljprNZlxWfPcPo4XgtUkrmPFehHiPloOiCXH5PTMPXFj8EXJPBvu
xqVjD+Ai1TtE5qogc7D8vWtlL5X7ajJfSwrbOES7RqTRS6PxUazQoit+c80ynNkB1a+8HyV8yCSd
f87wISpq+L05f83gSf1IVLpjqLF+Bb415yPS7cjjvWcz2hV2zo/fSKw0qSyvWY3DTOzlcWhDynjC
urfh+ZoTIftXlDXY/Vel29xqCfNCGWO4dp+eFmSUXQYxLw+2nWt8zqgdkAELVKZJ3YPAvowa8IPP
8GElQd3Dv3EBBsYIz8KsS4SggIxOPld7qyAPrZ6j3U/3uUbm8MlZ7aJM4oDmS0XbH61vj1EhSxRu
zotBDQtu6AnPz9zJjdyN8PYp8nHTFJjE0M5TC60c+iQyMHb7sAljw/jdYwxAKlUM9I6cqBdNTUUs
dKdEPnJ2YC/sDt+1Y0kErgTx6RvuL0k/0cvnwnjImLl7bqGyfh8mct3aWpbKiHYuApRl/PE38zEE
roZdEZsp7kca1F+mFLtyPuIcXftTs3P0ua4yYdhT+mFHpoTsaInb+52UJQ+9mcSQS5PEeRCmc1a6
ftW7jA3bQYaqlC4ZV+m+pKNZix64eTL81OQ6eE0gl+7YUUtXul9K8QLv5YgqCqN9g/vVcWx/fxFV
7Xz7ZrUWmDo8X7vSiG8STvwmmQlvsJxH8S7B2w+7FxX5pgLugJvVI1eZGaLpra0ZYvK/xKrbablK
BXxeZrHT/X0goCQLtgOMF7R5qferFoshSO+pM1cfWlgN+wtpNgblSz6x4GQq579IB2IOpHZoTw7k
e3rZ3/p78mA1B+qxSdEVmcqELd0ALFI5LUPiiGGBhjsY/iCrSvV6BpGNm1eCTjlhu+t65FKUihsk
KUII2FxMGRuXUWXrpgO04ZEvm+PzWQ4RZcZR9CXUJoI+WDcbCdnTvIYB/Gsls5kNkfy6xMAMyoou
61yJ44ZCxiPal4lZgamcveVUMMpwWCLVClsol6aSM8HWI24++ePvhzVSt8TWloqL2JyEtsiUqGxR
utalecAIrOyeh/g5I/hgt/K2MH1QD11YS7LJK0OqhZNd47UU/lBWjY6iQNTMp3ZpYMhhiW4c9/+G
wYLmAZeo3CBPjt6luhj4wJjbS/KqsMI7meKGSoxRome4DHIeKexwNLhtbGjJaPJjnDAP5vVOZYO3
id8XLEI165nvi88gvo6XuZHIKKaM0PJrMf72KqpwQ3z8+W8byH9UAt6wfltPA60W4L4nEhQjDqxu
3OJk1DqV5+HS8od8SMcPheyf9COHGLTF34cfCHTJXNhTKdJiJwRpwkD8ZeFkMQcZ009DPfAicO3o
uXKOqFEI+bE4PPGIpRGoSgbiLCDPN8D1IBV1aiq+m0njvnWuScjGxMNM19XOWFvbwd6DVL3W4A7v
sJgJVIKpzF+3azrniqZWqsU3S9DapLK/NZuSgEZbRUl16eU60Jtar8mAVhuJgF2Tvy13GJeBj3di
LrvOWfN0+9CRiBKrdbu3d/FrrLeBp19lsIDpsm1vBj3LgBYLrNnjecG3MDX/Phsu5coZwil4Xv94
Jh/jc+4b4h0zL72P0eMr8yDAf1G5KdlPwYGugKPW6eYemY38Bv4iuIRi2Q7cYS8sbEIX0F4nDASW
XEyV9+NgNTTQ0so6MJPTcgVcklSGdNogwc9QelQnbDAqniiwXTnX9LtEY4D+j1K8J9HRgV1oOSB+
/f8s73bMuxZuBcu+qY+kEwsgzsv1A7syqjIZbe7RVn+/OBfLKYgGdrICAQKdXaFX08HuETP/cPyP
H52dz2CkpuRbPHH/4jX6JKsEVHbz18HcNVmtYH0aUiXrteYHi/sm9hqw7rr/Fkco7Mq0OTUgzISb
OH4aKZnquI2h1qh+RKsO4bEZONhDA+NPqLVLWYV4+enYTEqUWMWJaZrHRTDuCqDPi2hzxGQLmPW0
IZ4HKzSgHCLWip1EG+tKQvyYr1kfuqbz6hlg38CS8ZX3ll8DYdxklAIEjroQGvcEP5f/KHfP2Fn+
SPi27XofwFxZiVTLl3p5PLiUN5kHtEDz2BHnwr2qN6UcH5DWql2nETn2GlRgtpDfdc77nBsLSNR7
dt1yX2wU40J2e4k2yVY49c34tGr9OiDoHR768lYJo6q6LxL5hAJQxZukH2gzgoK/TjcGmhmV5iFE
xuUzBi4JqsPzJxzJJnYTtBanO4lfYWIdk/pm+4wStWHRuxDuVCohmA45b7IS8gM69zKXXZJBcqEz
JRKNlV2U3U54ep3YY81v3f7cgu1Gx1j1v2xIrt3MWD7IGAHhlvzhpTHCliiQtIL54h4ngff+4aRa
BAh932m0/PweYZC4k/IjrJ7/BDTKo58WdyK3ewi1DwkOIpCldya0L8wgurypHPn5CZX8atKswDkA
kxSuAo1W8rqaaPoPzI5nIkC1U9xtf5lWHVtd5LdXIhonoFm1QiSS/xKhx7SoCrfSieajQMCuxYFm
zHmCY92/SjcmbPeF8G7nXfa7Aep+5+oEw9G6K94yoV3CNAo4y/0cSCmHI+y6vcdfgeYA5IHqauSs
ce98p6BfiMyS41QOCmenUZgIWu9iZfqKkrXvd3Gj9jbu2w/B1pbWyc2zj15KQQmZ8LaQj3ta7bMr
qkPt6YqvBof+wq3AjpZ83u344dL3kydrbZGttDNc2edW5O5Z2XeUv7oAqO5d3hPHkeKmakWmFtLn
c49Vnu7Z2ML/FWr1kEObnT0SGb1FhKyRj2kuG+sPhd81S646vZbA9qNQtcBVmS1Dj0sQJnKENYhJ
Y+uqMtZICoqqythp5oWhXj6N9LCiALhuBzvpejHDKz6IIl6KKWzxTICALqDCOXuFqNPmJphHXsF4
AYTbXhsxiHeftDG5S2yWRvmZsKLQDhaz1KRtlLs33eB6N2SlantMi5MmYxh7YOUPVCNyfyvy4GYT
73nbtB82j0JuGgx9S1hNw4oMIdxkSFrdetnTZwjaT6fRWo9muf6m1ytAfaErxGISTl687vdARJQq
E4P0XvWjFPf6aI78qEXq+6ake40I5QHqB51Yik7dOxm+VDc7F56142uY6oxL+7IB1kEN812zWspZ
xKuj7jQr1bUNlZ1coFNoFp/VrFolmQcRRYHf7ZILDShjW3mJNn4lkOgDb0Wmqfa/WHtCQ4VQTWOS
Pk36HlKFmF2Pl58eFvkxKXym5E3cw0mltP7AjH2+d/bP6uGsC6CBdVl7vjH4aegx2yzFN7Hvaffa
lHEv5N4bdYPbtPjKSxI4LbPCO+mscBKFD6NYKb3/zqk1+Qww5Z0htdZgvhcMbRP8Rh9fsDeNKu99
T9mtwZSzhoE0k7h9P/AAKMEuJIWtMI+4NYVZZ+lNHA65RI2a9DCPoQQ/KZM2DE+k6Wq/GAZe2ZH1
Sm5kH8+oVum2Q0LV8uX3K9cWWLUWDUyn0zGgiNw/5wjp4mklkZMNwCDThI/RLRM9bZ8ND7Jq4OIE
khlY7YAU4nqHVC/oBTPAaJfhvfHl3z6CceiTQ4cCeSvPCG0mHv86Wzu6JEAxjw/uJZ4sO/R+Pxfq
haWWO6qZqzco8XGv/KiYHnGMAC/fYuwYM806qtI8gC3QjWDbgTX2j8nQ5lIngv75TXTP+vp/wP3a
Vsn7pUYGVtkumR3i3jG8rVVAd9CNw2a2M9h/hbnLcecKZuKvdmWempZRgd78oMmqsgLQfxO6bo/y
Rziny1w3tJqPYkz6dq4u4LGPk2VfH90uuigFSiylToYCemc3rZLZVlEd5+OPrr2jswjUMUBWZraX
sJL+adzgP0PRIL1g1ormZjut3Pp3hzZAI56igIs8mIHIDITUqeCxSrEfk+JFvUnOA6PWoZeR176c
AX7D5b/WRdS+6amVBvyNLhbxjY7WvaIzdAMYnamMbQO+NXt6sVkYJUkp2/Ho3eIq9VTKCvRZAGm8
+3f3ImGs4cM48S4wRUQcsHEwaEGIl0Pux4ha6MX4zNEIFCG2zyPLXMkz+y4eHfpZF7t87BoGwxW0
Q2lIjl9udKmCA3d6zxj8nC94i7vYMBwKvw0yzjvW8SDBEk6Oha0/dh52sYuDJkM56cOmlyz4fy32
kY/fZI0mqm/jZ2nFVU7A+or7JMiTn75XPbxF5aws6D+njpqRS63Bog71xJNfuQup30pwSGQMRekc
S49H2L9yrU03cmJ+oyWqb5i/0gb9Bbwt9w86hdCFn/P5lmvnLlcRfo0/TDXeJHzITXQw/gtw9cLF
4VfzqyBz74aLAVuSTz9W0vO9YMjKCbC50FrwCWPmd06uF1iAFKFVK/qXjWvSAE9fLAqe5rwBT7bW
hatkZjXS96r62MGXQLfqWz9ZC8325n9DG5vtA1OlOqEFOY0i474nugF3Y0ZehZj3R85SAZOhPFnM
qhpDpfIZz/LCYbQD2EqxYwgm//8aqLyJwwYUb/HxLeXYT3u2VRg3Z0Cavzi6bPNX+idvnyyUM+Nz
mPCVJJNNBurc+Ctf2sNiSmR+nTJab0v9wNdSh/ci14KveUVRBt0EWDz5u8TH8TJswBrOd3k1Oa2u
GSaXpg1OyvEDTsnSdLKMF52/Fsvf2+wPH3ucSoH8wSAMOaM1degfjPsWZjZ2enbBtd4oD9ZdMKdS
VP6H1wyoa3/7lSLCgKypKQM3moeUthDykxjozLbGpG4plcVzBXBizpZNr0YlNH9a9fJsjJhzV1cb
fR2II+046u5JTDk/CGkuVMfl/KFjE/tkUSq9edJI77huuvSsQd7HBPwQNMPNsRAm17Nv7sOwJJ5R
yRM5XPjw16sYaEtmyk6Eq8jowcJC2kqf5uhuKtLDt2qDnb/h7cuZCM7BVmO1J3aydhSAS2RZwEbC
seEmsi+M7QlaKVCqK0gEPKMjrA1SPlD2T0UjOodf+P80V1htj24bV+I7ebi8/EXZBIRufKPkf4xE
vsJ75iHQ2OKQdl7BeC1gG+H21QJlTt6PwP3E62I+jRE+1hy2gXVpQBMri3OTqZVaaY8Fu68DWCVz
AKLz3FqChWUwNhFy8hGNqzRt7xY73Dr3SAe+anHmp+Z/vGsQqnOTv0j1q+FE6CHG/jChuedzF0Wn
BCCptamHDle/IQek2Kh0af/MrJUGf+9M71pNz5yfjRRlOqyy9jf041NHI2fiFpd8nrnKOcTpBagy
+AmU1Hy4tAnO2SZwBeqHRnFMcPEdzIyR7vVgJwasb37D/nlBvqdk2k8Lmyu8i9SQXvvyKbvmrUyZ
kCO3PbcolWUfFMTqYm3ouGflPvbVF36uasonHUiZ67XJBtlfOMtIGJinNY12uaIeVV3dFVkVZNkA
iSd7CQWn83cA+ERZS/SnHJx1ebHNvPrkwT2+TvOL+3v/U/65q6vCrehX6LtquEVc79g1Q4yj6yqz
AdkYBscQnfyDDe6mOsmJFqDZklve/yBav0qO+1ArydVl4qFTyR6UEkZW4NqUPx7wKwGhlwDgp/Yt
NnGYV8r12YI4du1mpSX/6L+kDVpZeDjjkuvJNRl6NoaSR9aPVW3oDrHZhSHprcF4z7ofG9TtHHie
9gkBCFJoFzCWN3hqTY8EMdcSWGsw6WkUAVOJ5SE+Nics+sfD18eB/GCM/c+K6P8FNUPsX2HbuACM
fCjWEedlhUA2mDGLMeMUmBL8fW9thAAa6xuABAxwcXRNPbnZTPo6QaFQ56QDeIR6659TjNZKIjTk
huMV0mvrO3zvsE9dxpYQSoCFEXTfWXBnjR38UnjIgn6/LDRXWLGepkX4LIe9zdB7gPpY+snAht5z
y1xSBeSD8ySTjluOJvEvNfmIlc4G6r0JmI7Ta/m01ZgW8gQqdXwayfiljQHxkTen8gRHwZnV2f43
C3mTafP6MaY7rA8KLtELKxkbiJAJ6CNXnv5+DdRZAQi/glYbV3vP4DDh3QwDIxmX6K5EoHKJuyPj
TTT4P5XXeHFAYhTiyIMTJ/zmWa+iHG/eyJkDNezWaGxGTTSuLL6ynJtHV4UK+X0X56gSvk2BT+OZ
acsX2g3n5u8b4savr3WEPZj+x+7qiG/rP38oQ8WffC9ypuabXXLpBt1zIBPP45w+IcCxLo/W/Ztd
/WPyskUGQY1pd6QuLV6ratpGIQR0kZhSQjdiNodZMzp8UjG6Jmmhuqq4Rr4MPDMsRBZRDc7gqQKl
SVwoYkf3qZWNUnnmxlrjB7zxY+9A+hBEYh2wJp/BLnLYb0NmRegu2OEyT8DbwJ/tcp3rdqP/2J3J
20UiRlDytEFzdf9z/Ss6ETtWjWgf9Hp1LUmY7YsrTnexDKSbEyXzW8vOhgeyfzAm2L5jX5a2PsRh
xM/9xzKlsGb439/XLboaXEqdhTmSb6OL+zAtO9imWPBn3iw78pfa2h0WS5LubJ6tfBy7kUKTXCiT
MZcYLXuvIhhR0JV53Q99MLderLqTta1X6jAV5S45mcRXGS7CsQi9YKLVahGYqmo2lOBbBdqnHDhr
ddL2+M26F4yRCIWcZfKkSsjx82wzA7VJx0ZHYC/Ur9m9d3oqabETz/8vKOU/JBPfIzoYAeLSWQj4
LqP+Tue50ZMkYdR67VKqPS4nKtaMnT1eCFFGsZS/V7SSqADnP70d/kJxz9E4xCUfOrys1Z4LHkd5
cZYw+RN3hMs1rgupxmEsxtfQZkjwWc0p1PDKdwLGZKmg2IGGLQAadNP2NK7Py/tEomgDIdehabmL
gK6SjQYLHyHTOcPWP3caGH7NLM2A1xEG63TeX1FzpIQGJN3Re70AB7VkR4cZg9ZY7Lo7kR4J2Jtq
V0RYAQPa9SiD09hh1IHh8d9ZrEgyK+kQtocthH8jipmdCxOmuW+jtjTygHyW9U0Xzq1R4IHYJKmI
TLUCHxytIL1gTtvV221YbWvB0J6YDvHQ5Ef991TFEomdYq4ShHX4R0ViAmfP9+55ciWFR86JXe5x
KAPl5FmEczeERFAVikfr654hLT6NHiip/UGHWi57eReR141VFu+wdqo3vQ5qJBUkTRCL+gOINcjp
nEob3zTvqv+NSDwHqPrRsZrZgU6z6ZH863JF0/i5G5OlQlN+/fsE9wuUqfjEmiEW1X5IGeRsGapD
Aq+V5qNLv7kBf+GLZ8TqPN6mrL82FLA0oh4MFrxJ6T4w4Nu88FA7uUkZxHH1hRgdGp8MFC7FDSPj
Gn3i5g52Pd4fVvRXyyJYJZmYHq94NHzluah5TVp0XYIV91NNbpMpJjy8GxyUoYDCA81xsMMnFXPI
IiPxFrhRiqmxd1LqIOjUoQbbo/KKtav4o+qos41XAs2pJngRX/NTMMCYl6rQZEKNYZdy6tyiEE41
oHSg15eUUbylcVADJD3VfmPkTjWkqOFzogMLg2yf5qWnyCP7tTWpbtKXRi2DqDYpAR8u7G3dtOyR
8K22kkt7F8aRNj/HsIXSr29OKIk+4aT2Y1VGNpQKNNpW+Mad0lzL0FgGYPIFRbtDFqZQyopRUCVi
95CEqsTQZ7Nzng472rmN6hGOgT+Ce16QJby4by7PquFfBYJnoMJzxJz6OpV6wP/d+q9xRLnPA4yf
YEl8JbbEaatsgrUtihVAh0r8K3p/DUqT9A4JzypjlPqwudVIvphH1+Q1+YL2UgbjNH14lf9Tdaku
mr2qr4BrMMCrz8koshsmQNuqydx8PUg2A1kW6arLsJmyTSCAngLxACbTBurz0BATLuzOk+Oh+7ck
hU/Oh9Xcr4ZLXJ7CWSJrugOA9eg8T9WiPdu3jxtR0mzADdeCS5kG0UVfw4wdCFgPriczRxCzPydJ
jTMZNpKC15suQjLvyekZu5+Wm5c0SPxoC2WtedHvaPlBUCPAInhs2O/Vq7mw9MlOOx3PbMIHz1os
r0FPcad/MXWQFF/U6GKPuRNec30nhcErxm3hfz/HGFFKZ6TThgfWgOgwO2qv0zYtjkNgcXAUEvMm
16BqJHNyZP4krt3rup+nBOAAbPdrm8rIz9tL9A0IOlbG5yAzsS9YTIbxX/PyGd+BYkWmpgNEYei4
+d4aJYvUOS6HgY+vAsL/2YRnEz2YijZuFmUOePpVFHpJ3vI6VHm6w+rsK/SQwYINPreSkGGAQrRN
nxt/U//CvS2QTjhxN9j9uFcan1P8XoDIG8X1xpItMGWMgNuSZA1EDT4o04a60zPiSJ3GSpFQgLHQ
KFFln6aVpReQPgOpmGZpAkpfe0OmDyy1HTAVD8EqNqjNwunz6pXhUayygAx24B7YVRRv1iiZYSGZ
kh7FN8FyffNc/plNPk17/IM/4m2D8GBf4tXsMg+jRijD0ksKUChpaV/M7jtkwZUG9fpN/e76AK7X
L9NEge35UnzS+wTpw2XxcQfEKDRUU2xsbAtyDqtD9W1+CQp7ILMC1gP/ssb7eFQgcSFuMekZieFg
SY7nu6cS1R8Z861pR9OuoAW8nHjzv+9soHKRH+yI2/4qczesnchX6qLsKdmvQ8uXCUWaIt9XfcXG
SsypIK/GJ07DaMGos3uP3RdGIm4605DYqtrBBTmvVnyyy75uObVQCEIhvxZRf8iGxWattuY+3MWP
dbk3krtMLtwYcXcpX0srT1twLnumAvHJHhdAaZ5C3owaVtgdybzXcqIph2lrmCdkSbTB3mqXO+Q/
Uqv1ENE9DFGqDl1WYApwEJDhBj/nhISjXwBFSAuf2/u1iJ1/n4pC+njPqLuRyV2J5l0x3lyD88yk
obIRyT5bgbit3sRIpPooUA1Scjug7vU1y+ybUvczC7jLr1jzWRhGQAMPtMI+iCPnNunz7Uf6cbRo
5dtGvRFRwkOWnlU1eqHboVXeXLrLQqrZTHHG31IifbuCG9TlzoDdesg6zYI/ItqpjnBMx5ds6wj0
gPh4YcbZbuCns7e2ut0NuFy5tFxHK9PS32gYmpnE4Jl65vebIkCKtsZcolm3JzQzcQyg4xnmxr+G
YLBr1QaaAS/59+6sISUgspSgjyFHnFJpk4nSpmQAtIT/7/yrUeUQ+R03VIB+5XUkux4YPaZAAbN0
9vwuooYazU+Gj1UbsWdxmDHEvnHOjzAliUxKV09uScr5iYh0BMTMOUveDGJd2u8AuPdk03D/4o3z
5nvA2gxvT+L2n3lvWvPdEjc0P4/siye7kPp96lND1HOsYxJnFvtaQ7mjUhtMJGRGXoeWEOeE725b
8KHD59v7YzgIyTfH6+ZfAM6O4au8PHtGz6ZngFaXeyA1Kn9PEH356Gn+0EoHKYIIZpO76Ez05l/s
/JtjC6qHLWXICX+yPRbM0/HLfkneEKy6+yFHDEEaS6VqLA+dVHHL52DiBNuS8MK7+25E3Y3xl3XI
WLxa3l4Ghcg+mLER8LyNMYVKK0ezHE99dAxAo5+qF89qzpq/tdpo/U/CF04VbxsHYnHvMt9dmadX
IZIacdCwBThHd+aB5TwtMJ3jc6vVzT9Th7pWitynuEKWdjbQsyHIbYdexrYa+0Xy+kEAeSinNF1A
TcCZsRPjiGmtl3ChvbBpmjrN7zWu9yTdzDzDiC1hv0wChS8behPiW6kBOg/pUw2lsFO5t0UfdtMr
NjN7qrnlsRDb8UCk9LRrv4UW07QVCzGF8y5lsNJdqkbTCFw7Z5l4qlah9UfohLicfK31C+79B3Ai
ZJ2l7YLgg9Ml6nWJ1ilqzqsO9fuB0qq6LNybsaRLjOyk9bVHaXtsJUR6einoFULnhUQzireMR+dq
XdxrdDR5UpXkWkmLR147g7yWuEey/TeAV/BdNFdWtFMd7hnLMUdZsC0itRYypw8aqlwtGpWcjPXR
omqUu/FWuJDLDjirBdWyDqG0YUSbdR/c/EuHzx91kbhDbEBVZHzpWhsrqbF/5SecOqzrPbKxcGfr
CTd2OLYC5OvtheHL+IJHYa96TofiPZc5tGBplHy7tXgZK1sK+zBkmF4khdDpMk/Pelco3ZY48SeW
pG2HPOAhCyHNsZaPKII3gpA/7RHgTcQ2D+pP8SUWqAvsI80JmtOtWztEPM5evj4FM/4MK5ZjEQ9e
NAPB/FvGFoylVPm+WX3gfXSYyGnTYEokwkRRrE7wgcP8xlDG7fhf+BNiD2hfw0sJH+8I+Et19JAs
Ya0uJuJtmcrJaqrYBJ5TmiZbTLGrRCyNvj6fJ/rH5tON6WjfxiRG4hDpXd9JDWV0YkeCOT0JzkMO
0+JYSAiVByVhUMtQJgExqJaJPWNfOwTv1R/2ThbRahPTs9HcKvY/Y5JRr9PVlsaBKnhh45yAzrMS
tlid4IGYZPymf6BqjvtVEyUoXYUtiD+xs37kuz8jZ/xtXMXyp6WoFz4W0ia29o2+FMKtCNAGoTOt
tVLTfTSavI5oIv7qLkUxDrpwdvMQOemejm0eJtJCAuvUx5HgnMz6VDzX1zufCJcjRPT2k8AE3fTk
xjiRBNLf68TMgfdwFaJgzwwPiYZCV9EH/8HUEjctbMSHsTX+DBWsaBi8e84mfDJGD9vYqTOS3ZEF
Ga862/BGwvjXT5kIHPcVb09RG6GGoBJjwSZZY6y+ZRNXKMoUH6G8vZbjUli6f0g/0KzlOPEo1+6t
Qy0IqH0NgdVetjIZ/ruCovzY5+yThJuE8OjIWNj6Bh04EDXZMSxa7KiesmqXonkk00o45AWRFW9n
UfGKqnWBvllHm25Klm17/9ALgDnKnnswmLaIrwokPr1PHNa/+Kc8V9AKDt7zeyFRUb4xRxGQfXw3
Q8dw3bM8VQdI+yirCceiE/sF7WSGSNogOkWHkGLi9gwJjZ8U6qUqyVJARUS7IjOnl3c+h8bX30zM
x1kaW1aWFA8i6qdRMKHMC+55GDwPfp8vShqsgEJYKwUbmjqDZoZx3dTYJGttaG7VviAC1sxrQ4Ub
FE8M0GoHyMUsCQxP5ZDYJXajoSnHr5eB9no321u3Sh+VkaaZ0PimGzq7WNwLbc/JDvqypwwL1Ub5
k8hxr+NpugzKifudc3Z/tv/nLAsUwEwWp2tjVhSaXTOQqeKiMhAOL3IRTvHR5+lvTGRGbQwO4/lG
QKHiW9P64w9YN09NJbfpWfUGNAMbUUj9ysIBVHWWSwSCm/UhWCmAEgB4YRt6NgiX39If0W+DSjus
weWlj9HoUDj6u5LXBFR+RrscBQTVWsCey68I/kU1RisFExn5vtBSpkl6HGK/6UZ9Tbaf2uMEtdtR
BU1y0MeWs4e6DckDHAhbyVhY39txTgzC4nP4mXS1PERKQMuOL3evvdxQnUve72DTibgQ+CncC8CM
b38iBYdxXlk3asiXzKH1oTD6IlOfODWWSTi0D3gb6FlAtBIyKP6hL4TV5xpc8Z7gacf1uTvQIzOA
2Z1TFSt7MQI2ERn7U26x2yuAoCMa4hiqTALkd3VVbmPPb2j0LvXGh9M6x8GQY8iTcRObiSh5MIFK
K+My7UBWqOovugO83yt6aWW1I+CWru7Tq5xJ9xmAdzV79sD2Jt6dqPnfCAgUQ8Og7Kr/xR2FnEHJ
U5ErkRQ1c3xNYny3bs3axRtrQp8d63CXJEthoYJYBeltty1EzVYr42UaTlESRXUFL9IFwL+SbxiN
DMXkQXfh+KJkaFN0pXzBiGFTvuRCvP8Hy4Z5/MVImzNyd18Qd7JerNnyUI8KPjHDXQAjN2I9z8Vk
NgOJGmrCJws03idKMQoE2zP27sjyWi9fyJlWSw8Q9MZRhUL7hXtNj7ZoxfhsNqR9TGlBoeO5xf4N
00G3q0YFNA4ageoUlMKhXssTggqE0YPzNra9zbWmPp4gqOgyuvn9AWSDS2iwrfjVLeWP2np/DNFe
8l8ZZ4xVYiIk5MywPKwY30l6epUzhjfiHxxOPA0sqKJvdTSxLi6e6iHMXpRYGWQ+xwW8DVYWXa2Y
YIrC7xvoz/Uc05JOT8JP7ctlQ9doh3hBwMZXGWkz7uxERbyhIR+vD8CpDV6QJG7HQ8n127FbQ4L4
z96SQPKCcwVB4CeLv/CLyOWCyK4AAdJ8nXPwSg91HNLn1UHoCaYS/p+esTTbhAg210EJDy0eb/zU
xYnsQK7fnvM0ZN7PzX2aT5DM6ZjUmMEeDB5Hevh4YGoduKwxho26H2V9TXlFFYNx4jS3UyrtjKeX
+UowPy5OZOGtbPlLhDrohgM8xwsh8sGunZmhCA3QqzRnkRAy2JfQOoBWig8lSoB7qddoQknAtwZ5
JyUW7X/zD+QrXznyqEBI4LB2suVx8sm+KK12kakg4sCrEinfrP1Ex4zs4dTcBEa4sgGSh15WW6Hr
S5rx0FyHrkBgyBMPR5aPT647KsM/ycYj9/WbaEvRckRJstz56bbu6Qb+OF6I0MeRKkA/avMbtew8
5EPC1au/GYZKkjMLwy5cAkWqY5YUXqHW/noYmQ3tUzNLJyCpQ9oQK9FmqcBduC5Jh3bfvjjkO0qd
bUelRw1+kxgf135Bs3uU7MG7TfmY9gj/9WSYhRstaoQVw+RI/OxRoV3LPhc5gi08p5RiQzpRyJQT
X8myZ5K5+ALexYADrfbLzTWlTGeQ74++5ZzeiKE3jVcLLiPRhjzNUTU1mNVOfo0qSGixeITsgxcf
nGoPMRUHYmo+93RgigWh6IqP2lyyaFkzMK/2Sgio+uBO8YI9ZHgRhDZ3lfTldPowT9fjM0/rvDyn
EHcDCZGQS7MM6PQoSOAH1yuzXQNMsL7sCPUppQHVkHtc/C2xxOaJpsnLpm3G8/tIdNYXPdD/M9kD
EhtwGHu4BVaIlpoSNPlUUju48+dTkWXiY4KMneRSz/WUxujQMHJBI+mIByOPhwt1gDdy0qh0BaG2
CJLIcVzqpfcUncNPHY5RBVm4cVX8TZXPxc2ZhLWDijzIEgRP3rrF9r1ScndH5clU5XuW5kr8d8+H
Mzl3uw1vOGrTWPkIpSzFPU7Q1k7qwMik0kb9qNt4gWjOmO2vCARbYOWGBpEjd7GlUs0lMZVl2/RP
OTxq2n8xBSKxxuKp565losRYrj3tB4L7SPBTvkR8aw7GTNU1Uq5cxYJOw511/qxKrIffUo4XvEW1
61Uan0jwnEIc0USWa3kOoSxP//Y9q9aZixJ5lr/YEyaOulhSUMrtsxf4UBRKvmjtsVZU5qDQqpFi
IMcgE8xEHUVfltYUqJm3mYHl/Sv4lUtsjXzbbA7qjOveGbN7zTIebLw9LbGFjodikenbG4cA8y1T
gantJousBqbHfr44iNR4Q9g3Wy9FrvmJg8phjPEL+lHH1xUuK2UzhmSfN3VHEsCES6gMyNQH4DHS
/b9EJYyVemhDepxmPiUWEByrulPWccXfoCv5LYDA8XGHLvErmVNHkcyONuD5IZnw74XcwEK7d6NN
JbxT3pLYO61GTHbiX8tsnHslkq0i4sUhYX8Fam+OAAPyosB6ejKqx4hGW/FaSuzjIZaDEQPG9y7z
LQZDjmAXZcPlWHIS60fIjmB7wc2zJxQ5S7E2p6qPAkHhZUdvjBj5jZUne41D7XTBkLokiPhYJDPi
l4c0kS22EI+jcbk1Nuct5Ndj6+bqpCeNVtPzax2uE7Ps6ZFCSqC2xN8P07B8AVVJOZOwtC8p4hF3
ClFWu1tATloEW4717LAWBTIK18VEiGUzv63ha8n4IvxB0mQlRUniXRtPXmymNaeXxAQw2P2dtYjy
cK42GcmHStctdqIavHGlW9KpDtuzoGLgy+9Z8Aa2ORLYTntWtm5RvEmwgCJRmnJ4YKbPf6J79pUn
Fs8XEusU9bJyMXAO/Y7TZUhP+Ct3QD/kX/lB8gXTD3/xp2AVuatQ+QIroCL6rWWIYMh1sKQs0Q76
K6l68mtKq+l1NrpUQj7FIxrjlEr4oFal6fsfi9oIW8QuHVldeFtdW2joR7+aENEzwN+SWm4KPFcQ
N2x1nJy9rpL403+Ol3/wrlo25fIqFWR+7IlV9FeBYkexJHnwc6C3gDpC4QAafyHp1s0u6mj5ouFl
x9APj36djJGk3wd/oRMuuxnfoemLRmJnED72L1vb2JvEUgdKl0sqZOY+yPK4MjtJhtnwX4zcRRRD
ipaiVT0bbGM/pOtyZNIhblj+Zl/x8ujQfnTXktlWMHM8IEBwaLjskDsNvDEOenrUN2ljA8ZdkTP8
hZ2nfWyDJWuU3unrQ1LJXiaQwLf2Ch+BGrHFDGAjjZKsKt4+3UUXReJaj7ZCurAprMv6UJqDdyNg
fUjG3mBh6WiHR+xlz04+6cG/Q0EkVNj3m4nuolar+AYlR7taJjuf2J/DPqOyIy6pVh/oWWJAxJhR
Y0PjB0eH6auZz5go3GPs+eN1Dg4EVeFnulqBtLWvdbgbKMebbppO/Q3Gsy31+XFBMS6AJIRbMZTb
5MgfEjCSiCYuJyKGhfXULzYPtBb6pJRnxz2kHzBv4KUt6TeqwdV3lXdiaVH5mkCCXW0XdSVXF1VC
m1Wp9Snl9Yq/Ulq/i2b0A+53WeoUrcv0+VX0IrE5TiBrNN6zfC/fK62zH4ljZNVJRXoNEL2s2LEa
caez9COofAPi0cPa3nrMslxUoLIpP1uEF9sd1tAhWt9t2DOUIRL4GLWliOaSGGJ/Rj4WKFcba7eN
xrdFxh1poJ6fDk+6BDRSQyxBvxNd0jOrjQNCbpQsQtih8t+DP8t1TeoBAasj8OmyX+9xKwr5fx5h
NStMiPeMJfyRVsTxwgQ8JuOftteZVT4fDZHHKUxXR1VARshHe5Giv/F1D4i9XweQVMk4Vkc6stxt
ddGEtmmNiUJkmetQV6khDJaT9VjYjHsjz7HFp9EXA5HZJALNAjTQfbHeMJDjA08m3MAxz0USXH7u
Nc7MBJ0tYgdVtFSLQEhUkz3Jz+QiHFHPoGY3VAR4Pgb53jqXxFQyXuuwhE1fGI1bkMoCw3/7oq6R
Fy1Af/a2VjeG0l+J7tFXSP8XOB69JoEw5EAAYghIK7OG5vW+UcqE5/EvGTLx3th6uKxJ+uzQcGib
Kf0Pzb8gkV+a6tJ6UHxhbp1114zlsWlUjW6iJh8w6/ctXtCMO9v2vAtnRDLoK/SZDASm9fnX+gvO
M9toya+1J1E25tk2KQH4sQomCkuOKz6+6MpGnMhZpFOziHE9nSo0iaeSEUbKYsN0w533D+YX8EKn
1jkR6Az8IP2p7crHjt/1PrLj1EZt+pq9REk07NvsPC6e0QY1DoipW43VjqttBbobB/SNqyK0OV8q
m+piUm1EdO+Ku7BasDXfeef1/B9yM0VX9hHOnfVIUZ7oPDfZBlGpkRmFCTYlPcCQEwPcbWtahl9z
Jw1D3X4TgY4hHE9LzPvOr2tJOO/vC8HPPS5LK6/h0898293m5Vbxea2X6m2Lq2buiLr7SKm2mJIs
quyVhIuRxBz+f+jGb9m+cZWYzkes51b8PcXQAawuQNCq+Ka1gE+zDaSiHXPWRIUJ2r8eUYZvfQ0f
y+ynGifYWPFsDWZyqTrse8DoEU5fCgipBYtvH6o7gCERTbGA07CVXG7Amkm6hCcvOqxmtmSfHgD4
YJ+Zc6ulr4PmpBXK9f36EJfrfrGO24bMK1H/U0LTi2qq91cdtNePXP7IPfdZCsUvnNvn2ir+wEmm
QS/SpgXSAnMDN1EmuDLvWc1xckKA4BdBoAqTe/ivTey+JTtoduVaXADaxs83tEbuuW9l6oHexcOR
JldRDrzwkKR1Dfs7mRityWIWhUw2mqVDiwdpYzhmPN4PswwTdxjqjK/FWv1H91Ukv/kPiXxMO7wK
NhiiZJfnBt/Vq1xxMF7/BA7AWcdiqfnB+fRi6KvQ4wcsW0xZ4mknmFkvVKRDvrDAM+KWgf8sNnyo
ybW8SxrcRqUuXYidll9+hH+dBzupBR6V2FOSimRU8z6XZS88weGC+rd0woMSQsEKyLRyUaD+DtLB
VTAV5XiH3H7ipd+1Ffd0m6gfxEtV5KlIu9pmbc7rqKEvqQLFQkan3vjNaDdwhpIUyFpcEIsM2wjJ
XGom7eGcqmCV3M7OwXKxA0RpmuWJNx+jw741rfgGDJvwQfm7yZ8ZE6PslZYVWGHJooIpGbtCfYzb
ErhzuIpqhIfO+iPUSCWN+nHkmBh8QiG5OCISGv4FxjPPuSWQtd/Ka0X2bXkRaYizQnrBNfEGkjNB
oUqqomex+ch4Yr6ZnnnErFVn5hxFssZI+O8Rvp+A9Xg4iGhH0Xaj6JdQaL3bGejKkJHoEXSTTZJ3
SJ8fdLKUu++mAST19BWOR7kSovZzQcN/PAqmaDPH5+XxqvlfqVNVVe60HBmb18boxbC/iQgr6iz7
4/bXUkFwKBEqJG8n9aNh/pSEU4MS61WFVmfkZxaVQvtCmlmFCe21DLs6AJhNxDi/Uj6ual4mK72p
uwYbvC/UZNZu/fJrSZSxJyjNEMJlZXs9b/Ur1QuI9dMnns/b+pG95U01iSLkdUYM78vxtIFGG9DF
4Jnv12SiEjg2Vni7WAlCKBgYoJ7HKHsrwqw5BI0g1PEIIqlQw9Yp9e1wgXr1jxMHoMo2t8wSfioP
XFxdRKt/KrxNz6u2hZXUdpK7aPlmlczq8sEyJXkM5NWbrS1bvP+eTDO/2orbxM84xc2NOkQgEamK
h+OdCc69nEwp3NfH0np5iKvgq2wW6uLdFN7okv4q8yMxw11xHun4b3mpf5YEvNRkpf/LVxPFkx9f
BFJ0e9aR9p/ELN39NjSrtxeqXBMSFoYYxGkb39ERpR++8DnHA2Jw1h2NNd0Mr2YCBhoZGcWFjgJ5
hkRkVYqURNYEgkFgqnHb2jAwk2sccNwyheo8qPhjIDKL59BrgVKjP4YuPovYmPmkPap3AZ+LZ+BP
JR7VzbOFAVFxkhMTXC3DosNgVv7lkqE1KTSXO5FgeaioQvzN3x6bw0Dxp1Ir7yNA1d+kFi0Z9LZ0
LbVzVgwC+zUlq0AFv/I53Ctepc3jbBlH3hJual/PSebHdlZ/2Fz07clVbddjQ9wZuSQYbu/i6WRH
2mNxtEilH6/Xa85w401oE0D11Vqvl/SM7NaX9P3Gbi/T9ywIyoQdnBkcuoRCzEgJTHflVtLsYZDN
0amvwoz5n18GEtv+ymDS1ryV5YbjO+GQHm36T1F/Gtch2GEoAvST0wGJAo1NdxQSNx8YI3cPfzbO
KpzLJVZ0IkThtuNhXeXZRTsychymn8X8OCENuoegAdqvD8yEXkMLrPo0l/S8OoGHVcE4ux1A37QU
kiXrmeAuGC4SGIslG/rxYCkIoLN8pwCWpiDcXe/9+OekSdlQg3sDHsVTRhL70WMi8ib4g/ZHE61q
qdsLn9JwwICKM96HyGZsBxN5t2sKAguR1kMlNioHUKXSS91x5zKZqPHAawSiDmGyItYPAfW8fB++
fFtkFSjI/x4/PzyrU/H9fL4Wh0DsOxlpY1m9usctlNUlBBh3wM3BHb5WaIIrUQ+TtG92Wi1p0a+K
+vhHP0RPgnEu3Pp9o7mV6Mxq2BEtWNT6mGvWuC097+coPdOQ4JjxkjI5RGqiIitr2/0gw4B/urK3
ZLklo5Wy63fTStY0tYTpOueziRpYlZtnOF7qlidhvzo3yMggcTm2SkPMFWGE8xLU2FjOuviqH/25
scuSi1u60scuqy7IDBbWNLHgwIK15N/aptW8oMRywF+znrayV2UHAS2oi1Hdec4f9xTBIiDDkdld
t6q6VqC3UbwqcpCzoTfv3S+1BnJv4SUzFuVLgTf0IoamzOie0QQ4it/7o51LMrIeZow9p4pa3B5D
jqYdFGQ4maeYj9EwdU10T7bTV7pNZuyyO0GfeSbNsFzY4qmiD+rYHDZjORvSYyMF01l9FTt8vcDl
GnznzDOgFz+piGzZstyHjoXM1x9Tw/r6p83LYwWenNqKmwHbRhV51uZ0vPfI53JEL7CTTGUVdsoE
rreFtg9C61hquj+DyCS8S0zRxjiEtqiHsBXtZmRvJoJOcFAOhyAxTrG3sdWMfhqBGYp6bCGuBQbT
tQQEQwWgazBVFlv48dxQp11EMUzCbZizp64NamxtZBKc0EaKF9VRUXQB1U7DakRAYBGJCBQMzVCs
Mtakc84L9RPgPRdcamRb9nA/adowiCbNSAP97mA2zJKKGkBielU95oRa1YFzUOQsQuyKpwWRYmd/
6GYkU8MzGb74l1xs1Rm4dfnJ9Nr3AmPOGIiZkHJN5wq/KL0CF352qydT7DoIVH+CLq+GsNYaeX/h
54mkwCI9z8aooIMGppIOcvZwPfsRUoSsZRIUyZ5+50XsLNVGNDqUNaU055TAMdkoywBkg+XmEC1K
GuJB3nSk1iWDfVFl5KmElONnHtH8zDiaQ1kbyngGbGNsezP/E895DfXznLRH94abpi1CTqW4Hq+z
7WS1vZOgvGif9Ln/OAHu0a1dt6rUh4i12QVU3YA1P2q1I4lBNItB8ioW0JT0EWodv8A7e0qYftr7
D2sdckJb2J7VLPcLzorI+IgtJXZNqQ8WCWNkEU3ZkmOZognVk27rpnRiZkiq9JRJSH9rWjWEFS8a
E0XIGNxKRXGXSt0eDTrcZyjSp8Awrg9pntvfgoqT5ZBxpL1SC2gRuqbPOcN3PZBqc+UORK0UqB0Q
n6wMZMmldeCGeiDRWk18C/GvBsPLezc/f0uUkNTgOuK29zBuYE4nCtTkprqvjxL3UvStxmtncAYq
SdsK8jXwpc3E64673HWvTOCahxRAIS+JyALkH/9HkZSjpbggfI/x0Qg/9ZU6kkq3LMYLNnD+T9YC
DqVZKg2s9ixhU6/0Cq/DVsFt19t56OFM1kKuR3pfJnq7Ir4KOOPcWuXxGuuUU9rzqItYLXgpfHe6
yxNoeJArJ/ikUMr9TqR+SfJj01b5AeVzzA8SgrFyWgEk3wZBKiBzvhHQy+UrGD5lT7XRCjlqialP
B48JTXDYLN5tUWkNd6kYiJVzJ3qBs//5TaRHgrEsLEOMGUi/afizG4cdaMnOccZvDOIeI0+HV7fA
ZX1sul7vIFgeXhlTaatP1YFqxx53TPO3E4Ln8b4etMHG6aq+21j5xlZ0b1saoHGVFgYbg3KkiqvJ
yeiiiIuEWL+4jehFabkZgHcQHf2GQ0KVSWUWmNftJk2FZEpd3wd2KEhMZTHIKBRLXcxV0jM1rdwh
wEPNEAVf7xrJ12iSd18nDKKwpjy2CqeQFNAzQHqxbjdtoE7jPyJZ5nAzxBElgNBqZZK91k0fNOwo
3ymX7dhgIn8U8mNUHIXd77ApJjfIujz5owePdj2Utz4NvhGrWcI/6K/CQFVKmyGMMDPAvbTy+9gR
rJWRSXgaZb+oa6D5WKzEA800Fl7OxPv5hTfsjnH3JYlIJ1QsVEbHdBVT3NvnDk2MdKDp5Trdjvet
Qd9fEJWal7Bug/6rT85RupZcOxqiJzCrFs+skUu2kQxRLeTEdA3cJ5IQKmKc40yDckzloXr6Yr+h
rx+1xVLD9JkqeAB4b7C5ebbkQdRy5DS8FCjs5maKwprstQa60gdDZa2fx57VY5cGscl99C51vji7
ATCidGQkHj9vf6laaf7Jd4Fa5ZPbYnfWoDink/6mmiSpSdnjs8uFa6JvcEB4gCvEDFQNqEQV6BAd
ML4WlmEIF1InEjsf8m432Oc0muTiFc3eLMZcpPiP8nTy5N+5Trz6hWChi7+xfd5yX179Qgr4+y0H
Zd482sN7lEBy+n/f+HugdLhSsxT2ygg+g9V8fxYb0ZaOlK+M09V0ou/PavVa3+BJJMbFezsY3c1d
RdoHehsLoJun8kdy14j+vTGhHp4wdnPaIZc1zFHzdpiGDwslDVhE3wz/FYOUTP/UV+2S487lNmnr
yN1n4LDXp/R7VpMECIpOcdU+RPrl/sdyH/foeWp9nP4GcjWCHXSSp1YtGkoKsA8SXXgvgTpFT6MG
5qou0tODECc4XDcdw8ACTwamsIpfsRAtKSTxk4Od9CRfmDEHHvizzugxGECaNhCTZQyffVoqDVxe
tKsT0wkNRDKy9u1SAbt/RlHRKkMxdZ40+DmDucbkEfXEZAfqgMQRX7GA9SMwF8cRA2WDlk29ZmMq
b/9UJbzR9Q/IIirs3yB2/4uSDAGg9tC2n+AyoM105KRC7TWe4fYWmBfBcHcBi5DxVeED3hMB4iED
VssSB/FLYWoIN/Y56IT6e8Q8S8h9frRgY03JMzrjqWUGQLMrLchlUkNrZxDE7NZJjYEiiGOKSXW+
BFLnBv+BZBUOl0esSbd9gJEkiwWihj7vgOTGzIRXPkeFhd99yUbTvEJFIkt2b5uiDlAWyyVztTrT
NGt18kbpWNhzPww0gpKWfJYGqdE5GWK1ZrOTtUtNCklCKsduiPyrvdnoFm5wC44FmMRuEmXjX0rF
U4KNVUdqEwl9sNkU319jvCBMjuTGMZ717pZTJ6mLBeU5AGP9XA96hnLLgw5uJBtomTnZ9w//TH76
qckuz2oDJmuEJY7G9LNSGDz4Q0HB0PJ/Ucou9JFeeOAXmGsRWMBn6KQMAbO7zVkjMXReVDGWK2rz
Zt2ZOKU8R6ruTKBV2PCAtjqvO0G9dz/qYLl5cT9JdocqiKlm11778zfJ+o3d3Seju7Og075Y6AS8
xZ/eEBhkwVkOo+GsNsMv6WxbDoyfZ+iQEw+NbTnr6dLezUv8VUkvmIcmiuPsq7tiRWGGv+dUKWTY
4bqGlfhUGsQHWIksKqLw+9cynajNcNuyXbCuxIIXxneX5GOWJCwdFvWd+2uO0h/4gnTRJyO3CXPn
8fLaL+4yAned8hVL4Kcr+ZGzXm3Soklfjvbmirp4rCnxgt/+g/ynsDJHWVdhLw4+N39FI4ggTulr
yKRlTaO1NpcV1KuHDYKPVDiAkdwUJl7jZUQWJDUzSsQsWsGH1nDNWw+m++KL7g6J/NVmzH8MJx2F
AEkO6XuJuFvEXrItfgIOWyGiEQhALC0o2i0mFDGOjfacouG3HtCndY9aQMUhgXdIDJlf7wvw1aJ8
9vhPX8/PY65EcPzvj5HccUeh5Ouf2f3jEl3uBoWZ+DbdNXBwvxQSBcHg/A+pL6QN/kS0UEYFGjw6
Q/qzbErLr9SJcfkIe1ciG0CzhW0rnd0hCNdHp9AhIsoEOFFMp/j1u90VdHwvePzFgTCyHj4sLspT
hbImCTXEvG4yIWV9/Xb1UbI1JGSxK8ieA062cC15uBhob3U3JPaxVf9oQFGVLSyIbcfSespxeleV
Tf6h2m/FFR6NueaPIs6sXwoLWHtJUGjMWJXr2JM9PZcqUt3uFqlVeDMAAH4S56Etv8NmUTrov8UL
+xu92Vcs/EZv2ZQvuxOocf9b9bYsekgk4I33EGjFv9JSLYBi1b1BkaRY4M+E9SpthPsD5lGkEKKi
V3WAcXk7plzQ0hy7rOwCbEfZBkms0fPZOV1e68R2giTTAIeKR+LBGOuJH04EybFJYH2QRljX3uLY
pNSyzUnfhCOeOw32yP5DBF/YvQxSs0P4HA08PCeOq3g/alS43+Pnz3M/ldbslCBiC2E5pDOiAhQ5
CA42sGiy5ZnxNoWRgmidQPDtn89Z0OhsE1/s/fBM0axky9Q1F5YKAiB3n+nNzMhuVy358fLcZQA2
Vek/4rRr1Rsrj69TO4pdd/dTe21DaQsGjZRlK0CBMw5xueoJdfpHUlNa2WsNN0aNshtcnWyVr6z3
ij+DwsY58BqKI+CXyd/Se7SMftduLMgf6/s9yvme26R4k+AtVxC0nO1wwXyTLca6P1VNNq070Gin
M3RB7r9CRM46U5bxd19qHr8lykH3j/5qnNxqUYTriQ1W+2PZxSGl77GxSYkTESaWlHbaqJSkO7ut
CnIRkAb3ZPvLULWE9lTHsHdXdzq2P62XFSc20CBykliKK8FvA19RL2eCG5vIMxF7QeRxJ6cx/YWk
47MraMZ7Tygkc7XuqYDSykddwGqe9BHZsnMISr+0GaMSPq3LsADPAVrzZ0D1g/hX8+oBy3k4gDk8
Iiz3Xj1BzLqRnXPSZyH7M9UY4DDjBrfBUSTGjMYb+C3Q+dBXQqrQpIiw6JTYXDLRB4VyW7K8cpgc
IxwhaA2KpDL2ASUGNz2//i5IoM+eMjSX0Br+DkTYb/2H+Tir6E12eS5zy1BBTCY/gy9AXkOEloOJ
YcF0/64nka9t99rUFzYI40MoWlCYIkq6ZB4Y/MhuIDZ/GncAn2B2oMI9AmpeuJHTu6uJuapa77Xh
YI2v+TEA/2vKchvcmpLwsoOy1c3WrXtAOz/f0kZkNxPAqx06tAkY1oPCiQNtZ9ryNvAm/HTLN2/1
Kkkc8TY3DT+cxRkYSrrEaYAWg1jXs09lqj41z/1UB1DHwVFSIPv7FaBi2CezCqdwE+cwTKdaPdra
8rkf0j/HNZNILo8eCSV4a6zhE9qaFxAB5uACtJ8hwZeMT0cQQZQ8FFPlV7HbPOYJJ7MfnBbRKc9t
C7Z1hC/c6DK07OlFXnQZSg+j3ZY22lM5bGSto1LfBDpw1M4jzJNr2XkA3AYN+WSpZuvBwdN965lp
9JsyMaozlO5DuhDofMtOV40kdk6jFS86vMyaDI3sLKfiUJaS+jA/mnEsjmlMPhPRDx7GxAv9Zezh
I7Ow/rmD90Hd+ngVaKDZw2NiJrrBenJjnQl37SmyB1uKdoRDz/BfuNP+teamEl8k/t78CAPJQ5xT
YNhv2TRgIeSHzH0EDxEdoxpuFerD9hMg3/KDoOCYeoXt/T6Zcelzgsc1+1Ip1w+Is9/DEF/Dpr8K
U6KPsPZ+rzVImd3COGdtQlDsyhvlHwHtJFWGKV+TqekxKgKdFjtv+9U9M5lwusbVUOgmbPRvloNo
CRH0VJNkNfivMBdeLLO7ehf8LmPHVoN25+n29KknJC3cO+mlz+eq8rlOuY5TatIOUg9XlpESSf6f
1r8nuwHYU51SS8RRcwFpNu7eQPB3Fj/tNFslMYs/zTZbjdp4dydAVD/LtqH3h2ogEATseSO9C5+/
GVqdfhBBYw9eHO3adRL1JM6W0/ujHEIgYhfQ/4nO+fIG5meatXUM9aEYxwQYx3UZq7tD6yoqzPsk
Oz+9JOm5NuAF0P5qCDYMd0p3UGituE1/fmqfDlIDQGGTsW6lFn7OcXo/YFMBEEIl7dbRlJcPIaiK
M4JbId8xy1/DmM0TU/ZvcR3qzmLPCoMHtaP9B/ksPO++dG1cHXW0C3xnCglhy0a/N6cfpR7bUvLJ
rLKFFs6cqOd5mlaGqVvsKViDjwb74rGb1MMSfcba+7oz91o04RP0O01S8fWKHOOjapGd3fXrt1Ib
4Wu2/yV2rCn3Oo/EKqJOJf/MwU09KAlq93Wnr+w9frTZodDNVVl4XvsxV3vE6oPwcDPWAcdQKVTr
hdaC7NvABxzaENzPqQI6000j3X468IwD+z2vIyn1bNoDz9MVUiSytYLHz+3Q3bC6tTUh4nUzF0g3
J4OsQBKu086a21gn1pH2/A9tMnUiIcYGUxUPBw6dV1OdEjHzT8TYVzOp+HQgnEGggGuR5BDn1s3M
YmKDEIVnV423PXjgq8JoAMBEJKEjcW2kN2/a+DCR3MMtR1JI/W/lZQ/RKk0XYFlOA8wkCRyAu7rP
6P8bwzgbQVV6CcARYC9H4iglzJNQXth1yVS0neh8pDBzxcVzGGwMSbd63/cBsYOYiC4BRbZ27kZm
g2DkHQ0odWMNgUfjSO8uwV9krq3L4zqcltuZ3tqwQjzXS9/h/MnaEd2XmCtBepkXNn3GPKTqoXhK
UelZFyW/eK/EyHYF408dN+2Swz0O9Ma9Yz610/E/8Ye4fy57nrXxTIFApZxxO9SDzFyuntCEIkmR
SS15Dwq8kPjxUGzipVenu3E9Km08RO6x3vlyG5t3nqq/rkElU1ETP8M/XaaODgWBnvTGZj4a1GXs
BDkJy2yBtPjceYITN/NqOxMWJDbbgeVwDiyWGwLWIYLRI9xz1hYmhAUz+tBK/PwVwvX5qauhhbw0
eZNiPi4akTWlj6vFOX2J2Ttgyb8rvjpFDSS9Qs4Lqn+YxU+/EfaEfLyvUB9ainUMPVIQ9xA3GD2i
Prrb5Qw3TRA16Y+n0ec/xgv4+63dnR19jJPU0iwokKLKyeIFN7fr4M/Vl9l8A20zIZebN21q9y7i
DTVEJX1YIMWtnUhe4WQXKt9y7OaFn++jeyE2dK3pM2ZyRdy56G/tOqaHo/v1Ov6UtN/8r9lqyMDf
fwkoUtkL8uPgqHn8EKlF28DIypWarRjTPrW5AIErgAmMSwOHp6xHjvpvzjYAJ1A8Q8DX+7Sk8vOy
WnFNPh2uHH4pdWeK8THiHyEWu3/yjDk1/MDneK2b+qpQqH1mzyTdapsMjcIfMHVZ/r6ze+eHdKi9
6dft+UhrSSUBerL5QjBYAx3YmWCrSWPWjWDx8Ns4jZYHnQM/aCAInur9oPKHbw0dpMY8QSB9Gbos
4Mw+0Sd920Rgf8lIUVrRGFeYdXRjt6E8wzU8q+pwVI/vuK0WakbKnixWi8aSig5zb4bBd/ZOOZBH
9IqROuLPj0c1mEUA6YEzYuMWCF9Remsvq5Qnfyoxug2lls7UXoIvs4boGoh/qCP1SG5aJCwlzi8h
SJLcNhdEF5Tab8nYPcepZoCg6TP1u1OgSqIoLxK46uksCu8zaE2CBlHna5YApo/l4oKgEARlgpqe
Sgfmmf/eZrklOThXel6+fpHjMdIn7L62MDjkHjlMVCD487vORx1Rmx1Y6zbsl/mGRoEcMAXCdeNS
Ck572jdbBKrfwBjN6EAx1AljzKr1Pk8Vlj06HRNTDccbW5Wz/heiqqw7yRj2hn8rF0RJUvglatGU
ZA8MrBW4bNkuMlrt7jNQydn5E9Xne/lLcPt/DSAD54YPtreccdbSSSacbQ1Pe7pgeLT6QlQTFxEo
lSQ1TyUzBI0laq1HVUNwyVfzitrgykepdM4rJ9qpFu8tJWHL0JeWnz+0Bc12BRH37Qik9WGQ5E7j
wuX/t16BjxotPUFiYC0baIW43gDtLHPyKGgEvvNyngcfFlFWup56O4JpwcpfsrjxJ16G/SOn8rU3
z0x37gDTIa11fh99KpGUcC0jAbmAHLwQNtSTMTsmO3oCjs83TcF+h9TRVJ6TyRitsuZy4vGdG8x2
b/86czE99pPB8NDGF7BNaKiaIaGjDcGE1bUxAspREUwP0uo0P4MBwBi+7OZf8QEw4Cmj9NOo5S5T
volMxJ9wvlNEMnCx5akvNzIWd+Abrxqo3062q+T4C3laeQekTXKuUvLrbne+geeM33QeoHWWBsFh
Nw7x8Hau9D/h1iI40KSSMFXf1GJld1pLo8H4xhT3wyMuReMw/nGZyG6Gl0DKw6p0m1S0USoYP6Eb
csaiwKHGuC0jXJ8kpY8LA37SXhJikp8X6r8YRSAIxA2s7d5eeJVt8GrqqdOHprFJNgH7osDefuUc
pohacczAb4m9FCeGXRKhMSnVEz5g5rjNiTNdufbznkqGSq+qgonb5/IB524NibgUcgEvlDcEEiAa
F750iGwSupPEiK1+Pc+lzlAZ669aOLA6Ol6HrBLojAOcchAtjB8pCnQYT+90YalrdEXdtQQjATxt
H1R8KLuPZPutOaFJ4fsgEJHz8aviD13BioHjB0cfTg2v+/M3FnXR8QJk3WFQd/5MU20aGiqMB8vb
MjNzUq5TVWdcPyKGuOitHSsADPl7krrW3f0HX8D8VBcNegDZ/Eozv7o5yiTflkh09zZJ2ncJslRw
OqXMc3wtBzjOAJkswjHNO875OvmKuN4rpVbrIOjVJ7Fl5eUfX9C1jkJk/I92QtESsp1M6N6+n2kG
ttbhJo1kORJex33LWXi22h9eUBQDACPyMTl3GcT/EgJdqzl9rBKwlGJKRQZhPNpTEHgRykqe115o
hmv8wXgoRZs3TR4D6kM7tRYYPWUCHWzWb/6JVjJdDSdIHHFWuJOLczZWASMGRFXC6zzbaJXl6nUc
2oAFoC0PZ2fPY0cGIq64cxUjjeWvG+DZJV8Fs0vXrM8xVFiQQJPVFtdgri0IyV501OhiVi8Bj0CW
Src6XdArNMBHi2GA20m7CUNAVf4Y8jpvmBQ1RoWfRhIqe9NRPYVbJ5wltJOd2uWKySDi/76R9RAa
tsaxqMHfr6dm2uIpHTaamuQT75xtU34TomeXmWjvyLCAYv7owvWiGI2eOozrfy0Y50psRmvAETWy
TdMoU3iAK0GXOsJwwGHhMJNULgnkioJ+eQ1gNXkRz3N7iMSyEmWAmc537O6/w4xk/7V38AVlQQuk
1t1Z5ysqHH04aLsQOUA2blUV4hbS+T6PvqQqaAcJGDObe8qMLead7Sl9/BSt4PzzftPW7mWQe2Gv
KpLHgVjh0O2GuraTHQaTaZXspgTLlVcPu/idE5UDB9QuRjleV7dpGAxhKJvk4Pmw0DlVN8w35kCh
BE09Y+BQnCclye0sq7TURYrzvbX9oZslHtmXN7dAONIClhZ0zJN7EH+yNSAr4CrJ8f/j7xRjWSI6
GDCQ7B8g+wk4Q17rHIjc00UPVEdnFBjBMaZiefxMC/JlYCsOCC+ALaVHvQzpnceRAfUuyr6AjV+w
qLFkaaB/mBeIy15YpdWgok6MAgrW4BrumNxgPkP43VbJ860heODrvklGzHU2ZbE8Pq7ANSnD/2Qq
V5BgXc1jhsGxkW+X+Rp6GYK9MCycz9jGkZPwdtUppr2/kC6ueA8M+sXUiZoPpRnQjhBVMvQ5L227
K25pmbnPGNNx8OANSeMu9xAuh0hZnUnpGl6g/0FNBIVFPXnw2Mn2lOGjBojQHBKujjgNkuqKSyft
OGpRv/1xW0g7zhxORiF9eXtPJz9nXIqrVsgibVb6rrFrOyLtlKyurxQHModXOl3lMi4qZflYa9+y
jgZFTPgWRccdO7hyZnWv8MKVb1ncIavFHNbCbphcEOcqdBQmW/+MZ4XxdXfeicbb6auqHvKAk5rG
kvbVX1Gy8trgKofWivdvpDqBPqZrXF0MK4uUt/ogb8drRqfB9t/Zbn+oBdoeBB764ADwKHBeQpw9
gId2gc+pFS67lAEZ7WnkmbNuSmvgxAuFucgkiFHoMGz80hq22dGqaJqB4xXfAPQgOhlETR1hqx/E
0zN96C/NQdPdvmJoJcqhiZkMlbHTqLCkFMNtAvHV6cfgSVCzk0wNEZ+or+vPRKZqvKQmHa6/0Pg8
a6f/jynE6mGbpFOgN9Y5GNftH66/0xl89g87nm/XTm5uIwUiKjX/8Dns35SS4daPquqzpfybxB6R
qzXRpgLrcVZ85/8z0e535+Pftes0PEJaH5exwKsyGOuxLHwYV1fI/7uChpDLYS90iFMT33IOCZMs
0Kg0l2Kc5ZTMspndkxeZapzPtZnFVaWebWv0LptM+29MKC87PdqemfgDi3pB0D7hycPaMg3XVbUA
j7RthJRnzdzXj/cmlUVEvU0qjntHMYzLYHO8qtMHPyt7qjlTK/nBAvEdJQs4MLG/DJg5+2rp8CeX
87h35V0FpyK/V4HewaKWv1Gub3Hz2ExL77iC9QhZqNZQpj9sYEDoeBJHRxHdVbPGqlkDNwfO3Uua
hBNsuq4b3qB772FDc9QAwKPjO1Oxa87C++zThRy7Koi49I3RfuOSZycLevl/F/utIWiWw2/YbMWB
6ukl6Jv/5JasYCtERSB3yesROTKDfpGFDsBCzVy7JDAX17Kl7wFtv2t3SKeM/rMPEL1Giq3X1/K9
mhEmtiUHOjBW/Jtb3VIGBSnZzoLB7SSmKsaVz4gShZ3NCc9cWLAaffUQpGn/ZCUlGYYXkdpaj8NC
jroaxHxmMznhGIfrRv3ngepM3wNP73fNuDfV13O+/1EcCn80ABWhnnkxHS+t/apJXkD4K32nEeRd
exiXWnFlSdV2UMYeqHk6wUokOUv6hjuWmDHwIw/KTXhg/uJTOXDhq6KucCKkrK6AFMeW/rYD007t
OBK2pXjNh4EFihSVqo2TdKlrNBy4gz2siG6eVWjtM4a3K3gWvW4mrgKXhSAW9NgCagbuLaoKeJv4
v7pOEgvRmpFGdcsuOnP/7V6Uk9dSmA1p6hD4hJ2zrAo8Wga9F3NAsne6gakONn7YRPgZ2xl21VC1
Rd0CH0fZajgg3xScEHT1QEypTQYOC9FyOOlumGdPC9peOJIwDr+QelP88ecl5ekXemNcAOSMyMxF
6TQHcZdRbxHt6jOFkFIufhM4g5PDKOknuXCUykpWxLkpR/CypXmWqtq3r53eNCoYcsoRuXUqduvL
inABlJuRJr4lnzeV9nPJ/NUvpYOM5qyV2twSTjsk/W0mqbsSY2FD0UrouH/jfkz1fORTLEqk4gBl
v8YiAgODpoKV815pFu352OG/XFdqSoKeT6F9LwNSQslk7kPbhmxzLLXqXKBN5KCIKwsMDLIz3txH
c7S6f1eZYP0cpMsCU7B+0Btq155lEf0GajEDzxpNxyRkl95sv4co5kKJCqub8FejfmYA2v7+kzX8
WTbeCi79szkaJxg3uqNBrKGcDfm1rL/LvQnFsQOFUxD7XPavaM+U9MTuMJELTUNUjSTptLlYCeoy
QSJ/PeLhTE95Pg4+ciVu//EaRzDpyPeYvu8SyRpiK8Mh49XgGl9KVKv2kq0aVlyzety6BJdS109t
q7txEKvwuO9NTTdDkuIopUtQGLCK+Jw5kPwljqiNBgoouTQjqwC6TMH8v0bS3CGKXkoiAjDdH48k
45JX4wNC9vij3ESY0R2bH0kYupoHfyulyPVDom+MRlBHeFZ7bF3Ay+OwKq+IYfRcbbtw3yLXXx1d
6U61hTeeGNphWWyaSoOXKZchi2yX5cobGYql++L2BHJexmRgIzIl1fhxVkTHERCF4KZzUoal7MF+
9Qht9s14z/Z9r24I173X2W3Ae2nXisy96DYnrPC3QPZ1UsRXqpV+6JBG3cU5uIDqwrzhYV/0slVJ
JRYcZBDfQUnAhMCVrGg5n7h+Zm9EiHUvqrtZKUL21LawYqJf+9di16yG4Uk3js286fLGdS+mdSIy
W3uF4U84AFYxf3mEQB1va3onb/5e5A6fpbkyMznlW8lz1JQCiNYBZo1JEAACLsF9/MRkQ6UBT5bG
9AC8CBRhkTtfYignrftG/6YBeMZbJL3pd+udtlVOC7mDkLTZxF5trgooGStmbbDBbkgA2tvJh3Kv
knX7GphXdZcVgAX+awspX6AE7v7CxhfIqltnDCpYs/gUeho285Vf5udmHE1eis/jj/hGMuf5MHCf
VssE78iRgk1tKvwQD08RX1BRrDJuJ4VYiw3bbgLDGcW27oCmXKgNCzf9y910cZvZc0H2iGw1bydv
+mrIRKADoHXcFckLgmD9NnDCwgqi7/ujM6SAnlBgMwL1E+xdmMbHtA0OI/Pys56xLLGzhxijfM9Z
3DYTBMweqgUeQA26YxfYMHjF9SWshZ1taHJySDG9PI3RZORK1S1qR6T3lnPVi0WvqYuE9VARIyX9
HGQM6Y+5G2v7zlGoRcTv10HA3fyAf8XCcdjmG9b9wUjg15aDYqX9ACIVZsbA0qR4u3UAnubFHavS
djV2DogcDZ2rkd7j1K58xyt7Hu0nve7KKpIPKMYeH7j4giwYpxSexxtOvFME9d0PiSKbuvQ/FJA2
6Y1Vi75Bu+i+n7SfngEMaL9hxQ2Vp0vdi05WMlLCi6m3GnLHyBfLsI5JKzkx9joeuOhSD4sKtNp/
54ohcK+1/nbNgHUbx023Oq8yQBlkNgGuQG4it1ZFxFSrwatpOQb3c9NhhEfNLaO4NAwW31S6W9Hf
r2A682PHViVGTabprFhNnV/848wshAqw3fD4H7IHajky3DSAIe8lmUsyirRg7hsQ4s1LIvh9v/Z4
na1PvIjsWEIx7dFyBSq9eIxuPZW8pPRcSqTJnxX0PEtoswHHSdxMKkKnW7S4stg8/VK1HAkYBPeX
6STawQsM4qMOjxdjNVyHP9CaIaDJ5Vd5YRrQ3vB15tR0YI/zqZ/gtB1AfY2UGABj5CgdZt1V/nNP
lTtjuQK04gVZ/aawhjlnvtlCSwlgqgIm2SfSrHQ+KtDUYsmNO19+q3jVg2D06CpKP7MuHDPVY5dJ
J/LyrNBwOI0F730iodwCfuFTN+TN8CWueMt3jFfMXEavVREMgB2yMPfRZL0WvKJf+KiapffxH37N
+nsgs3ySdY6uoXagf0cJkJN49QBngJyjoVhVnqGCk9vptgigsWWy/twEZq6QExFmmsHmzpVL6DPh
kZpvwSAnf9Jzm71Cj8m/0LW8hFsuwpAmE3a8rve0GfLq3Be4WQIorKyfnpoN5NtrZpt06YyhOsAE
irmaLNadNeA+P100pvDnq82b2JIwzwaC/xKOO0mgO+SmEQOHfJ11HfyZDo+9eWcfKJfKy0QVZZWj
iGY2GVBqkCgW2sZP8NrGxCYAh/AS96Yv1vlQCbAOK+Czy1gyskFKjaA+tV+0BzPvQlFAKsNIf1AN
obLrJLSApRQU1dC8G2rgdxp9qxtmSYXOvjYuBMunWLV0UTvqXjE4gNCLiTrcTVWXpUxkSMhZHAoZ
tijjzBAMtCiFf26elN5iYnIIuaqEIp7h8GwQXWwO8ofwYaE9Z9hvsvkuVEw1n3/0rjIrhYj9hXo7
mLtnGjmfAmpLYEA8ivn+H5wJbQnKnW+xOy6aCDlLMNsyNDcBRorC7jLG/eVTiuDyBKjLh9FCDblj
clEmuzO6qTw204kN2tOH34FH/45HQ8oYkeIS7RnSr4mP5d6Z6NUhJrabcg9zyacnRe3TLc4X3SVd
/LGRPQI9zpVycWEe83XRXh788M28LPe0SJIXLvEgUDKffqJHtL6zqhP5lrXp8IU0XCu6XhVXEZnp
EKVAG2IqpWl8W51a/n3DYoMWcK/l95S9ktyrMJIikoAFhiJphdMK51q0P3XPDqQXfu0nSe/jdvRN
SCeNIdniZCx83nQkVGXx35B13S1dNpQCImmF1pgy12wZM5CQfqF4qt1XJTMkGq9fCnpI44xBvnEP
f1FHqDSgKSCiMm1Vuo72S2iEp6C8ZWDeaj53zFHE910Q/jb3Iqr0H/JN/XGW94DPjgcBkxxrDlpp
LCvkJg/rv0gTtekMnX+1M1YVgO8mHPLBCPbhZSPYooGc/0QB6yEZ2wIA7Gv6kNqxVfT5uXnMjJK0
gyhXNvFJAULCsCxqmmAX+GLUq1YcXSrprw7FoKLYA+/PJvpzIyVgPjCsb6d0UU80YaGq1T1/LzpH
dQsuTefk6UOaWq1hUstvL1b0AzM5+tTKjDwxxGgKUQrBPjaOCVGMwvczmUta/SCyPyKIhXxg1zGw
wIHe+JqKYVhx4ljER8jMGSBgSUFRFVms/iTPX9uVmVWSqtyIRnTcLkcnLxhYvBh4XP2fWrQTct4n
n9HKixWeMppd1hOC0r2nw4kw8+piR+iTLX6o6kxBvITix0WghM96Ud898VxQaHlt6hJOX+bNgL/R
wE+u26WU2RhIvjsc4c4gzzIM1tyylunESLrfwzgNSkLaeQd2dXwRn6CK1kKQ0wj21yANAmAQ3Wz0
VyOVClrdfdQsjBEWyocxggullHwxCbrQ2TM7qRQQ3+Gisk3tRy9jYpQvlJqmTq4zi0WyU2gSDc2i
Hde45qGJpsAaUxyJdCSuhGhUW3MuwJU5N51c2Npmnxdfx3P1HlgKgIGVsXVBtKeB7P9swT0k3SOx
1l8XTOve0OBAvMaF1w10shibV1cYpIV3l8Zdd4aP46eKeAwogvQm+NUK35CLwsIq7Tx8UxU8btOk
PmUKdLlbqOXNuM8m1TYHjI940nzWOX+B0YfLzvu/NsjXfRoAEqjp9Brd8aDykfTgQKs6r6rYo3/2
ejslk51a3CrfwLidPhXptTrD4zoCyLQ2YaW0ToS9orQm5uBYn+iM8cqpOddJkJjU0V13FPdwtBKx
l2Gjrxcm0yei/7PDmnO9Jpi5ECsfqGb9mCRHqzpyUKxFCzTUunvliWwGfUpYWTmRC2sNK1pbcWrv
uGlpYwYR2z1oy988QLQg8Sj3yG+B70xWtAIWX9hXFCQKuyzJ4OciusHO0jpQG5EFwz/FKzoL2SVk
6GLOSHcMOr5cW2ud6mV3NJeBXZ+79UmleoubV92QKJ4hp0VCp7wa62vfVkD27NAfVPFhATQMMhBq
kycn6j1eysVDEVEmInPN8vOK10NerZ8a8opz3Izrsnt9KheuYquXHo58fsTxmyvxLnabEblOyvPx
6BOYflM7Cx3sNK72PAYDV3bZXb6VcCUaeUj9gqI4+cP2TQB6HmsF14NrTgrFWdMu2Lwycbn7Ttmr
y4nnaogaQAOCGDmlIopEO7byck0LBI7WEAqSyroLUUYhy8SMJjOwOo1F5MjRx+VlmYwffb0tEeHO
BALjziZ7daA9MV1FOIbz+aERnmxwTXhv25JRdVHiZF0ELjpbB/DUWiOyyJ6CddNFhiffPfPplKxP
FeEQMPs/U0Max0QxtZrxAD35XZeVvO6YKqltH0IpkOJUpZE5RlpG1TWpJVmx5Gq96imxrU6/uuOi
eg67TZUJ/8AdnQH48tPwqa//Rq+tF/1XO+TQLG+/DmeuJuTp9t3wwWuu39d2FzMGt9TKlr0N3p7W
RobcC9zLo2o5D8AcSCr3XreY0lYrur2YhIZSU+peJ8Ekh8sQTjWpE6mWk/PpNfjdPJ8FUVs2v/Rr
8S5nhSTmkjG0WfJWw49kyBPyJL5h/42b5NKjTAxOEgrufW0kY0/2BOWpYeyZqwv/Uk964gP+dTnZ
S6oSjXulK5Wh1rdrMF4Le8i1hITYE5sLsoqQpJPyLWtHZv1BiMZPJhLBzEnkQq6Syd67+G9fil+c
pvBVzbxKT7Ywgn1x9vQZd5J8Bg1hBD+yrzsKnVNjBhkTpx0tNp/TZXyduYvJ+Q8dKId2eNYURcTm
UTXfPfNAf97wjt7FivKHf/uuFzs0cZRCuDe0GxNady5BPlDhWTT+DXjUJg3i5fMAQvlKW4uPgsZL
SbQ/11XhnOsheDQuaEgHKrLdz3XBOgEpGI8+ZxjKtREb+RBknmqWSIgKoV9aBhdnbxWdZbxmAzCA
nUxnqBF84YXxiPTp28vz9MKGcLScTq1b6NxUjNrUXIegs8Mq1rXbMyTw/vu/ogj9bMWE6mlq0AQb
MJBO8xHqk/wwXu48FnhcbZ6J0Afm5rKCAUeslnqAaGHD3qqBCIoPa4UmjC6tN5TqH/JSI3FY8Ys8
Kz7HFfKOhGWOHiCzE7jHKKKjx1qpHp1jVVCk3BjhEEpd0avt/h21Afns7sVuHi+ebHPs0IH1k2kG
lQIr+2u8OPkyyQi94j3zJhvlCYLel/pNv8apiPCwpBtoBzxNsCPo4gucEVo5LgU0XaYV3lZ85teL
erJNzVaqJJMsRGucID9ywG8bpONNrI7+t5rFuWpqS7rWfI2E6DahtVNITihRQT0xj69qs9sfd/Kk
OsIhK3kOIIRqxnLi3dK4JpUkrw4qRo8v+F3BlpwnCNVYKWUOSz1McvQ8/bpEGrF0BOVt4WjO69He
lhV8YKp2YyV7Rlwd5DqTO93CREkyDBIgL6NC+/p5oN0NOKzwXfggTJLlVPtuTZX6Yi8LVLxXku5Q
jNHDIutSCKdhfnFzrZME0+VnVt1cMbIFe/VrS1attqu6tAvcrEoQuOMVwpk0KSr8b7hIqCPD9Par
9PiSbD35z2BK7sr0ewjLq2kGbkem5s6xhMZ4XOFSV5UdlfbUDwsCprg+6S/kfzmWh+epSe/WtqWI
cr20D0aWnT2aywhgAgY2yeIYXQW9lE+2p09cbK8sKXIF05y+2xLqxtHctcmkl2Ba6sw7/SyXatP4
87xS+yh1CjVe+PxWkoNrzZ037UHY3MUzM7A0G0U7gbvMH/ZbT5MCuMIfm21HhCeulAExfW/vTdVo
IhgEk88oQOCqzCrTd/nlPh2i0Rwo4OllqGf9t0tyxXxv65lLv4CoQXDKWDbiGiVUiWUODhPUpjp/
a9w8IrgmpEPGwK55tvsQOPSGRJIysKnMQI965TMxVyhzguVrz649Mank4N2tNQA5dGc+kBj3Qtwq
CujLGdDeoxcZIiA6MLm+0loqRpQqEMynh06l/qX+LvgtK2q8i4vvYrnSyIpEmL5SzPzOuQiSqGey
8njoE81nHPSZQjPDzg9N+UAAMAz9aDFdL2+2+lTXocpKb5iBosn/LGqOsiHZQgL7a+cnYmWi4VNC
Vl9TGSHCpaHstTYArfuMx8lerRXRdVvQCMJj7f6CuD4YC2SyzxkiTCJr4f5ilKA2jyCO4gtdYLQ+
v2z4mj7VCfmWMwbaxew8arMTIvfaD1iApwp+IhMGjbmzHkDV3igFxaLzLfGayxRQlF5qBSfYKOXV
dRN/urfZxxTn31kdG8rqhp85vlAJCAgt9kZlrw6hQMk8So0VmBrmW2Uenz5wbZeSfTIXUe4iJbh3
qMhbmT3oCVPPhOhQ4S8e/Vehn/ibXOGygDo6BWLyPrkV4RcW70Zv3eUA1Iap9QjeuSMUid0+MenA
UV1znp9okphHvJq8Dde5qLOxtJku81I2gJOVImGiLfwqLhRZKN0iwtRM+VljjB4aEFIRCkDFmDcI
PLyfDeiHc3UZYx6vNH/Z05QBdrwP+C7iv9oQuWURwUE6GZ5BgVyY3fqbuOtN+57kAK/Tz+UpIM/v
MHK2adrM3tozRqv69ZIoj9BcUnW7JlC6SagYBHChvUkY32+ANXFN9gQivC3/MGY3LjUJvxed+pav
CFOouQJ0yj7uGzWRwyMmfL6gdbA96cGUq9EWIgBmLPRvtCZwbs7Ea9QnPYQmh+PVs1hFapdxxL9+
zeEsvVqr8+fzd1FoG+sDLM+cudWE3d6myoloaWl3dCGMAuH1Oeokefx8fHGwlAFZtqABrGkzkALe
QOhmI0pciJ7lZOb2dG/UMwmy7TzCB+qTUmT8OD4eHfzEJu681ZnZ0RSotjbKRNuM10jvyQE0SMT4
ZIasvRnq8M4Ql5FlxjriJQC1V80vxovkFP6gcc7d65CsNrhILq3HtWq4HvxFG1/ktKZOPC8ALqbj
m0r4eLKejKxxkROWTIKhVNjzGC8lBYSH/zOjFHbaXWzgnmGhqOoJyLPC6qw+kvWoVyrYj6SZtB8r
VCOGmbX04cf193xjt79Px7FbcGUywf4O6r9tVj2sz2Tktj3D4g/aw9vuGoQF3lt5dnnpBDYm3OHW
XAoE+CS0//JSjzsyditSCxZmKQxz8K4naZMAVVMH5zzQ1R1eFGXDuN2P9qMj8/Wk5RXfKg1e+008
RNYvOUhg2IarfBnzV9ObGvR7qxhL96NmB5mog8fR6mpnuWNuEiYKyrQggtfbot9s0wU4fTyzemjN
Hraj48TyO7PDzQqvmVIgPbvoyjX5EC6cYRDO4lzyWdbRT+UUePpPhUB99XzmukfxY+Oa2DlT13Pu
p/7c4pPP/2IHFyVPqOZuwgmqreavMXrHojz1tkJ9jt2o7KJe6htCVabnvQO+Tu3ZLQdjFxVOj53s
4up8V12m8hIjt65hh5c4loUcyo9psD3LnTaQmgvw+ps/ifpIbjTzVh7i0//3r4jRWGB8Pb6f8/pA
lRAtaGMMNqpIEtD6jxG0TJ+JGxX2JXcaK/2DnTeGIMX6whfpNyUBQE1s/3YULIsROBGHoD9DS/pN
Ha1KpbuvdC9CNu0JslT3Qh0th5XVseOJd/VFDvCbsg6bmbbJSrj+GlNPXNGcwO1BcqZzcS55NegM
KXbVvPlNRYRGolw3Uh111W9qIjgpekD0GzgEstiDwzM/nmCQlfLeRXReUSi81Ky1iH/cwoAL5CBC
xBieul2IFmbFcCQ7tIXN7mgplTfZbeG+kJidM94tLsaxlLMr0i28RjAK0LCEU1AdGhjAJBWkKqHO
Qaxj3sNfh4vieHUUn1MmRbMOnRbAjUrbzoRf7s0rjq2I4gqE7mS/hs+UsWVhHVhOgXysy77P8FLB
bKk/U3NUufYzZ9pFQi9Zxas0gWPkDtBXYlQt9gR0R42x955J7WTrlOFcqmovchhVgRB1RoSjuMlQ
5OLXQ1SbLHujoVnkLSXJzL4xKMzqzjxj1WpXxUKiXV/DRibnpIcF2DlR3WYJfiz8KY2qbGm+Qf+p
7t6PrVdlm9XaTgu8XqpOhK+WDwo+faV5CKje4V7qp174q9B7gRbYgCBGroABi7ARMlADR5ufJ/hr
SLUhPESr0EfnSMSO2LOC/kM5J8zkhppSP3lyh0qkz+115sVDCdryMR2ejkIDXSdxU5rZtC/goYLC
akoi2YuCb0fRj5R26ZEhQmw56PXxhWn91eCj1cayXYWEZORHLMyuu9b9J1ZhX2vnS4Q+q8OOrujS
lR9YmxRZQp+voKOrTr6rNnwoWVX8uUmUgbVum2Uosnjw5GGkjf70b9QjSqhaDnrTXjmj99udrgNz
wjwihRZZRjH+nlmL9IlzzcSCcvqaTwQtLInSIsHU/iBqOJLdirsfKq4Uw2v4Y13UvCM5Yiqc1qB+
IUrf6vMYbxFIuhiZ/1SzPOv1F2lHeDgPPQisvSj+Iodm93a9oqPYvLGJmIrpP2Sm7DhZBjnC+DG1
1yakp8ARQGyYO7pGW2fJnUZOLFlYC5Hth/NtlFpS75c8Mg3DCiaIK57P2pfRrmwzoLrgcBemUAWb
wrkSkOMWxmXyHs/2g4lMAuvip73euZu/OiBBJGIOH4j4sm9W85CtDCQgqytuh60219D2JBmQkGgt
BSaQ2JH4Mi2NqJCiiImkeY62l2iR5TyFQF4fZZk1aRZueStT20sIXiTdHVGp2sDgTc7bucwLcewO
wsvX4UO9Q3fFzFmQmCGeZQhgDinojMlYcV8ARPkyJacgdVoE4E6C6PgITeYV8MJQvpdR27bge0fy
ar0S2WDp9jknc1Exwfrmj30eKxEL9Ppo88oZqYnXUDQI7oBKrVLVFNbhpu8yyRcGcPp06V0euKw7
nMEyqMe71VY/Y3bIOItQwBWvivGT2M1fJj29s9LaXS5vx5bRwDXc61k8eHSoSuZmkpb4CshUlkFN
I06njgwmranjfiaMuZu+UloRy6CqmyE4qefjXDb0q0Iyg2J5PuNLZ7uV9B9IKQs5wRz7LBT7l6rL
JcMf3FSfaxbOwFHuPIhY98Ec0j7YDgcX7fkadX8BYDNu2cDcAMU7XEGTSUZv5mdSDJyXGa3C/nr8
fXw+GJ1SbpSnT1gfHCQbD7oUcjWI9Q916I6tG1ohZimmQHO3iIchn6N+MCxcrgevWTPP0/rRXLhc
Vczrpkkw8o5PNxVdEVfDSKKKfkU/3RsBM9TVmxsMoPpcoZIOFOaOPjVWVPI1cptsPrbpw6vQhgoY
pASdN/hdkBZLk5YWdt+ZQ4e5UZ6vTnn1EAcvBM/wLCcPP6jYsUd23t9q9NVHFM0PGbasK6GEwae7
wZjPQ8dt/HL6rbMxQLhv1QldT1GkxthRlBJK+ozPv/VOTBEj+MUepSJ+BzCDb6ikd+kaOlLYIawZ
Z3cvht0Wwc/M7IB2bDJCh0E6oxlRQ3fQYLdfOk1MTXAkxoj8s9IACVmyTOtJlxsVf49oMRXuzPRc
nPXLS0uE4Yy7G5pamP41YVoECGv+rAKVS6FOT5bRJOwy5vQb5vWJ5H/8i7rtteCoIikhgrXJwZy5
IrybI83lKTOt6vVpXp65kMfH1derB7zGYhIGwHa0zWoO/c2bMDxxp8BemLy3DWwr6VQSVrbofeax
FGhiYRZcZHA/uRr40wfNblS53o71LBURG2Jw3riEMvAEKkeRzR9ZON775q8jytx7G/62DHc12W1F
v0HlQoJhrp5tiIly+Phe4g1/aaYY9+asuX5JEEceLrl9xFMbi/phwJl+kFcf2CzHWtrwnXIYHr1c
yf4FgBv2Lv71UBDSetWllI8CBxUmd//mOhIgGp/MA3hAzTq/ngaqWEcgM5SxqQU4YhifCmFJgamR
Fo0MLvMeZMR3BMeAP2WbLs1g/fGMzCzHk1Y4xWp/2SkDgb27nBD8osx+EWy1eM3E9ZWdvm44XvYs
sLtOg2sLhGrfY0JoSCGuVludRIXyasvbboJQlnoQwJPHZzEldDuab4T6rD9DfewL67mPNypaFA3g
QpNoQ3VOqkZ9ZWHRUCm7tUMDbVET8zRenOGHZjBEN329hd/EDqKZmbpVBdPcZIHvDF4VvKAs0YP7
EU24ozj09BDtnnGGmHIU/wbsbLv4lApH+DPK8Qdofv1fzaZFOWMgzlsDurj+4YDVgY8EyBAYk2HR
2/hg0zGzFlplQYN0Yo/tF/1z+wYmv06MEZV2eC35mDAWwpTHbOgQhRE+EvvoKc2Uc9sqnYCTSrOO
+vGD5cgS4ykXvIfWV7HBbmwY77+uQFSEdYSwv1Csw3ZpAmusGeIUGx7/5HQzwrtaMaDmQU6K8CmO
V4iMnszzeE7i45qgNzOGj9D0sr63h77VQy/tXG6pDWtlHGHkLzlfQ2P+EnTARLNkBePtcSdjP5vV
1QEsaq/xAkU5SW6lheVcIdsE6QfiCjkfCTk70I+VyRtPgzGEJCvoyv0vSJvCEbQzoAN0D4SRVC6I
0Pqzlkm7mnjyc1f07CeJGlgg+pe2cESS3dvKiWnC/QhE944no9ilx8HjQqG6w9y1Doaweg8bf0fT
jgvJeTLSfr7Z3dEgznl2bK0ucmqg47FunRq6rHvyR3JRXN3NtEBBmrBbjV35ikphC3Q2qYFneoDe
gJymHthp1MghJZfDTbQpP5fcfIHo43PJQXhNviCHO6kabX69uMqPPkwQkNL1T5tJVpRcpY6ih0ff
KOpTDris4LcRHpjMOa2k5YFfJWDFwboP15h0biG37bOhOLO3gRA9gKNMuqNB2rBk6w5Ui/rxP4r1
WkMJsWRhYgbKnIP3+96q+npgF/MOmFwrSG3urXqVINhi9D9Zl6EMWXcD0a57xlwLqMtyFp0lZG8Q
vUvQk0Sj/2fZMgzA4wzLozZsmE1eKWqqomgE9F3x8x1BdCMBXZZH9fTNmLqMwREKG79zMzUvHfJF
J7a+uYpx5lahpeCwtSjfRQMw/5ApxcjuWOTwAkn5peyNtIQaGZAlAQGFs/8SNej2atZdJ8wOBmWG
hfVniX7GrOyMnl3FLi4DhdJNLfMEepwJQoNrjLZP2SR8AFVS2IGjjUZ9o4bTidjpXAE9umnH4UUU
oduiz6PlGtzKrPkI7D9Po6niKUVfBDq94blL7eNbSeL6Z84x+Le/krnTil+OO7hX4piFpV4WUjfz
I94MmWguu/neFDhW4I56wBQd88Mz5OrFgFy8RjFk+D2NpEV0SWSwcHMgVddg4Kho3a+ZLGSS6wiA
3Q5zpUivezM7tQ2Gtwt12VU6cKnZ0ub5wm8Mn3WfjegKwcIN1mLnzxHflwpAqfKRGVysf05xRHPm
mercyCDghq07vP0EcbeefA1Mz8SqLp2rLdCtpRaC9ywF0PmJd0rXt8l/GsGVwCHQuZu8PRdG+/20
0S7EFQjtFabGgjd9XmI0bBy0rcZNd33hdGVV92VaeNFU9w31xVZntr5IW0KwP759uU66wDXJLOxC
J/xirt+hRoLHgdU3SGsLboK80kx7Dp4UlbFcRC1jwGK++o/FPpinxpicU7yzOBtmHY3Yod5/wUtZ
wghXQFJ03pcOyvsL8DVwEV1k53lOIyud2fC3KCG6gexxr97j2/UlG9xhwStpSlmABzP5Yl95rqc5
6LvAeHXI6+9qpLEJ2EZ370lfmNI6voGgNhfAjOx8dfV8p5JrJKfCwJzTwc4ZLY1l5CQ/LWOxHP/Z
fwm558mPaOJebV/1fyPIJ9ZPrmDtKh/ocsf2tkLC3YHcTck7DjnlPsDXU4Pmux898ObC0cgXssgz
/wXZ7WT55Crk/S8yp226efNmaZXBEZtgKjGy9UWAOLSsR2fL1fsAtcYk56nl73BhK2RI+rStQbAP
9flbzVX2bU29URATKroY5ZzA9E+hZsKFl6QXtRRok6G95P/LhZF71yif8FyxKisva356MhUQGnS8
l+uYKk3DA4UGornvmOQK0Io0jNvqdCbPfkwdUN+pcM0rgpar+2QtBb3DbggAoNdF+QStPcTB+N/W
t/JbH9CaTPLs/cvblbnTOvXErZ2F520YOneKc16WFJOmzRkAXLowWIWfFEcRymYVBSnSft+Mm7NH
FM494iegP2RGjls60vhbnQI9WEKJQsBU2v7SG6o1/5c12w7HtcxlFpn8fzgqEAsZUgVdbfplKlQu
XBMTGn2EC74rcV1GapdEGK1hZqw3sCOeFcg581q9LGNvW5GwjukXzTOO30dMNHi76okxAeYgkkPm
hB+5v+PEy6YQlL2CEfKF91U3ya/egIps2mCCetwZPFWWyiZAbLAd4An1kRhyD+7cI/pb4dATKjia
dV2Y8Ltq6f0ZAH0lBXeZu44HP0SXMwPo1QsB8vWJoDYmVaF+W4LEKMWpx6g0WGnkGxE+8W7rFQTU
7nGwH6L4qRGMeou7WQ0BsLKXARmTpv1m9cIS3neLqLDI3/Fr0S7BkwW4sWfRkqU5ll8BJpEM5xS7
d/6ox42xV3y600B2aokVyl7vamaiopqq9C08H2YVAiZXPWlfmAn8cpZHFS4btcKnNqedNQPJSvew
japY8z/Cm9bRjeaiCmTKTtFzUaKh5OSe00Dn4GGBgPjff3q+ahWajg+Ut8XpqJEjiaDOIvVVu2FN
gGrsUtK7BQPy14ri2gmewXsWtGmVmhCEYN56IWYfdmM/+cD3LrLbldPYdTwtdJ/Oc2KtCVtfqX7c
/8r8TeyPYyUgQUSti9v6dcq7pstp1jFv9n2W8lD7dEHa5Ev8cyEio0Mb1CchL1+PPI8nXdjg2GOK
nXu0ejvq4xwKdzRiBBJOqVXbTfbWEFYhf2R5w0wOC5e9XKrXyzQlz+Btgsd2keSbEdYzQ8vDIPCM
N0hggXIkh2Tx9peluBmf848GGl7/FNCHGn37xzGlUo6j8NlH7h7m/LLeZf01Yb+qdit1nP+46ZRI
EScuuxGbqzMlhBotucxRDesnqJvOmWR/PlUABOnVIuizcjmwuGj6siwLNjMi3mO1lLzMX9DBLa8L
H84SLY4LVGM/iNX3LdAfMkfRABTHUhnCI3fUSb5/Dy9Hi37T01D1eo9oOnmis4qBFAGzNz4tnclo
xbkDzPRoAG6bLJOcLBlWV3VVbJMqatDdnZTUwTEPBgqWHc8oVs8J18PVMcb4/FAr+cK6IAFilbNf
8mdcnfnNyuYu1BVdtjXY8D0nWnK7e/J+P30JPCiVl/20+dZboljT1IDE04+7qyOLlvgrDJCRlSno
FeOdVxYCnrHf80SKM14+3i41IUctiP5yDKeyfmymN9Qu4wHqqg5aOrgtSDAPj7hHRPpFibhTfPaD
QDTHakPNbQr7hZ+8LYLPkgEyG+B+TtwO7fPwdp90j3tEE11kwksZHpcA2NFA+1Dgu1d0J2NgDH60
IIL5FsxtSusCG1zjCVF0Aj5bKliqigIweJN6X8xAa46DDRjiPa8FzlOU9MsEqVSerbhpK5Ig+xfX
XIL+FzZYh1BYExJiDktG9xlQ1d6F4PiEAVNV8C/Tfwwfuwnzca4+4zJFZ9CNqF2RqQhRTa9leHfo
1vzaGoWnD8sRDe9yEBMU7Hk4LiZD+loOPVSgS/CCB1DIPOUWduHeFASqGDfeutC07gMKA8P3gjR3
P6ohusjVOt8i4qi1UeR7lNULINMVbaW3cc4HcU5p33A9zSM5F5cQl2EVDlZ7DaPcSet0kHJYHVPR
SxbE5+50sW5PgbE1qKOjb1Yfs+nQS99WefKcRnZRhwXJFxOJDFew5CDeT7v3sV2l1YmBaToFbERe
fyM8qY/LEqg8ScEVGPz6+L3NWbAnz7Se2HooCjsS6SjV8mQ5BS2WGtoQsVUi+AiZ3NFXR21W75jp
F7oFZhaKaWevQyTEb8SgojlCDF65gkzBw66bopsbNG4doCEnzrqJUEezhjz4p3aPnQhwkd3ouK1P
A+ubezV4a7xb50guhjN9Z9pKi1mmDqs67uTxqudGaU84sb58bBnsMijtKEGnvQUkNehfJRk8DbZW
agr1SvLzcAXoEdVu6x60le56IyWYBkJjgFcHdw9ArXbQGFb3OnfjBlCOxp+5bPKg19mc1Wm/zBT/
jeOH1FQpl+VqoIV6ZfCtqEkp5tzQZj69cQuVk8LSkAPCbzt7kSJ0XaOa1s6Di6+tPyIdLk9N6Ci8
IbVeYy0Yo+lTSRRCZEogd6LP/PS4s1YspSUo5skxHRDoWKd+pipEVV7wzPrkZHQga+ZXrembO0lS
9OHaTWS9C9JCtL1jtfX8yUaZAa2Hd68cX8oCpRedYUcrL8Iw1BRJ7uu6Mp+agkHtYWc3j039IJXv
wGo4lghP3gydTUvfZTeD/am4L295VboPRQoYsZvoGfIKJQKELaj6LeqfKr7e2jTPkJw1pGy8WSqy
wHuEiI4QxQRob3ZctGG2rkbAbfl950whVsqSO8bs0i94z3CrxJfjgIfzaeNQ9PaC/8l36AwME97G
Lqh0lKBMbrbU47zZUVERderbegKjKKGbEcFbjfH0kHa9KS2jLjcpPloVzOthC3Ul9dhC0FxTUBxT
bVU3J2jBixxOt0leW+B3dyOzV5ORs/spdNQMWEvK0gr6R8j6Sto7a+jpQ1HrQtMuSfeqaE6McUGU
g/n+kxb8YT78nVyNz4WEw0BgWpa+a5z02DHZAZXQLNnHLAcbtA5re8iZmGrirxP0v5jFZHEkxoLW
QrWY3DG7A01jI9RFWtB5JZDO300izvbqFz0DC5H9ChhKQ72QY6mNLVa7g3T7HyFWbX7sgHF5AvaQ
PReNbOxBIkMX75Dqh4ytY0YHnfBdx7WB4TbzWv+IjHg64J2+JrNsvvpPSz67MJ+8GoyjhKrq/XWe
zS4eiPalm1oIXOP5kj8dsq0MWIKDs/HuWFuMP8u6H4S3Lsz7MO4cLHf2u0DTmdyXtBRBC4m9n7Xi
VPOrEtR2EO56cNTIQHAVrWxjEAzmT/ewi+eQJgqeEJzN2Zvf54P8mRykJm114OQPWHYuuMFGtk3L
IXIkpR0qhIUHG2vEE8KfPYdt5vLe3XqX9FhXAk4O93t5En8Y16nAIUfLZ/AqitRj2F/vj8thjXfJ
DqBF5IPlvs+mr7jozfZmrVTNpRlLykcuXDLizyQzT1f83D+z/pu/J4CmiFtxr1IafgOdGzujndF7
Sfw57V/9FmdOBzfGzgowU+Or16We0BKxp/lsOR+1Uq+A72pl2PYv3WYTXydYbaXiD89rLWxqDa+E
agCaLADE/Y3Zp2rUw3+SwXEhqu2S3Y9V/I8vk1GDoEGTFFboCgVOMIQxVM0GRTMGCqMZAS/b8tqZ
OmNntJNwanAhUIgDxszfswOl++T3xowSkk/wCGQEqnZFg0vNP5LBAXa59RMCZoUuM5zDI3va60id
vHrcSoUi4lDLBckL4/nje6szkPZn/hSVy4/p6reN3zwBhawZV8tMLrTci7v5UqbLZz5qvQNhd7Ka
F9vSEzu5Y+xGTO32qoMgGi0cFBLoHmvCe9DYhO7xn8iBNFxUtwMSAPJ5ZKSnTRDXTUxJoEeTnCSq
ORnnH+xKV1t/t21I+kiPkj/29xEjPjTtvLQn98OUJdMlapl0wvYUF6MF4v2IOYJFWad3ExOGAOXQ
7Yv7heuUojmRqdsA/G+GYrtay1GdzNYqsTCGMiWs4hxQyGfJPhlxImnAzFr3DMWic+kCNmrx6Pha
kUFkzGeckCsp23Ib10Ikrc6/jTa8xWFyRzq4rInuZxzUy8CSxSHo0lLMDncxPonUOOG75kRxmfca
xgF0+aZ/ohJ9l+HZ3e7s+fPnr0qmXkzFdC8TO/58mnzWhWwmWnPTh7lXubKJoNFIOZqNI2xBpLlU
TB6EGFOUXd2T+XTc36FrEmmm28pZr+Cfyfm7NNWp9yjMP5Pz5Hj2a7IqOHD+LMiCqe9Lzw+MwQwG
NfKDzXhYoY7uoHCt6YGrtdChJKsOy3l+MLx+aUoBGnj1tyhxmLa8UgrbAkZ9DFUZoQHeebsjF6+K
5BWng+X+ztDoStuWa46BqNYpjKMYL/piMH4bgUE8VeUzDfT9UNkEyLIdzkINlbt9k+V+eANcckNl
qeuqMpv8moUf2NrerPhpGtFDzm+KBCrCjWkU9I6N8sWEaSxCkdrCq8kunEV63OFf1eUqKmx3C6rT
GCqFd//IUGDvd8d6w9Ra+H+AJGtdI3jhrqsKWkrUqAWVBm2S5f+dwSJBmDI9TPkmuN0plaw0dZrK
F0/xQ+Q1hYMHi8e7e2mRpM26x9qCnRyTDDUTYzfwQQYSmSV12RRngpoDaqTemJkYis5X93F1661V
nuJf0HK2XmP4AgvNL7JK8VR6+nax17IRCpDEw7wl1dVaCFN2aXXimjozsEZmPXVFxZULSig1mDn8
g+PhLoED8nZ593uduitW4et4c9XnDCPMtB/hzFg9a1zCsJOvxnaaPgIOZ+Lp6DH1QpiZGCSCVH1U
Y+nRaHoZ0EMSMKn7AyTQ4HSan8YQ0zWXvzMCTnNOXFSWWYyg1XDbyqPeeK35+3R67zTKPzOogeEm
3l79n6CFtLdzbj/su18AV1nrT9i2NulrApcFV8/ZHD9/D+F6kZTslZe2FsOJxZTFTyTqBNctcj0p
M+qhpib83IxzgI+khv4CHKJWHo5Mss2ZEEj30h4VxtYp/67X/QvefPKGdT+UV8Fe7wGQiY2cFryK
ljRfS3+fIhhhSmzAJQr4gwnWcxlaU5eXUcOLGeVTh2NLYNN0lcP9fokD23vHZzCZZAnKEW1DdGzX
gMlbuUDwdZF3gick1a5rIHcHKiErxr3SFOr0OdHYkaORnwCS9HJMW9K9IcVKy6F+pyCAGonAZHeM
Xp7oby9gOVWlB/Q+jPFRu65QTRAjka+4vTjdzCtwQWR65/58hYsYliIMK99FyCOltuwpNRUCvL83
tEqgQRiuvR7+KpOUVhGiaoO7pVRf5LL092tZjfQ8pQDvhY3NBF6TwRDyIq8P6UxVDLFieYshqdkp
ZoYjd+LQs4sx0ksvsWyi5yiHKaB6ECpuUCWGdShEmf8yraDbXOe72whIZAhX4gvzBrBR7bLnBAtq
7Z2kTzVPId9UfRi1uohFUFlZbmyw/r7Jiiyx3Vv0XCescq43XAvhrY8VO6XQQE13goHuKJB8Lgfx
3ckBH/2j4+VOP1gSYdvRsX2x8JEF47yrHnqw07Ie+cBGcYlqjN5QGhsHpah4Jo1dVXEW+CO/OAym
r4YJ33fYTKNCeb5M6vhgHDANa9TZBSqkWU8gw+rar87ROjsMORva5ZZCjlgSxZp+jQIzwknotmRG
Kik3Fpkz0w/81CdCjrSomwGC4BFJY7Sgc5l1zJe59oezlbuC91wT78DLDI2Wqhul0o0OJqJEwvgA
043XxRoVS8rkNOyCY7lO/ajwxXlqkCDGImdkvLEGZnmlIIxzx5ZtSHiuyIFK1ozdyHb3MhtyoH3/
ep/aAcIZOE4h/20oJ2t3cOpCbSLQpO0mmnlipcSOlAh1I1RUBPIr7Kmy7MkREP/Q/AucFbZhYPoE
08qq85QEr1eSXRCJ/phQJ0/Tl3KuWc3eS+1iKtCWR0pJkIXhEh7abhJzYRc19PpBQSiXCvC+h2ok
mgGSWlXiNk6iMuXxdTtkNGTk5o/8KsFx/odAyeLvPmmAzEX0wjSCsY5JVqQmerfajGW/htL9WQ4j
Krwj1WuxdtXhob/ugh16qNdtLDvB3G92JNnkgbIOwmNAVDS9c3IH8H5T2wlnSsriKFa81Zeb5N47
2PfLMUuyqpVP/VEMGwJxP5ygz6HLxk0S/wCsuKpz2t5bvlfTCaXElayPKh5WyQ7PJHkIDdq5OigH
PznyFIkMWca9/0DcE/3NZhWND0EQYbfy0SNvbaq5DdeydQD/hX/JLJr9RcSZIWB63I+f2YQ+0K59
lYv42ZDWZnRGbFBhzXGBryny2HO0HEprxC1A6Qugt6z3l08dm84Yrgq3HZQ5VMQtfmTHXWcDnT5M
V4n2F89qqdzNeWOlT/aQSFKXPq35lzfHxzPzd0VL/lF/tiVtTqzhAwvUkB5Ids7CMyR9tU1gVHDq
u8Ee1EsknmI5dhDkQwbVWxUeQ56vqpqf5qYImhNyqCj4gWAW2V/L2mK+OkIDNKNUTh/qYENzYfPy
TIKiB+KBHBHFuJQmMYUF36ZaVczOMj3YGN4cU7zrYSHGQw0y/6CK3r3lpLeoqqqlrfKhLiZrg2Vg
h9vJccHTcWFHIQr0tGi/OgqXYbX2AeeU3gEmcFX30kstNSFcjVDLibY3YnXiS/9pT+9b91tGeeDV
LjEgFMMQE1kJLucrQ/0nhdmlpS4Ze3tOuehFdKq4n18lBBC6cfWZqdAOOWyxkwSVpzB9gdn/tTCv
2R0m3U8jeFpYUh2DfAdJV30M2UnhfOkADbTI31VbWGW/1vTdTG53euHogTYbgsYurB6qAqxlDobh
+PN2WzlRqicY3owvEDjqDHK4dV5u98HZG1UOvy5tdQ0xyQW3ujwEKoGn8fnO4cAEcyCiVijPycHd
E6i/DLdp0Qz5eN+PupCkUoUxNUxHeNH43UpwidAC57iZju9mIOU2oIBu/UErpp2f6352EOfEroWt
KMSGVn2VM0Q3jR0lI8K8877KgiK1jF7Hb6U8ytx4jq88fEGzpZJt2a2D8/0TQiKNpLMLiRhocx8D
ba2kYNmew+fktx3h7FONzuzIgNKIrFVrp1u13E/ALKyq69wXg2/p/pO96irTKR1MQieX8Dj8jOmG
hYSbqLVhlZTHESbYzuq3ZcHFTwcE+oPt++BIVtVdW6f2JNF24Yf3G15lSNEnoqLtSm/fUIjOjTfD
LZK0GYG1kAbQwXXfyOlAQKpMrZhw18oSHC9rIDa2XEgYtrTPJIoL6WBMGz42v1QyhabPqosdtZ21
BUIXsOOB3memFHeXLWy0HcctCvNGsSHQkOgoLUwzcb+QrI7+FBIXCoHiy7IdhDwhVVmKKzK1pf64
PF/2Lp+H2iHOgyqt1wASymgDKohY3AYCAaxeBpvv0CYsNHB/J2hjDetmYyvgqctiyuzurWRoahdz
bvrRNjT3YLF/JEeNDtzISjgNZz6JdIpEGVvpThhxukHPT8r7Te0lNkPqpK0UXFpZ1HiQgMu0Eba+
Xoje0sJEeoY9JbuT0yn0Jss3F6S+vACBCxsOx8vEUacCXf4ujurycH0MvGRLr7qjSUjqudh0rLj2
NJjNaIfqesUunj6qQuzyB7jcz3PYySl4qBxnpd/9f1I9tVZzqZhbdXXGQe5cwOOi+5PV+TR2MEva
+YqnSpSVFDYfc/AvH2hjPjAxaNed7dJgbUH50BksGTbJ6ws7TpCH8Su+C7KTlZXEcXO9cF/ECWS4
yTrBJStD7Q1VN0+LFVcwAR191/0MfVKT4SVL6CoGqnew/z+G1cH6Jkg4FQpG1IurnwlK1OkND9PU
8/2RMBqBuTHBtR+o65HivUTVyHwC+0GkzY9CNtUKipoY2SNGAn8biIkTQ759iVM+IcrK1hKTx8Je
ALuRSYfYj1VRmI6XVOv26jRoaBZo09+tVgsssqF4YnNgXiQp9HYUwdZ9TcavGwtwE3KhXc5F7T0y
z6VK75j04KB2lju1aQlXEVkNYt3g8q7uUBvjQm813+Jzzmz+gLT9ygEsb1KNkWwcpECppRT+IyY5
UcXO1CjIt+lSRdtrqGZiwugBN+wvUncyaXwT8eEYrQSLxyBujL7iKpOaQ7A++W3ehs0WoWXl3Z3N
hveQKr6Z8cu6oYAHb8JfLLuA8TRnqDCD0AtR1CXaMlT3rn0KXLY7u2A065vG9rTeW3akZbqSVd1t
6uN5yoQrDZyRShojaF1sd1MHUQJIy6o97wTzgBXW+xh2L9g4lDxjKott/hAepnRoVYbwL/f6zxpv
UA6liEDLTKP0+XWPP6vhQup47sTabZCtbomO8Gj4Tu+LVueP6wXVh5jbbfgABI3P+As+VsPhuEII
bi2hXQ20RZIS7tALFwZZXq756kmDjYByv81xDh3tSjzOptuJJlKxG8zKv4ixn82eAzBOebCTlQIy
ISRlfPQkjEYIn8oUUQpm7REZbGTqmERbOHg0ThBWD+J7jJFmnq2XLOTNqDvFZEIKdtwiUQdQVCpF
EKStFYXHpHmGaJDxkrsGAxShtQ5rGXOQUEhZkrJrOPFesQcOkVOXfgMp/FIdKvHiIicUPCnFmtXk
ctfwyD/XgRrE0zHznr3EXCEz6uUuBf2j0a9Hz+HIXrOESaltGlYglBewfMfO36r+U+mic4S/1/5I
Xpz9/iD3+DGryhUDNONzyYIxuAFPyM1Q0f1/pzZknmxVpXGzzQU9hXJkF2fFHa6cyfhrdCWEH5BK
Loh8cy3UzLgwnLktY5ZHj/KSMBJO6j+HQyJPw9FRaP7T8GhdcoApd/zs3QhJ2zbXwHtRHv9Aax0+
TE7YvPYnmsD4tO5R6CJUoTlLpI5rejQe8HKGNaN0NYW5F09ld48gmW+wPu4Nq27tHc7Q7+Aciqyt
cF9HX0Lw34VqFDhFIhLM8vCbt2qzsJinwNHvcdUVH040z0Bk4/mI1VFhThL+nJloKibWkBA+/YWe
AFJCzW+Juo0nPYq62YcUzL/V/pa4JjxDnR8FT2ueemIS0jDihPSC6XCSq6s5WGFfScOaRU7zpufZ
wNeXhhDXzUou1TH/EeUycew7QCo/bBt1TPD7a+1smNgT59/EF2N+k5L6VFgIZg8HNzmQ2oebXqj4
IuexPT5/VEdfcwAqG4YvPBcrN4I7wxlMdthVgM9+NghXhNEpy84Wpf587e3BM/LCa1rzPboJ7Fi0
/qXfrQNZyxpZUqKYut/BbirnOUKAxvWCLwZwJhX212z7+L7HGfB/auq6gPrVONFQy50Q1EaOD/TA
YXvvJS6folKKP45BDpWlawwCtWlBWCleH96i/Ywcccjvruq+HIl+wHr+bpIo7apCC9LXEW0mZlOd
68kLIgcts5OlhBEl2PDIKS7R//vqVxPNmoRApcqec9scehnOk72eRHdlsNKptpMfvB4Kz3cypzYR
j4OvSj7mY1wlFhbUVNyQxEf2maOg9V21X3gbtzu7gyGTzOX/FeVFnMfNCuL6ck+6Fs+l2HgOoREj
zCanJjpkpFdSiyejYgjgj8e9gtuy2tCBxc4XjkZz9xgVnnta1EewDKEhHsUB6qcnC2Q2IckI66U9
YgQ8mmR4fUZfLN+OiarZZzvgm/ph3mnt5dRtxgqz5s0Mif4FVf4tDwJx0vv70l9FJ2jKYEPAd1Yp
Y9f0BBs5gjIbcDz3z+50CzjsH7mDE8tMIuPflm+9QE9ghfjhtTFdJZagGFLZr2GXwBT7aGyNTYB/
qBbfpFX9KqGzAmeMuaJBlPAq2bt+bwnpURnUOiZbWy8Hw0KKbt/KwOQkMr1lZ4ho8tYvWPnw6Y3H
7mdn3mX4YD940tOzwymTvo66pT+9sM+2S0TbaPSn+bMBqSeEmJjBGpL05A+Dy9Aq1v4l1I1rcIS1
HEggkCOvTQKNcONSekvZCk+V/6mds38Nhs1WnKFK5yHjNKXNyGf2zAEqSEXNdqKtAPRNKNmi8C/J
1TDz1J2xKWCn8z672mXH9I1KHVvlt29kwLl1ymLePDExNszUUURMRd5NRVYfCekNB8lZOTSloDf2
geZuhRnDUltoBQNy55A/5Y50elGqUvecFgZvP7EmcyP9kP5yOqVPtU3B3W8hyY0sBJ6nzxXAUAa4
s+0kkOgSXPWfzZiuWi7uHUlOrh7i3epUJGKWyKBCXIjRyuGgO7YPn0eU+WtT4pI4y3hiXKeN5YxT
HJZOc4bwK8p4bW+2wuYgjDEXbIdNL6+7YBI1Ot0au8r9IDazozTM1+hZI744UK7RIVgVVloxm0Co
3qcr1WTqB4zYbLrj46vfBZutwOY3P2quxRrRuTk99m7HujGaPAiu+IsdDuJzjdrpi1NVINiQ6fy7
IJMDkjGyVAqXQD/ou0PCopyR2I/d8hzTDdd+iRbwF6r4o7VFE1AIlYE0ltkgWaK0rxF/CKq1Mqb+
sd+mlMeim7mUxn4qbEt6pE1dMib/EcsN+T8X3FxkWBuacvjhFSNEB+o1N/agj3Lrr8onr1UGu8ok
Vro/FfAYlcz7Wzl5jua7p4SNAk06lwV/NQ2Zfp/bwZU59G7U/IGp3x5A53uv3DAUUVGn5xhcY4dP
vTWtNTP3HlCqjDPldXtjOuJQCcynviuz82VbKcmodZFWvsQaR0VQ7CxL8uJo2IGltpsQRpYPvDzx
1+3ELHDl9WxFCB8MiScfCEkozbbBaP8gP6Q72oThdFEiJCbsSC0/CE8RNKXCVSlAfK9A/uex84iO
7UNd5szioofkFqBDzKf87pGpckOqYiDaglKuAWSP2Fpviy5BJIuOVahllt6DY0wkdplw7yMXI6jv
BzWAIktHS3oRxW1XrZXIr4yUz2i1aXrVUeOmf43orfBjCcUNN1aPPD+i15cd/khfY+FKkou3EKvk
EsrA/tBV8igpP+bqPIx2SZ3L/OxgIuNLrePildxburBTwhaBS+NheKqG6aInMmPpgK8O09ilBnvX
sQLIQPycsc+H6YFwXk2X4CFiqKRJapSuRjrml/SKLzPf8cMkn5NaM7dAJ3WPXZV6kvKd6Gd48thm
/ImsmnsUOnfpPgw3G2TFRpoEAN4PUjKSvAoAkMjfd7mIPhsi0yk2Eo8WqbmVHNlURZ7dr/gYlqyT
okSx9Jz0LvKyyInLoZB7PXuLAJxa/D2KyXcwOVZmqB7gwG9aQCc61smKWb2DdLwzLwpqCh5yBb3S
4OX+3/3kssTLflUabUn+VwugO6zaij/2cXEArq8gYP9fj85iprcmPIXg1l4BMJ/1YFTd7Vw/3gat
2l+gKCJDC0aStCWOZH8AhXHDWfkaONOCgwUSBLBCySHKa1ytkCScyblgFpRMJITT9cEh0ysgXoAU
TpSn2zC10klPeqA78cHOZQ+gvSYxXiKn2x6TIs0E4Qy8Mk4twZGhcz06Q+9YQFnOMJpRlFQV7BeE
vZbMFQ3JB0WfK2GKNP0WG2Us1IYfNAKzuDUJIZIoR4fPlNAFwpG15vAwA0V/z5DJJ9jNBveGa8Gg
gqGDky/qJAOkBisNH1iv2ugAcdWkjPZtaA1U6gCm5piHhv34bKV/SaCGlFyUHEAjfQT1Yr4YF0Jc
n3t+DGNzuNZ9V6ZgpsG4axlB+1B696j1OKcU4VWNBqOYn9Cf2FiViG2SdH4YXtsNENbU//qTd0zH
Zm7H3HjSDf5wC+M8CKUGGC9DqgooMmdCaZCcnYh7I1+VPZJyJpsPNh5z0rznS0qypUTkYSfDuR3a
1YPBPighu3D7ay7igVSFLjDfiScbztLN19YTDjy56bKjPCt+tKn7K/DGY7GGdFN01Ic77lqyPOlm
te9O4WXYHugOnAf/Gqrei41hQC6zQ2NCYeChm7uT4Br+J7JgHl7CEzb/2OBeTC5Nb3NuRnXzp6hz
gZxwdl8TVJPeEQqYElaUVHtoAHh8C1EcmNHebpvt1hkx81iwONx2ABxJ7AcW9DfDEMUfj9UR33io
q7rXrM73HafaBwieI9xwiiPNNRhXeWtPFzj4feAxq+5i5pxAdV8fcXrvKbVdcVP/0s1gMe/0Cgdw
XTrvh+5DRn8wQWEqZGNjkfK8Edj84xjUzex14kDq4rZBaLBkvzmC4kM8cZrDxw0866G/Qiazx2gV
rX+Uk4rND+I1L6yaWXEaFitQFVLT1On/+/tReieoI1+MwVuKmitQldp14DVKW0PdVADB7bptVAsj
CR9jL03RPk4eguVSLwVEv4xK+n8vRkwdvZI8pYV+G/TLIExfsC/cN9DdR8xuPn77P67KoYVcO+W0
pH1hBiLeJ7aO0OwfLwqnK3Vmlaz+cOMZfP8iwQe6x1atKbpB/jy8wxbofQ9WauXZCqyN1R+twzDq
j0JQ3AIsNA+bTuEscvxtz64+OU877XGIt9Sp3nC3iRgYcsLaD8dqBjaa6uZfi4bX/dDbbnwLuLFm
/jkiz1kliR0QgXKX9bCbTcFUGnylk+UDaqf1/7/rPdsPL6yoga7wsxhYEfYCOQiu8IXDU/5Ks2ZZ
bm4+newzHAz6vJVX1eeQcvqcD5floE9NgwPsgsbHExcePTwoRO9oxW6G6UAwRfM30dMEtG6O4lzQ
7rio3rhprF9HbBZZ3k8Ihd23QTCQ0ql4FwEOK7gT/zw0CT5c5LNXKzchCLD1G47Ne/RMwMZHqkNP
iC8kWLa/R1Zh7ZsH1PBTI22aHs5jn+T6qWkFE+qcnxRBl7ClramyAzDThpzMNtCx6cWJw8D/kceh
W3kcYrg6U3mnATv3rmJB5EtLCx+yGylzxLQrdA7nGGrefoTmydLbZTG8wqNn0C6YU43Ccq6pJXFV
0BD8P6zeF2zYAUU/o+fbDvcuaQ61NdeKG7ShYZ4hHTgO3hIlqGZRuJrstUGaOH3Ef6XXmx6Tbav0
3P1uRgO6wSM4Qn6Q2wtvKVAxoeDScmx6OR5NNrvG9FIFcm6Tniz9A0VRGcfguQKdl+wRFv7qJPwv
/PhcQE4n2oTEMDhQqjf5pduPwi5HEF+g740QBCCfmoflNLG0gsAKDvhyXMYHHiRFmgNr5Sw38COL
SQNuR2QJjQSf5D9E3d5sXqUdOA6dbo1E1Zc7sh+cYDwBMUFuEtcrvX6m53qBAomZrQqa5jMS9DPN
rw82EgvXHMg7ZCX1rh8NtUO8EwjImM96fxbZ2TMJrzjfbkgO2I1HT2lbNsFOfk19KSHn3GqCDfk1
FIQFNDKr+F6dwKlhKjGpi/xVsZM64cov2puPqRaSalUr3/C1VJUxLDzzCM0A10zyNw3c1NDhdWoD
6zP1y2oEsx2MXOH4V5jPbdWsi8ZoLmybw/F0tkeHDOdA5LJQxHdwNrWw7lBhKm+USSi1OzYCvKXj
JIqBovai9UBgUgW4XBnc5PP3fvNV9wQeDarw1bjD2fb4hnC6D6hOUJ6FeJMfd7k233/n2mP3rOWK
/OBt+QG7dim9N52w4bG8ng68tgqskH5rj0MfiPZkqelZ8D1rGT/dIx0LN/G6agzKp1ezrJeFL01s
6Tz/JrVObcIQBGtmjgnJhPVF8syMc0B/CXEjYm0ot0zWCRInqQzry0ArnZ55IxS7NmsMZRsSmr+c
L8RcKMBaLTLHDEZjSKKXLlOhw7GZOL7w4PI7j5B9HukUnKrYm9ovgdfAX670LSf1aVg8z7OTbWri
O+t0NBfbjyHRS48ieg11UyfheJ7UWvTQNDemY5/FjzYjWQXgqBVsOppvqHlWKe0xdHsRWwOpww8T
cg1vp45qzXye46Wjlf9ODTbMrKNdZdfLAdKKWU9Uu7447CBqrjpTiwI2f7tp20y7Wm4BC6f1Obvw
CX3pd7mVyKEKXjZZxdER/TMusmGNR2WII1a4g7g5Af1w8AnQlk8fn2mCEcZUlRjbaPbxSHve2aOs
pTspYbE6OC4yF9L7n5d/vAK4yF93Cpc9Ns2GDgQA1jM6CLvJjHwG2SVudNS2eDEZcF+Lwlk4ztGp
H0Dbnj/uiemVJjxcQ8mDH7rm2NOuCss7vTtVr5l6oi3wFBKrFAYycRcWJ4FNPRZ56BetfjvcU5Ef
W+a2+9QXDNawMo/Ul24avhRgbFoPJyohCiAiq1MVuW44EtF0BXV4C+MLAGE5p14xNGw7MG7qyFxb
bUkUVZL6PJPdnhfUHQ5dFrCDA+gSj3e3kbHJI1Fx7oNdRcBAlZ1SwAoVA38y5+DqjvVL75RSz8sz
aG33O2mR2qDiNXtfLlJMHAXQ1GOzFU4Co2slNYMgUb/IH0LyM1z71e2L1YAdcBv0iPaJQ6B3+zKj
s2pIhBAY2J88IMgI5BljomoaFWrywH9MECpcKkFp9J6RE5VfIV6fj5aD3rsI70LbrnHIM6eiSVHi
SvIGIQz8P1gvvyNKZAaWjR277UEv034hCymZ5rlduc9MkKoBEQQSVBzuF+G6JELRMeVYIxVAPqsb
8U5T3rFnE7ddFktGIBTVglKj6vqiXYoqeO7CAdxilCu92yBKfFghgzFFDgCokZJ2uiZfU9HT6v3m
YF3bbx0OGoXwZbELUKkrxgxd7ircUsUXaRlb6jj3M5XRlkq4cCUoQhqBbKFVfAR4vFGyLxPOzrOd
EyKjkMcugzCVz0kMb6W35t6O2gYsTbG3V8A15U1e/eWPC+25rYcMl73GMUGLRUhJfOQQO8ykdKq6
bUvUavsbjyIZv84/gtQSNowrvD86qKZA8pc/CIk9z4l9uA1PG3e1mH/CnZGf5WO/jDJMC8hjyZ4L
5566sQgXXJy4aD6udjcUcSwfvO4UMPpMGog3lZS7/dH1z1cBlN56AQ6t0E55ZtXocN/2VehESqzm
xSYEl9U8Sa55MANq1QCr8ydRvDjWzyEClkGoiO6rdM6m3h1jTp6jT6jqDUw6HN+/PzwfGbo8TamC
L17teiNMxsOR9HTIHzVCaiEZhA0b1kx7csHdTsRXwRlj7mmdiF9to86RhSHIO4c52WMfzaXgz+Yn
TdJdGKiylfU7btU3lMYnFiIX8IV2bHzOvpxHfsk62FlhYX2/8sND43uWpzjonh/JMIds+EsPmdAu
oz531/eBVa8GAN3k1eAf4JCO/N53PQo+nx6/3BVPvX3Fm5H5u7LYeMXjiMWkFxwf2FkGEUokgGvT
BiOzR7Y01V1buLA6pcXFN2AB/i6eW7yNnQKQ+sCyHEVlJgreWCOCpaEO5l82xE9wtARsXy10+XV7
VNA2Kv0WqkX8E4sjEasrRRiSsVozWsfjDw8kFWKPs+FwQZTwGxP1m/gCfYF469toxg7+e0iLmGBl
9GW8+YJa0ikJ/vBkaMWLNKFSFSPo8q/xVpqJH4ZeQ5mVn9Dvj0N22zifEipJy3OiY5Nh8uvvvW4Q
v0z2S4XH02w2KKTtayfAoeLHyWjKgCSwhRHTzvDvqnl6zg+kjUbJmcsP4afY3ZG6sVGOwpfIY0+Z
GqG5ZMq2aQLvCJrQufm9VMSm7Ts4O3/bi/V510EMjJJm11PWTi1WfFpRrWVUjYUz7/sNZpf49iV1
bakuKFUhAgsS0aZj1wxAucZoW84cAI3K/Z3cLUTXskAFbN6S2xBc9dofJHV8mKOQ+rr7pFWcAvhz
qq08PIngoVovd1JIvSYZmwji6W1rLfZPvtfSmUtNnGPYh6Vj0NX5iUg5kYo7plAoR1tWfkkKiYx/
HrLfumxIufrh+KO4eNAWbYBVST+MQL8MjCBf3+WF0lP6KV8c2JV3nqNKYQDvxB2+b+TFPKkWjqFG
RvvqkNRr14VG2cE6l1/sUNjGa7MEwzPljxCcFRTWvT1OG2e5mfegaHUbWDde3arQ40q2Ne0eb6n9
Qf+UEKkxCvxrTtBVVrIEb+Bd9d/lupU4dFfyQ1iFqcU3w6tbsWNP8a7Vjtao6VTLLiWjANLA0Rxs
OD+CEzoFzeLL+O7CWp4f4WkNhFwSmRSESFZFUvwPWekJV5TaHS8oH1hQqYzwdtJ+RR8Q5J355J8X
vXsZb08eGkILmU1+Utz2PxasA56fjWo8b3cd/hCigi91MlHPb5kojj6BGk76TAZ0HhkH5Cq5aTKm
tRpa/sakn4rmaVME6Hif9SJFr+DZIiaMGSXV0UmgMX3cKSNuz/9uBavZ80+KWf+tBvA7Rx6YQ5lB
oBxpP1otliVtXz7H7l5Q6StHPwEoleqrveEpyFCM1kRPhGcC3GpoH4ti4XvM6k3JvNTdtC0ei8mm
wvv4rgaesMxnCdu4X5vo5X/VjJCWGADm+r/wNUP0aYG2h0of19zUo9iyrWeMsnlLRXlu3LYV8IUa
fMEyWt8m5KKLj8lxFw9eSu+4ZKRlwo9ngwiMhSIhURhYI1eNIKnuyXYH/qlhr+gWd+3vkwDaOsa1
MLMKjTu1RcDePWbwrhTCR7iCHwDPWFcRXsUQpbtlKlkUGkLXzVRernyLX6dJMEK4x+l1K8tgCoF4
ofg/+C+iXifA/NugH+Vz5X/62PA2EvikvVXh+IFgX4A0vHbZmfJoQWPmdikQHqGu4mJNc8TW2syh
xz0QvQFZTmGj0gMiIf2T4zfXM6Pd4Oy1xDcV7528FQFqMl19POz1f71LxI5heHfPsvzKBluQK/hu
5iSW0PRkCw+ZZc8IJLoRkuGqXQmd10RWgD6KfmXK3X0k1AzR0QvduJ30nrWxBbfB+VkA1+a89OHb
IdGu35PSyRbRt19uEM7z5cd28U3IYVFzQgphNmM2rvOk0TaGEB2xQGfMQMUFTL3GsLAIZr0VTZuM
Q+XcvgQ11OsSun6K4tQNgwjCeMWwdaaTujyVV4oJOmE/7892IDRkv/yQkjHhldbuA1e9E8vEhT3E
zGfOPv35+xhbfLJHQynr+5kgn5gIcZ2x4m6k+ZMeBnv8e0ywuzTJW1KoUeryrdNFSqDf5y0cuYnQ
VzSqretvRO72GdhHeMJb8X8p8soHkKUzpiWQLVawzC17+UyWBdwlxZAvo3BAOE/tIuyivFh21o1E
jytipPNlWqoQ2v3ekqxoSbzkoWdwD+EX2raB/OjlE6SJvfuk+k8PVe9x5RPauTUzPlHcivuUh/Qg
dvhj1sywXzg7vR7zoJK4OQU7A2UMViAz8FiHqcvIRx+2fL2PSGqywch+xyfoeWmFUPoH/il/nOQG
xTNg3FuZ+0XhDZCPASetJmvnNmChaHSNSrRXjCEGLAKBri2mjvFXTU5YFqrkaVI8y0kH4xMFyPLn
ou+kxtIB/v3S/p8q2Q3UWcVHdlNKJ8usJuyQ1UR1o2ePREBwhmaKK4jNavvt8Pc+yaOdyVCN6Juo
p57uWeEzoEkzbpFA59S6ICEaP439ZZGQ7clExy6T+nVQRNGtPIcj3+mg72KHbccBiCuWeupDqKg/
hVUuHrGoATo9G3Da+xi0Aj5XcZrhSVIhPUad39JVq7aKfiqXbfRQBJ45k2Vx9ycx9bpE3kzMXxAX
kLxdCgkgNzuIceIpHTbvggs4buoQeCU4m4me6cB6uWYP5l63o81rMY1nHOxZ3/LS64ZyE/sPf2wy
TyY/xr2bkFhosA6nnPXcx6pr/NoT+G3n7CijxpQFC550JLhX5ApVEkFTnZFVFM73eeW7DJpPInG4
lAo/yYG4B1AcHkGj9Zjl8vlVkVM08tqEG2pGuqrHTb9ZS8wSx6R7CMmHbzmHHNANW5DD2az3VKIG
ilq4HvyEz+0uopo44HRaQYfZwF8ZIpHJoN8//y4Fc4SRakDb/k/L7xhyZ4JqUapER/20hhBZrBmF
SfWdu3+FL3TCPz9n/NrCSn7c1VXjmHqu378ZzihW5jraIusLGcxDQfvypCRXmx1ZEKdOSa6fbL1B
G7D6mPyJhQd10xHFZO7NoWIn30Vksjk6Yh0ENaN71rqsZP2NzRexvdftIgewL//JBpLOwfSPsf3j
fYBleiwN+QxtnIzjq6vr6UHKpAK4gqyAV3gFDYDYpc/unRQatH3nVjtz9RLtE+lhvrCUKYB+BkNz
AEgF2ox+2K42eiQh+9Ooio8zN6899K9FbAHkaxUes5Y8vp3XEce8i3MsxXwdyea2a2j/Wgc98wkI
WR+byc1NWVjO+KgrYbOiqnm0EZylzV8r+N6uMW5M/szrAA8lWGvIIPI7dLBcQOIUAo362wfUEqME
bU17Jyv+cV/R35MlE71rMZ4MwD7W+A6o96thDdkbiz0eeILAerEVfNFdrMX/568xRD3axU5YUFWT
EFJBC4kJl6N3MpEUT0O14NzN1R2Ld8vfxnM6tHW3LYsu93iuEH515paDjAQWqaD48E1W7Dctt2yd
s1iYFnJu+7ril2WYqxWALvdv7i1SmQM+tuZgDpoWCQxF+BgrqMotUX9Sw8QSOcLinYmgefwHMRcu
Eo4mkjn7NoGp6pGadZuqJsOhXL9Wg68k04V8uRRe1W1Iy6LB6cF6EPHz1dcaMERk+HmwhUpv1MQe
cjby0MNt70GMKlXFPAjMmNeb7Ju8JjmhmbtuWNP0QqInS9aWnDbi25rmbgMqra9/TMPCan900LvI
h0aFNQXbLUz0j+4rxqExLvFS1mfRJCQmbb/dMtWO0xoeXxFGqOB77EZGur7S5RuvaUjcYZu4JEKm
hpp2BJW+KQayJBeUKpFLc+WMjotZxHT6IB6sQ4Ag26RCthcCp7Td8OWdOB5qqpE0c05Bk3W+SuGj
X+blt1j/fXWKZ+S2eDXAqqgLrrad8kpLdMDEqD1lHhTwv39W52rtoZj48iHhBRLLxCRosFaITOfG
iVjPHdqslqL3Dr02XrjXsWtuKxVLh9RKTRjEsbDaTgLAqUSG6u8ON3Gf06cOvANTa61eG7+SEXt6
eDC+IvQyQEG7DqHBDLVZoL4frChMU+h3SrUl5xxqMWapCCaJ2PprhkcgKG3xZZ4fWaYlG4MEjIsO
VW7k1Kx+2jIXQsl3Q0PTxFVxzbzPKSfDDsBlQa6MNIQr3gsSlVSHKHFwoy90j3EY3RnFXztUntps
fSNUig/KuWWD4VyjGhMu24DK5jcy7nuaurX/vbL4388h0YDPkbR8XGVIMiwxezpwRgnygEihhYep
RQz1D7b2spsid0R0nOaldal0K1qtm7puOjGspM10p/FSRHGQXQ/OSs3b2OU1MRtXT9EbEFProju3
h6vTXYejlgJzAS1xChp0U3VynPY7G5AqmMgh8MIQ6PNTziil+/ifoWI3h6M4NR7lj6ntWXIQW0N3
pZ5nSAHAUEZZBc/fHLaOHIatyBGRCaQpnkSDRjSaVyIJ+NJg5GXGRHzA5len7ABerP92NitXABON
IAB2aTDfRW/kIx+kVF45XrNMTV7Q7Pn8s5m5/Q+oeOCz5S/12yZ++089uJ5/vnZiLACyMDc/eMCY
SQdNsBpuL34N/3K9316tsowRdBpTPYE2pdR8erxl/eUmJNj/DrP/a2lXPKUoDCyJZuvCR76Fo73q
egX77m3Igjib/yIzzE7zpVRPptC55MUowbsQvpdC5+DHyUf0LWjQAHkTpnnJCHn8Ly0+RPJUyadr
IpyOb2HJ81smS/USGB0z3fxwW7bb6IZ89+57J2Iy62Y+a01JbXvC0fDk6j5IrfUxpaFyMngiwJbU
5CrWawHD9qZZqyJBIOG3OXPmFRgBomsqJiclWOJGqVo0OvfVyqW7BRkSEeEp2GVWCh5tkxBpYZYw
c9B2hxarhwO/D/9hI2GtzoQLFiyLGhxB984CqAZ2QLm0Os8wz80UUPBG+yl1Ss3bFOMPLNqP0BRk
hhlBF8HCqNJtfwVKdRAAb+B9yqGBPn8vAJMjm8Lk31ryiLLSj8A1PXXBu5sYEWW0NKKXZD8sKav6
MsgvX0VLTYWiaVNxxfmDJC2Epn26e4J03kFCv64w8kl4NwpeS7kXEHfZ9ASZNXGcSXGETNy0gkud
z9ftj1akwYtNDgi/oBaJnW4SnA8Tb3cKWtvuYkPicvIzoM/wnwIQgMfk63aovjgmwNVxcyya1VQK
W2qFq1lXiG7EL3S2ImoBZo0Eo347yCuK8ZDX8iI7jHNpeKMRPEIqXB3JOUZs7xcFmsX2XErbB2Jc
8VWdEacz41uTZIqSc7Io2UUtyxTm5w75nKY/Ejf/NPwSfpJKFIgfmsCo+dO2Bn3FHYMdcle55/gh
NrN8emBX/b45vhRjdEYEJ4lYS+axX9aXUXHIXcJkIgWs9ON+M0cil4CoHn6cGFq6fvH162jBIiwc
pkdd/7g+9hZxrU45zYVJV2kcBVZaiP+3mOKLze0aXOrUCN9/6SUJNMt6AeCHAVRDM5JjSA1fKTOy
0ljnjTGdN5h2B+P9A6X6hMJUnQMZ+5oC0YZMAgbgF5QBrHXhJBJY+6h/qeH5P/K18/uqLwicMdtG
i/mSuMbhn7DHO6EokcG5eyES2KUt3HPfLAI4SRY2iMj28J0NuCz6q4dD9WmOCVyNWaY6VD5sVT/v
WRaBCu9iogKi+LTztZtZun+4ldQ7A1GpaOzh3Zg03b7EtFMQr91FdhROiw5WWHgO5n3xNvluCFB3
7jiMBr8wL9WLB4GRTbaYSRw0gg4BoN/r/8dBT7ns9agpPHr2WNRiaZ0+m66INpBbKLRl+x6py+W1
z7f+h9GvV4wvEcUIHa5pF13TreMIom+mdMohZ/ZF4lAOm9a2vYIIhyXnZzfrj5Hcs/MvzjrPG55n
3/S7Op0KdheZ386AbXFYRytukoZlYI/4wELHfcD0tNGpuDB47QrQDv1rsVnaHmyS2395uMNZEYnf
qM61ZZdWic7EonP6aj8XqZNGdbvcGVpuC30XPKcnSIjpn2rKG/xwWOABDw+9isMO/MjyfaaI343r
9alJUpVFrcbjXcNgSDo+pKG+urIPxqbWmcdF1+WmBB3ZwE8vgyhqBcKoKCimummZSSrDthxEr9V6
lLsHJP7de5Dl1eiGV19uYZ1PAdW95jWponn3PTyr8eGLlzNij2H+f8FBQHm8pGMk77gmdYY1KGvT
zAPeYGB8qwsWuzZPsFZCm4OSynRVRs1fCHyh6WP22mB8uXKfRyFphcv5zPvWtxRIMM/WSY+oOrOf
jN43CkZ38t43UXdkiWD/jXfhfuQaASyI9N1mlwjbFZCsG7fbg/mCgqdJPZv77PbH2PDs1LZvoE6o
7LH7QhAvBj7PTcLvohp7Rqgf1MpPOy6oRZbK2hZ572hb+3Xbe3cZLpNdeM1GLcaOqkAt0hN0MOXx
WfL8Ts/b0p3/0kC+EqzDd6Y8o6tvwbjQrxpz6dR0cA51tRrdfhUZUQbGdxwYDW/TKIQB2ZYqyWTe
2KKQoaT1+uC7MUJTuLqTqi6oOA+mpZGoRosToqmSxpbCdTGyk+GWwNT3cASnkPnXnvm1W18Pik8p
bHfC5JArt5ZM64d25NZ5f6ZDkRdAqEBlFaVhnS1JxJZd+UbYz26NQAJ+6ClpBkFdTCKN6WJThp8T
/MzezOau+lpubvz3K0kG5kUCphjbiET+ADYfuyQ8mpQaygAee20829kOc49te47b9oSEx9gcBCHC
OgOMB6OgKxb0SeCv2b0qlJzGjjNVynVfEQKZGOFXoDR6m8bbjgl43ctz7pr0DS6Y3XI5Rh91pNN4
pPAFw4DQvN5ecEvinFycItzrPB5GIv/jxHPQss3+0AO7I2jAkfQoIGYGBX72rOFM2V7YaW5zP8NX
NfPRVFF/uvWYqdHFkWKOwllNK3AIR1P+4dQ5ZKmAHE8MlkyILDC1IWTnKN5XO2aOgz6ErPZ+LCf/
1dWEuM7VaeujA5GszDe30+KoIXuwvrD1/mWo9/ORnqG95oHTPNRpzPAqWlABIKx+7ia07gpjVcA4
eP6zHk2GcCDuRtX/79X0QfiW6wI/i+jYf0HrRZp1qmBhv5FxtI3uhBUcJWmlAAkSP21hc742tgyZ
egzYhfyGatbf3RzLNu2QPQgkv4RKv5jKcmxodfJZ9HOr4iovfApgnrfCbTrPr18rYgsw9Fo2Hfc1
4MaIo9+WH2KJ0AJYmeATMFkVyQF/JhB2o+/gPpo1iB5PZopfe1wPXRqpACUJHLzho26vdxr8v7m3
pG3I3qFlMjY7jFfkHZ3x66qoPN34KSWuuz/W1bCHh6fgIJNSrdl2sE5NH3hSI01C08TBzZoAns0T
V2tZzyrzwh/2bgfwoD2U3IrK2DNXX7KgRyJY8y32L+2pQ2YdjJ60wtznzcTU5BqyXjuzcJSNiw+d
62E5LUzNsvqTYY4FnAGhTuANmcJ2JyclO+p5i6Rz3p7Pl/Cqao7pEDY4jvQ/smhByH4PTfvr/kvy
jdYm2OGr3r2jtFb9YMu6XoGhxwe14RRqZfZ7K+W4UI5WLxg3yDtOL1g/fjb+QnFhft+ouwMlCL3B
50i38HcccQBk6bwZhYuGKvurppd3lehnP7JoO4IwWtpyKIjZYscDG+Zu3OOetJD5xCEu0nwoDqK0
OXHQDQAp8lnFl3UHDOVR0dUJHU/0IjSTqJ73OgLcjXWOe/F3NuzD4PN7B1lhgD5mTTJu2RigQLaR
trQ569oj9ZznOJY2ChLGMSeKX3VOkxKp1EKIA3Jd5y7pJ9EiDNw23flhD+Xf1L2AgZOtpZk6ZBVN
clrUeo6Camksp8YrbQeBWDeOD7XmZzcgZz1BXd5hlTZk1J1w5xjW3wQVZ7VKy8654y2ZdaDEd1DM
7pni/AUNfrUYlBdxps6JUal5CIQio1Oo4kIsDCJUq35jV7Q9+hgHct55dnWrnGpQAds5jp7FkB1B
2lt8RkhK9II0sms/GOCMt6y87yJdZwrka0amSstqGZoOk6kOxeT6pTjONG1/3q3ftF+67MjYZO9p
htG0yuChYUjH138YgUMcnPThZk+yCmARXhk40QrYtdW8Vd+F5liVwEEqDDUja1KxJXgjEJp/YT+q
/Nx9wYbywX9r0fMS8m1brLhvuoNczsJPNytfXGadllnFlCaDDHm+/OheepxOUl5Ulax8sBNGDaoV
pp13UOadgGLIhzrSKCJkIFnjmnlsKzu9fEyYrhSarVPj2eLOAei3tEJPwVo+4ToCQbRotWIiLY47
x5DKuSIDV3UyrpqtwJCe3nrFipojK4rczx4KGg0Uhtidw39Lq9DRFhWxdXOwYijvWBNRCiX5Fhc5
MmUGk1mM1Pow0dwhBVdzggN3RFbKeN1AVuqo1brOw5io4RX8QCVg0/3MY2DDUBCgWUhXGgZc4Dqk
v4yDW1ZrwEZCcLugiobEzJQPJNSKYjoGh73PvUSeWpnHFkTVF6c7WLkLnCfaYEL4L9OFnPJ0td6b
F8kQjOSnFti9HjuAU7KlyD+nKlIO6P5eBW0RdAvdqumXF7CuXDuDipusksP3hkGvEIv/PaNc49Wb
Eqk6FOCE3ylxU86uY1IdWf533uFaemDJgSFsLkZFcf1YLOsSpAnRJoSa/nWVOd+rAs62xWn/dk6K
eb2W4DbFdE3CayHWP4sPhyKY7jxlCyWzZ1XNuVQ5x6cafIqhqBB4OMxHOX9pJfZY+VP8XnYyrQmP
jHgegu/K7qD15sGvOLMM+SSO9y3aUTqxheWLIGMA4Fj5JQah1VGTI1pvZ2kx6lzpt37w7dvKdaPO
pGh0WbIchFFt6wowL9L0bjHTqeKZVylFcRuWfjehbpiukYzVdF70IdCGLcUb0ngrHHPBLZU5IplU
bknh6gy5/20G+ZtRrb3x6dMtGa/8S699O4DjcbutywUQyASxz/yHRfbVXOgJSp56POIrTQBBX+ht
ZR2msKpGOoOILmqYH4b2Z44N5iSeAA0TLElln28rxQ2QfMCT00RTPmbPJG0sHNZPW149x2xXw1iZ
MvWnvLOaLZL7Suh6rJdS51G47xR/XV+6amRaK5ZyviCdove4BfF4BR0VufHQ0Pm97v0t/3+5rlAa
avLUUDi4+mpnXP4joujEPEhJOkDsEuAo/uBN3nTMfPx8fulMVzApyDWngpoJvX9O7FB7x0aDV6VT
KAAAaK7o/WcxA50b/H/pbPkN9rNldmPvJTFyHXdKdbmr1eckvTpDwV+Ci2u+680+4jderFUpv7hK
Ce3plfiFFdyEVGTSdO7/f010VhY2KJa7OAZoMkEhhRd65Bmp+FQgbNqmjdhXUCQugqxladNJpQvU
hqYQQSKDOZ74RS3B+dYq8bg7VP7IRg0CqhKjJhfVFIhOx0f/M8LjPz018br6g5jAvp5kRVN7jmiz
pk8V5niLYaMdLhj08d3aoyQmYoYrTxmuJ8CqqfyWFqB/LkHnu69ePiyD88Jd7AlVhIfXoIPJ45wI
T3pTjiWWSR4FVaD1RsEK0aNZXvGwXk1Nhbo3MYxNMh7h3PhXEPgCT99mjfcbrk/olcF4+V+mgdVG
4w0BjyzKLfDykeQvmcwERxQMkdOF4EFC7IYIMVDKkp0meZujVnbTet0O4aXJs40BdVFw4MC4YRVR
mNh9YmAIc7yXcJBKsp+BJJYpy7WFx6rOnkPI/BzxA6RpymX+3PvUVr9F646OFft8FAcrevLv7ihu
6kh6LLNY/kvl1XH+MBKvYWsMWF4R+Xs6/89Tx7Hc8bYjW2Wm+tZjOel6wiU1QBOnxpAsVzfog9C/
6zkjwR473y0+JACLq7fwjxwNOfsDzeuaqLG4rFJRMViS07hsgNRTm+kVA3SOUNatebNkpF0WzaUL
M9dtQCO0rNeyBaZ9QSCOK7eK/Hl3i1ceegNLmCuAzk1S5vRdKoFN2++NF+9XGi1ZEN+/SG4dZQBH
NN5nTy1Oinco3t6j6HoC6XZktFqUjGc2icwZSJ56LU+QY5w/8HQOUdOARdQ42oYBBOLQ05ybBaeq
mCqSSq8RbVD9E8kv+3fwXz8r6PEpneuaA0hieF2JbkR/Zqtl9X+OlhL6OnhDT6n5Ds6YANpEALN8
H5HeN7HHcMHWXM6n2LNKLdNwuJ4FS/hxWRW+KtF2GNtmw4g3Y4WxL4i97/8I0FrMJeFvrTf8PA4Y
EoqbYC9WzyEu2Sz3FEq9W4hNSAQBUN8EnZSdfg6g3jJ1cLBGieKGKHx3xcAbGwYJGuqZy/Ci6pyk
O7xcheehAXIZy0D4bOD23AEu+38t5FTV/DYW7zqlLMvfYK9g9cys5pN1fYSK/vCcNpRCprw9/Eer
QyJhTiM+UTU692JJOhMQR5BaWPlYCr9oBGXw5UHL1b64P9cpUMtEzt9HGaMoBqLpCV4Jw7Jo42mp
a5kZ6XKmlmHW7DX9ZBZkvET1Ol7Wy7ZRp+5GAbYXsIlT1pP4VhA1LRCt9gLOKqIhreRkflCq35EC
jPOfoXEgbDQ7WkXK3/6g82lE1cEYxXkaJErlQwlRL5diTnAvM7rPB6fQqPprlGuVi01EBJjcnglt
TwC3MY4uh52CUVxlY/j+SDGP3yYSq8ixZesby7x3YHswS285PUTw96ROt2JBvo4xIXGeFevVqccp
qmVypq/cBCWg0GFSIzjpS6YOLnfusBfoHCFTNenjmv5TOIL17SbBfE2b+YX7AoCinPQqJM7EP9uS
XkkjYJMd2eM+0/yaTbzBN1BXgi1d8NsaEUDh8ITesOENyFgXNBZZ/AtbAfM++ev0T8YqWcmxW5O5
Qa1mgQuHWnQsrRX0LPpkQh5PIl/tv1Dc1oLl7lZerrNIDMR46bWYfLNNWSgdjgS5r1maqy0QOSBO
z+OFFwHvFYfEY4Q2QLxJ/lplh54cspcQpqkqZ2zA0/QSMfO92vncGhze1XNej6g7iCBq1gL1C3uP
Fz5nPEGG5QjZbE2mk9DCDFvK5gPBTx1Q1MueEXgNTrzEFZ5ZC3BPvt3WvWYK751yx7l4MImSx4lm
DeNMHjcPkGmy6zDkpOdfsDe1kuSkWsbYUjF0Znuqln4uvp07G7RtxhCcfvEkqyAqycYJtP9DvCVY
fEthcLnJuP+N1zU/YcqBZd1fR/KgX5oqKxNEvaAUC1vQbK2ULQSoXHQG9aoGf5z3oUtZuu4M8vCM
Nzr33gjvWSseuT/c4MtSiobeDMSzCfgKyj5Nvvk0VZihdi0PLMK9jLTyTwINaKzGvHNtekI2elCt
/6h+SadxdOR5dW6EI36v1dUZSVvfxgT6+5UZZiGbbnjfV2Cr8q+qOxI/bkNvrH0aC0R0ErtWZ5xv
emkfOsSZyQWSksE/cmvm8whZ4rFHqX8e1vAI5VR4V4T6lwPWml5Rb7USZJpQfMdj8XCjq8xp62bJ
PXlTtaPPjO1Bx6JA0BPdeU006nF5fgUs+Loe7fBNhCoBEAVts9WFVyg0nhAKhnhT52nME9STWc4O
daBzrn/UG2RY0P7NDBfvV13KraCqxLNIkvw5bAUVy3D4Km79yhIJ5bYWzxyh2CT47eLjmmGhXN+E
RGO4+ZHPXlH8Np1cELO3Z86AJFf9GapSfdqEFgvr/371lkPRXacUCf5+OyiPaThztx/E8TFU/6NV
U/H39F1x6xwvpKBQq0+1FugKmwdEjIzXCv73dtl8Yi4n66zmJttvaGs+YmSknHH8FDaHmKCMluiR
SDIj15F70Pp7Cxk56JGDTMOnLXxE+P01pieEJ0eV3t5+mEpMkCPmauxUbpyaRzsMvWxdTZqjhSZR
lg0jrZ4qA8ncYYKKMnJSNd4h3A1kdffQvo2ODdlDPmD+mdNbHLm84gBwxIZM63TmeUVki5LHdQ73
P/Pi9RlooECvE4XrBCiicb3z5CrSWutkM1InVd7CZc5y+0kMEUvoqUsQH7Ss61ZKaxeHbqPeBm3O
q4Vxy0UBiKBxnJewnB/PqsRbvqOtF10dSA84ZvpEx+aEjIOUdcnfzVUyDiFYLybT1UyTc0yMtpOI
hwx+G+tavAHcq7RUPhl4mtP+TdWHcXztJmBD9L670SjBLnn4jEl8hVajjVtkNl6Bx7ZIs8HoBgWx
Hgiq9j0ms1kkvC4FYcajSghvY6WzO9/gS2UTkJmU7JsORPOSSDj2P7bNVQWePnUd9qBpX8veOV91
aonOUXmTI/FWNXxELnxC3BL/nrhsMI8aNHzkxPzSO9AFJQKS7BvkZgEipZ+iBmj4m+Eq0sw0LQmj
rDgte4C8cN5qM8sgfK5Hj0tHzuKWGTsKJA/TUhKmD+kI4+PurzPK1/DhaPjidZMVIp7+VH5KmjxB
7MencLqkMElGxumC+iFXEkt5O0eCwk8PSrjErlmpnJupAWDXnU1csCa4ZMWeaYGLcg8l+wes+h7z
Y4jxwSomil5mC+yNQxtzRs4YSQQdMb4Ci9qVa1tJ8yJxk5LMYpwS16zMCPbrJTA3e2oio6i4Dc7o
VKGUVaOp4lMxWnk9hcNNTF1+XvXYX9b9sh2byZChMJUUUyvmzNLfZS+gk1EftS//VZZA+45mjQdl
Vc0zJIunJtIFwPs4rr8iiKdzheoWzRo8ZAREuHtYmI5QyrX0K+TopKijNdIZpgnpNNr1o3LrK4c3
mUjjcUUUEk0zQpNZzaE5QPwWPtxlqEV5hdAlHoHQPt9/sMH/bR34//HVFll55aprUSybgBbxcomP
BHmw/gbwO8vS4jOi+jvLLwkbJ8vfv0bCwZfPvPSrIMhjXCFswSrmYl1Z9Jseq20yo0W9dQwAPjYb
vq2DQUQhlQQEVpOwq7lfnVkqmClj8BG2yTB37h3aoDQxS5A4QaBZy3xPHoeEGx1qeomYdn6x0Ki+
XW6HOTQj+nKqoSMUHh5Xwj3u8QuxgfG2Vc9ATadOwZw1cYl2dEfKHWGmzVFcJKowijz2KEhNykKO
8QYBDHJcMAoR1OX/pHvIUC4LtcmJ1m7T9OyKeIpvg9WxjqNEFnCnu//Xp5RVoo2Y+I6lvsOdhLLy
1amhFU8TiQgMQg97v+JoCJhez16Jth/mvEzMWlDIFdprKY9QUwCLHX9JWTJVRWfYjDWRGfmThnqV
1hFBlJxXXFULa2NLTXj1TVqpNuHief/sy+R1e1qkOAFHpOKT14K0Cj3+l/haj0+5QMJxq2QiGs4t
n25cig2XgM+KDt9uK6r2NoxN8F21kKlBlw2uBz6H6qcLrlRKMOHovkf9HOX2+5KTR6FGJtQKCJgm
C43lWJ7RAfeJNXK/D0ZYRPtSDrTU7lXIfdWztdnq61LZVxsOdNpD2bxrXR588DzuQ7dRvak6avAu
reH5C8lfbiCoruBHy2SeGqP8SQn8LFdmOSwxAWWHZG8DFtlEia6c2DUwWG1ejtsiGHbsEgvkCgKa
mfMMqx0sz7bvF1NNn0rm168R7qEMpNfOjCQHoCLzQXxosF2oX3awBpi+MnahZfKzOB1z1MAS/tgy
taX/HKcmIM0X2F3ixf937U19s3Fm+v3nklm3G42g4/EpK8luC1jZQLcev/u9GtUruob/hMqXEFN2
RCz6CEF4URGoZBHnHODa7u/M8zVXIEFupangcJ92OVwXPd5PK4WcWuML1j8RPRHlGBi5SHEiF62L
lNdgrKV7BIhYnR5zKmCELlyzaLiKJ0NQKcjRXOT6QFEJUTUEvYlgruA6ZfR3aaMqpP/JO9Yb0eFS
8awgFFVgyRVKDB6vHfrf1VmzD+HAOZLf8lVj5Z86G9p621eDPHBfuYLXUxJjpiMTylXfGZscmEb4
b6DU6Zc0JyOWCXIbbURa53MQhnFQRVq48hjH2zmAoTvu+54Ytm1VV14HkY1XE6lVjisb0tJc5JyM
bvf7VLO3CDYwRFTFA4wMuXQ0y5BzxVhyM+7ucw08bohzX6PDFjd44FMZvKgsWR5XtY6mz/L9YEIn
RDZmc99nqW0ZIwR+LvjM4Esddg2mzOQk4ERbOMib36E8iRq4fVBMs36RXGL2qQdy6FVuVhefIEMF
GmY+Q9lq8TQJ74y8CcLcjGh04kSkki9hGXtddqfSHhBEPHD7iiKaBIohoVk+W9MXbbfd9FxmfM1E
WjVxdWq7DRnI13MaDwSyO83EVqGns0HnF4EXQ3QmTjMR6M1f/ugzNblECaX0YN1AdhflH4O2c0TI
VldYZJa4fXwLoHsAnnEjoDT4eHEMsjmUGmWP7vcwrzedIXA3IWBthf/wWTpVU3SVFogCP6T7rZb2
0bbQOVkOH3jKbzefu/KbD/6a7DeNWUa7or4ll3kNA5KiRtFB97ShpXj9weH8cbR4iVFrNvo3rEBw
hmh9ZDtcZLAhpCMMhnQxoXc1e2qQatTvDXRwicXtXZy928Je5ID2B1h8iK3GJSxaWumHTEpRgP8N
/kKDfdXw+oZ9RuXssdckdZRg2D6yqWBu0ty5guVabSLxZaxgbmfdAGRqpunOAftH4M7QKpvjyB/h
ag/h/aEwDVbFlvatPAg9pXoBe9DOczuKx0qjfZ8VVTnCD42mO6GJTfcE8veJSdIYuOetXer7MF6I
O6XIEE0CA5guvb6MxDZs2GsBpfNlXrlBjJQYYAy/wry4yarI5setpHKRnJ4PbC4mCYTiZOeg7Ni4
Ob0D5ft4T7/uEa9djuDfkmiVAmHpIHAogyyi9hOwvQJCmOn0/2svMS/H/7XHO68U8lXXbek/7WaY
gTJPyrdfZwVc96WAsgNu9TvUUkcz+Cx4l7cOt6DliltTgQwJaZILM68CU5ylhjzjWuN5FiNWk6HA
pzH/tJciCatwKDUX3Uq6qVatRa2e1vXboQ+LAGEgN4djGPcWTWO4r7Uf1GO/X2zOrJUDGEB0hZlr
1za6PqLEZUCKxrQVAzIYl7M6/Tup7ibsMJllXPIvPCjfQfMKpZtodUelKIUwyj2m/lEzChg/MJF5
LD+hHvLxqcXFk1HCyYTL7BvgmSxoiN5pAo2GUn6dog6H56/PXlvbJmkNBX27pApXrtacxziC7WPC
4sYnB6fcCpRK8czCPFTDpII9PfrUK1eSTkhpCStuzFWt2dTsTpMw5JUW1Bf/0KmHM8CTw17Xlwla
VUViP2dW6sXNhmZInDXl0XO2QbLg9UyUg/ingbrWu68QrOLNHBS8TlS8qUF1f2517rcK9HvdX/zY
Om4TcymDYQKpGmz9J//zXHS3VXQtjvpEXhiu35ELkj8gDDRJYHqHY6kA1Ut9MTbk8e9gaM5aWTKC
eOGZxEfJch0PMaVsgjxZEitCpa3G35v85L89AGNC4KCor/Jos+USMf7bN3+mG9vLPEXr7ePEZgw7
i0ljuWkTHfTAw1rjQ6kLSUX7i9eRHW3OzJTmokpQvHMHgoZwrikBU3F6gWwwCMG3Sn64ZiMFJegT
xI+MqjiD6IjQjTZHlfag7a43Nzsnz9S2wUd0TyAU/b8lmN6vqpLRa1l+EFwpNKwzrGLGTMs4VD9h
tvBwFg8cyj9BKhFNWmutFp2cJDTOewDeSW7iDp05k0vlhd2NaW4dKf79P31hSinbPVq4t9qnvcXR
BVpPRTmuMTahmuyEfzY1z3rzZeOpfaUgJR/udFZ7UmuyRNTE3tpbodRByrLTURpPysPHGig1G+ue
aWd8rjAj5OttIf8LD5oArKzDPX22q1I+2kAhNS2Ok08T9/Uv4Fkn7WG9pXJZAVDxU8W1eeSS8LUg
H1aRqSNf6v08eqx8Ib4ZP3HqAWH7lgycawR1lQYXJyoOelL9sealyIF6kfAOQ2nmOUFV/GceL/W8
OaQscBlbPRAonYvXxJEhUuIu9pKY3WY8VykDCTlMdV6qeoV7F6gkQ2FhWM94rp9zXepqEdjpKCeM
USuor1ZxH7zaH+YR9ZKesgpt8zZnIF99LPdRf/wz6rwQKo5XQmGUbmNsS8xNf2gmWVvx2cI4NvEi
vKrhZNDo6Zhf6dVKtHaXn3uT8yO9Jw1sG/j4eGWXhV8WJZPMLAaej9aqN18+vmV/5B61IMoHIetE
bKpqWUlal5JT/39kPVwhqroQseu6y7BiqfaE9vDYtnb7sBbSGwAahYqPhXBy1Q9QIHN1sJsKxjXx
2Ah7YAo8fhExSAlK8zmq9nSLM9I6aXvIWKx2ERKPuKIFNX0HlEgrlm5F/6Qu4v2+G4nCDKO6LXdk
pOvxviPNnS7ebx+yT0+om8+osfu7KA2jaM/yrp0P0V5FlrJnKJT0xAeVfxzcrChxt9ktzqC+9bAR
TvpWyWOjyZD/k/Py1Q5yp8BkJ5tAv8eFZFjrRXf47EeltneQR+ABt6aiZE4KjjqO5xJvNwcpCiyg
oOAP4SyY+FCDm/bkfKheV67RrUvZCCFyALKkjRFdmywuIoMluhRh6qjUFo3zT/R54FqRiiO/fPuR
FDDsDNSmZMkM4h8yUyIGswD8O8SWCRq2QWTJN2WT/zWxUmjW1ABYdPG8ptaA9tfWiN/PduEeC9CV
y2k7JaieFMpOKwEiXjka68vro2XYRXU9f7kJiTll17YoBRfJmiGCqcQBj3/JdSYZSav/kdpjqS29
+Vi1ApXdn18YJjXj6qpHp21cqnbFknAfEJWYXNcapZiJ/y4YkgcHcaR4Ww2G9hm3R8qlVcBJ7tgo
KOYzhrM7bBBuhw6TteZfvr0hTJAGuJYHK06OHl6W/D0rTzlI9R9Cp32yhhuHF4J9l9v0bqhPTUaN
W0LTf1oDQZAiGbL2Kz0zScuTHF1jHq2KTBrFvEJvgOtvtCe/VxwuUPlfZSVJiXRfXdoFYSsveC8w
c0O3nfbdCZvz99E1Rk6FtqVMTur6ZzY+yH1rKE+Dq8k2tBptol4Yox7d9jLshNqpzN8F/yvNP5iH
ODX8mmGMw71/SwEC8Byz5iR/tnxlGAUmF87edtJIbCIcdJ/PdKzS1OtdJMgQla7d+4H2/QDh0dA0
5c6xHdXI6jtCrVZ0BAgG/z9bYVUmgp2G501wcBcnGBFXCC8rGRXW4WqrKFQghxNNzdyukgrgtZT1
WCiQQ++N/MVU0SiwpR9/Ge8J0nr7ZrCpNR8811Np64mYoIQyw+pdzMwmhqK4TZ9VQd/yg5jQTe22
cjgqLALkdj0CKXMXq46Gd5Sm3ygkDo0yCA3sBHk7RD+KhPV15SD2ChWG0wIQUBWtpEYNgOnYMLks
hvsvoYjZatvzdYUUqgKjWaValfzIsOkxz51KxWJ3D3Qd8qvWgRy/t+NICB7H7y0W5wghOqBOdtM8
FmmezOWmlhDYzMYFKADw3O8T/n1Yd4KypHp8lNTJh7zjrreWYEqsJtt4faVY2e48Ns393uFISamB
9BvKSIhqoo5AWUjmq+q8oIEpPFQR1O9A6Kyj6TI7ojzFF+yqVIUDCTuRzfUuz0SMp3pO86KqB5fx
tV98HVdonw1iT88bQxpPg/SWdhl+x5okjAMIVrZi8IXWDwQdf9toaJrsqx6HPMb75bOiQEuaCm+r
xsNpCvJCuxxitFbA8l/XB7AQcUbY2Ee2J86X/GIUC9r1Y/o5iMlu28yfh5dhJjMsVLwBsNskTcbv
af+NI2JSQBKqs640kJhmG/edHhJ2AXtJrUNd11iQGmMZOAlcqgzcUeMrb8H/xrVhFfmwDFHm72uH
kWd9Vgn+i6vAMs/ZaCJCg/2F/PhYTTwdXHmNQARqAlEmM2hVXd6ZQQkSpYCpKkCZinVcN5cgucqc
p0zaxWAy992GuV57XjmmJcAzXdsbXgS9YlwqB3CFwbBrq9FIDbh6Cbi7cQB+3b7ZnXoa/EbGcFki
4NMQ530YblfI/cVTAjWwEmHH267S20hcxG9YVXTGkTPjeiDlgJe1wdxk8le0ipU3PXifWrIPSpHq
Qgu9oFJEned7DNU7im7xpk3e/vk2ySnyYwcwOrRBZ9SD3Thqz10Eps/1uanMiStmYk9mdBC4YyvL
ijJwrXjHkIeEdDzJAnlBMXxVNXr0hFT1NEJrASQcjbyxvQAghiqkkNucbPV8K1l1ZfxbyRahupgx
8IDAZWeVWL/XN1Dg62VrWnPmkLV1YtakLMA9v8GRaEnuG9+SkJlmpgzUljZehF+CkJp2wVjx0YW2
cQ2kH2g4kjCD9WS4wouHkOartf2pYhgXNUCe5xlhuMjT+jOloojGMyRIk/lmAUMxhe8YU3FOzp4K
NEx9zdVReuko8hbUw6nx3Jo8vZW0DuNAqVJvEdps4IvHS2zA1X8ROKlnfs9CiBZckgOQkDrJFM1R
NNiJuib6WJjnE3/9VHyYiJbUnYrExKvG/2imFqRg9DWehBLss2gIBJct1xDVpl/O/JFsVYmMF8UE
LJVJTdUm+XC/aHgnaYJ1BbCK5/rrauWIzjVszDOfjMGhkaq+pqKZx04U5gM62zNsH1KNKNWbGPg7
/Liu0JoMz/v4CET2WRP3pXY+oId1O7u2GvC1tNtfYJtaUcbOqKc1CC2pNIi46JN9kb+IKnF6LQfa
c0xqPo0yqyViLGCDDP5xJiq+vBDwv9dotzsKVftRjxmw3QRFV2YvSK/HFEVQmS3mg1mF2b54wpr5
Sg8mNJWwyHaTulHpXzjXyxCbxd6+V6BSjnOxRsxd7E4JVcYusP14ICWX8fRrFVpruMWvEOPLtj+X
nA9VYSDhVqj/ihg73rmKFVJdUoDZ7PgIsv3Apb+iGAtU/7jthdilX1KofQcX2shfUBEmjjDcFvSW
xvx9zVtuP1Z1wh0MWXKPNBS13Jkk7iUXRVh2gzf5UzwEZCaS4GSuSbJSQZlN/oEDSU9OdJSvcaSD
zDIGUOlA5X9h/a5tt+pYsWYqspyMRkbm8mvSBjtGiFVVF9wB/EHwgU5S4xrmNhX4kT7/s8svMXDC
oJNkD2aZb1rIGyMTXQSHN4CxgaqDiW+p++AZCyqU2nA69rJJbk0mVyQN+Xu4iH5vA7mBHYfwEl/Y
40FVYFyZ9p5W7BLLcaN2D54aa843jR+lveLyLrEl8h+zE7N3uRP8+4xRmHaItpnhTDelzq+WF7w+
hrgOn802fg69TCt5ax4QpYDsk+popmnxh5XvAAdYn3BstAwVlXoWToc/rh1RQN1QnGMC8fUJwB0v
NyEWbVCqu0thn0fbANFmQRjzoWvP5m7Y0tRlTcLh9KJ9PdwMkLlRAGNiuo1VuCnLj0yRNgYCfRYw
Gi93/Spkuqh8GeOIUO2Qvnqribmrd/wIzGpKk135WCxInFAyq/RpKpW5utPFz6+sPIERHF7Wn6I1
UsGKiQYlpKO4oeWKOA+kDcJQYg4Ljo5j+Nzb9hAbNw4DnRIejOxETlKlIFVGES4Kw7XbKBWfsMJl
1PyvBhVfN0gC25Cvr8hsWpUAG5jch+awB7R7BsYEEzEPpflDUh6iQ67GuAVuelRLPZMIZGqW3CL4
DEEqSI0SFzFFbMTamyEbWRpT4c8GXzfYKtNjAlu0IhEb4EBy8vmZ4wOqDRbF2eCHdMlgUUUwx7+c
cNazharUVUtmlOgzIR6d4fikArKLys6GTzZa4gVpHDmWwEksEWujrJTwPPxm/bmugXn62huBbeEe
5py/Yq5Q5xa7kn/zMte8A12gmX8J8JZI923045eoCMNSI6hJZPQU0OZ5qx1ZVWEnu73N0DsJSpRs
NrFORUYAQgbbuTB5rXKU+85JILu3Uttx8nkODn7s9kQZie3TgTM1ekiGTDkQxsVoWmg1I6NfQRQN
lb6nWrxlmJBnugtUU+EwMgOzmXRKseSMd3AhvEB5zWXPSOVC4bVuB9JDhfuU6Bv4vC8oNWdG3cNX
tMGFrmZe2Koe4L0SIxH6Jo7ONYxS9CjCZZwo5QWmY+qwMAAQksy9PcwTbyzE++b7NGL6rvTGIr7F
jRAX+pbNSYvtU6ulLckyQE9vdKkBKukpKK+bvXd3VEmnwMMiyKW9w/g2QCtqWGrgbxea2jxbjHRF
4TIGEk8nMDswgEaGlT8xViIuk/NLcCGgEhFmzvYSMQivOzFvl7JcHQeb3FC9XMzCNR/w7GGYi5AL
SiVdzNYNnFiJLWGYvKrXnwVT8me5jZBPokLeshEu4f7Z094OxnkQeZB+cv8eHNsiKAmViYmCqasO
feM8VIprZTPsu+KJP/gXRu4T45LGkyDlEDUV8Sgg8+qw2zaam3rKTkBvo6s2+q4WMV8dYUO0QHM4
cSFRMtdCy0yXhYlyXv93hC/A4n0YgNOFlUwrD+5Gasxif4J2Oqiet3IhdEJE6mlvTBXwRmZXT8ar
I9wIAUuqn7UwnN1QmrF7BxWntByyUsMdEla/ztow06I7NKu6/HformcYaF+31HM911HInDtKDkOV
SmIwElzyb0RnevNarUDVD8EzfGPPlP44N3XtE/YTJxkiKlHCCRctu5hZiRWYf9sLXMu0EHSeRfvq
n5YqdMBlsPPpr7BgpZPYlKE7DLd25IY4Fl+BUt8mJwXdjYi/vI90vGUyokwlglJ5oX9VdHnAFlzu
w0EhS3/+N/+nKEmeOPqNMs0IYRR/o7dzkgnJ3kPjZeTUdI0Bv3eipwYIz5LnFfMdHaB0UpQuFvHk
/ad0k1mQx4lM7i+JCnO47qTBalKA41RSFeu0Onfblq6g04M6tcuC7NFY60dBLpERlSxMC9SD185C
0m/MQvI6BMgT8jLDgEYxiKiDPPFxXRxfAy9cAlHtNGrrhMK5SNxImhBLVU3Y3yCcKuomCXS0+eAB
HCC4ujkuBW21EKVikcgA0K616+HvcjaIeRb9f7LnjbNhaOeQ1iEd4xsKpUJl+fG0Fu7pZwnLKRSx
dVZ7rTk1fQDlGYXtFrPv4vx+lE8i9yrdZnyJgDvliK4wdi2ac+KFKqdgGzNM0/dW/7sWiGzWWDZV
tl9wKpe5n+RTAnNCzgPSR1a2UQLC3uDzGwCfqGxoTMoalOzzCsGL7e0G0Xdck+rDmrfW+rRj1AIw
QudNrjOxDEKoHgtY7IkqTvnTjTqnh6mmBMf2HUzcMc0z3cTgtYd8pgDVxhY5AeydoBmMNfPdYTGO
/lM9J/wNGZ2YxozOStftJFpdK0gF+6ZVFLxgdA1SnUKf5PX9Xu3Ti6djoiuM1XEB1BOLI7OzcLoB
sPv4wKCC8Tq+P2Pt30HszP/oXRL3moUfZcZqw2bpqIgqJBM3/mNGAzl32JNt16IofCn73ZH8k/eS
kwcQJSeSVyEPlYQPny3VUDg9ek79bSNJWNlvdpTPiXxvHNGxslN8GectOGkhj2ZMcIw5fHsn/UHE
3bLcdM8D6W2DtCEa5VGsuqMOpyoY3PNrtpITGISIbS7reKkBVLddyKPUBqYRSWMetqmOVO1kX0Gw
Se6O7nVUT6D/i4oIkk7NqR39kuUzbJm1dteWCoish8MgtHPlHBOVWHi8uD0XkbQP7bFZIsTR6UHJ
ZiPEgrb5LUEihTRNf3h6fZAeZ5KP9C+5bS/y6qWvqYx6DdE2iVf8vRn22coc2PCQ1GFTt2OoXE2b
f7VEGBSdeVu40HmtrubsxXQvBUXBVeM7syNo61K65LETPhuJlg3iD9qPcnSGvy2vjDSHsgcI4ary
pfZUqnlve9ys2guUXRxI6Y2FEjus3e+wE84srfFVvkujlWHpr7Nh8KmYCNw3lXjkD22cw5Qdb7ZA
yUXUc7cMles59J2cS3PWSwdDfMCgYvHOUzG4OdhWopTM/Swkr+EKqHbeBbxt9J8EfGX/oyVr4w/0
w3ivTPipL1YRsQG0tvA3dRNCSs12+DCrDDX4kcxBI+UqGGu5HjR0EtXRI0fMfMRDnxYCcV5xzK9U
j0TDq4GZ+nn1mQ9tle/LeznBpEh32Wg/kDh6ViANLpZaDoVg4MttukMotIV8J0CcN2OXyRpt7Tn8
N8vZVvsS0JV+3MnXDLSo54drwRexDLzomIu54WVH/NBdz168g8/cKzcMPnLyvavkLE3G6ahzYZ9e
HGqkcZobvEkUC8M9S8bLVe6s9Ig3TmXFkJgdk1AZUrIeeqiga8EW58ync4EPYRo6bKwGUmF5G54R
uPoNJ/sUYBn3dpFrN1n6iROHqBMa2cYZa0Xt/OY7EEpI0FJFEi/jKh0x81Xmv5xyolOYOxQWRCbd
BVlq6vY7F4nHxFnBRuIOWKIBsbxuC8z5r3xZZlvXg2TI1wKiQGItcFxyspac14XHPKBiD7FQEPb/
wyd30GPTE0XCEhEtF8L91xc3wKN7yLUvaFXGAOOp8FfSvy368AnS7VRhLxC4aAD7rfeYdqmFacFk
sbK+UeXj0y6Un8MdPDZ65CTn5/fgKUbwgc7QZJ+2xv96M7twcFs1hgoMb0CaR6CbEUP0wvZuBsMg
fH6H1mLpqdvP0D5AuLMfOUIRa7j3SXPW7rHfy6/PVNsOzDU38NUjp9kcG7Uk+gJ6l2a1lPc2XCTx
Y881SiCAj8WQAHEXgIQk2t27eNKQsZvqCrRxizWQwFniXu1Uzo182+/zw1ZvPrO4CXVU9ZiTiOdg
+CfSSpeicYHMbHy3xElJ2qrHPHYwqX7KWeXHfxqpo8YGprDm9HczmEbeND5J+pZzUMOGBemA603s
mbasir5rt8Amv8HiJhkFvHAaAr1Vx8QnxLucqCGqN6HnjPl+zzQcYwhobQRufeOOXEPGlXu/Zo5k
6Exonf9imBrkwgHrWeygiFQbhkKViUGDgYxIRMYduGd4Wpd9k7q49UzJXOhbLQ4LwuGu+P6lTqXC
x3ZF5kSsziqymQcBB4agtvHDlg2C/iUfwlBfhLXQkoxQP4d3Lj2ZeuVTzi7rAJpgjKTKUJHxDX8n
+rj12c6i/lUl34k2xOYyMhUS/GIFHfy6QbQNgWNQQ7xR4Oh1kP2jkSD40bguayEtOWDqDyj0q2y0
FHrbbUVVT95QsFfmeDodXtqCWPD+1jolOeCoVMUnzmVeqqYdjOv/YlkBvFGUVzr0o6VnRfLIgSNs
1iof5plsyIUMGkwYcP/KBRXa+CNyEasGlu9F0/d271lGOjNSTNVToEeX9gCTrdX+PGB2V8JRktVG
1YoylYlZjJ0Lhad02R7OiE17xH2LH+TeGLf6tfHfr2JXtspacBaMIZA5YD3WBr7g64INt+gEmk+9
1+5mrrVIvIYcudvBoxlcrzTK2NkaQVh08KKzhV4d3hr0T27ZeAtplAXhWZjDv7Pl74Z5va4FeLy9
0Vuv9yP5NMeE2SJNomAMBMDmwONU6Yg6x3pThBxvLxVJ3ISC7TbdpQPPBl9oeGuyK+adaoJG7Vux
Z5lwX8Vu/FiVxulxj8Bw6GC9C80md3lRiu7w+qCHlGj0qGgFMjHHs4vQdnBucdNkY4eR085LP6xq
xklc1M7AaTumJ+8j5TWF6vGmadCOYsWefv4PgZICgyJl2TkCTKFYMApsLYJgzXDqcFCaZfekeouq
IrLTqZyyzKEY6kkHvQ6YxDqejxSHlyhCObaSuIgX12d4IEsIWxJ0ieJpwPjBvDxRQMdCknOO9t7m
zYZtuai7QGTh523O33KbOLUTi5iQ0+jkH6Kih46P4wThsBcII52S4c5F0jKE+JSxAhO3KCtNdSmQ
b1/LRfLHCb4lWRRI5edbz2njShmoes02dclnWlnbW0QfNcZKzWyWuyPHtewJji9XZOWJYxEObpos
n95ab+ZvYDaLVtnhQAvYnFFgeaHruR4ghaHU7U8rAXt1Q2EclsH0HiRkY4mQi5YaanwSA/GyVwZk
wlkr0U644Nk87glVOr+wy7oVUb8UXucpMr1mkFjm5tTpodDzCEAvLNrVFy1EgquTIRWhluh+QlI1
By6JUimpAPZ+ihj//9+CXhKsZyBwmlEf4KO2ucQX3pDSh9eOnSN4BORm7J9iy7tI+ZJoi1DD2fGv
nstBSbT/Gwwxa5OJokuoK36Om0vtVqc6D8x3S7+svEV8Nm8/dsQSbTNwWeaThkANKWJyZn5j4V2E
e4wSYtzUg3T5JhfpQ+4woBnaf+pd/W4ZOnQi32BoToyXWKGLezQYcWPu7vE5nNjxbOODtzOJzCS+
ewJZlSEO52I9Kg7Tr1bXknFGPU+PrZVfEMWO2oz0h++f1a1y+Brsr9esl+wdtZZBcNNbFVyXoQsl
eycF0rgJkZRJ7S/2l33dUHkHIfVhXZi2XeF9PmXdVKS/qbATrrPa9bYLSXBKXtMGtCHL9foDb1Vf
3XyRKb3vCpT+l9bjYbQh7KU5+fRYJATDtRciWhyWjJROh1X619r+f9tUniKtk86ZmrEMTv46AeAX
kkHqCE9DBKfyYnhsFkPYgNo2VNCuhRNjEDzNVAwRHeoNyE1YlcaIlrf+NFUI8ppb9ElgB9al5VzU
F0+rmI0sG/Sh1jqX9wUx0jPr2h2POeWO7UbMn8uATebfUF6fi5T/KCgUHuZG6oeZWYucxEJdNgtv
OTBlgY3HmwW5PYa4pWFiAy0nsZ2LWir8tKXJtvbe3Q40QD669A4A0O+waURe3LqUcKP+vjm70jW2
BZ9dgCcxyp8ZPibKTD2qb3UB61VwESPB3ks/lqZVzvKbLkM/INMG+mBJ9ZAFWF1E6r57EQXWVpiw
EnqxlKfB001coDXG90dDgYAV7rvz/rIOjdVtFX2xlyokWhzEUnSU1sIBU1+/Ggx1eg7P/IoyiQfD
939PYIVbqd8czIt3CmmIx8iKRl2VYmrAyAgw5Uw6y1CPiUY956OxpmCrjnL+368nyTaCNnXun/Wn
MSDJlq2cAdAPP307o6VpWie8/pjjaykQb1LVErJDcg48ZXFm9ZmxKe9ocmXfPFqTEcoyM7fivYbX
oJsFYIqb18YtbwozhXDYlztjfEyp7q0MSyfl6JNOJYpxQLlyZ1+ltWBkWvyj2cPnEFGl0RCev/Zo
kDQ3A4UI43GExjSu9Gu30mS+apXsmFjjOZEJUwVSmxwOH2njHfoVRTqs+JY9WseHIYc8aUMdI0bt
qaRzII2+wZmAdWmZTb3O07Dxw8IDH/Oj7Ov/rjNf4y4MYhgWP3vNbkL5NIn2WP7T3dbb0pJQo2f3
tCQOag1mwtuywIEVo52RYDWHW3TwmGwGKRZ0PnPsZpiO34lDW5LvjzGjulcSfJ7F5yxYQU7StQdN
+QTMap186ne8KeuAt2VVk3zm/gWkvwmLqBrMoeYbFGpdPGeBaSOKmiwoVusX3KrChS29Y8sO68JX
tV3mgsci0qRbNL0iOmM3k1DUXrrRdUcqTaxJnCKhJCdlS5582/xY+oxQ2krrUCf9GeLdAoq20CVD
uPAM1Be/XR3Vgtt+Rkyifav2JE+QeD9EM16bDSI3Ca914ZuJ+3bR9VZZZQnPqRaGMhmKAfNlG47V
e6Qjgm8Pt07xW4xkC0CGYAlqs1wxHqtuS27b0T7uzoJwzd4D+CcabpPMQvcv0Gb/Dz8sNUTfKEYH
wl1Z4rGdlxkrnEJMqPZtaLLt4MDtf9PEVduOb/GM/3tHrLZB/1JnNScgwWvtj3/YQRwkKQxPaAOe
lqyDrzNY1bbDGKTZ+K7TNlTrM7m1+Xu+X+oH7O3X2oD5XgbtgsvR3QYrVtLfSd/wxQFKWM/LxG1U
O0BixWvNi5xfPZ6kTAVitNdUpUJdpOIjIeUMkJWdOnagzaqRAneWylv2eVZk41VUOz2UZJ8mnaS3
uEdAFcQUJSShMoohMvJFL/HkKfBliMydZ/gkQSrR1KF/KKBunHAf22lvGrCCcpodHFnjQwkBvFm0
zQmRA+4y4KX3WVSZsGu7Z4spfSHl4v6VQvxN802yCpi7tZlkjGpV/QD0jvebZWrE6rULEY6tVQi+
+RPBuZ2rHmbvDof+0dgXTZnX+REtKcc+FxMZfGg6Z8YGysU/z5LqDKieiR4ZdZCHJT5V304RSzZh
AcfMZl8TZpF0AsWkpqEQ3Dytsou2cphHuDq/B63mETI6hjIcURqJviJkgHpQC6ouTnNoCn6xfJQh
gN2w4nrzhNR19TMBk23HgCCRncKpgoP1E4DJ78mNCqGKrf97X2qXsNCYbfqvrGXHiNQknEGQfZdL
ZWK7C7fqJB3oYHEgdxzq7h7Dpg4GRplVbFgg+rywpc6f9z73Osy9axTfx5IHHvHw2c2uZ4PBPGZ5
xCkQ4NCxecmFNUc8Em1/wWkO3rXORbpoMyFkgl2bre5XwxkBi7/7mqFMRff9LOAPOf8vQPJLYoua
MrUpXSWkaIzgGFFzv/IsNWpZ091+pM0w0XbdO63PuEoobnyPlpmM5VYBXuv9KzKpF2mnNtqj+HUb
YIn6u78LWRbEFhlQ2+mM6nz3bQVHbmPY3yW8opaaxQPKvSxMGVJNSot7WRyDUyAw20wqNLLYMf3Y
zFX1hSpeB6D71pzqU8qGtFRGFIuIIt19Gr7Y/xEby5fKEczNGpUViQh2kfCWDkeXyawh0Zb4vqIq
9/sDSyU7k5yJgLDvH6X/85jU9KnQ4Aec2HiFCYHFTMolWDdnLPugEZEW4YS2NH5WsgEZGbLYmLRM
ZzusnezSCyID+oDHnPnKIRSoq/Gi2t1ZpesWlJi+ttybtdKaFWvZgJa1vRFSFF5QUjiUsHdYLPw7
hblihcjtgQOuZUTOtLtRRCk+IhmJSuBoWoFziAIuUrDBLzD3m1xNqR2W+5p6ushZ9BzRToHE/Wo9
SxkGP25XA6+b2Djt8QFMCuxWzSQ6iEcmjuoOKqEJCgR89RFepu94pIpiITD1s1XLYZlMBc8hLuAF
RySM/EmrhCSUESSUCpKIBRzbNv71jGzEI2NkLHP3Y9lVNBBO5AwmaTdIqjRoJMctZB7M0AUou0Sf
Y5L5PpAn6CvIgT3ATtcSUKt0OjkozDVKR/fYCzhBysROOxNQILauXQsiN1cAF7vZ+w/nR8V/JIab
bQVaMm/enQQOhJNdl9oQsV4P0uj38SXOGE4Fm2AqaKnpEyKoveSiv2s2xRZVAZpdYWTFgU9OEKUI
feUKj/sMwUNeaMNG5+OjdfFPsfOKxsu527Z+r/pBLZEn1Nr/XLLhNHQf1XB3uWtPEAQnf2nqlm2I
kgxLJ4Viiw0aZWBbuJYtzPF8lWZZVqWojAmHhkvAVL1+69BeCbqc6vfklFlRsKaOwRi/ieGYZy+v
qBTph1bEnKi25eNe9fGWOCTL0b4+XdZSCxFAh00EbFgwc2QX5UFL/GZSOYdr4OpslkVFiFk8J+hK
OKtXUm9vCOm2WfHO6DNdgYrS08oxxcUALK9OOOERJWYAfg/vg2UKGAZKbBEIWU5MEwJSnVGP5ddX
hBvzZ2N4XcS2BW1IW05wcFNOnxHgT7y6wmDir3qwgnGEOE97+ZqQxZJ70XN7++H57raeOq21vH5A
9cFkZt5Lt1nliap95Z25nVHFVTGr6G/d/aqOeki64OsGhXZ/FipjEbduloXDL9RdzQH+EV5BS5pQ
bBa4np19ekuY7f8wLT1b/MAUdb4GNlIoxOnhlMVK5jViA0ucqInbuOhxmDwI5SRQRhDFiWLMN+bb
VHwlDbDgdYTz9sKMMc8rGe+jb81NZ5Ctp9PHuI0wqrXYBj20V4liq46ohR6e0YuIAiGNMM6ueZMl
3jR6maKdolWvPlPr1NnKr/EWZnqrN3yALasKBNgE/dEj4yM8whgmLQiiQlx4ifV9wW793vKgcGf/
G1ik51mi/w86c3DclMG4HXoGPIMlaT9EeJNeZPTqUAynjCU6I72As0O2nwrHr/+QdbU4bRLf2lDb
lJ7eML6FYtvhkZriKV4Oc0DtO6In8CzBuKWgfoYp8LWUV9CzyXcEfP2dVB9VtDhko8zT7L8Fm4rj
aCOic1WQ02LLDaFBmN7qROU2gzFqdlXPzEMKPFKc9EDgqqyHvVXZ9HaCFXyzff9SB7D+jD3T+iG6
PrdQAqA2WicrGO7iFuafwXZCO6MwGnYFjO8SkUYt3uBqrAstTeqH3XeJFu2f1h82hMzMNNtVbHgJ
lyJec2svQCLo9O2oZetRJ5GeXAQUooZ1sm20EQ80vPOvJh+xQKjggHVP08v87viZG7wBm5FtRwIt
Wxrqz7LMjPvSP710QoH0xJbkCQhvVb+WTa+DrxnNUj+Y+Yt2pdoxrDO9HPxajdon+Dh9AEVu7Vr1
29pVnzGQCUsxARWf6DIu95C1AGQrlQP3pmDjswoxJreIzASLSVHEWbHzInj3y6p127Z2X4dNtijK
9E6+CJBWsPfecl9GV2FjY5CDHqtvf5/CLzZoHNBW96CmOSk/Yr0ASNaziWqHmzgVOiOKC4uvo1n5
lVp2eiBrOa9Ik/8r/RmEnGa68PoGk2TQqrVwdDf2JurWMHtJAXXVihpZ7GlRZ0kw9/MyqBYUloiV
0mEzznghzf1LjDpOaSBsGob4w/n3SuPQWpMis47zAKf6x8l9nUGxT2wJStqlv6+VrE3jqMzfEWtg
NV4BFo24R0paEPbM6MypNmnVojU3nt5avLfJSt/nibT8RoPI5XGGnUWeIeCSph+e0RyOvQ4QKv9K
ma4dczoqgvmgiGCc0a9eg9k/JbLOjUcmzm81AHBo0Hs8/dZgqu2IDmKU0hbKykG5RxvKNyWk8I6j
x0i99sKxV3iJV752tqNnL9zlzwTbw02vAEfgfOblu431xy/wYi94kPZRvuIgOoWKtleQv+eDyrWq
ZppNDqT6L8yGWY6r9anIxhJSuJC9ULv4ua7PxLah8cD2aRgnXLctRH9ihkEAtz43qVRbdKg7AohY
QTZq4MvxJFNw/wnTAOpWtd57xkgYcwDRrbv2ZtuEmB0NWXu98Sx6WYV0J12RrmrJfAojg1t9iJir
SyylGSgqu5hdUR36++XkPQdT64L11ZiSuDEnNEKuVMeSu/7ct+GVZGkQ+oCGrIAcWq884xOCTyKz
rZJrPWLjyCtqp3meAkkoawGAPLhtmdrwxoXpuPgabIETJQQZDqfi2DY5q3oMhF3hWHithdJvvsAu
+5g6jaxosrPmsBY8zxY1iioF0TWN1s5f3QkhRQnj6WukMOC70r15jxsNzFz5BOCrfD0L0+WUbvKa
jWhHgyF1dE7l1dQHMc2vrT5x9ZFZ41nowxIk5VO5KdyrNDCPZIgT4JOEC2jHN6L0UD6TQDPYHvKq
XD4SFGUg5v4WFKYgT48p40C/tE4XKl6DBGULq2A5JDs6rKhF3eLGsDhTQ12UbKyZTrS38F2LQa6t
qgzfQ5Dtmmxfkcbs06qjQ3iU8aP2/SVxb1iOCvs0MWRArqJFYCU6m1aHkyuu/3wTYzSj2BboajLX
Kq/b2GtyQSvcD2VJ8lOcUuhfCoevFyBV8IlX5uWEdxbN5RkRVZKUyYuS8Ozx8V3TqMtIYoBhdpVA
JGLBFSv45wrGGgIWxxnZyC+BvzxQClZsm7zEctqWKFkpRuPd0q4wSVEHqiueiK1f2jzgS3WUWfIS
C9GjPwM90FQmrfqE+oscMQ5xole4agKlCXaEwEn6Tnu3iq3CoAxOH7dFRJyZ3T+N9wR0CNPNYu5Q
TBPmpAyJAS3tawo25sv8ssuTnLHqbyBuCaFAUHPxvVHCkMludGdDBPbQvuxLWqrKi/oHN2bZB7VG
V6W0uhlIwF2zSar/m+gyN9Se8k52aV4jpTqd+s4PhY7VSNzJqTsAPbQDfe6hGxLU0467QmxEjy2c
iKIh4tm/KCP+zTSMJcIroujWtVPVnhRrc0Dd1zNIX2oOxV0ANHsgcrSNqHI7QnJt0l1xKxy3w224
fXLUi5UxPhZeTGTqXzwn9Culc0nCI49593n0phlEhXYZ9ad6CwTUJTfNOLbcb+chOr/sWcNYlcY5
XOU32e2SlwefObBiTtzHrFFl04MLv1MU7kTDdSgeber+U+2emT1/iingi5eMHrp39b7Z9KgQPZVn
NNvPAPFxWlsVsdCVTVpCrOXZ7K0UMPveFx0rkgRL0Ccy9I+Mbfx4MhCfKBBILe3ioGxMjy7xmwWM
8KO4BAtm0dVDELnqGHtC5ZPtrpt+yZ/AkKXtPp1fLpaOm2FsAk0/hA8zsBxOEH/HjftDsHb1U70G
B/IVcosKfOD/kKX6vNHFVrAJPYIPwCy7Hm97WsLhPmk+cLd9QeNZcfaRH9+vgslSk+uPW595ot4S
lzefo1E6P46ZLC3fnMCMtDXSHqXbtDGRIu8HjjX0qWe1U0DqktW7B1zSnl5x9Qp2Z6gJC9ScBX8N
lypzgZEbwlT4eFQsLRCWoQnSQtlAWYSqIj0/HouBHe7BX+HJ4zMF8yl8kTbrM4buEEacMunst88J
LeD+oWZI2Hl3YSRK/WcQhIIoBLXpthSeGhqFwrtKDKNfyBXQthhadhDlSO+sz5PAuM4LmqGcM4VS
aUO4CcV13nWW693BvGRyVoB1Sr7QlpNIY/lwxT+LC4+FFFuTT0cSwVpRWAY8gw0UBe6C3bs0K7II
HYWkM/npu1+tKDr67lTkX9gdpWJD7bSpdZ8blvjwlKnX/Ee5k+HXuTkUuSBAE9b/JNZ1iRuTgvAa
WF9DBw7noxfd9RJxuASMmO0PmPEmqTf/IJVkvNDjUPYLWtyjS0uo+IV42QmjZ7zP2DsyFd0GZ5vH
XsfI4GYiE70BnYev7DjhgK80q34xz4vAfkCQ+yDPEc59sj6tw5LeMFYW8CeuZOEfbd0Q+gIoqPLM
bFUL2nJBo0LXbmD60Gyt0hLdrSLcPpCpIysNtgy1EC0S1KA/7f23/CoTGi82vNlkitFaj5/XAbmb
dx3n62cvihhTqMrlT5WhvrJZGyOrNHx6DK7LBJ5aySJG1/82AdUJBgPUOMZqtnU/shKFiIr2+a5E
9I0KIpgV0UGB539Eeq6nZEEWrYUPAebK3/ekUCyDGF2aiPPTa2zhkdeQAtqSgxLAIooDQGijuc4Q
TZjBFNXc5QkE608k8qiaEbYOlFSMtICJK0uWCguy+4qI4WrR5zvHBw8yodi6myzWocArP0zF2TxC
2Zy6ZOdxuCw3tiCnNH489sWiSQLRVeikZ5o7yHn/qzDkRWC2S2v3CDGQUIYZWQc44FVD6EVxaais
95wPbDIrYOnvAuljOg22GIZSFSw19ROZ9VN+R+HJhuzEJwCPm/WMq/TpJLvW9TksZSWT6CXxCzVP
pft2ww8ZWr0UTfkXnTxks55s6AV6OEHzn5tebPi81lZZlYCAPowwk93+osgfboVVKOCYcxe8pNGZ
Rm1JMVRxdWQnZ+9wJYzEy9MSTY3s8m2kmxIY1Fk/GVRlFknWP5xgNTnLDdECI0Ri2XuFvu7LvbFW
fmw4PgOt7B4FGTxqlEwnd63/SM+FHuND5cU9akkrmUiMvxLnF3/RvTQdaRW69MSgvx9bjYH3parV
IDq3AbVwki7IP2imkOCWFoTIzR+QyTUPBSiaYMZW2RovEk9DiK9KmgvwQr3Q8oXzEaC35V+DjB14
F8IHUcg2LlyKDZ3VDMvGV1t8iibkKlyjebUXX3cdgOvk/2EL3ljdEhrD0gBZx7WdGGYKaBJxXPti
kt2NjFj9Gy+vhryB+zwpHMeyNkt3u77/8bqBAZuKodHV3wG3fJWjer4RC6gzR3Av1TPi6LQW3T7F
ITH7HcSmaaVtb1tMkhxscnvAcCDwxnFeM+/WuW7eZn5BMJiXD8HiXL7+AbRuDWPhVii8JeBNJjhp
9HOaAiWZNt6nqknfZAdHPJTk+4QpzvUPNxEASbvpVu9W8ZOERGB3zAd99UIIth1YYK/WRF8X6Lz7
FyAPYdbF5XE9vBiB4QRQz44A+cJaf9JXU4w6QtunDTTEeKztoBrJxgkoK65RTsU9HCm5gAOmk5o+
mMZ68nByu3e2+5zamUaBmDLyqtvxTcy/Rz5jxOGHlK9QYUqXEb7G1OycIgGu5+xT1JgaHhAnuMsM
9BgA3d6/5bVUr14x9SaEuHpTR1bY78oSErLvMy51o3WozfGFsRCDfY+6UynwlBOeS54amZmDY82u
X5uuyysdpi93PKkpROmgEkGGPb8Mvy1OjNhV3ARsEyRKpXPQ49mpt3jbz9TkfKRq8Ub+uJ8Wk2Vf
Eqib1B3whEhYIMff1nE9YIeSOS4WkWsc427GQ0sHgwxQqDJc0KXtqC9yeFrk9V9swFIV6ZLl0K5X
AAamA7mHwppzZQ9QNZlF1SezWND8HWu5R+0H609NI39+0LEUfqYo5DW8C96mQqJzKjp+29nkab6N
dtSkpjCKLSpN4vaJy+NSbcQPgyVMVrQB3mcD9QnztbK+pzVEIog/vB4LgG1BpryUsfelxulXh/3V
RNtll5qExA65B2EvvC9sXMCJ+So5lTvOM5IIMEMsHzYUFlS2rC+l3igt+U65yJSl/LW1I9Ue7IOS
t0SnZju1KsORZXJWjPIKz/oYyRPJzLkGLVgylu+Ejmj8wTuyFOqyK8Z9kFPhg3u0HWl9bqoFvJTs
QMim+qWWA9RwxAs2BwAa2W1QtZcxQSbxkos6z/Hlg344X2+ZybeKkGgUCsH0S4mrXGTNG6+cCKhT
dX6JHOmk33n4I6q+yimAHTc53tH5FkYLzK/jj8WOwKNqeEyn7hGgzb7lR8zoecF9UBVGWhiR9FmA
l4o11vhhiAxH1qitFDVfK1PavY9KUF9qk9BG0V66zISv9KKMfN3s7uetnfEmgLM7waA3BT+A/tNp
9IHYq/ItRr7s5TMi/ogeANFUtTF7syLa7KOrApTrLA+p33kf/k/Biyb6aZ8zH/aFRr8qZsRLdErm
d+7wdKXYvaad0hwX/Yz21DM7Ii//SdIUPxk0M1GgsyBu9rFql0DMLPLIR9g6Xe18KA6eyttgAupO
odflagczk9m/tG7wXlFzNOBX5iWz6bFCgBsNpjPJZs2I6fQG9fQtf8ZnNJbVKEZsaTbjPBu9hxvz
pav0f7HGxrg1Z3Csw/QVslgHs8QyHvrDZG3n2vyngRADfT49biI0Q/9ywLWAy7gm4y2qTtCQXLnF
1r3LCA2L6/EbdwFCALkMyZy2QEON6PSSSia0Y1+7rs2C6as6WR/TS15nbQBNPJbjpgJg6nXs4NG9
Ekn7bAM1a5U7SdExBH/SgKqhVYvmjqqRQrOev5fiEyVo/kvAzjzmUIHmU++6X7yjeIAq+FvQWkGa
Tv/1bp0THzvOJoIIY8d+zdOWy78Sm2xp6Af5U7AKpEo5Yp9SWjSv4ueOO8eA0XkulYlefMIoYQZQ
q/aFtMESaQKOahkIvfDYo2RVZ9wcl4GAh0O3kjpPydkhPFI1g9QeZTc9Yt+y5kSHtoXYdm3U5rAU
3SMmRlvm46oK6SQY93rfYjRilw4wVVRhFm/IFdqQuS30BnAsBFMJnQbsAkTdgj0szCl5/UWxsdHF
2sAcdPuichJwQHsc7xzFFsqYPavVKFVLQuiH9sl852kVicKtvWoy2NYOx6s4We/fgwUPx/vdPiA3
dKb9EWiciX6GoiC2OYtCZYJzKETvqmvgpa0KljIor3nPv5ZmOUnjsPiJbvsDW9CFryGKYBv2+SPw
3SsFbmx9mFHVwLBCLWlDI7IoMn/ydFY/DKln/fzzuNH+AbwnQCxOXWZl97yWsbNogw3F2y5MpfNE
WrYt7uPVz1n7TcuIxSw+xeoHOojfKmoHLj9OdsTiAQtdR3w7sSTUibxPzR6pT2swwb3zDbQFOPMa
/fI8qfS3+/ixwmxZK1BVb6bWyZNQENPGpEtqCoEBRPdySY2xeoy4c/X0JtQqYuOS+nBe/FrIZBcu
pUyao8KREhFuA7L26PnyHlMVwaBUBd5fUkwXoBqE+4b8PDYJ5JUeuu4ExzKZi3gHbhk1PdmENQNn
km/lU4FDUxnbkw6RebHqtceH4N/9gazD/rUFIkiGQDzneuVLzXRd2G3EbWHyoXQHIKPEEc3DP6Qu
Dm6aCHngxUTp0bgWTPKdA1ru+DgR0cKLSl9zQ8TBl1sLjaMbhmGgCOH4r01nTeeuHZrF0XqwRsCF
P8HSSn1k2r1cGldec+nbERN9Zh2/l1nwULJSXmP+uN3bY2J+oNSMRhq28XbDPbcN5E87d3i69aEU
ruAY+UMn9Hqnp90DOKNHFNol0GkbQWOL28LJ6a1iUtF1HNFzCps2j8pfDezFmKMYC5UIVMWIqysf
dPjWfyG6IAxJoAKgaZx1Qf5LSqIPLYJhRNpwBFYLx4/fX4tlAY6jgXx9dXfx3G2QvcFzD0BU8flX
ifMUcpPCzFSctt0tUiHY1xH/qOQEltt+I9SLD1wRUf6QrI5umLxIESQDGmKrXh/ysciAzgCD8bUm
McTunGMj0B7drl2+PXbMRhxdT6A635dOAVW4an2XtwsFEn+0Ik5Z/SJazwHfrFxJIJnsIT2P7y8E
GCY/AWbWdbNDOlOM6MG7M3BaRQK/nnEv50grtIoJyFtDPaWr5zg+YUYwsTaBd6JaxQ3neeRltpRi
ogL9l+zEoBbZm9udOPhO/l6NQNZ+30EDoSoPejWuHssCJZNlY5Ibw7aPoEzfi+G9G3VLIa7qJ5VQ
FoAS2Nk4UKeajABNqPvuKF18dCjngKF2TMu6l0+nUMqsDmFQLJbjsUKeAAH053Y4IGvxdE+r7pyP
WmFV453YMHa9WhhJwHJdd6xq3wj3I9YJJm25R9zzGIE3X7KF/v5f6xHRpyha6H7ewL7ns7RoNFr9
XCT2kJJz1c78yyHFb9mrkhH2xFLNkmfu/1B+H1KyphN5vwzK8xvKJ94YONp+QqfQXdqKLMPBORlU
6LBYl3hfzXc48TPKKNVCivfJVJe5bmSMMhUlSdXVn63mda7MiAoy4UVpdvW+aC8K5CiiWq9BP287
mfH8s2D+2ddAoZLnCyn1Axu2MSOurdK/88s1FGaDJRIOqxwtLVqgGy4JVUbjv61fY6ogm1jU9J4R
WXLobDqGAUNe43lBtMBNT50Houup373VbXpkLg/zaIy4q708IXfb7BKmn5T+Yv14nNSx2MCTLgHH
zDT9GxD8BFM9GaH+S3E0YIjnQGtbzg2jH8N0JCzS/NdPAV8Q290TA3NAFOUTPkQQCXNoO8SXHoli
iyb54LP2/DryxL96tJ4vrYRhF6UtdSdF3Eyi4yKdkBab7DZWl6cAh0oUQeVjbapDPORTMKUsOU69
hIXDOCOc0IeeqyAupJ7214nJTrEZSBmZcuxlluMNJkJzNvzQfRXm3epxCoZYz1ExF5JO6S+9G7S1
ym7z9M4fV/u1voqfM3e8eLjJ1Fm9REn4PYzUTLxpVxkgKfJkVEmIq6FdK3tZPdcCHooUziwHNmOm
5cuFVXDk7jARCRGlXWI7Dfli0pRoaenSGfpeWOudVEQjDa1iTINGusJUrArvhdadU4uWMf59zjQM
xKRHTrodGblblLdJTYxIR+eVk2vu6Ekz+y0rc+SqRx/PNZcUsyd21G5zMdMlbskpoM6dMmVdQJlA
0lWqb4i62+JguEgDyUwaQwwdSvAEanIHRMr0xBj8DMRIPWo6XBHpWJl5exCgdRDuHk3EMWGrBbfq
7JmXiJafk77EFqt7cdQgxRLtM5Y6lsP6j0UlIrUbPx6riVXu+34IJisdM9p4OZSDCHHBqpSNR6EF
IboC5LbtDENcppgf5j3sjLJpGaLlAb9Nybr7xJgJFKdaukD+GXgL54LKbdh0dWWNeLFg9ZOUVUq4
ZHrBmApIPZLIxrQ7vzy/picNfakeVmCtfmvG/W36C3y4k4Zc5UZ42sifdGNG779dvV8/YWABjmfH
tssfURCNQ43TkKHI3N+esLevEpFoe+EXdhFNZahrCfG4ZllUTfM4og4Ialh2ri2FzmJlcltkhA84
y2qI25FwKw9IO2v7Ib/Tf/O46Xe/gkd0rU14f9lwNbnmDmxOP0XtipIHuU+EuXO7gH69R/78mmzo
/0gEaSTgXllqVzuDcl3f7blIf1kchLR8U1RynyIZzT6oSLaD4weUF+L6ggaP6zZ7gYDK+nZBKa6Z
9IdQbY5jer7QT0naX0tIj9oh3RleG22yuZZoHf8rbOX97eWaaYLROA1P2ll0l8617ldYeFhLQitu
p+thGb98AHYjDrZdsK1m+kD05DEUPDxeAasOL8MdQ34hHsQAxraWC+7jCDZSgT4iklwX70j8ousf
iuXx8g4rrlvgPQyOWJlIBvr1OTr9abuPmUR5XXSvHElexHaUJe4Ky6eMV4fcW6cGas1uZVDEB4bg
k1sJHCgovSNB4B6yXimNPp8bc7niEWk+YAtoeBtsSdFFc9A7sxN4XSYFfIv8ZWDgx1OPhYcQmpcn
uHvomLVPqSfV2/0vs1ITob9f6M18MNhs8yKZqWS0NZU940ufu6xZ4Dca+sdl7DgG4wPxEB17GCcw
JZkRJiZ9cThE9UFfObmMFC0adA+I+quBJrkNEZPe+KYbawl/BuDaAac4GWcZpncnXqEbsy/0SZyw
8PTrIQ76lqwaGAFgl8zltPDV3ckR60UP4KNmIS73YBQ9MFifZIp2P8i20C03qXM/eC5Pq8w+kmp5
yYXjYfm4j4KBOC8l33rXKuP2bcp76P0sIP8dBrCW4oNXbGFCGILLxvGUqzRewYH2H5W5Jvm6F7LK
fpBTvHAiuxMFeMCzCG60ZzyDs0OPK+imSfBEI2HoAVmOmBNiXkf87B7NM548yPRL8FJBZKWVxBLq
sl+32uWfw9Cf3FoX8H3SMgATX2phn/+sYr5U9QseOELVqAn4ZyOPjXz4QxsgbuKHFYDwzjdWbqbu
MMHk/thzv5HQMWfsC+rUG5mpFDP2nC9MLRoDWKRFhE4DgdN/cEH5IjMx7ng2p4YxRmD5goOzcNoq
e1SPLZv0CJX7x82RXsghFj4Rr963MKmjZvBb+JR3N7s45Auj2eIU8XJtrGi/PeeaPhWA6HNPTKHD
raEbpyeahjuDtIkTZC9GHrCiAIh+9LWZqxAe18dH52qBZiaqE7wO0dNaO1JDHAgmTluXuOAiEZAw
c0dGfu1YnYF9/hIk1i5ebzV4V3YQNPLpxMrfZXaJmoIJl7iKmyyITFt22I6Mj6FZktL1k4sIXpG9
zlP6Ebbg2Z6aPIAy1ds8jZkfvfmM139sjy7JON4JKpzKibsMsI2/1uHFGiNvDN+3VzxAOS9z+Mms
Hra/sQbZ6D3qiLt7Mh4E0Xtc52oHnFrygOK8xp9lkkNHzW9tMYzfU2Gz5l2JZIuinP/IGc5tJMCG
XvyQTiU2ofgU9BfWbjLHD+drtC1nPserN6JLyd9hrRIIxg/uG5IMt6+Dz9iZuMeDDJkXngTu1KIv
wuh6e2f0XYoUa2TVU0gKVAtf5Y3LYHHwRWn0bZzSzUoVzhorz7MmtTLEIMhe+a9sWCJUvIOQIo72
BdO3WBP8Qm9rYz5lE1aha6zyJFL78k1OYX18KWGRbfaeZR9fLw2YEUS7Zt/J3bzYcJ/CWeB8IXJH
v7vZHn5aEMhq0DRJh/VNzRDfWjk1zKL6dcM/b8UPNWTe+ooBO9wlsRLFzWiqrPPriLQgcNeeze92
UsUMPgTlWsFTXgRJekxouC5NVlTjABGkd2+GoUTcY2TAKOI49aEbtleuR8o7M2tuGIAHblND3//V
8RTPxgrO3vdqqL8uf0JLtIKuyc40GWjzBgzlrDce9qBELc8f6bq/tJrFscvU1G5fSnwRRTLahgyf
uuK9KrEi2UVuGLaUZzZeFP5A4xrr8atBpDpjeOkk0X1hr8/gbfKVfGHJEaXsol2quuD1LD1JkuPe
LHozH67ZshPD6CiDkOkVsoOdQCI9uQAS/Wy3eAFYoijMuaB7WPpfZAoZCrJGwMPphFWspuWwJ6Hl
f7lnd6VVrYUYbpDtACMh3HxOZE1Piz50xT340qZEKwYS3ENgRipYtyDhu9xKJ79C0AT4m6/7Cef+
yCvhxNjHknhQjmwwvyrqPv8w8XCdjNCDOwTQmF5muVjxeK2zvREuYLROoN3QLwZkYdI6qK1BFDYH
6hk2c8F/jGXvCWSWdRXYZ1dO7BBFgiWMgPLKOcZgWE2OCMxd+ScTbCfdKyoEqRAtuhe6E1D6608N
4pSrz5ksSy87vx6i2cZC2fKOSn/wImU0+6mHoxMYv6KdHeO5V/a6dbYqV3NTA0Na7wL/bDmo7Y2S
O9Z+LYNFehOy7M3reOE8kQpZHqm9cMyKrlWov22JJVR6jzyxjg/4TPyHQ1JdOTa0k158M0juj7KL
ijC2Li5nACYhDVhUp25hd4MzhE6KsZW6KE4Z8Au+CAlFUKcePk/p0sGDJjTt3jyHWsh72qKfANtH
dITu36KsEVOyddwmO96FCrzvv/kJ7nL2mgGVAUVYK2JIhuqs54khDpU8x0jLMM9dKCbYdNLMf4sy
JOCOm10+3OWhk0V4E0Rr4jpmhGK+FA+fPlf4d+sDbML1wL4CfjX0NktAl25D+a87PddEBcsY5y4u
oR1jkrZVFugXC320LPjYqZoTAwGTg86A31r6b0uOrZ0ElIK2I32Vr6iKK4uL8Q+5aWs4WpSgDkZ+
Y0Dj972gUsQw0x45VWNVraYzqTnXEZK6Y6XBYg/BgD7ynuIDrblAzB8UXwo/pi0YvA3aNl8uygfw
SCMkbTZDBwA/Wxh3NmtcKrTyrK+YTLjLb+ITvH+aNKyZhZwRwAC2fU2jFrjIDtF49D9D4vRONXMy
bRTHlF+lqJOOuUqrGe9VIPDWjvvOZYvpvMU3pb16uyNNBSKoM49ipSRGvhf+YLyAq4Ikci/IhGBn
jD87hucLDzqmUX/RRAgwj4M9cA/bbC3RUfaocILpl7X0vAr+I3ce2KQ7rSZd1Om06n9Jyq2GLwf0
K/gDVj5KWCVbZwCV6NI1K7X7mxaYZzPwKIx4yQ4aio95gCz346fQkFPvj0MnqTsdOF9kAiA6LWFE
CEmFgRGagyZV7ZfTO5R5eqLuc7uoFOoGBk1c6F9uV2NWF/K3oUk425BzJxgmhyq9iFB53tGg2xUh
18rdLPzaBYMnCiHOIXDXEQNbepOFKCjcZgh7e+l6DpGkJBlvjk0UwUUTro7CN43yad3+L5IK30vK
y9QzDZ9Edh8P5dwOyYD/OQf5CeIkGFzfBlIdBzyVTvPPbuilQQQVU17k/X60aPv/6q2HPocMtdrQ
wA3JkWZAV4KAPrhN4ulElTdHW6ebZCsBbR7FpsPmJYF7/WkGtZX9v9is3yEViNdqSxIJCqmoDOIo
iKpMwH4NJsQmrzlNK5BZAKdnEljVZfRk0EXhS0f24IYGeP2r3BWC4SxRbMdT8e7pIdK90nqC8dvz
CaGvTp+ToEnLCwmuMD5HU7zu+dOsog42+ALoW/NsxlXLOr5Z2TxD6ZhnwTau56jw4Sy6cPCva/SM
fZVAJ2D8L6rPAGTEdPeZgQFHqPaz9oKOcurWMO8/enznH6F7lQhwovO3DvnRYo9BGicx3ZeN+Ads
illGOnJkf8dtEV1rPpSmG4yK6hM84AvfSJE8Nw147HWOEhw2IbNOBgzPlbwloX+DB3VnhWBlUXRZ
CXvurBY9zozhkJmUcOXJUDKS5cwcY7cKh0BAnThYfLtV9KCdBDI6xYGYZyASU0JNymKBVchCUFa1
ct6aI/hhNBWSwX0VbwWrvU1hYJ47kLgvTKMJcLEtJNCVQl2rMIrAk0sSrXp4vdVDK11Q38vBD6XK
XxFn9nZDbwaCZ53dcNe4NCgT7loVoSTbYseIYIfyh0vZVMtuWpgqjktcNlZySTZnD8kJfRrrFWFx
N8Xt4Q1aKN0H//0kF5IxsUR4gxM4WPvn6qlx6xzZzYM2yqRtpYP5RA+uJ/ghXE8mF2dJwNvIau1v
/NQ6bMIam6jfYbmCzE2jJkJrnKLZaUAaAeWasvDZpawA/KbfkQ8RNkrPO1a4QYoExIdiqLdcZ8Cr
JcmHyriCU+K3FuWeL0sURAiPti4DIkAcKiJoHoAXu5KNhRhcaURX/HxqSzzSO1inWRKtr7L2cOKS
1h+Z4GP3/X4MO5j3rolRcDtNDsQOO284hSjy6ZRRxe1PGtpGK/72nvPt8GhzwPEoMJTsJ93Ntfut
ZBBta2HM8KdNTNVePAjLh+sVFhHEPlM1XBbdlo98v3sZwewjpnQYkN3gpUvlfgtdX4UUVrOL6+7o
0IQ4U53Vlx3UYL18WeW5qFAssRfaCMK1JCoaDgMEtvFl4oyISreiHoKqquKpxvP2EF2mQ1SW/84u
NxM7O1DQoOGAQTBL55A/T/2S56nIPDCUF5VTjRNQOHzbZKs+xIH1U657+AJNbwqWtF0ph8JyXO1V
rrHHDUJDhfPupnO7zgFSS8cR7lLIq+EDutY+eAxRGkWDDqg0SkAKsCkOPWdPE9IC3NdR5tDyre51
MQ+ZaTH+2oorhku4RhYppJmsKwmSf+2HHkuXcVU+E+a4DXc3zmCDja/Ul62aTaDVvtFtSU4PkbLZ
JU6SSBLDExN0KlBCtQpa5ncvLVKB0MflmuiizM5LtSyVvFmODmFdfV8tpdMhkRm1CbVBXI8Cww5k
dNgjlcW+94Dq9EQqO7EO7EFSH23to74GJzXaNO6BIhlgPsmolcPFLOO1C6YTIEl/7KOXAYo1J46S
sIK2ARx9IcZC1MxatSJOV3a1R913lmdkIb017Q/4HeU8le9jaLkSLUK25zi5VY1RzAItw1A7T1TP
kOADiG0v0ejQ84rOvZsXhmnOJuNZPiuwIns2k1UW47D3VTmLQUs0BZv3r/CyvhwSszlNyESg6cuR
Z8ep2K63LCBhgERUmCReLtOPRHXNx8kq6dLLWJhCUr3RJE3QPqCU1gJRRXpCklMgT5wmHEd7wAqc
Ne8VVRKuUzgyTZPzFk4KX7kBhQSKtqLye3HdZKtwB8TluqqqiYHDd7M8xIkC64bcrWAKHxCatj6T
WTLTnNc/6t1FOFM5cFFkRwzlzAJU/cUJ1dHhYAsIcsuk8FSdEM08l8xVs/2AgKgxFiyp71rXrzFY
dorAHOyr4rbcVA5IeGaL3D0pXEJJjNsvsvYjMtujqiqE0cgneQ0V0MIqT1uFGTrn4sZyRfCgfFx1
byQwBFMhgQOb2gKwn1k9qE+OMfNnPfR/WOkKNJEurd0QWhs909LOp52Wz8y04EVhHLnFs5vjp4Qm
nnjNZYPjtJc7Y4c4a3r28D7UyIbXVBuYtR/L2aIszbwBbm/MvCiS+dyLFIxzjMdI02D5i76GNP7T
GhQAqSpocceZ7f2V8ehdzfhFCECRKz+3CjBybZZq6rSA+wutDF2pejMFYAK3Bbviw46M3i43oY5N
5BOBisM2pCkcywCLsLkTk6ZiIVF8bEN9WhFucvguQOtTcRB/ETV0UMN+70F4LemrOnKcWaZsxu6r
HARhtSyDfrFkNTPsSxEMs0oNcAHur5I5Pi8SKVdjJJsD4YSeCoGk5K3D1a8bRH8BL2dwEgWmpJhc
A/ZP/glCS7U/g1W5wKoJPqCh/D45EDHRMz5jboIGMxm8kYVmJmzImjlYsr4XrMJvckQ2w2U+WfOq
4ZEbjiGxI6G1YIDW2EMCaYspuU6dp+y0BDFsb/2EQ+aOp7Od5Wnh97HdvPrGXqS14GST5avoakGD
YfEi28WIizTg3nqxDMjP5nYXSVA0h7AVzoy9WC/SBM+X1x56HKiCIw2PrkldB64GKOv64Ee3xzIi
C0o0EsKVBzelhyHjCCh5Rdi0tWYxhyjNeXsruH85M2xzJwoIWrRpZtsYlQ1aSFnIp0uyZI8AifLV
FzrxXW9dWO2GohJRGBABS62+ku6ipsV/5/hYuL+yFgmUzDfnUujsFhWkNVdjyz4ThcPpHPfXpBeq
h06vn9wVj/fdR+nMjhly39rUeIYh2u3BmwWVkPQEd9Q4F/jNbkBnYDN+LwRZbNYmdyevjaFXoYOU
LHIdrh4qTzzh4MlAqPUzTxKV2ZkydqfNJEAKl9lhzZhrk7335/ESkEM7u6YAILQLHvOLMSU9jfyA
utQIxYzdyrSrAAUEArIbP/IYtHA5fkLgERfwhNjIda1EdTYGNS8Tx6Hs6SHdXakDclL+1eE/RDs3
aVskPVaCaW4zKDpROKStbRBcuuRM5nFbvkLr3Fb4N72a04CVe7NZW3zxz69Jy2FUaPOnu/UlvE5u
/C1tuU1IAdsHgtA9PPyUXGTR0Bi9ujY2RlQ3ogxrmqKd44dds1WXLVIDN40DAbpPUjsv1RRW0udj
BiLw1vuuciM1B+AWuD2+1+BcTEoflkBLh/SCwdi39nWomTRa7boQz7AjrlynuZy23yCJstkRV7bi
U4V6zmoTKRpN32O6IJ5hh9Ufok77g9FagxRX21nPbZeeroXYPFNnsbXIPuYRECE+0vrh5drLpXYm
8tNEw2WoIMVvFEMJfD7LAwP96YNGjja6OXaZ24qHGuTQHp35fXW+d3MXiutcxp7Vl2MD+mjIzNny
00DNbXB3aEEBColBygMBoO2GdeTIc0jNH/40rz/ktBzaS6GITmOllhkctE3LkiHaLV9t/+CO0Qpr
xW1nD4LuFPA8j8CEjAtcN/btaZvVU+FKSE7xdchFomKdsNvYzCuzoEeOaV6lqg0uQTf7QVaTws2G
bk3isNypXTAQj/uG9r7TxNb6zxO3/tE1vD7NXykvCuKWGFKMqXcWTPdvGXeTk9IYphUf2yIPXRzO
iUg+EwGxCg/JF6zSro2bSMD5lpmJ3MvbP8uk7llUg8I3YxpdX8w07oSSmOSwfH5eGg4w7lsJOGHN
vKwZZD/wHngZHKCBtfkJLbZs565xxudtkA/ATHWgulFhF64gbcj30kShPMEXz2nl4bexDADda12u
sEGazjiJlbultaVoKvtrsm0VKDRF+CaF9TopOsjf4vKVxxCBjuXC1Gth4C/ZOWjXLO4Jeeywtzrx
epKFtcwea0v9NdxesRFv4u4a9+WxAwUcdFM5fsf3HnsRTJN2SaW+1pN3PFplQekkKTqrUQ80FZVW
4GD9Wso3LO9zuwPJQBIGzWOswozJezJyHH5jFL9ZEsczzB0UeMNPeqRCZCHblv4VvQ7vvpGeGmnC
LsxRkE5K8exgj/E3TAIQggh8NfkZibw1WK/gf+831LwRH1JMUB0WA61RrmAtUp2f1edHyfAhGqnm
Zei6f0FhzgI9yQJFTJ4YAhAZrgdjg5K+PNsnDJDn93iPLYKHLpAZ3eB874c4PhOVeuG128Vm8Jdh
fgCXegF2xuqmTJP4gFkqfnbUlMbPFvJ5AsJL3KR4rn+B9epD/RzE+8ym5Onsjg3M0HJs+45PrSzP
pn8mYz6rHiVQnD8T+J6KDHzyEvXGROZSA8cR7oaRUHj1lxJc8hQZ3Dpd5uIiqs+N1XnQVdRpUssq
ndR2jD5Gs9fmmWVRoaMikoy0uFj9Tlocwwy+/NrQbaalHGxYvI4jMI1ZHQKup4kPC6TT16Uk3a1J
fen0pSGrJCxX0CmD+mZMaKX67C+eX1nW6xogAS4bhqLGB21uYnHsEtJ3UL2laNm7JXgzG5/YrF2H
Tp8BQe2MOsJCVuUISTuLj16BwKYRBHtRXLm1JOB4TY2WHy9ZGJ3uSU1yZmJI4iipKAKYV0d4Enys
Bq5KbGTOawjKzRy5GwxTJHgfAQkki0rHojAJZblhyX//EnEU2s49524iMmTtUwRTpLKnGAC7EW8p
+dkDvgxhASbdYZBuKdbW8dKE4KBkBg+bwPnoSQ37N+MVKvvVa7Y59vLuYf6NlqIkXCwllaQkPJ3L
VpSr/3mDHcnFRXjC3c3MRauR1RHJ+9SRPvpdlGrLRTavmb3uCi+cy5kX3vO8y5QE7Gx12cfCPGpa
XqnPKr1S7Oz9///Jx8g4HXIDGVu6/Ba6rvCZLnQZvRNk/gUyl6mrIhsZfbYIPAAK5AxnMN/LEkdY
JGYQFzwuprwwUMIAKAR4f4n9iKXK+2d7Ave2tKVwu3FkSLJJ+Qt62CnK9iywhvn21FMvKR+AEbwW
Bu2cwq1I89EoqjGGhaJ2qRAoZZiYcsl+nCsaK07KmanfZGSV6y/vLQIoweX+fLf/sAL2hW0XU168
AZu4n4s/9A6S4O/x2/paAIJfgPLPQ2xWZs0KGiYAk2AA6Yu/0ij3cZdtWbgtSL9A5h/1pzTJF0gb
s8Sis02np6WcJwNB2avbi7nFueSYX00Ct02xKFaFelTO/qYOEWbQkzsyKOfKOvsEhojhv6vCe8hm
iAYfJ0x6UCjfR9qH69qANbTo/ZcyrSt5p5tGgLTpp9xoh5LIV3OvWsD6P5Zrby6RoWbaO6ESETKK
cRx9IRNrPn+3pDcIhmvMcaR1wnoQcAYR1lm7lMkZvwkBDnM98bQ5tjR6gHiaKNcNFTbzO3WEHX5C
iTO2D4T1A2Gv9I6V77QjUpMNwgNK/m5cAcZdUnKcoFHKvdn5yID8RKWVitbOgx7VRjk/5iA79dy3
HFUkLRh3aWTRMQ0/rKspAMgZy5BEhBGWVBBH0DpEPSye36BwzTixrJTShgekER4K+FUneyWzdh1O
PwSSO4wtMIIVupSglnC8/HUuqtb4PE/0lIufSiz4Q14/ooyJwCkORt8JV96zLvkwY+Dv92Sv1396
1MeIYTQu4cI/vzm8Xg4j9Cr1ynMBJBnnG9p7wDsPFx1T9qVMwV8p5vMlOLOorXKFz25iRgfipbjY
D0HicnAFOLZwrl5KB8afqartkylhsGW/eEPUOncHRl7DQerR1Bf0bRN+2J8c8zwMkfn65Lo2vfA4
LApkOc1ogMokbiW1D3SuM5JOuYz1hrf3PlFzcAEWxOuQxOupHEBxfIc42XiX9twZ4UFaT0+jT2cQ
VKHQLwDGAatMtDXIkX6dCEnEHzK2jMBO7j9KG3Fsp1ifgMZdH71S4rQbF5HAeqhhCVRifIAt83vj
WHtDNfNMe8/9EcDDBl2eqczeQP13OdK0AGcIWc6YNhcO3NLHyA3t4lrokXFpRCJF+cpht0VaADkC
CAPNnzDQmq7ee5/N9tWXSE8lietFQHlAU0BXrwT9y1m8IYSQm2sG0MjKudxblhlfuAZDF7XMa4Dv
GYOCbVSiWx7OJdqRmsEEkmAmrhshtdmLIOSyrfsNtnSpNc9rZbiBa2PtT6MQOnYq5ZcB5s6vnWyv
wx/UxRw8Im7ptOhiht/+PpZRlTWB7VFRe2MxqizC7B/zOdb4LXUqZ8BglCsvIG4CBNzmcDB4Y5eM
xUotzfqMC3AJqY9vZ5i55XLPCCPHiIgfwd81q015o7IJWcMuKOwY3HUTWEqC8ge5Akblu7xzwKJ6
6pjRw0jib9a92MU6lSwIdbDMcmChqz+WpLLv/DkgaBSRVlV88ftpMTMFNZ7/A9TqfhwXM0e+6O1s
q8mol9PeCZ5rXA8ccsr2BPvsGWjnc4sbyPl0smj8Vd2uA1evnK7EdGPmRa0Bc5RmzcPx8sR/oIKO
mSbZmTrY9odzmAeJZWG/qMoIfbygfK7v38OEQVL4jUn2kJr6mr78QvVp0HJOs7YOe6ZWZnA6uMbJ
w16orMyc/Y2YjAFZBue1Gr7a7f3UBiL5vUMZgJmzXkCyE/S8kVlvOrfP+c5AiqgJrGDHhvXTjeaB
Y3zzPjpm6svmTFPfJ0HPQZps9JFiLanAwfvFIIay6a7qOe3WT/ktEF7Hjxjtrb7k9yMDLq7DSd4r
JreGkyvmgT0mLgIw2wnWwJXjUnKq79tV7yz014fztNrA4M6Xv1t8XKki6Lg9i6OucYKzVDkcD1uD
qDQnrdWgSPj1tz28QcNB+9jPhhEbFkv15i7XAq5Nk2DaMiZbvMJYcodOWKStpSquXJBkcXgkqwYH
1AAkmO36GSNNbDE2eBwmmN45bz7P+e35ph8PleuyXCD6VJ4uaaqxEUKFZQEMwlfuu587xgwRILAo
M1RbudptW/Xawe2sbTzpqpTglFQo1RdbMGwKG+Cfx7AKqF8ZpQqVdPRBPPfoYm73L7VLqiN6uPUI
tV9oSjdAE4qpNLsqMW2QL0V7sSMpXBNZQJvJTfbzCocI/Bn2KyRtz51fe2ago0mj+LoI3oJpraYY
keZ7TAr5uQZ8AC/8xAdB1VkR+7ulAIvsfxbolPE7orxCnhVfUTHm5ixO57D4eccdjXxVuBizFNrE
SPzjFCSePFhGWISy605qzmd+teVExYtbKWiFjGSr8u1La/qzXHI1RE89Fpy+wJ8vrpqLTlSBKzDA
eRQ2CmsCi1hqB7zaSQRYuVTAY4ovlWQgaBIWl3YObGReOzMUOKMaiINSKhrTM+5t70rfC0Ge026l
vp+w0KFiBpOZTp+KhFj2p8gHvCKtut2RPxakil4HNIDYllj5WPv46dtvPBXxd2yR+GhdHprXTld3
q6+SBTuQXSWJH9eJNllsIdav5eq5sXIZStC7Eo2hRkBZqYMdZ8enutF5aFNBxswgbJ+lJr9MUwQ9
wyG9FbqBrBospBtwB4ypeOFx4EAoq7t67Xx3JhLqcKigtTUMxmicSJFE6RpojEbV8q6eoBTssM/u
K8SnIZDYg2fHOjYrBecxFzjnhVXtEbimID6mF2nLA/KCtuLKg9sd8uUZgeTbQzCkU9QzfJYBdpD1
lJMjDpuoPGmWsKNJ9KcX4JMWk0AuyFukwyWmwGZaCHxri1p0GIE4xN9mie8LfammVR9562rFuYuP
cDN6bEEtzTt/Yao23HV2X6covVOCE2HscRUPvun6G3J/4zRF3YxNQpX9B8iIBha4HQJmATn4cXbD
SYSPaftVoos5jl6QyyOikQoOtgh9ziTKVX6zj2OztyRCjPbaBQK717bAj9IvMVar/b7i8IlIJZka
huGV7/jckhKCnHH0JRCv/sELTbA7aWVN86+XdOFFNCAovQ3bmP5yUbtdDuyVdBXEe7DUDm8nsdhg
kA9/jFDeHnA27GbRI/5EHPAeMCmgu1wm7UOLmxL3xc07dMFZJpzaFvf3y5W8cXbDzqY0Pie/4Kwb
Gz9EX4ES8gQ2BzKvHHz0dmGp4feqvp3gAn0ICjAT/wYUttVcADhqySvWh1HeAUiJg1cZq4KhnHYh
/+u+Hg+7hHkEiNbcBh8PvKA9b1Pl3CFin4Zihdp/qMooqT9NwHu9hQ23Go61Jgz8HZLSS0yY4iFd
vUEXXGajHhok4tX+R02brGJcNOxFCacLewFPT7/KtuTvZEt97KL/G/Aq/B3i6AWkoBzskQ064WL8
kwlL1+O3xWaczfYoPwnw2GQQOBRCf1SrQEB6weZMJ+93fzPOL257DvI1ylslFQovoymmatBJ8loL
5a1wDihiPHpFMY53HkbvmH7q3R59xgM0VYA1Mr0Mc15iib35sYp0+gxRE/29DG6bcMudiOTqbad4
bxrC2Mallpm87vP2YK+le9vIuYm9o15MXpA8qmbFLGCGt49E1uVlRC9jkzYcoaH1OVfhD9NkwwDa
eO/cuezinIS9QNWXEsWzZxnOmfT702Eg+3QdeZ1zSh6CmX5A5g1CMS1qgfwTAVB1FediH30noV+M
4w4XC1zgV37q1PmkNNc5X1thMqcUT2qY2m4r7y8fbv+H4vP9sQCNnSNcMGXa3xqS1fvKi4Qrat3e
DMs3nqae+jYmwQCsFs+9ZviwTie9G2EIkLTs925i+6Ez9oQFt6OVHr4L/GRsoG0GycSEcojZzBJh
C/BM2hf/8SpatAlAXZiO2dk+eYjGRPi4tJGHdzA1LR59M0/mNPWSpiOmhGIkh1CLUZGutkHALjRm
iuFqDRH7stTxHeoYKF6+D/mQanK3gawE9JP5zZidDoDYEGlMov4W+Mj0VOLhLUKTphthHEZHckh6
muqCsjhZOreqoud6SXeRDBd80mFP6k/TBEl6BqrNu7oPhuelnOnYMfNTGpTc1iCj5b+Goa49Lup0
pHN3PrhR8B6IcLIoa7hS/XfARcbNzrV8pdhpMeKsueRdOAapPlosM+B+jUkjv6Zi0ShUtkbEu1VP
Ba6jIDveZQdyeRaXrUaaLHvx3zXotxLI5Se78HgXSOyhwYF3fw0iUfjo+88KlGRokAZticf8K+FV
oO6aBTx0poiRmfGcLBlvZfKdZxw4Rx/WrOC736212O3B2CX6lgvZ+FuV14FtIKKiePZmqhBJddwR
+5oEXO0etmmkfH7d02rzKdsnjYWIZ0p7AA1TpXCi0rWb/eSDR543vVEcxBzDUlxiVRw/I730yH+7
MTkWxG+zBR9LsLy7DHi+qheVjIlL/XLiaYRDZiUGz8tbU3zk3mdT8yikGy2OtE0V11HbvT7nMH1B
he4qpX+b1mYM7ZwZFnvZ30triDg9i5zjkHOxaO0VMcJNUoWgFdlGFQWq31somj0kCMqZd6/5OauZ
F6rRggCDYT1AqbXwWTW7g5UR0btTEoQgn+wSCGCsxjdlY6E6F3e7qrLa0Jbom0WnLUkvGMtDpM7H
t5s7UihDNAQRgdHzTj/qLGPcUsx1LJF68woyHxhCGL7Vrnrtx6JBkTJ5aWitbkKcn8syQ+VhjnkP
t1tmlywlttOsb2zaBB235IiV6I+R/Ovcc4HJ3PwSK/y3Ws7VGWlfJbFVIqbwV40SRv8PRnK3EArl
5S8eZHRmeRU1gqwt1a1GpPROPsaPkXg2DAyLdDhTFah+pPb3JfPlqyjmoVk4u2/q9rYxRxezr0e1
Fb6hLc0Lt5u5DYGaUFUB4h6T7B6F3eEABPYfIHJ4aN3GTLH4SFMyTRoDHPP/ZcfLpjK7/tcSY4oA
gMWFrszNzd0dbcb8WOrUR2rTNjQpUFLsgbz1zxDP11rsysdFX9Svto9VHWL6fC+1YKnhMBEkA1JA
Xzx5uZWF/Xisf9Ae+Tij8LHWfpzWM8kZNc/HZD5olgEgCH0B54rb9PCMzMRlJAZZATi9QXXY4Nze
rZTUspj/iSkqYCDJ03ZG5C2aI4FC4G1pNHQ9BVvE6cNlz/i9PBWy9kW++8Y43Mk/dMvmXd+DCvDE
30qxibfFjjFaHkQNILeXrzz6qBO5bP9D+XCrN39ZPpS8/g5lmPIqY1U3yS8DAVCWsyB+GeLVAsLy
VxdoiBJe9fwpV48q/d82WHqIxz6r3KIZKlY8sEPfNqG/JUdsIbtQqyqlifbMJx0meSGcnrgQEemz
RbJzonA/xQYP3Du4OswonU0v1rmn5nJmHrJy29AtfkRSJ5fzy6er2f6rZso+SVE50uh9wjeYqlxX
lF5l1ZuD5lENkarrgGxxjr4spiv5ez5fURTPWa4hBrFwneQ1Ys17QXd7TUHlcHiG71OZ9lh9Htz4
QKpjpLBy80InQA/byWN6POwXP9PrbmH4AJ8eShnOgPp+M+0Xfc+ZkUnA5mN/aq+hAVaXF7wo8Ere
XhEMv9DJDupQnOTvJuznjuYpQUOz0WgJY/+VbXr131y31Uuv3Y4Ab2GQM3RZLbc/cLq3VgUle4dW
qN6uNWKC6RRjPfJ7QBiVhQUzfv5nW+61682o4cjNqAmBLCUZ1LfO6lnl+sNhFyJ+7Yh8kKMO7wXI
0eucQzrJFZw55TaIfXEEGs9E2i1cUmf7pLBwrfodq3QCwXyBeOSzSEWF4YMfO2I589OCGqBRrz08
MblZ34cxKfpPeQVwhU2bjx6JMH9DthLonKq2blgsIi06tK0rT1l2u5M8CcWDcq+cLfXpyqOr7REy
V27vsAfP1H9I0mxrYETU8TtL22PyvFFx9BNN939BHPbGokn+9euwGtF9keJiWcJAzF4e7axbpQNM
qU9I8HmaF3BJFS1PdnxZKTiPuZyaw7RVKGkmwfHS570CR+HHBSB3GOwgC2VI9t+g2XyS8HSqXF1H
VgctbjXyY9YgAjLiKlFazy60ODW9SwwuwPAedayi9cTg1Y3SFuDVcmrlOFIzLHO93C9M/aClykiO
k+MJxKbAmAz10IJT1/QbXsscUhaLXhgFRYjoBoQkC73se5nbicVijEHJLwOqsuvH7Cu9qqV5lMDq
uyDNPUyupGlB6UjqED/hLGsudxa3U9Fx8+Z+2SCV8uAVVSqgbe6Z6WyUGq/rkpcuU5VLkJiAzlWr
ixQCQqwPKFtP+BoO7lq1FDgKr9GFGsrA9CYLV/1mjb+nIGHuSFvynEOXgq3RQwlH5G+ZgcU824iS
hP5EP/qGhOJI783jMolyEpLEZA81o90Li/pfhRRdzQx+//n6TRfDtRlzlFZnejH9pbw8rOsR2Xmy
Jt1mkDK9Vr4k9Uz7h/rmiFnyWCfxJwpF4yfroN+mbpoi1PYofbfwVwfG/YxWkeMWUW5eiPUSyIx9
ZRON1SNy/VqlNLA0uI5BIyNnUUnRmBgO1ibBpCZHUrUROXTZNK8fv8/XJsOq2wCIcbmOwhtNoXl4
B9QQS6ZkYx2q5jtvAyZ6mxh5+ml251u8UBde7kLNJMKgxIiTGifpQxpYTJOjM9+k8mklDtWYnvUn
MdStS86rlP4f5Fp+W7oIuaRcOq9LtTzceaVcUsMCBDUIQ2iXPjruRfgvm4I8qv12kDUyzlmTSZR+
W1dTmlRKZOQnIO92/rMb9Egblxa2zh/BOGK5ToNGX/S5LqyY5vhHib0MwJ0sCs6x2bYFP+oqABpU
AqYe+k1hoU6mBI95kMwFJxd5hFguYPV3Gljnt4ViU69ypNx56DNR+wCMqJ/+GWjrjAfOSaxlwWeZ
ag/HUUjRxgcnTww2yJU6YKSnbO9moxLZtjz56LkU5M9UOzN8DAa+v9xiCkcrvoUXHXINAuEb0RAy
wRWVPKiiuU853IGr8CV9XWHg+HXUbK75jD7gG8RyLGvDvkeY3tAIQrIJJIq/f3zZNuCGljaBs699
KqARJo1o1xAif3SHpdiVMQOeAJ5F4Zx/UjiwUlJ1Q9k5DuqaP+It9tDHDInzzoeD5TLrZA8LcahN
8kHsGOFsruI74XE0yvyArRrjhnrYxjMDQ2CiqC5N2iGBPT0WoOcQzgKOdSOWMHAIRlfqrhFRb72h
16Vy0tZixkRB99Hj2cUqb5Jj+wX8OmNeKEMUeIoZM5NVOddYTnBA01aseP/EvAnDW/5CxcsSLciD
fxMAWcBgeHQi1P4iwy4oSJmlCKS1nIsaNtKmL8EExvSPGRhK/E5wkoufzfSqFCfsW7J9u0lqyH9L
mDu5AIxhl7ggfC35unwUirOs11mfJsVTvSAapP+hdtX18DmoRMyWumMbKgW1DA58BWnIcTpbMu6Y
GTOZWA5fAExM5BsDw9NNjnzkhPnBHyoUJx2LhazxDbJDWEHf3oJTn8JS7xI2qqFp4AvDLbQtCQmv
lUdACa2EFqTzp6UHIVmUi/AAmrfu4qrUDmyh/e1S4sZ4BZNjrcf9DMW/uIyF5lXPUtQnA9JGuS5m
wJEdIqZ1PdWJfzDEOnfoOvqc1D0T4sjT9ajXP/T8SrtX6wPZ4HAl3u79+JJ8t+JEOmb3gwLNPAyl
UinBglbLT92uuAdYFbXVon9ivPeSJaJfeMfZFHQ6SI38MtwpReHDR2PElsDf2ByLmd7Lwz5BpPvh
WMXM+/7YR4Br5d3au5QvKJV8gtHeIqn9uaV4yMIaRW/TAfK6fd2ZzFnFQlTVs2Mx4ORaRKxsbRFR
04eP7oBz+FVb6zLgirYQYzP3McSDs3ULajO6PLAisnQBGfUilqHoX+JE5vcTPsVbl7P6SZfZrCOo
+8wyoodEOqyjmb3OtJ2nhJAHEzcOOGeybFqkrAQw0+keybsCyGQBXtcl0JoVV/yrEcC2sEhtxLME
zqK8dkJZqtH5XRdaso5cOUjO314bn/TFQIpETq1v4CIqGwbRjE/vLwzVdoJxrVP8InKjVzACzdXZ
gAoP70taA/0NP/L28Q/xL3+IkldULL2J7Y9Hn7Yq22iD0LLWmsmzWqlT6HYygikx8Wv/olc+eEPZ
YTfBkTjo7sAhKcngvVaRfD/DCquVJeID+8XZpNSIs+u0DKEPdZbhdcA6A/cg5id7NTOTBvxU29pt
VdZh8UIm2l2j0U4SFxS4gswcSYp6JXmdMsuOZHnP0oT3J+qEtAb/fupTBYe1MiUFoROrpyTT4eQT
WaeODm9e+dkt6uTAQDrSvQ2QYut6wHa7MsN3TZr0VdHnEWfz7/DGQJoUuh8JxyfTIeI3wXm361KA
KBeRa13Z7xhhVWCbKGidkRprTmLiAlnVjZrQBVHqWwoRICsYEKzPBA9/li/McMa4M+qtudwZocWW
7un9Y0GYwqMEVm4i9Xu21Y4XA+VrwVgJ9rdcHHQ5kyVbJWzW+/PHYTQeEhXxb7eMN3kY33zSB5ga
DJWjT3risvJMRpZm7nnVwNkO+at9zKGRxz4WHH/M+OhBbRqbKco7Zex5VnVSZYhUgJ4o0cAl0feA
ceajQi1xG1Udv3Ouvi5zMJKJ+zWB+5v+4PQwXZ/R4pZkVgHze18y3QHDIAWDRpZpLFZsGC3S9Stq
ZDo+REw3/xkrkaAcd2JUNmirGJ8oRCxftFy//yamQVjHcGdjDxfST/LsjSCLaLWme3vXdEhb86UZ
LNqkrh1tLYj5LpV0GPBCgk/2NZIxiCFtbgQgI97SdoKjgI0gBuX2dpuFxAjqI6pl1Hol9QHrUdhR
OQ3RCXgHxAepnkKObJEfKf/4IdDQtlZHkqxQkG2z0UKpFN59dMawS2dSJyGDrNvpJMqbO4hBBAEi
H5wKkS1EhTPHPyJ5/BegfqgcsYG3VEt2gVtPAnAcyy8N97SvK5fuwzfFSI7rp3U9tclUMLkQ3yod
BlHkeiKFwoiS3vCB2qXl85nGQwuefDXwQyU9ptXS1F6F6qRzaSveOMhSystVhXzGlJPjlG67qiRI
5ePCzWWQ2sApWnAZUcfsW7ebXqY+jjBp4E0UWZqN+2F6fhhJpzJ4mX0oVk9xW2zyA9nCtNSDNEDd
dBdQsESm3TZhHQNpIJ/NgEerq4a5aomoxHbVh1IUkcrUBB7pyD2qGVAA7r91ckQ9qjZFXRbEChZN
uxVS9Bjckl3QcDHEA7t7nbIlA+GB8NkFOZpeC2hxv82TGWBAGLFl3vSDoAgrnknyHYyJevQkoUhy
DlxFCfnEA4uhs+HpwfgT1WOyCJsGAa8/RU6IT88PlMl5XvfCDFrkk995xaYtJIiPvAhngiep44Yo
y98rXlRo9Dk47xHqr9jl0Or5+iGl7KMeA4t1yS06UTZJD9rYmGamt/6JVGprE07QvUPCyu2MxIHy
TZb5eNR0gmKyGU3Lsf3AUZeDdzE2s1C1ZFHWeqUP3S6kiMoe8TUHpUFrCMj/ytP8RidGsOqJ2h6l
z+Gwi8kJDVzaVTNEJIlLtR3yGIw3TfvB48zOCC55WZaA1QSzXTOPeV/q3TiuarEm7h4rHmIqTRNS
/Z7qBXYIaDuHy24x7C9T/WASsoopIyVgCoLwGORiNfsUUW64H2253x1Zju9yjPoKTLZbeTqD8QXW
hjb6pOFM0iaBLK6Aq0uK5a2u3g6yEcRYGoXvjOXb3XK+tc41dRHu8xPwOi5BBKnuEJH0BocaXTOM
ExkzLc1HFhN1j8pYjyt/f4muS9gcTpP1rzX8e7Lume7IzgqQPGt2Vaz/8kpZa/wOPJHSCrTr50Ew
ftls3CNkiviEmxiNqMbliJINQjDoMun7z+DNT6FVCJuR1ZZOxRuzmftcbTtkdPEg/dnitnUJYpHd
S/fU7LSpynj+pQwWdJny7xQKPucV3+SxsIC73rlDPr8XCExNlJHbQSUrmvMU8pkjAqFVmVpYGhyQ
4rBORLkc8RBeH6Hbq7CkjQBTOgAAEVX9dBW+bW9tQ4EVwJ2V22qFv2V/g4QFCxQS+iMTaN+rep/v
JxFduyHIDGD+b11eUEVGk1gpL+jRNAwmhzUWS5Oe6QcJ0ZyfVQFINbD6NtOLK/70gBJ9heYkkhKV
2t7Wl5cyKqNvF882bGolYcNGfidY0oV3WluJL59jLxUIAXxgiYkX1yQhIc+q8xkmsncuabyiB6l2
kFWwM3jtuIj1zpaKxXNA6VKZs7Kr3FsL/RS57NvvKGXyG8M13vXm6TC2ggmK1Sgj7PU1vo9E4MeE
lSYHDpzMS8YP5Y7ezUKSsr2toqYbN5ciZo1Yhx3ImCWbYLlIOQ/HyGuJzlUPyh+NCNr7cLAr2+1J
5CMikGiu7aKH6jdcLjfDQ17THLnV/qEDUqOfXiN/Mm4v3pdgQ/nJ4qPqZd3Jdnb8/Vap/WFc7jCW
g40nD0ocC6oBgRRiFPMnrYvGD7Ki5+LITm0UiVZpaTWPa1P5OjXBT4MUMYkmJX3i6tqETR5D54Sg
Az5FvxMPB7YqrhGN+xycz79H1PU2yNPI0R2yJmkFpfWdvYbNnYQfZU+3+3Hng+P9ulKg4I3gKMtI
w/3KTppmwAdEXI2kiQVMmdST8exQD/+HXUBsJ1T5mAr8MbPfRnBBt8KZwkz1RU13v1nfVBNxwBof
D/YJjjZWITDTxLCk5xiNKyuy4HtM2ECJtRX21NSkWflP//xhjdmcDIEZ3XP1B/PyeTljU/3+UbHx
a4Jmv2TuYkGItsTWms9WA3JMrwWJMs1Dc5MvFFrn+Zcz9M3s9vTBV0kbTFfEJjPpfYPbqiiErKCS
NlydduIykoUEAKGP4pbKkd6sAXuASKEH3Z1YE0rJkDTvA47EJDbXK2xVh4tUHfjvx8YVAi1c9fjn
x8wVkzKqgaPobFZvWk/s6PAr7GotQS5IKoNfk09MRVcLRFuGzpgw8ITL4QWrfMCC8SxLWKimpTvA
IWSs9wEHyBegQxtlZN3ZVFeRXe6331wRPVCPmxKxMQtQO6RG/kdLSOcnlhiDbFzeQn3PL0i85e6a
tnItElOtDRyc/lBZbUcXOPfVdP2B0rnqhcBisA2r9pW+W1xaMKhLdDeEONemoW2o5ev0uWE5/7av
sObOO7egTBiBrnM7MPXbpQlJZYn3zQEObv1aFhKZEDMI3Uu5GRYa78XWbtGQfZd1N3hM1ESeETdh
Lenlp+ZV9igdjcXZXQ+ZYdcT21JTVLzR0QF4VcgXH+6e9IZh+iIsEwsPQB/PYTcG3AX+f8ItM/h8
IGa/YlXRLerZy+tsf4LvQtGiuW7ITcmw9iXv8TzdwmylL3A3U5ITuZhT/GFsBjbuthmih8e/pbOQ
0Fpn4YJIn89iHnu+fF8RCmqiu9cVvx3iS9vd4o3D8vHp98gbFxDi2lgXkt3y+qg1iKdtiLSzdBeQ
iVbdsQNPeSqYG3nLhBgu8Cup6S1mJEvvYBbAGkyPqI5UgAgYxhjxDl5nQLvfe8sD71X8LPurTwtj
5SLC/vmw7o5hqjTrbthlhg4jxgSLZgjqW9sO8uWMX0N42RbIv5/pLUC2ocG4L7ckzfTGRkEnhAYI
9wjvPdMjvUG3F//JXidHwaoJxY+d5Bv+WuSyUIoiKnDJiQGsNu1Fv836j36wRJ5oBSo7lSXtN84O
C3MwE07VnjIgVTVo45JGve0lVrLOyzQftKs8+KrgKshbiqL3twsELgi6r5vu/j11LGBbiZ0uav+A
cskckP8UzATDDnrCS6zxftDf0Tc6yhE/9ph2cDtzl34IZgKAMXJDpkBmCYM+B8whGQLtzbJ/ZHTM
BegqABn6cG5HNWw8q3HkEUFIWrU9QWA7dacI3GxKfOm02mziZY5WGu99DDN/a6ieu/QSCh+9Ob8C
pSYh9gOsRmJtngGJS/IQeMS2AULEcCCHSLs6Ra8kuc/OZTS7G9PjuXgJfEzztRINZNSBjoYz9ZEG
LnjL4WuCsLSnN1r3XZkD7My2Yw7mhSQNhZhFLW+0ePTxRS4qA8GLmgtcgO5pQF5+1+33I06ahPkD
LZIdYuGdLQ9xgCoyMMzf+u1YraXwrXP4bLnqusAVvoU9ycwagZg6vORzz8Vx2FwHq2ZhxpOerdJj
rRFHAzDoI2pjd6Zve9W73S4c1sSdIRTKUeMTSkZ/Ct36wclePhkaVRyj557r6dp67rsNxo9Bhn5B
EemTREeuITB/objKFQQK9Jj6Ci20P6MonrE1Bub0qxWpsa+QUqhgBpfP0yMIoUbkbcN8ktZnSu//
9Hg2Gu9pPrB6aI+akjApL/vOQ/nw2inioTdgCzdlqUrqiBKarKVKbQ3p0bDhmqv1v3vl881PJaSO
ZLwRl3EdAx/H2ZlZLydDVIUrhaB/pvdfnyWqKRwrucBAgMkSVDU/bxylRUeXUkx9cLjavhxFk868
S33NUVHrc4Wvw8bZUBlKDfcoVwjpK2FjY9DEw4IrJ4pHIfCfK/gcxdbm86wQOceOx6CXNN+wXRn8
BUAlCQlnU+rvs5jcsA9TxJLAZHFwKX24+vAIm8H5JG8DcQw0ZdNdxsLTama3ZeNp4RSb/Yd5/5a5
52XCI5KVoMLtWjljTeTAMRFgSx0OTPxxEjcDBwxDiuxWs3l3m9ZuDbrhFKj/X15E4EJCPrqFKqx3
Ec3atP5U8hftP+xK9u5ztXcYfO/2uYqTzmGrYB+f22+psExEpXVx82DFQnnAWdmFKOioX+CCxRzd
R40/T/vAPntUgCV7h0ku3DHCbNE8vjno1cPc8xIL5k+SD4p+w+F+wSpAr96W+zNcMZP1Jsw0NFSD
vn6gs0Nr187sds2eWiRNFUme/uxYWb9ml+HZf/t5dcxWMBt5VXDLoUHoIe6UoPXRZ2QPIH3pK5V9
xVoL8MCJzDvijuSmowCiy0WuVibDLngfxrN6BdOW+PTOODPOV8QU07ux1Y+UMAWWOgG7dBr5Nth/
3DEaTbECsewsBpGVn2bLsmzCSc9T4mPBAvCS2MzfDvdhP6V8NFNoJDdQRx1aoecAxmD9/U/FgE8k
HpXWxMUsRTFSAtbwiYDRKDSTZr1000r+o5/ej0/17yqfMl/rKIf3OUOPaFduBrsSx1hfVroMvTOI
oXdsqyeE2X/hRknOBAKobWTSBzXfmnxj/ndFpRGvaVc83ZW0CFl2WkWDNS6yj2JMY76LP86/RN7P
v1oe9JUagQ1i6Qu3cwD2gucGVu0ZWvpHRFduH3ramcNSiqUJE7J/uD3HsK6MpRrM4q8zr3AdrLBn
QyF94wX+Is3NPM4bkVbQoXNL7smNHhb1HHcKILzWaOOPhjirSNK444qyQD3o9UBC6MFLFPfreeIV
VQIPeNQK9cCOisY6U8+53X6uSg+rkOIXjCnvvxOKLnWCFdp2wEVNkyYvLHJNnbrhx41fWogJhfyC
1I+94Eqr8VGP+d9SyQe8YpLr1wDW0cwBFsBp6DjNqgvvVWOpLX5uCI72eCZgNp47H7CwCIvbs0Tc
hPT8NddPUt4m882Dfzvrqwr+q0s1nllcDdICTbiKnJV+7S5gONoR1C8v0TBr1AwAxbCuyPRWrlC7
ouez/rbANNO99vT6AuPGzOSc4wh2vFL644uauPct+3Qs25OEPL5oOod762WnY/+J0aivcm0sZ+px
fGLxaXjlHcoSiXAeRbSOdBB3t+eZ3wpGCSdKtq2aFZenIKg+zria9jgw+7LFTeCARv/gFKYDnFBM
Pjc3bQUGNYA+BxaUZoMshiedyrToiu7vamkE52BDqL0JHKZOKBH4BxUnYXjF6mc/G9IvupykcSqG
l7kiWM7yeNs3kyLmNuKTBCISILGZddCg601AJoAmy57QGK0sVFlXJN2MyyZnLCiCijdDivfTlgqY
eNqfu9hGTRc7hA1j13DIvp9lx/5bCEz5175r/Rt9He7aVwgsPXmZ0wMEU6DP7sBhAEbGAnZ0MWzm
waqfzFjo6Y217iJTI0ppXSwc7J3pDJtl1/2iafvwTHLaByHl/2cKK72fbQ6967lMzsmSWt7muESU
oBrpAAmrDz79nPxA6x4uS1JxO80v+y7JMusfWfMPM+Mf+0UfLS2XULSgNDc57QHRPD6BLerykWNN
MwmrP4DySsrY1hVtdWEC3g/bQKc9Vmg0yb7pFnPaXUDp7sbcpArX/7vhXESBW16e4dGcCatmzmR8
jppI3Lrj1V/AF8qPdXQZlMKJBgdkag3K7KGhnoX6jLbF3bqSGT+s3BlkX3117QbIlkxdfd/8t18F
jCmTX9ohtMtCYQWv5pZOMBiaVzsAFbkj7vpXwVgQpUdbiqGeft8PpL+eSWAADYlb7qcjpT1ZKPaW
p5FQrX/UZra4FCf8PDt2Z+jGh1X+JsZdCpUChdWeLN93ELAZsmn3n1oxBu5p+UhpJcARclXZ8qAi
C6xG3XxLIEFzw5p6ZvUo7i4EYB5W2lytRoUtp3hHX7CdNcw7xg8deUJDR0pjkSua2Z1edxqz4+L4
cW2c6XVvkGnpEhgC3yKSjXn1Ufxa80o06ysMTewH+YLNmlaoBp+kD9wat1UKxG+p6wpvTeHy3q2y
2/td+YvXbE8GDpXjU3tWq9g/npe76a74sa8cl0qk3TW29pwqsQ9dm7dvlOg+4BqUTV/6YmoXTyyx
yMdpbxGyTp0hFNPtPaXVMBOOi3P3duPUsd4BvskoHAICnatdgwxxKaTHkMUOOZSBQ55Dwnmy/FQy
9B0hoojF4259B6yxIZaFEfK/ii7/sTZWx81q2W4QyT0r/eOYcqdL1xLmmS6p8pNIef+C9EBDidqu
jRQTLq95HW9oZTWOPqYG0yL2JtxbLIeeebq4lRXIS32xLCooseQI6Mg1jHroTy8u6JzFWt+t1sdo
TI0fyG9CdefNibN90Un9c0a24dS2XZK8Scx1ungKLFVlHRZmb62JiBjM7HGRSRG0ivBVsZ4mpHg/
ZwgGeVjQa3Pwr+e4CGpdnAuPU78j6QuSB59S1c+Xo5BuiIsdMrDg9KlARZLyMFUDxHIdEZVECGqR
GhAOfjreUSy50X8n5+Fnomqjhbyr+me9LacrNrHVT0IEC4LAnHGB/YP+WCU7ovimYrjkxpxZYM9m
J8HPJRMBSMbIPKfB5D9MgRd/XJQpyuQXbXa4h5cbFoiEMlcsjAmkqM21Ockh629MQ898VXoi2Xfs
iOcWplSFi2sEcbOvWjletGlNWsQD8UU4g8oRPgtV/QyDLnosu6kV2lVy2Zgp8ct7ay7V3nAmLXXs
V25+KzoDVpKExtokWM043lae8vSiWP62MwvPOifLexqWzvHaMBNWT1frX68HnLYWSZ/rGmok0goV
9SHKX6yNs68/Dmww4fWKoNsR5mhtI5CdKVICFD+aXbWNr+7bBfY06Afb4bxyiBlNNqhAKAujq1R5
BQZ3j3/DQHGY6hBh8loWe04qXgBasR2OZkpRTlPJVcle+GDbqZ6AdWMUNlMQ9pSwnyiqGxoKefhO
VQ+WijF/o8GZy0m5kx/OWkCnC2kAlLXe/1Lj1BjbtzT9ri4XKt2DKQ4AOQMwCC3r7+HS796IHpwW
1MMK463swk5UR8HtomUzAKjw59PRyN1NfkrQKUrVh7+XV4I8NO6Vh/qQmrv2k0SLyGRQzOQoycqj
ieg3fZMx4R/vIbfjmkB7myCV4N28AzbQn87bVD4Vt4WXd40NYxS90oucdkmt51VhNoiwfLxsXdfK
dhhO9tUgMj7Y8cWQ5CnU7lC4sjQBujBRMKhy25xaX1BSNHIHZmMIXVLbhR3THG6gvrDhsBXdHPB6
ffG8QXhDIKnvehDDnDruLVJd4mqwwxchgx+HndhsBgGkdEzVroEK6/TO1fZdJfnXmcbLSQB7zeX4
qFPWY+njDc+JApzHZ7GafBCduUP6BxtQT0to3qQ4V1lcIUXFnDCfzGb3uSpINn7Md8qoraYAWIJX
bWzFB8pEiY6nFZPbA8UNMKWCBeIIb71Eg2pFfPTQycvlebcN89Hx5piyGJDCb8UW9CaNO7DBDz6w
AnMyw3vtYGXwzhQQlbZMC5nJc1BO6gwFCyDTDqWsj0xO+wz+RI0ygq4+gVwgwG45LuHnGu06DpGs
AOYXntXByhf1p1KivWQmLJlbyxEmfx8AmSDVKiMLicJwumyjmNXIkLq/6UWjeMjtx3JRGvtdusoI
AiVBrbyEbaxAe2456sFpzLuGdSRT5t9LhhldVlNl/G5vh4xbNtr6a+X8mK0VCiOJa+ur9CZ+Hkie
2SIP5KR7qrjuX/4NhhVvQWNVTIcfbtJLkPdBLLIG7gergjnV1JrcKt6VtiTcbvFCnWGCZIaHg//1
dtMiabGmGT3gXB2okUbK08n5yNGg34zduqlnJQyuLbfVsIKFaoakBWTAEImxxyApxf2ZSsjaHToH
cwJYN14e7wJ6+cXbV3wXfgGvULqa5VXE62BnrkIfk57qxNYxGa6+PExehZrMIXx6Cxi0fvDajgl7
svw4Q4upcwvE7wBcpc9CvpTZPrmLjxkV6IJRSZGONHTsg4sS45OnIEtIjIkQKCRywrFDi0xNMH0W
tGA9pvOyk+s6CoZeUCq2QaVqTRtEh1A69khr1mZ9emiZKw8fJON5KoCIICTk++kD+LPmb4IyfE57
8jsTLw/jtSKJy9hIyTQazL3jlNhNnAkhcZBAa07IFHyQ1DmQ4sWedRqa5UzQBBW8hG+TRkWcQ7UU
VCvS4VJ/Grwh0EfkDvZdEDPZ4j69paD75v+Ms7R2Pv9+TJHqh/cZ73H7/TCQi8GQt24Y3gGKlObv
/Vbq9qllyLoV59XPe+JR037yjOjK3dH5enNr6+culR30RbIL9Pb+Bl5g1wCJB5HBYJOGQQeaUahV
17az99h6r7L/x6nE8XCgBk2hk8BdwwlPTC8j8fUeLOLhy5vRdjhmEW0XJ/doN19t8fE+QUpnJzPj
ErW2Gb/xj/g79cVvXIOgB+DNNdjkE1zQJlWoMQ4E04BuWSeV86EHsEujyqbyzUiSIjY4A2Tsp+pk
36uUKY1kS38CUVNxL8VlNXczVAIET+3D/rx0Ful1J1vg+NSgu6xMyh/FyG5jL2P12JE/0NzHHnY/
Mv6yQ/fnd5xhirGjtpfvLl0fkCnZ3VWMLPYV27QrrU89giKxyO4T448cG4hpQgKZ502huwZXHgj7
reRO4NnfBpCjRh+ECTec5EwtYIz5EPghSqamWBIZHtGKG3Yc28EPcIriO+sr0vtjOV2QulTMNp+D
NJE45pNnViruLtGn70xlATEsQed+ex0a2OJ9YKK+yv+heUeRZxHAOjpN/d7nTrTEdkOMYkCbJZIK
YWBhlt00ZQ8Zv1C0Gxd+zaG6vHXWLK5/0ohVprw17lPylRTAbmFn18TFQkgqPmYSe+JbbymtFa9F
1URZj7Ng+imcxXEAjlLKopQc1bhVnjtFYNNOR07DxIrd57sMXaELAMInfvjfuZo6TFMtN3tmByYs
rD0m9l6rpFJJrnZ3jKy9ulNUjA4O2N2JwCw6Dz3PC3OP2zB/7uglmoBtntDX2DNSBmELa7+BKPxX
f9bl42CBJAq4LkHGlChkeYSbX+KzzWyP7QcRvzlgz7/a7GAvLmaqkZO4gBWQ6RuTxT9ef7928zjj
vpqwjNDycDMoAzHIgnXB6KBHtHwGHDWgM3oBEORYUo2jWTuUSbN/5ufNH4h5JV/PV278/PBvHrEf
yQARHmQscFMaIijgH1inLCjTHlDbazTUEge96m7tH40P6kSJN2hcJtwxrKLCxhKhy0Agy2wPzYlY
RWLaSsz0cFrFlwhvf69XREbkjBofnARYswUmsCqxLamibjeOwtr/O3GzMK66B0eCm6ibnqNRPdyb
EpVeG+pahEINBrXNhna+zAYWYOSbnS8MS4Euh+lQIgJnXRFJamoiRKS6lLMZOe7ydUCkZeZvaZtG
RaTah36Kil1mig64q/nbT51dPPw57ni8r0Bu3b4l3rJMGWi6iH10/lvj5PpMtzd5VInYoZiMBUvL
17mlns5xuYfxiUdQSyRWoFIsKH7svlbp47asdKRFRgFiS9/if6hNBuExaL9kQazprUnVCG0UL67S
4MkRoAt1kMBExNGohGNrYc734BJVtAn0Obk4WxFc0wdJDi1IbhcdGlt2R7CDwqAFVE7EVJyJ+p/N
FCjhYCi5E1j0N7t39rbz+oKVvilWza8kIUawTsV/sfiZCMquWhd5nOOORtcYaQkQtAHFBw9hYClO
Qm/Z9+S5m8hxFU3onHhOodNSqKZl9j8EqwrDJA0Zz8elM6c7iV0+6dbQlDM3XgeE95qWsmHAzzyS
nuY3y0XGykWZPnO1P2WhBf9Ph0QJJWZ6HY3+EKyh2kjIFFdFI+ATzrMi6KKCB2+e51jW4AvwoSup
HmWXkEL2p3PtvTtu9xK62ADaFujueXQxCMh4Ui2b1Xay/OG2aLNIwMx/d8NcTni/9brY5DipPaoq
36r5hfOICZ4xFvZ3fB3nUOKkRq0oEzf05IrL5UyInnAT3q2aAcqwucC1ziWbYy+HTpiFy6T999qF
GFuZb8quS2wXCltFQKE85HMq7ykLTguYSXVr1vaprQejhNkgGvKR+ByP4Ma5o5swINKUt3GtllDW
sL7+Qtt5V47fo7NGnHSPdw9MqnBjPs2C0/i2hVL6nQwcuFu2PJpCyjhkAOqxpzWokGvMFvyfmg68
L68gR9FCy30i4PAdrWR5K2UFYMyieNgX6185Wzup47NNmN3BqjPzMay3aemzE5gcCQR6+dKubG0J
2BB7K4xhKhSmtnIP6DX/BssfDSIwWoINuSbQdXapF4HnEN+43X459FaYDxeGxc6IMTwLPHtlNjrL
XyuO9PYpbaMTonoQ115CNzV9ailUt2WYUYEGQRcBPOr4gziu8hGNmFCRCxNupPI5URtAoHyImEnX
ml75spZNsgJggVKG0qhoJgCe+UlnPsWHiqfQ/I4SwDQbbgc9rIaLmW6zmpMU24xpGMB/oB/zMvhi
j3v9xrTRTiXakROq+ozs9QPYLjOs4of1L10KL1NHJyO5o4X9U0KAMdpBMZKpDFo527fLQFhjAa2E
duNuOzPeca/WhJSrdLHMCeEZ2x3nTMrwzpR1Le+K7pdmnvKoBKGGv0dfnjat0pA3Qbdb0NJhZUUr
UO+XQAf+ndGTRTj3MRwphTgSprmg7ZAZVpMyN9h/SFL7gBG0NmuEZRnS3gTZsuEbn1s5CsCSt2Og
tZhLmShxLz3vPFQzgfAR5NAy5G3oh0N/emSddLEcP35vKDn4HnCacnxUSiSTyoDbGAG2Ep2vRkrU
vZF9tsMvT8mP62X0UZ/HwO2gpbaAHEBzHyO4nlAOrPp9qv8XmBbvA8CMGVSRgFFJ3QMjOkS+8kJb
TXaRdvcR3NViEKUfy8cTzH6hU1BLHFaQAmiTl2GQf4/NJVbSE2tMK159BqCwSDPB8BL0wc/BNTVI
lRbggQz3my4tMoCdJGqvtf/ygyWqtLwY+inKzcKg2SNTQx43aX3a8PNB9unjhnynDG11W9Yf9Mrw
Fpj/Hox8OM+ODZvhtTfWa9XTBjDLvsempveK9P/JSePjuGkNHE5xRpJCQtYIdMVai5r4pRm2E4Ci
18K1IBrL48PpcFzC0nmzAv6QQXVLzpEs4BvhyGSGg20FVoy8Sv8zO1PAa8SnxTVhlp/HZiDs2pMB
AbZfyJqhoq4pJbhLFFBFpUeG0S9C3jQPAJJ1mvd0EuiTVS9OknYdQgemKKJKqh93qUnuEtAfnBQW
6EBKy+luv3ceNLf/FMjh+UCaRPgqq5qvPyqTbt/hj5hJHR1mbyzlshKZK8Gp5KsSatj0KNMr9BZc
ZLdgRuwQVCt2BiQZqe1tjD9VhUw2c9eCycv108iMPeoUvrNw7j3q2J5D7fCobTzuuktWlV+CF/Ks
j+c4Ms/3IiEDI5foVBG+L/AHry8OTzZR5SL5cicEDg2D8jHNjwW9neVDSkFXQMC941TPQE4deqky
pv3m/ijwl7WS9t4ZSsTYiiqLO38tYEZTrFs/Krf2d6oAfPItjq5ggPHVhxXsKqjEukikc4jJAcc9
AyBc66GTKsO5R6M8MdxKrT6/DTpdGr3Fn5RHEL6DlJZnbkUB+Xpjg82U8EJFgzYGMEBc2A97oupp
7W4YDfzJisOdLIyLa4dwoYpu5F8PdGG0IB4iuctZs9GrPDT7Z7rDZ/lzGXB1yfwNRxJAfrCyXQJ/
n61rS8ursHTefDN0tNpdn5TStMQxsjq/YO/xkJtqLvKBlntW5OzuhgYYo1bQycEFz0mGMLsO2ce5
ivbhvNCC3NHKBHfV/2FNSDosvw3ukYUvNuCO3+ExIs34xBgRWS8oA1chcvrIMhVhIDmfB/3PF7BR
pkhKTUuxp9+uoYE844noTE9+yHaKqRDbALYVtYvDN6kNT7iPGee9qNP8vkdWvEMln5dI8Cz4+WIN
UuUxAd62UqWap/7Ch2Uuq3E7LQFSMdHSlUumEsQPmYeYh2GpSc50MuOx6kQFofLNMMwNwsrwjncX
yLAQ033O1ijIauXj77asxwIbx6NS7glvYKpvfDV07Vyz6DtYrv+7IBe8/FBJRnZh9RtfyVDD3bcN
0/WvtyCtXODWS+uCiSpHtFGBiBI2erA77oEGyZprw95LHOB+DFS9PwAykXC81DvpfyWmiqcfoWSh
yIsvu4vjWfuM8JwpIHtoWC3kvlaoYv1y78UyVoiUVCsGw2uh56paSBH5FGNV5Fgg7/85gQkn/Ups
aWYgGswPTdOZ1gqp5Ro8exp8MNW2AeAPeGCnX7lqM/d4926Z12r89W0hQCD/bAPulgDyvp5Sjkte
wBU13WoS3sim4YMQfr/qXbw/YezX6UEz0eneYPHwuJBBonXltmynMh2T9HdSCNQPULH20Vgkkf+V
KCnHw10fvne2te7S41doNCCHSfVCNyWx2B1opntqvf9IAEEa4vKaB2JCMJfnsyYXEBF1DUo4eB4v
SLkHoikoZcrYtUilfJjMeFNlKU2EJgn4jMhLyeFR2vCtpPGE31xMcw0hXdwYD0OuvOkJXHpZrFyH
sG6cqi/jJmx0KNbLpSzg+UnHD+c1wozCWYK2fqTl7MQUw2qlUZqeR0Wb11mkFqvOOMiMcGZDtIle
ecq7N3fc+mcCxsV2US8rtsUB8DSIlxzdMOUFIoLDau8t1BARSytUXIlGkBebHDwfU2S9lQgO2im7
QWy5aQL05vxbHb2vbA102mn+ans3tezZxVftwuewtWSgRExBqgPgKfc4ZcuIgCC8DGyQ0Li+dNIH
bM3y8LriqVaE9w+Akm60L5a1rRzQsmAnA+ZxACaMldgp3M2kNA556zvhN2zEstRAJbdrI05Lm/Hf
D39rd8PDg52ClvtmtDOYG8eY/BrBCfNyrsmNwYCo+YVWCt32Rmn51noO8dtI55hKQrQI5tRZv9HP
tn8VPCj1/QFJ3h/4rBZbBPf+ott4vrRPPDCQK+0Gqjp8BWbniHUJN/r4GOKQXO/Qmbo+4usOUC8m
8jaJ7ScTIFcFKNrbqVAXsuJE3te4URFlDB2qD9/vU79m9UfRoodykiCHFnxX/H+7T65y+mznrkVv
L3N7hHdGGgVLp3vFquy73yDBJudl4hMA6PmyKy6T8bupa003LrWBj5wUsLpJ0SEp/gcybo6FADHQ
7G9rs98r7YvtwY7YR1hpU7ZPUvuNuHLZacRfbVCOkP2uAtpxg7KlhwA/yBbPkJvcIVn46pF5NRWK
MGYtLt1BJJodJnihOLiaOTI6DMPgKL3GMGu5BoI7fRYClSdu8805UNHRWr1HY0uev4kC9Klkmvhz
UwPRPx8Z9EcfGX3CgRHSnZPVY6O+IrTkFQLGCBqqiMmma9mg7ShSFPLz739bNtSJUop86h4PjjNv
kqxhgzEN8dVQTy3NSCpqlPWSTn60AAKc1vvl2SzPxhoJyQ7PYbOBEsvUksGhSLXcWbzIQf/vYGID
5KnjrFqJbTeq3aiJ/wv3HfkpLYj801mOeo8ePy6ZSzI0DnynbPIY6DK8u5+eU5qQ4bRFM+d5cNis
0mVpVNYXdy6wvCegY7MZQ6TIeyk3nsY4SBclYqmGPfQHbxtNessx10QVnfhmcsQpsxBIF0nKT431
Tgk9/TMeOcpXT4FlHSVfW1+Lo3/k98DVvDN88z7gIquXdBe+GYBdHrFSS7jyk5Dp5PV2Kis+7A31
GyxkFfmEWpw5XhhopIpQATpQq3hWJltKcSltLReWlHkPQ8JjB14rmktQVWjM5+qoba5Pln9CODkl
3Xf4YCTdTkjKi3GEIqiT6nULjLnPa7FMwKEhb5dF4vzCsCN4UCOLKRc9yz+5nmQmtUeSLhqyfLDT
EsfBBi1DdmZds46wRw4cRSrjG7TlTytQzyGsCA2Oac4Hk9q5PYdLbkFymUuiSvm/g4HprSsALIED
532KdsvAY2arycr3hJIX1kwW2RGPcTmD71i5ZZOv3YJfvNVMf+7dqoFvayBvBz6Y1UVfF2ndgyvq
ExPjstPOTD4yHh3tetH+Qa/KOYXq9602xOfYyaI9i2fcrIzgdbUlR04j7pfL3nu7RZGPQzCpAJVD
YqeTBao2Q5D3LL98OpQ8ouoIdS74l0/KiIofHLb7YSUSp/m0n0NtdCtFcxdXzAtfa+BY/Sc6M1ep
bS5gsWPL8vH11NIxcPsSPVvY20xVleF5mB1I2Q+Os4OrZO35C9S5H56u0Gjq73EdWN7O2n1vtf4k
R3pabtRUbp57Nb7zzFVZIuyNDZ/1EMcY+8JNcTguVg/KCkKBIShM0yiy4haiuoI4Yj3Y6Kv1th5i
YvgApzHCCsKvXCaI+xNUghbOqiOnYDmwFFiDfVCvl5CyInP9ja8RAYcB+P3yLgfMgUMHB36ZZ2Jm
sD/VpMU77wBrkq1KlUN18/FcnsF2+pK67rppyeetvViLtAa95qrudq6/2Dl+UYfrA4mLDH1M/Uhi
I3yZW0iGGdZmh5XBLtrTQEqSsHI+O/sHNoo6CQ4TTfx6UlAsySb/xq2j6E6Aw+3yibbWnz9gCCZ2
Yl6eGPnVTYhP9rApOiDpSFdhrrfDfoCrfvL+N3helf21WhdtUt2dH9QJfU2d+EtSyVVWOBdmSTOW
vIz18Hjp5yw5zs5HSaiYZ8Zuk0JJ8tWOk+tW7XTPVm0Zo3+q/9mbOwMxfVhBBv5elSdnCd2TvMB/
kO0WHnr0ahDU95SpomgXFQz8PDRLb73B3HhfLWK806CMb4CsRV3SYv8F0tOILXH2LhLVaY2WxOon
FmiY6Sw9n9VxwVeo8TUVjaUvto9BtlZhir3+jgJdF9zRtTTwJu8zfidBkcRcRxL3bKyXw++SVQJu
45MyRNDcjQbOiYvk/0E+K5X7CCVurPyTNdlQOyytqDIS9TCapq1Ch1kHrGaZvnszppOwp46gEJXd
Q4946g8ojWPDWZkRWedyD0MZkVbaDfdW4fudrxokNgZoA7hE8iEADsA+8MX5Vz/siL9N61edafTa
2IvKly+b4sENocctHB8QWFcyg4jZor7+17guO3iOLoAdD20FQDfSKX9aIjCXjvH1uhFQbJXnlgpg
VIt7IDa3V9vYCGtwlycS/07sr60mObbEDKixeDYEmeE2OA5618v+3SwNGu7eKksXALea3/Chlxby
ZXxY6kXtHAaOhHJ8gbOdcww+RExCyEyeGq9qgp+l+mtfoI0AVDZlnmIOMQNPD3eI/YjbMPufBxiW
qivuS3SLGIw8FpYuRu1YG9zqSa9HDmUTeb/zkpKBbwvZ8bICvsZBjGR+UP1WWuyWmkDfDRaTTQMh
7tPUOh8As0Pl6mJJoEHiKXLjsL7D7xtOz2RxyZ9ybpb9YzBCaU2U0wQXtE3HRCyhCt9jx0p0k6WF
mEsIzX3U0w7Ml9uZPFL2DfkH8ZKJObBx1tIplKEv9Viv5Kw+QoC/qxPpFOs8zMA9xSeSiqGwevBN
9QnqhcKAqZ+FFD7wfONKg/bIhJFyUNDTNV6R7qpd+suabpXG8VeJfsjM7Z/RHL4bRC3BYxRPaia7
m7EhshRhqoi3VRddn5C2eHNIGiZMIOuVfyoL3qZVYCjO/WP9qj8enCdP/znugtbIfUkPLOrq9ffZ
8GCodgfWtDrhy1ARA4GBqlXpCamiMYciGTxc+7Ueqh7qOhZjRx81OLG5XfA8y9u1Ho+yE4sKh7ya
gSuagTwVAbaD13Sz19FcYbPnizvZ/dHQbZe7mNboStY9T5Igkle4DIv+d59tmsorxWhgHmTApIFr
ODgxr2/rHSWm1Ya5fXrvWBEq5tLWU0K6B6u3HP9J4D8/zmDEjXis+rMfLSwZjK67+DVBhks6A219
DJJgbA2X4YQ9NWXT2Xm/GbTcmJVgWbr7xF5AZA0uVVCQ/RpbzAj/dBwRVUFHQDtklcZ4YKa9N9XQ
GJOXXS13XBvuaHzAN1iOff2TEETyy/xGHWa3Gdz6bA0J+VnJY/8idGMC/dDmbZu/goM0FhQhh33u
zKVYoRYlmyMIEd9bNJvBH3Za70EC9myqON1tL27rcxbwMlbeHApDh8BX6z+WpI/2Oa+KwYcpoX3w
0HqtKnOsNFQFPuHtKdulpYSJRUwpBL2pqx3KREgg8AZq0XdAbOXrOhAiwZ8hW7XW7umS9S169J/2
kD+6rtKY32WaPWnmLVG1Yeb2eqYMvYJ5ZaNrj1wAcZHRPJDquqId6cWbYXXShkZRQF3o294J02+4
IdRg6PyFLb/n82PeSI8432lU6tfgg8C1F7QepOdEPL7QsRRvNPDxyypfeOEMphdaEU9IrURWAii/
kpl6at9zMLAvWc3Pn8KX4dhqWmWp0+AUogqlSU5yEZ+ukgpO+85idz11TWt1lOvdlCWLS2EM0QwN
sB32RR47qdWxLew0NPG3dS7Ikcau7ZCZFHF5xnegO3p+RSPggfb4QbQQYEOjLKpjyIezjMeTvpsA
VwvQt/wyW839leTeHG2hea1PR/V2H6x/ZGFAycBRx1FTUS9vTi7gyKVkZBKL7+xbcdTPVT0mIhlh
4vQd9PDsZuOfMvAnZYfzKAIHoGLFl7LJWEeEcqhEBgF0wXCiDFfwfG9kVqzUM+LCDDAaOKW31yfk
TioJvvpRCgU0lZmSNZkIx2aToenG/AN9sE5Gf3/T45nb0vR8EdQBg9N50noI68neJIGQ8uVCrtc7
zfofp1/iZoAk2YFreDNe1lds9PNDisa9yn4ikypEY2PKBuJ8HGSd6nGE4QUuTUD73jQnfqNlSlis
M5zm0v8/uQ5TRCHlIfHAoGvqK9mlPlRIE8YOAnI4o6dDBCjYpzmYSZvzzYo5/TJfl4CAgmky8TTc
p6wXI+J77I9rDqOaif2YOT6sGjCgbvTBG2AdWU1l0tBBxclGRGxN2YdVYwrMJ0oc7RBjTcIUQAeF
mPqhqYT1VRfLRiTn1ydeZpSa7/OucsyZZArjOjA0/lu4CyFomYGf3MPyu8orCzLVvB3TS/w4ab29
vHOKabXYKgdEY82vWb3IJL6z7IYmbraQQfphgqTf7r2SK91yc98s+UUAUr/NQhmw71Fowwvb/4oE
WocG5wAVB9zprHJKsu8hDO+KmT30M9Ls77+8BDpDJHIt5No6uABMkkHVmBEPdJGKmHQzIV7ab7mD
wXTPzdjeuHEaRcsMwv4wQymD1CKnKul5hNtqsOE0Z6YD9sj6C15s4WqVUqJyAscKfUpV6aSb7V1y
muX61/foOPfggdgpMdU5Yvr1NmUA/3Z0PI3OGtRc9CHoO29l8vdlJG5qwgb6PbuePVhlCmH9WLl6
jRjrVMMSBQqAuTGKfuXZ7GxWBXPlZDTX0NYc9BOVfecVMbdwlXM74Px8YRz1rbKtD47o4IlAOAcK
iqivHcWc8JnPjKMXUGMvPKGUI/9ZGXEaIxU0ghVpimA/gtUfE8ClMJ3fKS7IG27QLQzuupXPJ4dq
P+/eBCUjxppBYFMWn9SsOArLGJdKXxoGY8WDuYbS0+TWFsb9E8sRe5q0aXZ/nKg0omtDmIGIs/xk
VB8zGOZDzM6EgMkN4YxWF9w7ERoMAZCfA4BvhPUt/WjQGm7zL08DHMMNSlUL/IskPDrHufUiUIVG
3E8W5EDepJxJPQgou33dE4kton7IAbkvEY9mlYHTO4hik5PMdcgWEmIgI6PirPCU9oF2YskbjL92
wDxgObN5EGTIgQbSabd9cqcF6GIutJuZ0Wtcnj3rGQEMb9lJn+RiZC8lQ+RkS94lF1BmUHEFMLk5
zgEOkE8Ne3FJTHC2fWq6TBWNZxJDs1Nt63r4Lqpc33n0d4tIgSbDSvgVzmD7xgGCrr42XloujqGE
2HATcjROOK6lsqOHTHJvkKpA/VbAQBRLYA0C0NGa7El5+5xryJ1Kt2URY/n7Lu17IGKrdf/ERF7E
ec00P3hezzWc7cReYs4PehVMQpF4XaVaGYjjjd4edp8WQdi5TyO5bdhCAxYwxcZxnm0tSk+981Nv
tqkTx6T5ILUS424RMKKzrCpdNh5jolm9l0lC+RgdyhLBc9hYEg4N9A002fmnQf+xs92CKRBbNEWh
RhISAGD1hFQnXqDWjeItqVa9N2u2lFmIDWXPqgoHVzYUII8m5nAlwliuRNV7fsqwTZ/smtSKKO0G
s89p5x/3e5bhE1ZSQeUYM5pW6zTYdY8GMoQQVmT0MvsMkOTCVaAc2POmQ/wtAXYaQm5Rda7i8vtW
y1Km+Zly7klSLN+9cz9w1gpa+QDkMOs5q5QudEU837PbyA1g/oonJU/Mgh9RfXZa20VlaoeBkBm/
F/5my+e/bV7ixedQFbT63Gc3h+9ar6ndZ4eQQ+u25XPTq1VfPFWms5x6wu2UFEdsWcze0gGnNfe0
sTGV5H2yP0gWBFzIHW7szvb38tpuLiM9LEMRZYhQGOy3C64ZO7qR7qWHJhrpgDQx73WD4R1V5pS8
g9Whn9yY9Xni4KxLSWFD0oavJyT8Ng4YOFZARsLWrkp6rmHUqrvo1QJ8OQqJCxe6tNa6Iz+8HdbB
BvK7swTHdNCCg/L7N1mz0P4g48y+Vjs5EyEnIZoGLJoBdwF5yTC6InNHx+2+BDeE9jYAdTrq1H2Z
FeVuavDkuB2mrc6KFqf5ALSeItLWMcTMpZwOCe/eF2OFjiU2uxxRhaP041yRWFsu0PH9jKUX272O
CKm8DFGPCNDuSR8ekAtzxvCMNh/3kp1HiokShAEiz9lRt4ASJFSWv7K56jpPN7PhOZzQGwMy6ZZS
Z9JrbE7b4WK/QfGRpAmnGinyCGGI22aQOOEBfNZSThxTh/nFHUd2wDbPjMxZANFlMCj6hwrWCJ46
QW4WB+OUoLV0twldo9pOlxL6Fo8p7/WhFZ6UZhCLxbgzJWSYjtByRHHlT4EO/sCWRjWPi/j4kMbt
z+3DearNkiokXDsjaVxk+4fs2toia6AYHl11+6P6U7ByYMqnTKq41ujp7Z+jv2j+WVCSaX70DDNI
u5KuM2/iiART/aY8WMWx3Ws/dQDRKk9zLCp/w+Yc8a1UHcBcxOhx+9wSGD1T0vOvsgi303jsXghC
yziGWfRGB9dSq1gef2aG6dVzHORZDJERJr5psnh12gmbK7S/wFGRmqyHMBoaDxpKTStpG3TlJtpn
eYMUZPbgrpakrwADijkhiiNtyxl4PPeZeOmvfCaULwdRs5crvFU5M0ma8nw161mjeNO1vL43AFU2
uUyvAWnW4V72socoENQhxQlOVbmk3JBThuAHPCswLbJxYzRTy5H4xDi8i69zUBepKGQUjp+Fl6sy
bA8FfPbYVm7vZjDkmu3w0ubgyHVXISi51bpkFv9s+O+T46Kv6ZBT2aqTk0J16jJwNciyCUvJYqF+
GYFUMeANEYqKxDeBz2xwhSDVfFtyLv7uAKHzukl9J9TRE2jiQf5x3RrfftXQgTs9Hay7qsO05ayA
pMdYChhAuqnGlwDARe6SYiaugnLhjm8Bzkafj6NpqYoqG5zcoNyscXcGfTjAvTdfbLDF2WPzfC7u
nRH0zPaTTDHOef0hH4mEtXO/yZzfenMSbEUlodHqsWm/O8GaAqIyK2n3Bdg5W5Jsd+z9z9wrRxQg
CxbDQnNe/Q2VtL+AZa+Ue1RjVhZoaZm+zzaS03oHuciWHvrahIKRdS/SlBNh3s3Z3c1fluAFpMLJ
zH/YK1be6A6BTTTIPIohosF4b2L9oNu7eZUoiOc1DRNw+SISZGnI0WHC2vBvRJ5PH0oyboAAJ3f/
OO2J6/s2LQtkW3LX271QoP4z/myi7hbkefxKqutjkppp+PqtOf8FaIuA/Nbafg5K78iOQV7Ug0M4
IiiLjyuDAtUeY89iPhjXFfBPKYnicUvr52a+zTccHdmR0As5npZWXoT8k1Cyb8BbZlPSZHBxTAqT
n0sd19EDpOXCTiRQtqwt000rGQZ/BQefxpJygeqW4HrW6rqQXdyzOlZTKXZSkb0Zi0hXjGCG9vgq
7d002bYtiS47AbMpNnG2kmB5tRNIZyg4H9MxvXugilz3d8jwVF/6JXyp21QlfjBl0UopZcns/Jcp
qI23O/EDkNo/rBXqJimm8c2k0Z8UszqCBg2E1VW598ouRTnuNBf2OueiuloGvRdp1dJsB67oK1K8
gvj9bB26CRMklvgyKvjHE1A6PanIYPuwWIm43BWk5S+rnE6bAxi4kd5ag3pz2sKos1lgT9VzJYCP
inzTiDRF7Uy2Yq1mga+JUCdKyZqaYVjgdtinU1sFGsedpZuzMQi18Ia7sv4Km0VeMED0mD4xvx1X
UuUOdsshWq/03WNk5MKqcF24aMEFVekNFlosozcWZMokCuTJ8lw2UQMbq2quOvaODgzTfE2yNRe7
ZD6aeMI6oEcxKMjBjUtodafVlEVg6LYlCuiQqevKrBp1E/w9d0FS95vlmdelcSxNSixW2GOBqpQb
H73J2Zf5S5iAbQjyXIMo87T3OPfGFynN70imaS7sA0XIQpdGLDmxk2qcV1TiSH4eXxfycojwmidI
19Nrz+GfTie++a9ApcZTKOY94aoSPDzVi58Dbf1zJKQQN+RJW+oFpuCQETuLS8Q3+utk4vfDVHcy
OqFsY4HiV5ULytmll3TqvKkaqgKY/aBoxOomkw2LYC6UFgMSGI+HeJbS9S+TT8osekYchx6NlyRF
eOdIuLZure4naRWdlRJL6DIA8lAIAwjwsFk6B6imwDeaFpdkDQSYDIhbF1tIkncBfOPUZA5yv9ER
+7BiKbS24Gf84NYHW1KjnDnM+7FJxKf0Ngl0dINIgZiSm7YiaNUvBOvsMuL8vhqj8uASLRTyCKu+
P8CSyTlHbPB93KiMwmeWWYLZzwgoD9EpEszhGeIX1WNtd485EO0MRnzPs4BbsTqQkeJfqKraJBLx
TT2AEs4csE5xMDJwCxzW0DGv04Jpu7But/hgWUMieGsxHhaAhw2c+4qA5jxIKhs2ckphiY1xq2iH
5ZXbJYF+nCm6OE332bqYXt8VDy40VZoxnVNzqRUkHGOB73tnRenc4sOCDPCoxETu5yM7RHB5ozdB
VkidHhdHgVk5+5qyfuJGfXiUrsKBUX8XHi5svpufUL5lZgzWCQQ9xizj+xHotpm7mzD7EXOm0Wdc
m+SY3SrlhyoQiDrZk4Iz04neZRqClTqtz8vErTijQT+8+b2xQ428z4hiVCHZhq/aPKHNaFDKk3WQ
nS1GV2qagDkiy6ARsgN4YqqH685zPa2LPRE5VNv3rDrWjuBDYnXTWbQEmmGn8n0g7ZwRLI8RQjWy
+RUaQdigh/4Hd5HYYEwa2lXTLZ6IW5K8JL0yHpM/vy4ZESUIawWlxy1L9T0kVtgDrF8/4M5p6rxN
h5HzSc02qkqq6rm/BorUNxCsZfg1Axsp4AZ3ALXtzisysg+yBimgkZG9s8s7HOLDspbPDvJSzvfC
9SFMAUZbiOZni05zgcVMNSoNKA9p5MYY/TMHTZXpu5Ov4tI2YcjWFs6r8YwSXFi6U7DNsS+HK9Ng
yUM5VvO5H5udkmHtYUjQV+umeOVN8V1RSjBJ+EyHFtwrSUa1+bpCzOzmi418ZS1zU9mVPaRQnapW
BwuwRChVnvhJCcnKnEp0LO/19Vt6aKM2JNjUmgFD+SIkwhEf3hKZs5WuD7sfhj04xFeItkHLkWYv
mF1S5RM6UgEe1JI6b7beOr1kZImLUP46CWJfSEAlPEPKoYQ35+DR2DQ4FDW1keJVOvtNx41/3PFe
FTxCpy4oN/E3UcbTR1CaigZNYi/dMPQa3nX2M9bjVj/dCEDEfXibgTDpke4+IisK7OzaKB5zl8X/
biDgFFtybY7zMntxu2ZrY+RMHV+RnJ+Osnx0QOnvGwOqRXiQ+geQqHxFQMqJNs21UXW5eq4JSUkI
a+4dDzdqiOs9JyRyv4mHvlmPz+eZZmJUcnPJ7dSZevwu90DD77vwiqmLoqiMM25P80nqMGJ/Cj29
28IOCwPX36v1rKpce+Q3CrAwh7r77VI6jjMQqRsSKNzTePeCPCXpneB2cjvI9Soyqbt+5+lUtcCB
HT3qqn93qapfSeIuT4sk6HsZ/Lkjn0bNAUO6FPtSzT6QOGHoNmeIk6IDcko2i7dHoFja7hYeN4p4
s3NXjX4hnwH83lUMTUJS3zSa+v6E7A571wyX/s3uv6MeKMgvjtsEKTpD+PM3WhliTU/YyjIJ9WD4
dq+/7TPlQTxY/hitnd1EfQIPbHOjLXmJO81V/ID+SlASRPBmL4CNMAR5ZnWzz06hRwqVPiQLJQxs
9G9Redfxn14fPj4yt+29Ep9efJMq+kkJiyHA/o+PMa4GYoFlzFyjm4e6CrMN5M1527L39hEbZIcL
bOX2a3RjW6pn05h78/yH2+G4mnP8yb/oUKnNsxYBiox0iTX/HsFOMGCYqoABRjE1bKyoZcX4VzLh
g4KJ3956XbFFXPFynz2HD1z+sWZTohTIYn5S1wQzVrFO0IPccD0Xqp2a6K43yhXaj4zFZDQrRA62
oeRBxtZk48TCuWfLqehcxRkeFpk8WU0YdCX+6UU7FGk5VfD0w7sH1+xVxpVtsOCE/r4gOwtTL2ts
lNMrJRGGDbDXcs3x1QGNfBhWjMuDTfZvujs6cfA7ljGf0eO5+Y9M2x0S/p2kCaT6hiXC99F8D2nH
REyXiRUWhLRGFnmX04Il63NIvqOuRGD41CkKqvZIiT1BNzRM1IMkwWvXYMYPe2bSOelIp0rZENF8
+9Jn5usSUTFpdIx8EkcgEO38+1rrqAnHGxBCOCHletHSzFAUCO26aQUZwrwzWXc9ZWGqgGqO0n1q
IHBJXGHzb49MBKiMw73V78TsSTMM6pyGLUVPrZjoCm8T22JVALGmdBdHe64iJUuFRi7W6L4qH7Pc
DSdWhilAwv9fBMAIf/lXKf2X/B/QWPdZ6JJQ8ZWbDnTLbqpdNs1HL1hOtuFIBY892S9ANzvOH25P
KA6pxBRy9mM2c9VM7KK+53Yyc59yObjiUKhfzGqYN/67SDk9/JlM2Le4TT8Wf7HgUdhJGikYDUZW
9s5eOtHqIUJJVb0rp4svA5e1+mQPelrA7THHgolrpuLPNMjTfEhhVU4OTsPag5GxGR3XROogAQnQ
nG55jCjsXXnHdBP3UWY+mh/I7B8LnTnKvYaQCzzUbatZaLULNom5OWEa5sBfMX4iqy+/Cth5U74I
bDxVRKz2kUR/9X7R2CUGeAOamMKCmRirjqpv7/u3XTygtXjwPYSH8TZ5bCFSsk/ywxzokz78MQ//
Mh5X8bSzPIYd7pw+zzfvtG1GSXSzIUO2U/oeEsuxtlNPLct7V6B5/t7dZs/Jhb6XH+OrEB/uSoZf
llFTYBQBdaabWGugMu+V64CXkW6iQN6p1hYihana0hY0Ej5Djbq80LjLfhb3Z3lrx+cqHL9i/kK0
4Q8WbTQuKB38UgrWUBaYQt6eS8jMPuMbQqY8hAYMNStf3/SEbcF8qQCrwrccMDZRMytLJkvinwpq
65lIsw52dB516KmLsud/mmTynkEmta14/Cb0V4ed+hdKcXBkcREQ5y4jHOaIaI8cZ2yFjsE301nG
+wCXm4fWGNf61Ke2rkvT6PqOnRnMoKxrzq4tNl5B1sg9use060PmwqKAm3Roh6SYkUegaR0KmN4O
whhZxmrR/xD42r9KeiFInv/wW1ZqbZPLQIW6l35GmMB3EbaitgAVixrJzsBWsdKEFkeVtGkJSj/e
1B59Y9CQtLiAgn66Dgt94dv+zLUqTmX+HC5L+66JBkYEacTKttpU+mGOsFdxFskPYJBk2lLUDavN
HURos+fEHHv1hXiZSr3SqeyWUA6RzWytEiq/CUtiiBhNm/7dgyC1VM8ztruwui0q2pqeIB2UUtvW
MDRlPykUkyF7b6SASAayqZC9II465ig/IN0le+DSyXhlGMH3J4NAuzNTn6SwX5ZXC6nANm4IzLlz
iqa1yujIpuWQNrafaDkF/O5tiYt8c2wO1qH0CnvXdsWeQCZ91OCoalSLhKmkkFfORqmOqMVjvaBV
qEVXEaKIQgnJ/kuq1TwYroKfhSxwqfyqFlmnaksxjuYfhMqo++qaIXgcv7DFW5wlwTsTCiWl9KXg
zi75hsL9bwm4zOJEJtsnSb1mn7CnNNgGY2pVxP4O5VucL0RTFhKC2ND+DRGclqBMUwfGJ7zP6F1l
HNzejQFt6JVSyU1CmX9huMWcGXAjeviJ86JEi+9AfCKLOccIpkDoTJ7VONr7GJ1r3luJk0Cg+qRg
rRgENt/tnUWq/UHCv8EBqvH/LHvcnAXKsEkmRIqjcW1+T6XWLYEA38vx5sTBMSYDvQAe3dWIK7rd
zhfiSfSaBYJHxoZQNpk5Y9CARHgKkMfkCVz5v/6Y/EymSNwWzUv5sKMhaMzW9OEu7gzIB1ZDamJ8
r2OLCqOWddM4Tbcfc18FgTTS3Oo7FieWAyA9Y+T2Yt8yz5b7oREM/v4JWRLKS0kM7vf5j8MmQr5B
I1fkpFYGBPvSqYx16eaqyqTgnpPvWWfTGl8GlCSpYSM7ZQDc73KTPoLjz/+QMHnLyuD+cEZOmqdQ
U6Q/CSqOfSviNfRmpbUWvVqSfC/K8LH6YhOy+MNx02dDctbRjqcwUtaTIvxyJel6p/UczB6YpMub
ZhdzdACM7xF/jtNni4cyznb+6Ebh+2GQzGFdDugSwkoEtTTHL0JAvsDBPy66WrZ8PRFv+8AJdRJU
17hkOWPREQcYshslRc2hjTzHDm5VHY5DMTRT29NlwtR46WEQskmru3umJZg6khamoPMxCao5nHvV
gAu/MdGPNJ+rOxXcaIgJZuNoyKCgnzscIICff9kCIeWVpV+mO6fn6ETloOouzlneOJ+gOdEVjj6q
386rqblk5TbYlN5v3p8CrBw6r4Agos4f1tYR+KYxPWzTR06/MRh+ZyQemYekvmRzSrNg8vTLTPvv
1bU7EmQjg2U0JSM0vy16o1Ow1khWx+Ga5HXksq7UwQZzeZEYUIT3829AMzbIHETHxDjx9VDcoUSs
Z98iEGhMaIUZDFNFhcG7oYuThMyoMpZF5MW/I/FEVtWrP9hzIFQ5DLRHIILDqaLaJ59vUUjMr0KI
sIIae710cFgvR7uOHHhSevZxO0UmBox8g69vjpN+G1gZjt7jeiNUaL7D2mXHpEymJVvyNnxYpyR2
v4x2vJ4zHsP1g9KFTHF/lvx3H7aTt7IocWfZWCRdyCntV0C2ftJmIWqEpLvi1hBs1Ug2+n3oa/in
qC00msfZDHU14xUq2gqQ+X9sqLfH7NlNcQlq1J6l4xqqM65UcSSLEIx94/b8z9g9JU1S7ABqGUv4
CWSpkvkkueLI1WV5DTJxTlVih0oX23GZA7F8oxt933w1RYyK7z7DuneEDAeFT0+8NoodeEF1qZu5
3GMZD/+ayBFEO39hBEAfCaXxLIEatFtEZIvOc1yURUmPC1XfZyz+OsLwhUtojX5exOKKaDKbpLCM
zkzb/s/7s3qKFTNuZvenv4FPXeI/FL1a3JcOUZMZRU97ATTOTic8Is2YVkcpTgyVgcF4LJaY57f4
3DfGSzDR1mM9bEQSxsHyePHpZ4nIH8t+HmQGRzhlj/vGnLLI9+ayArAnrBuakuNeLoouZ7UI+AIN
KznfoW2/DxgkIy4AC8nOFR7l1X/7Aieo05Tgq0WK7iWH+BXB6fhqXtmUlfxsBVt8VvvCoRQHAS9a
mNqdr4syo9adhvSzoUu1Z16dxbhLgPttFLl452EryQQ7OB5pF9jUL/5q+yrQEaHF4TL6NKk0324J
C5UZ2BriEErowFQb/cDFaAGcb+qr/baPNjp/yImFmFBNB9IzaQdbIaMbDHxCsOpajtRQw1WZug6e
0EF/tr9Izwjydjuct1JPePiBmIOpvE8AvJkTWBFmmVcn/RLidxHgtXCoCFkb771ZzsTPqXEdQ0Pl
HlGM+Uyl4RTnbH7/EcuZ16f+G6aslgDlELzD5pybfU3kJ9W6/9SwqZniLzIyAS2N+pqmrqSce8oH
FVzeFcomjOP3KcF6M8MjqE7L6fNqnHUAfVCOjQLI1YaMJYK8Y4ouQhqymKQ+19OE+E+0jJNjN3ik
ztS1zNEtXVmLIhlBrQPg/RxuWETMHNrYgIXD4Ecubvn3HgL7cfetgOnO5CqPHwwiq9TprzUSyiWL
9Pi1ZeLf6Pqq8rKuJLbL0JY8H5M9b9O8MwvSoqOqMyG61vn9e5RMFfgbwz5pZ5Cn0FwQkyfUMH7Q
r0FMvRfV4nrOBYwUHEFFa5b2ujlcHBoTgEW4ysEfXLJlD0iYT7mazoAo3IWN7Xp3Y2iIduaz1X6v
3VCRcPSzIUiglW25A99waHCU/l347cWgOfHuO/opSCpf8DeohpaXHN4g0gabWkor/gHd0sYfiZhh
zqjbWlSFjFIho4EiA2Fbg9L+BBagPzBMss6V1WefQOmyE/QNIzGybbcvRdv/TsOctOVJPQHBXTsx
ZnZXaGSPWub/4oDVG+uV6DUbcZMlRlmENxln8jMxUSL40zaPiW8NpU2mqE9shW7CZHeYrZvPqpeS
Js+FEE/GfZ1kMiWvmiGF+yl1Qixzfp8RYJHXf99g0iFaF+sZaeNidR3tYJ+k8SFmD7E64I/GnC/G
LV2glBhDSYH50GgE3Fqe90SIrMJezNPIiVDAeQTkC7rmaV+8YDmsmL72jftLRxqD6dUQazf61OWD
1v8wWlz36dx7e4RCMCXZYPz4gEbQjsZR4Z4eZ7cw1Q1NaNlo5/DvE3y4DwrP6DDUIicQ1uKHBVl0
FQkvfw9a0j8OJyhBwR5VB8w1vfPcnLiKfrnMCLdTEY6Ry9J8mwDrQWrmv+gYTzSiAJyK+T3zYa4u
Qu/RCase7BuJIZM6x9WPZxM6/WT8wAmFTsYCvNcYnVNOpBPbZ4+XhVRuZ5/Lc/Kmnff1v87rRyVm
zeK05zW/N+rEZ3ojATjSE+NlIYkp0tEABbYnAVIlBYSRP1Fyj1iD4s1+W0Gd1u5FvPkxlrs8CCe3
478PiDDFu3GcA89D3eajDN3dqsGEDWovDFVheFP1w3FAJfK0AzCPpIipewRDCASWH7sx4OhLctmA
BizAMCil+p/3vzZXfFLowbEqwFL/WHx7bImyl+Ul2NY1JPLX6wk3HS1TKLQfwOh82tXK3TIik0wj
j9ik4HcEMgQBlZE6FMALEYR/AYwwxg195h9oNyBMjJA8NIIqgYwaT/VFvZzGQj/1U5PMVOE3IFcs
XFYHAkjxTVhsNhokDl1oDEHe1XASlWfi/7cmBV6hvB/Yj91iFZGQ3fpYvq55EDkHecdbYUtKrUIn
GehAOe/r4A2AIJNfbOFHhrn55TTaDHz1UjUsdR1gLM1Dnc3KmoqL9ojqDLWIMDnpI3WqNIHzyXFH
UVKXAKocKkSlAGHA/QFWT9zYHD350ScJKRvzqatXFDbISNZHpg/L8T0mnDmjN31bcJau6ItYlV6A
Rjf8BAhK6n9O1qOulNktodyh8qjnEdY/ndTdrZyYt9XrE3NMpwzeHFPo4m7Uw8VyB0X3yZk4wSoc
rgDmAjlezajOMbu2NiZNj6FEjlACpffB228KJmMRpt5+e0PPGSlhGL3Rv7u7ue2huE8T32jhoy23
MFXVOT9Q+420treRCl3gEy1dcgbA4BDDv4oPTgAJEUsCB5DtV4Ib0rcYiwpldtMvkfE26YMkp48H
w70ezT1XLjZRZ6HqLoTj97GW2vRluv8NDYqKeoZmLcw9FxCqd0vslpV6zh4vl81pV9xQ9KpoI0yR
Qt44dm7kbHlt/bRr0yGjkOstvRPhChcgFj5ZtB/r6AOeCkMoIpQQ/gOB1OdeSXrAfeH683Z+crD6
kAMETbYLKH8io1qFDfUxCtJGwI1EEjoru0qb1rFUUW4WVL4Yfts9IHGmw644QcXm5uTPbMM31Rno
DwFGEiozHUv73gxaUdnaobUf+kRoZ2kXxT+sN/v+Q+YYwxme13j4mXoBPiEI4Lt5+qDZNZ7a3PQQ
Uobpcp/dHVwH8pP65tiiYB7LTh2Uew2vK/VSrmx4Va326gp0nCiU4dLe8+NB2c66OqSe9qdkgn7X
0894YjYqnEmVc4wzEDfZvRjltGVWVaIZqk1xcWuBP+U++6JPFn4KspQdszJWUMaULs0blOq9DAVV
IQY8SmesIPdyAzqf+NiAe+8C5AYmDNq5t5XVxzfGULz1a98A2v1kEakSazZ9g44nRPKW8+q4o6NQ
nLLkVg6qScSz2PIIJnigIbvFMzkiGhP69LHCCoM8ArBQTB+IZ3nw8Eb5xir9HufbRIdBvKJMWeH5
iuTtw6JZN0iyFLtYzmELNFIEekojFb74zufSvfb3HLaC2G7zP2dg8EPLSaigQijSKdnhlviOFtJ5
84jjeRKP5otptrAuwLN0gK6jkuzYWuFI996gW5D0wd4FdV2DZ2DZ04/wCvuUiNA1cW5pWepkWik1
SKucaUMX1UKnWUuGVDGEbhT/dSQZ00hKA+YE3rp/Sax95o6NGv/HG0rqOQsnJWUkasiB6uIeiOYC
2y9CMSM23+HE94HaYpS98p99f4dc2iQ1hjG5R7SSttpj3lP4gtrAbTt3FLlRzLHTk1CTe4B1KnkK
CI064dCoA1Y23qgGx1t9i+c+PgpvMEm177qZzeg35O4C2N8gwcLtUIdyBqg8aZ8pQJmNQI/yAB5p
0SnMvW72XrTMk1yWnQ/7msONiYNwtS65Xkh+w7TBe6pYdZcXjWltxVx+29PpFhyXRiqtoXlNE42P
F8qJjByVVWca7M1UGK1yTPNLcQr96prEk26guJzMSU/EVYPiq0tbIEm7A2xkHYWQOKmxrwdfiiaY
dP+78Yk+5c9TGTTB5r9b22Gc1nGzRGe6qaEJMv0qojVNTL5GzXhf0ny+jxhhK6Yw5ARt/DG3QfA/
TnDT3tjekuxVEot9H03nw8SY2lSEgKyvrJ+0flQGswTxap02D2Hl4IHrp9a+I/XNVGV4XBq7gWkD
fv77xVJ0o0Ou9d3Ra/j3W8binYMg3aOIlahrwUUxcO8pdQ/bHcTOLGFL4QQuzn2aD3Y2Pgy6il8+
JuKX2Qu9t8HjJS70SZ5zdJYNcD2AJSyDyeD6LUhY3tcpmbfXTNg4dpI4shKqL4SiBttH+KjaRtLg
MhfgwPATAgzYJU5OXwzzz0VqIlNGMbVGpdAjl9kED5WrnQjh3hCjaYM8Y1ACNhXhhIaeQMgcbib2
tfrGcw/q7u8nzE65JZDMse4fE3cHsRtAqg9s5maCYOh5hPHFUosm8cms/GIpEdgHKjjbzRAwHi+D
0G1aDVvBUvRGlcjocN59UFQD/A7tix7LOS9JokU3pb/DX5cv/shH5zxz5O8KxgLeIVm/1Cu8gdmg
rPo2C3tOmvO13pTB1MOV0wLG24hPRPiQ2vXtGifxGxRjMdkPvY51tRRrcInOzW5DkYczD4dlxezZ
wQv/8mAw7GaVL9M1He+YHw2vBgsG7sYf3WZRoLA1rmk0HUNcDAV7Lk5I/QMmw6mSL+sKdoVW9Zd+
doyqdyipigM07KBcYsD2SQ5RWcXyHmzFlrrsQp/XVi3T16yfOXTqaaNVd9AxmraOr1U3k8aj8UvF
AjpxCIksv1pYNSUlbunzZGNsy5sWNsPs3pqOl9Veq+y5mkdhjiJe5n7rudR5c6F7Ctk7wNrsGepc
fsMHAxzAvOa/ut8q/4PfmZftpoh+qs6RQYNbFu9VvUUErFJxw7giTB7gwIk4D3BwflnlJMS9sRoD
+VGbVwwuG12nVi5z8x4TyNVjgTB9ac5fR7k3vJ9Eb/ks5KOptj6KCqNiUjK7H5LH0r+0YG73atqd
q2R+w2cTUo8X9Z+iShe/CTlFjWwYu/CJbGccw7obGZD3e8Ng7XmbfdahMATDwhtxdp2XNRfblz+d
c4rjQ2ZfItXf5MX/18M0NMw1YcHhuKnW+1Q7nEPChaMMuv563ALMMtWO/CU58/NSLPSip3qiArtm
1XS5/2evsu16+HjDGMJ0xbVrHEXiZrcBDiqn75x50w0D9kKfCA+Q/qvKZ6wnu1XE53wTdak+gNX0
BHnA2MPrrJHD8rJDmUzrIUMdTEjffcsACLuH/zB7Vex4kor2BeywhwO5h9fwZX+L1JuHzoKgCV2X
jkGwl4XOD0q8RBNDSVpv8HmgMG6cD3kJlyPmhQrcUqLYnFRu8oX/CFd6hzXJZl0XdGx1AkKDUp1I
QCRbBd4HKkGYmmMYZmsExs//fF0ub0IW+8PfkMVOtC7Y0pl+BBgJ6esbkj5QoF+KAitQZdvSflfA
octezVQLuVk06yJdiCTugnji2MNJIRYiFdry3bJ/idPW8Q2sHxw1+Allbtr0M+VEYTFlLJEN4UMM
f0iF0uzXqY/FQg2sofoFQ34EuTdmJJLbw4rVfZDs5g349Tkk65T5goaMRECePKQ+H0aHzlraNnIQ
TJsTtk7rXkp29LnWslJPayKJhh/wnrYK6fkiW0Hm2tWuGPFKEj5zWHPWmgQ5CyTqPHJpxTHKtb0L
er9ecqIdFb7MAgN4xQc8yKoFI//7ddCfK8hgTI2vKWgLWeVqkwnFpRauzjrpbRCFE804/oFSkrZa
/zcJb2PAsZYTcGS+3/orH4+q+8tqPgAQIuD09Ol00q0YCiRXHWowgdqTcfx30ntW0xqhUyPm8rEH
2K4O0sW2pP7GnHXX9/YUElv8btSXZGMiuqFsfOJlLDhYb3SUTuggL7baI51u0pFZYe3teJO7Ji3Q
Xrw7NSfcfOF5hcW/f/yWcbWUghXpwMr6armvWPp0UmlWpsQQsPmv6O3/fKrl9SubU9AGHwPs8S76
pL7kH8VEd/90QYETwjwE2je0n4HQLMVeAr/M2cJg7t7KBy7twec5WRB0AtS9jSVqVUh3oeP+Z0FJ
ZLXFF1KwV27mCQ0PZZI/KQ5jxp4bvMwoQLGoEkT2OBCRs9Q1p8VoAgXztWJP8u/OjOVQLawqA5Sd
j+SqenymH20wn+udLg6bDvSOHAGJPe2SQ7D1sLvvE5/9H2fu7jC0UuQWnr0PnmaGlCyFbjsV2fLP
a2dUwdjsxwF5tAOBRuri64obWZnRF0DLy0fBAhy2h4wBRhtMJ/5D0OGUPtoorbkW9AICBZncHwps
5EHQpGJj4DP2sewvsStBRciziLNR7Kix0958WuJFmryllST9pQM5+H674X/AL9luzuHatLsgJt0n
qhefjMRHo4PWnGUMIEUJj/V2DfC/wMJmRh/GrCHwappzrTz1uab0bt2HCHKKQ1zE/MBNCVIzu1/1
R/6XXQCTJnr6O7CXMPEDvipII2Ron13y1bqDlD26wHggjOSP7qxyfBkPLFn9WViR1+vlOJrKQGY8
Ujc8jE7SdbztvTHO5DWIQr3qz6K/MO+fAvnxfIBNG6gK0asGdFJ1qVi93xk3T4OD+1PLfFi48dX9
Vmyq42dTXirIw8s8csZoWlAFcIgW03I9x9iDX7QnQV4O2XnnUpdxlEwp/ZqISR+RERUw0FICR20T
dEJ+NYyVRIvgLppYRIukZVdDXnh8j7+z4hJm5pata2T/0diXPHX6eKEAkXnXeAdZOla0kK18f1wc
T8gJEVWtvY2r5Ofcs/8OxG3Hyc7/zyuxnlT/xQ35mZpOnd7X2yqJTp8bNn9xmDTNET2INiHBPL1h
rdGZrJCkrcIMTX7TQueRvryXZMwPQSyerCALsKpt01WabZN4igC+23CUVZmgmNFmFAxh7C1cgY4N
/lGySyxluW1BSKBUI/MDcrhyGNEJfIMVl+slWBItA38+JSJkFJq0c1OXDRTkZXWtFgHnf1hw5lFX
vmx8W4AE4t/8Xe2BRxAD5hEt0vs5FTjolM9yJVwzuLtlIFrxZvq3Qzk0XGox508WZ68Nkyk2lxpE
AkxG3cENU/ITHmKVrUiWQGQ2cPbQGf+Ho6FGhj2MWeh7lXzrav2kqE1npD1DJ78Ea5wkICgpev2Q
bkd7SlWDh0ktLOKe5ePyVN+JmCG5EEe1pEXCGUGIcMh/ySULdxrV/8M+/9WgB+ljRlXVKmfQX9w2
xh4/8iAvmYkoSC1BAE7+OHGIWp12C3qn4NjvZVuVXTBNQZL5htxOZOwMrXUIKHwkfvnfTvOmuks/
8ofYnydCIKaEcM9NL6QtaLHwXVtSpkZIyc2GRBfzK7Xtxaryfk/5y8FQ4sDF/r74SyswfBcTNk/x
nipAm2Dw0ZlDWPFHrgzWyGW7/fL6aeF7pSJ8v5GzVKvKtzqaI2uezmqqzAOCL9GA9L5WoLO9Jkzj
Y6U9VD86ngjar2eTEB73Jkb9KLY2qn9YQpEofVCXXcYAd5RBMuwFkoR5hkW54NRVF+PWTLd25Mhq
hl6ce3pVZsZiRtvZuuDnNGT9S+X0POG6Zz9hzqkHJE9Dz4KSGk+pK15mdVXmRsmg9H0DaNpf3CMz
KHmRH7hSNEdBjdcvk2IbYoGMr9g1yk+QsNu4wa5aEmA/Wew6sT5P6L6tSz5Hmn8fuf1ABYK/LjZM
BqpW73aeKOF6ZtMO0lgK/6EL8mej+zo/ro6x5Rw+aUj6rkV607yJYzr3u6YtrScnK+4LheD50WyN
507EVdwc2OhSHmLmyQK+Mxo2/ueufrlSwEyBrCgAVaYw/8u1hiby+y6GOiZDZym4lWmJkx+tocDh
B3FhRef5lmYnzoEXLPqzt61q5N1XcHJJUwjuYH6ABKsIoVfAF3N1jrl9TO0dCcL6JoD5pGJlX6AS
C8RlmKS2bUZBXuROYbUAOx/a3T++QSws7lw85STG+e3WtqfNqh6bP937EiC/hDsKzkDhS5ejrkN3
Vcztw7IGK2HiGmtSZoVwxDj9N/b/hnweOsmMgUV//3m45628kwMZACpkw5WnQtbbrEYzU1Laisi7
hOYa1ej/2DqSRjftxDf/QvoZXjqOQMq9J8xNRGBmIy5Nv7lxFgIfSCjWGsd7cU5Cf9tcw6uaPH5c
Hj5AeLxmOqUpAvGoFNdy64mjGGsoWZQv0txQ1tDSHN7CEPMA8f5FxCSHGPJDOmVi5Ac2W96+mjoO
wsjD2EWHrkIbfb6JNQ8cqV2zLADl8CukfcK3bV4Ff3R0mSxQuNU5LHQY35y61NzJLknqhjX7/QFQ
U+LpBjML3BJXKHsq5TakqVbyQ6d6xoiAfRJsWbAI97uHH2LXBiqWwFRptDHd94I4s+C5iXkp2NRm
x5R4YSRzhvzGB+2hSoyshCWzicH50ZDFgZepYURIsVTzr1ZlHNNWWqd5yQRenjtFDQaqrvu93ane
lgpTwGIjeKUlJHj3lKgvNeerS/b0qbejVnYT/tksFSiahLG6+tEqXQvnFy1ak7vidNyNrl7sd+s8
Z1xjvZueaCRBk93kubrN8s35VsMO3UHuaUEE8zf2xhE1xehrdPOevHLFzlYOxLxAvJAGYaCYfpom
6104ducws7eo+sz/Q2ZJ2kB1aTd7rYr3e0kdbOOoJaGCVXnJYSEvUEcfXpJdEbzmbDeO4BwC6Dic
/SXJHRUR0iVzE3eQr74Z6S8cb4etFPojRNFW0UHKau998R3O9VUuqCjVG7wzNF5MGdV+hO2m+Yl1
lF2yZ5H4Npxy7vweRf8VNSAzuYKuOqEu0ccta2E+8UabU51HaMUpjOfeK04IpTthr7p0SIkeBxlB
IfWXuXKz+ZbC+MJ3IHJ5BFJV+Gm6uJ7jMeunhYBuxeXmcDAaKGVUwHVjZvg6SH2RCQxFCbYlb6ps
8brD66hNM5eUG59PWQugBoiq0S0WIA4pb3OwwTG72hRsmianHp1CeNEAR9m4R/36zUSeuf4AQIxH
i8rPZA3etrkaSCQJooONJCDG23VHCChxuIbD9B0+O0ADKbIyQ2XJ/o0esv280AhnxhrSzknZYmWp
7j7MhKYpOYWFJWbDCjwjrMDvOftwnlPK/5ZcUSt2zGuDKEujNVMpuh4fTecy7Hrhk+qEG84KCgWt
YrQuAcfRSr1u6m2+7R1ol2sjLRLjBpUcfhbuQRRrZmr8QRjVDftZASwypD+zksLC2jYBdBergc0a
7+b6BI3pFOd0hE6grJFnxn3qt9DuxLUjfm8rRTh56eNcxzXzz354cKesyc72ePG+IkqVjVnAvVAV
vFVY+srmkO3QPSOMbbhpineX3fTLL30S8dRaBpPRJX4oDoYdzcO4DoMgj14EuQQGXO+czCbsk3xI
AkWFc0T2Wv3lqf9LzkUdgJqhW2T+PTtn9030XgNJEsMdKTp8M71RDIaRdYgZIQccIwJgacp2L5/t
ghhxZ2x5lPd7TR/WfcWjLyUqmOD02mopifzOFzFE3RsDqyPCDSoF6ah0aBwzP4fpbfwBNjVpu5XG
KHXaZH0aEoJ3V1MSj9rgIfwI/xQMyYVpvo2l6KqjLLvhH34zuGLbeRPxKbrzpIbo4/MVhx6Hcdbb
VIQg1eHCW2fbEvNYXAcMc5hkP8Y4+Jj2gAuxmWMmuBp1lFoBtUNWJa0R1sV7y4vM30C7tQqgF44p
Ub9A0S/wSurOlszacGKB214s/DWiaR7c0LxA7E1htNVPYNdsD8gssApOYjfXYRXscEWwpvOwMeN1
MV1mKBuTCb0YSGQZgqwD++2eZkGzuVgyulfIB+QO28no3E9HqmibU0JySZ7c1c9/i5TO590A8cmt
J5TuUbbG8qNmBPW8MrDbQH8kEZhaol35wTudftmggahaQbIA7RakMBOWXMg/7eHDe2rKz3dGn633
wXdZeIffqN858/zZGUPRnI6kobItJoqGR57aStPUyjLkhwd+NdMkApOzLiCe6ajinCRLDbOHiu2K
Nhwvec30hmvGjORauaEaB1khIeI62ZajXsGiyI7dlV9NDZ889A00rgGVa8LdPl4ZWRNBCmNpBzZd
i6TtIZ2c714nmezypFsn6JAeM7gnuoltjSn943WsTEmhnCIWWoBsiJu5s+pKmrq/VGOQsDaNut44
vgWd1virS7leqc3x6XVuPkM5N9KHSP+mB69z0CLLhJqX06hCGBdaBQsAf8DQ4u94LtyOBY98/rwR
VkktWFo/EdNuMukpbRv3eaYLQ9+SSbLgK6sbzMsmNbuHuWbEd336oFWA2Os7+5mwF7RxvgMTIzsS
w1EF0uhuucwlV/3QJG2jWb8V/wY7FT6bX5VkbmhKC41KJfw2Gw237AulFoYHwQK0BwtWNMIFaeCK
IbqHwt/1wczmasUykBMdXjE63B3Zhm84Dv40tTAJ0XIFSRpZlDtnfBkr7wcn1bZFoL3owOvSm6xW
1zs4cOAMAwdDywpRY8435xNkXpaQ2D+O18T8+JRG825z3gKvGTsizSy3VIHD0FjZRZ8ouHRwZmk0
5IiVKDh2LSbjlto7b1mj48S1wbRhdGzbdxDvNNyRMg/1Xfwj0YN90uRY5Yv4GuX0pvfCgQ41lIXX
yqZjQrGWYD7OmD4wbRxc+qlmvesbG2XY16deOKvNj2CVpCT4yvIVwrplyPBBolFLh7LLIECxQBXM
mJzL9rhTGtrTWWj65snId75jsP2D58Tch/St/yIsxt0inpyESK+keVlN8sr6WrAFV/q6x6G2dUfy
8QmJ/BAwwMxC1vBuP/ce1EQpjdGHLFs9/3N7AumZ4Lq+l0CkXcoSGBk6pEyB6ACVzl7/nVs9qrtB
Lk3zQc0Olr1VzWSU8OTrNtWruQnZzyTpTD5Np4GDY/dpPu55Z7wYe1HQm/JcEFT9pF0aKhBhMedb
Te0fMFQWgtRTP1MsdPGH1mqIvZB3+B9dTnUsYUTwe5sRncujXMWyayU+TXxNBu1mEW3yCYd7s1SQ
u8nFWGLB3jl9DbDV1781KVWFPBJFZm92ynk0AF8sFVRFgwsqsi+xlxwf2qpABS5GODecgWg+pl3H
QoMZqw0zdPlblMrRW6wJLRw0lBI3jHglL3FQ2MrP8Mydtbjq2juoPpPjr4ygdKe6hSdpa6Eu3fwK
r/lH+VFZtg39hjTdflDB7mKB7tiE2w27UMV+do5B20E8yMAxhUd3lk+S3itC9BivzJbG7zJWiJaE
+sO6FoNcKq+zlvR0VZNYoxx/SYN+dHuoCcBQ/iH4x3S6TLWTwF5FF6Zz0kJOxyI25H5eN/fW4zsw
17oUaHFfBRwHLWeWWcG+0bYDwgmlJYtnZNdGcporbiBYs4E0aHIjCMzBOhMEAKFjkT6DFhF8Hlxb
31EYAVO+S0VntcjlKLUoMfzyH3igD7jQs2o86loJsm+KOzKGq2IJCSLBIkwh7uQxW/u12C9KiHbh
DQ8Ep3f9bQv8UytPBEktRO+PbWkLUs8HRv3Gk+ZDjDt25ijXNt1RtfNzOmPYSVdq3rXCM8vY82mN
Tp+ck40dyNuZltqlzBUrhz59NEKsc64ifqrDC6mfNGExgEMs+aQ4IHlUzPeedqCGalWwdt8ShXcn
1dDA8dfi1fvArqoRNJZQO/BCzjdc0IpXb/Nhrw3/X8L1xTWt3b8kTc/3HGusAT467h9jMBHoaJPG
Qc2kmFNcqFFOYsuVit4kv523Q8M8XX5T1TwndhmwMCynzZbgpr+BkNqYZzcSf03vRZhHEV4ndR2B
euVa47Ju9fzHc6/e9fLwyCeqAf4E07nGVt36haxIlWyjMzEsAXViLx/It2065KOhagDzRNzMHxiQ
3JiX4fsIcJPYYW4Y8uZthZ44Q0U+aNS302bYJ3hGJcbUU0sP/tJlcdU57fBxo7yp84K71N9ze/Us
vZmWjpE0ICGX8LvCznaAufPKYgNaU1MEj02FkOJ5z1GPZBvTmu/Opbicss3F24+8VN9axdbqCKMH
XfJVsCwC5SC+bNmsw+R6U1Q0TO/FE/Yb4JeVwXgeXFAc6M+4IxEe7G4NM5SUuAvG925iMDayO6GG
7ORu45fdM7Y9G0cQN+Wl3UyRTrVxKd5tWShGAMycKi6kO9HyEAkCnVdkbeP4pLErAXESfnwgTJ7j
yUqtPSgz3TqpO8OpVGHWJhWStNvq/g7UDzH1VePjXvkh9T7zgSIkdRdiyIzyHq+RwXvlfYiwHxTy
iYjF3PpRffCWApYrjXrt8qhsvrPFgwG0ZpUU1Nj+3TPYAWXJCVEtZZin117TmrN06ME/iJEJDl1w
Z+4pH8AzZu9TskfL0TIuRaA4a+BRJeTx5aX3o/eWWV6ZRBLWp94Fb1nr57GlJB8lEyW6C2AWyjeb
2LhlVhyAs/RxE/m46Z2mWp/oYGTEYDaCh5HvJJnScg9OOl0XaeqK28dtX0xmHNtTMv6DYAHDJqwn
sTgslpqibXTFOiJelUmbpk9VPP1SfCjb3xlo0olW41B/vTNnxpKJ9i1SgpGfV+PFf3p/nKwh75lv
mLBw2RbpecvDcbeO5rLuiiYh03U13bXiaMxm1x9p4r6wLP4gW9P5j7I3l2EEdadcLSIlukRMWMPR
B9wCfyDP3HrwJNONzJPW9ZgPOhbbfMqEIwGBzkl//CPq6CIURs4Jr5Jn1Xuwod+v/A4ggwmI8ZrN
amxhWjN3hUUC9x9p8TZ+NUuz6InhIav5gHtVahJ3y4ACq1MilRbMB7Yp5QcApa+rkYfUIi4VAn+Y
7+BAZP5tzysGr26pTYHN2wrDIGzCe/Znxwh+WajAASHUNHHgAD2WWlu443AFCKg/8f9wwe927M4X
ixkfAWacr+kLbriHtB2Mptur8cCLi60mlj8K0F8nvQxPdi9rYvps2bfWBodBzeHR1cpfLql6oiN0
wprZSqo5t/yMka3CgiW8l0WRBy5GISau9sbQwtX2nI4y+CWGFrgYOneDHUlH1iOqG1M+QxSUgl1d
jcckt+63IE1YbJX5JUYhReGU75hLvMActByJDjaPRB5gb1hnzi/eHuOu2K6DukNVQOiN/KjrRCDE
iJenuunNONk80xfbJPX9BhWplPgun+CGwVl29Qo7d0IL0jo/uZJCwm1rU85p784zDvCSjRem52Mm
38mL5P74aQM84xPTe7V6spnDEh6Q0oNycN97+KE/CZ56TR4ttEjKdbZSkxOoAqeyBpTngtCJY9fi
Fg1SoT+pRc2E2ipdVzUVkZ8OEJIA1mJB9Le63fzsZsoTLXCLl6GpjuEWurXblDyGBjOiWbVPAoVi
W0nw1MHNmzwpTP3u2CMMDp0OH4AtkFjrSVPuwgH3POglYsLafdr7RHcBngGnVToC72C0JNfhbX0I
5/LXreMCRbXg0RWJGDcJ8Ac8UQtISr0nCGqh39+uFfSoznXrxhNNEOpzt04fCPn0JCvy/+GDaBac
p5glk3hgvJfn+HKt5ffULHsg5WQ50EdgQJwt+8FrDQqmRpj58p5obLkanijafKNZcNh+QVf/NPWN
iUn/GdkSzU+/xyCV5gttdgaQnth77UXcuytWpFucLFCpvkZMuRN0xAlEUv5S7mUxn3BjHkBNlYfA
RVMvFOb1uFQWrQiTKP1NWJjpUG2o8UyM+rjZRN0XBMUhEQ0Sv4E165N1MjPQzmF2t/ATY+s+bgKB
eTuMBS1i90SVyCjJhgzg8FS1lCdxEJxekU4nl+q5o+64dg5XClXIWNHsQy8VociTHLh2Uv7+N2oI
VlYpy+nyTJh9rS5Rfbm8I98NQmqkCZSRwFd1vx3E6BJ7Ln9rvTn396j9VbDyBYI5Xc89OjUGqkrQ
2/pME1VDlr2OiuLhf+REYpHXQVIhq+O6E7eNTPZN1GdU7If4U7DPrw01O6acmMUH8TaMcr6DPyE8
lPtXYhObS2Ik3cm4QCX4B+w03fa3g+9C0vjKxXYlpQ+SznYtewtIoPTyyFZUCd9NGBLb4Y12czl6
5jpWrh2HRzi70ys1C3ayw8fAs+slz8+91823UZ1dvaL8EWcHTcyfO9vCap0dJx3EmCRWowCg+juk
UTPFczXeqz8Zh2mcZ4wsiRhq6LF1JPDelvMS2GVg203sQoe3nLzGnnsZHqVVwgCk+rq3+NlZ3vmJ
hxEiebUC2jsfkfzTysUogCG/16xdh6Mut6UkMSX7rIysNwXkLM6UkGTLcZU7CNaZv+ZmmNuxIZkv
4eOxKcXgEjiWApE8idJXOuPARd7Ps99fIwBn1HkqmMHEa20TDT4bArmIAI/TJa8IRCtMP6gkVvgM
D0LSKCN/wYMOd/3E+nDjLhbbOWYPO2dVJs5+WP3sT8GrlDMv3BVZyn0stRZWYXVwehr/4lPisn91
YWjWIyNqpokhfZovykrqagu4Lcm56dCx7DnevZAfZVr3rx1hjfHqaHi3gepw+3a81nPSD3wKLRbn
Iu56qqau/tCP4J8zCsjdOvZ8GxrJHBev69fSHIkshgK5l86NgXPPrG2cbld/cT7uQEYPT+4YmUgw
IsXFFj7mAgLPv0hpW8xTYMehP6g/C58L4+vyP1Wvo0MANy7jCLm/Sri4EnSiam7Pxy04/IujBnAi
4KwmyqCyv9JvKl61CtWZH3X2P/E+Kn4sA4pJ0qsEDkkVZw+hT2t7JkbTCsQYeH/PdACtI4QCCnGj
KTDknZ+zYouUT6gFQKBJ1n5nnEAINXqQ8CvKrV/0w1a0O+Y6nFWH/qWzuyriqfbEB+TIUnUMbmKQ
wUif8su+MHtYn3Zg528cEDMShXbWgE/OqB/ihhKYLFQopkFcd7xXBap5DmKOkG5jcAtZmyLJ1pod
2dDyr/u8hqxSyUOO8pDz697iW5qQklRfJKhwOXWPvsK1YbAoLUb0Zub9KomcvWilZz0pv0yqmfTO
zP0hBvSRwBVr3A4UCzehbj+SWrB1MGA4wFQtK3lh1lOoZz7EQLrr14BdKFFzCt9d0SNaB0I8C1ue
C3XtiZvGCrs9kmGwKoVwgg2ioc2rWf3fLrXZjJLCxXjfFOPESGXIujX8tHwdH7bR828RsrN3JxKw
fDDy6v6ehCrr8cajPu9paQa/E872WfGtgPYC+FIOisB4Obdf7SojXeWFGz4RL9HTjaxgI/+hcWJJ
c/rzV5X04jP+o7kItXUtsdQ0s2bzTCGI/Oz34PIQeTJ7bSzi/UOGYgnEdbz6pMNTWfS3rtipcYaL
k4KMH5D5nT1dM5BtWJDSU8HiU9HmpFvnHu+8HxwHB1M79wfmCsAY98I6UMrqclZuKEjSPjtByvKO
u1GEOayG246XbAnwWykQ/tHvYKl7P6E0q/9u2V1Vgf+mJJyvUmoP2poROXgw9/tjX7G6YwTKSUoF
l39Kcyc16I7294VP7wWmOeNVKFJN7TNMnHaxwswwynhhxt+fjop2rafF0WWQMe4z0D2xwZLnQ/Z4
IwAsxivt7emsl+Vw8Bh0nZmbe3kdiefvO3anF46JhP3eAj/JUvhv5sDEka2IT2+dPyaju8hewft0
cXmEOc7L1ZyzXzJEPfDmOo3xgeaB0Z7jSsPxA41app6u7SwN6Gz+mb3KUAZK17gR1lxPudp0yWmx
bvk4yu8Ej97tuC5/W9jNjTVXnYMc3MGIh87Ahb5GFyGL4a+f4pkJlneaD314d60Bkcic6KSxmcyk
A5P245I2UUpGgPkxZr+7643VwMhctLfT3iYgAWieJzq86cMmfc/SQ0seU3FiHFibuTjQbgK95w1f
dRoF4Pf3drB8gj+2Ut3VSFmWBieGjVsIBPkhgoifzKtT2wS8XFJDPoLnJ0Rd6gUksp/pWfSLJ1Cs
7MJNCYT30iM20xJ755Fm75P9JU/8t0cYeyjFPYXZh0zgdQaLrMSRC+634llIqtricz6PFzL55qqa
fg2AYqoKVeWrF2YfAcJq0vzf+CP2C0wJp/K4IXzHpInrXFzJYl3U0ME2kvnGNY6/sFQM4+v7cV82
A6pUKmwS0vLZvPMEnf4aG6DJllftLCqGAG5kzmtTzJmclWUkQaGwc6EEf6Fj7U2+csthMbYreDr7
ZbFhtoGES0k6FsI9fOywP/vUSVUbyGR3ZIao9+XOO5XaDuQH8Hw3oFL5+Iv7poSVyE8KKZJNpdvP
M4nhVrKPhTvbiw2Ii48WIMxGJY4X/KglUhg3nhTlcYRNDPq6iFFrYYpYHV2XnhuddchbJnm8Vd+n
p/Uo7kM5AQSonHAMozRQb24OacUKWN6fYnUpkbixIDai/U4nMray0WoZUzM/CbCoQiRTGKKl2Gd7
uZAXx/nCTwvkW1TynPfbjko6gDt5zPvsFOFcw5F6/e3hP62iG0bNE8RF2xzpIw2ta+By8ifLjgHF
vsBBi3e0dBmGwHc4lZHtBTmc+/1lOXlK0tohIDNuOFPIq7dPKYWjpvEvbE5f6oC4bhDhw30cAzyM
Kc/2KdLA/gYXAugK+ujUCydJNToFkh3t75Z5Y50tw21yprjg/2HfUcH1Uxg1dhC0eC1Erc0iDFrp
xUzG2zJlRbuDDgAHY1WP47IWEJZ5/xQfC2cQrZecedc8EZ/44zOcVckhd8SRfhkaNQDDBUa43SH4
2QEnuyrGnM71BwMlMnkZVFoDBibdvQAKW+5MNX+GnqPuefYfLTqoerdq+JJ5SKU8bvfSIqIy6QWv
JeokfiQ1PdmyJFdFrym8byjLGunwxTC4dEL/3N/NEsm2jxrne43PntuBzl2Kp596QD1LWy/bWbJb
Pj0mByp5Dt597+zWqVOLFpv0JymyyxYIHShi/3xvTmKcjYGsV8N+j7u854DbndSFhmAQ41NHKYlm
TI8yzC/e5xNFgroOU7GuA1piWCH3Izo7MGBjD+cS7IQkc/V9+9Y2dU+8Qg5Xti6DjEed8jl198Zi
U7Osq1tBYGXmsIIUsWzKsssGn2rCXSFUzYvY3SYWf+NPL8Ftv1RwLgPe74wZugLZzfrwLpM0jd7F
SCoRs6e+DBTMEfddZIZGMiCvreZTsDo3lUpVgdFEWmFp7VavUJW42bBWAhux0RSUuKuJTfYfS9Ue
pFIP2VVPwXCXJWQXj8iLVzpb5Tz0NHS3YQDmCWbxmHAGBNZVohziYGBqsfK4UTQngbFi8mhDn1OM
j1iisHPpf0fsMgK3hrqAjsYF5fKEhBQj7ZOkZPIdfVtE+MmQz3/PH4FDitSAIIcl5UHHjhWUVmjs
VRMLgcI1129pEidsAnyy0yIcTg9UpWxXVtUMO5yLwNtbB1XeC3koMRs6w2Zbn1GHtlwxppgZK77s
UOaRJAITJtXo8q3N2UtYFj6FhQlWyKoxjxlyYOzzxHAywLpudxdOzKWmmT1Z8N7XHQrTxMEZ4/3L
1+Z4G9S9RauClrVNF26BvaXSQV5aiwEvON9x3XNbbmByMYf1fRZJR+COoLdgP7DQb0BZCfSGa2J9
NEtjL8idA1OnOZhdGG+UjEi75RbC1SM3BsJld+MatDNgZV7F2VmMtUkSt067NU2aJJdV6Y16k6CK
doWoZEtoTWlYu/4hC0oILQyeXDV3apXsvkAdkF1FcGjBGYh9xL0C6e8hX1mBorXztOqa3x0t24J6
7gXB8p+m+4azIWabr+RSRkHYUeLYxHgkGsBsVVLOnnCAsfKA82Aqy60HFRI2l+RwMCJa1bbL/Pma
PD4e7fc14RTnO31rjJddto8nQPNzJIZTL8mVdBvBzlobeA7WUm/ZXTFLy+GB4m0eecxUw5hiSEI9
xKgXwZFPhf2jfQyGV8+owYz8oq0UqILBCKI9FZXBWdD/c9KaNJ6t3l78x3+3sTWPtk3JrCvuOy1Z
LRPG1jpYbNZT+D1AbuRStwh4CEOYX+nZA5ebPzjBojN/3SSN1fVDXU4d56I77n4XUv0bk9owQ6Kq
b4qPTSpKoeq2+wqlRDUss1IuwWFLKXaITvkZkA0k82bJ2VU/7C3iThkcUGOovRuxxVMkZwQ1tAkf
znfDhzxznDGCXif4G39BCR31C6/ut+c2zYvqgVY4WLhdNgOm6MlfQYFkCuO+13Lqhe5cXNotsQ5g
pCGz85XH5u6YRfsWlVI07NSF8vjicYA9Jn41dl1eV40dumV5BboKr2lFuA84Lcuwg9XoiDSVHEmn
PrTCcW+9vkQRQOJgL12raRYke9PeAm0C25+oqyMJORdqyFgKJG1NX1qU6+xsH6dd71HaaOOsX/Fr
BloTFhEB8Sr1gmfsa28KkO8lFUYdJkdUDq9edDmuDAdY3O5e600clG1BZ10JnbZGKH0aP8fjXCY8
ncLq71JPxF5Mqlx5dYsftvWkbcR94SMjJxESAAh8BcOztEfwQWoLix9N+ILKRYYeYPzfWr7xlj7r
TqBXkrzeM7A6OTjx/+dZtsc2zRq1LKENxCMJ4L6CPbhMUqPlLYVhxQiDetrYELtJlnYsV5NHcW80
fej7HjjKylNqU2DTKdh52h+aHSr/ksoioCBpYpFBrMX1LQBdJrjsgqRw4zRougq/DFs9Hg6a5enh
KgxLodb0Oo0ELf3trXWgFHIaobvR1A+9/p/gubR4B9JO/2dlXaOoN2DL6VyH0p4+le/kRZ+jmg+7
5cAd/968eElA5ijoa84uMYlRWLi42OGmf/MDETr5xpJ2850d8wsvAuO8RoRh5UnFyvxlXBxpUUUi
SaRLFfFVdwiblwJlLcU6LbP6WI03qlCLTYWk2VnHn0ZP9TJiHnt/IiKSmVRia7Mj8uCjTxHxG8Ai
YlvY3gNsnDiX0UmHMcOm7gdsbCZ+98tY9NCCR5N/3zdNsnLJp75PwStg+QqxZPYJB4JlyQ9PVYQo
nZ7UTwRxoTf2sIaBLQI8mAhB908RlVHPm7unHUGW57FWiAyN/ncIm+NYdPTfZhnrW+tk74/fk36W
eE8ILAvSAMdb6Ndob3sB+z1g2VlGp7gFoTQ+Z246suL21ETRsZgMtg3ZVwUIMnpko/ea+A0zI+Yz
dUq5P0u3imviefIWTqCBNHDMh2iNhirXBRcsCUjoQOSoAOIxjHcsv4hh31vClewlfUc3FK3V2gu2
NWzrPLquo56i5WOcUkj0AZCaTHPa981CtdxDkD1WcFa2REVJoToH0a1V3jkHXbD0FB+lLZM8kjMv
d0j7m8V2na3s9wgWLGHgLLW/HwgxoSkrbhJXwBaDxwCgPQ9fE+LDIyo0H6i2mwYCPpeIKJF+lWkI
Um1GzAmm83iPu8CBNatBhDf2R19ZVXvG9FgdNy6C0dJO9C9jg/r3uypBSulP/GSOCqjhRt1HEvmK
+LJW8UZuxRVfRFvUcCW4+jnf5UWbxriaDBQNspL72nC1zBD8WXgYarZ9O7xHM9/BS1I4UnhosJEY
NG2heKTanyWfvjbJc9YrKjBFWMMZcXUpdvV63tXpL9yQWSRDdKbVU9Gm4MJbE1KY8DrShreCm6Db
D2rVSlSRh2Zfkq9Pt31J6wQAZoVJX1bC+BVZdcIovPawM73GXQLD0mCSR4VNXqeWs9NRSGM7drCL
vhqUxw1JspfVuy+rGZ0YbfHhoDlbZiKdFMBZJuGiYt1LsgHhlz/zDbRnJW0cnueFD7quw9e6KBVn
rw6gtKmYxtyLEwRgPbTQ0JMttf/zUPawA6Ks8x15qAuX9r1+a6HcvgS/HinljhjhlHEEabrftzAZ
pa3UXniRxXJRFPk1CSCtQgGyCiFgJ0bltNSgb7vou1dgiV4RRN5NFBn9KpJHgRtc4QkhOYuPKKZK
S9ySBph2TPi6iezpoDTpgRZGyMB/N1AIji3AFj3AHq08xC4ex6NR6JgHC6Wtow8ksCCVWPWDHfyR
sIsCq8Dc41qOua8/QnB4e6d6lPPGkXX6YeONJ2ZOpy3VcRqszJCOJd2OXAB+kMjG4TVMwXKSa1lL
6lSi4cdBrhkPVMRRP4KMH7mZ98hLyxHC/rYu54Hn+VXs471j8DsondlG4icWhFxpu8s/FkrxxnZZ
Uc/jz/RHWTJZlm0HseOOSFtiLnPI8YeWWOOdiNT5DapGvKtnfoejKGs2Yafx0VaozJTEQT7LY2dw
VNdHyhZLHadzp0aUJCf1iZ79ND6X/KWWB27Ue8qU3OKERaI4T3PnJW66jTiiL77TtARQdqQiCqRn
OYrH3eJ45TsrG/OpSAalwvHK60DXyfnoBzSm9gEfygwqYaNPYcn5Bwv4wQPKlTaHVfHzf7o+Wojj
4cfl6U8OkQOf/gQDAeUaZlXPvTicQuYtChIG+VhUJqZuPAJfXl6N8Hh0goroOrZ97ZYq3w9rUKSZ
R5CYGo9d9xkiR+/Eo4/HGnIIAZqkAbfPIX36B3Bn+lg8I3QXHF4MM7qMrWh9xTJgJ+sYzrVNPTh6
qnZGqKGPYG6qZp1ldKRKcGiJJ9wkmG+ZtIA4+J6A0qoRVARZa1yufSACP1fv4xQ0jKh++aqZuri+
B1riUZaz6Rk9kjmIezKhKI/9XHGB/EYMzc5XP++FVeBCZqk4Ga5ZPi2Zn9cz7nRFqyzzlVArrlzA
88M8OA74Sxjzje6BXA+tSR9gxpV9nXSoZcQs3cQTvD2slHiH5K+UMGL/soomnJnj2tXauF37I1Tn
8RK0IbNaJEeigdKgpdBxzi43Ae/y+z5d6fITDlQ/MJIlHm2ALMExurEnP4lsjARli00tOrrjl7tE
uGUfBkYq9rlDAJ7ojW24oubvQOvOfOxfZVeMxOyLnR53bP8+6jV/ahMrI2oa0fE8AstoK1uP1ACT
c1cdMsr22uQ69Uu/3fKBdwF3MvdrR1GAphbQLLoBs5kV40PtY7iml75PW2xvdylRAVDwKBvaVJVa
J0hiDG1tkfHsYIBGtdwvqe+Y1448pq0q+LYcn+5U1aYk+OAcmYpYig1pwgObuBJ6qdLjFNwOQGB8
aWAhQoiv5PqBSNYPcU3LcCR4+s2CH37Khvhi+2BZOkmWnqaOvsre+0PsP8kdLlwGVyzS83wUIO9y
OGOwrGZe+aN3Ox21My/ArA72nTvqXAg+Ghv12wbnZsnU7WrwEajah5YDuukQIj5aNY8IbpEwgsKJ
kjiaj6tFsy+JKFSgkSAGuIMFWt3+MlWjNF4NU1VtazpkcVLx9aUAP+3bxzDws2wuPj/k/dchBUYC
G63ERu0MR2Y638eio+Zo3u2n+Q132TWaS8QghoCnihkyrEZiwj80j4yBL2+NMHndvbfOfbKA2Ijc
YfKyfVx4AfQnWvELhlLb7SI+fom6MRCti05N82vzvW/0jQvayoi0APHxEJ5kC3ydUdNiQavy/gnU
aC5qroGRkrVk/m+ZVUQ0LIbD7LSppZ6Nnqs0nmKZeqKOVJGdrP/3P8m+/6WkmzVwXjGk2A9OedKs
fQXGREpjU1uqHj0SgpXOkUlsEjeZLm1QaqtC7b7icdLm7ArB1InhiR+eq3619b6nmX/wUp6I/Nuh
gr2GvdVjRfBnvqC9RcA8m5prULKFKTvBUMGpdCiQ5AgxioWvfDKQBkiO9uB4S3Y6eB39DwPFo/fr
JcNw6yYJHGwdvFp8JjUo1FDzCFCg+x6hSFBqLuReqD2KKMyo89/IUOaUIq4d3mo3pj5NKMeVYrQw
fQLGnRS6QoDttwF8ml0t3pGYTM3m4Lx1PwFJ3YU+jrULcd72tCOg4ToadnE9Dq9uXneC69pK3Yvq
oh/FSU1ijyQc1JYjJnoTUw70tgpV5cuax+kp5d/Z+WgwEAAJMFMHOaxNGGz1ulWmLyesvJPKxg84
6VSvIm5NCMdSm503CYjTxMYHFRXeCBcknvWzDp1y2SzPYdTyi0x2Y7XXOhun1ifu3YO9IXEAUOUE
Pt+QlhKRz/B0IRXPKIpp8w83nNfAmlRX/xPrvDE+YjelBSpds6sCJ6deK6ubARQyRiJhIJf8OnAI
WzCU52t60PbYJ42SNdf1mQ8vdk0jzWR88qfg5sWEe/AH/bPjEDCeFRsPN9PcSnXdQKGcppp/BS23
k9f/zlolIRoLBV9CVnLEjRexUEJqRqnWq+xosmQgwXFAITzDDY0ih+DhT9xPIKjIx9XxSOM8hsPT
jY5ZYykzz/IbUtZRyGvxdApXujcg+lDJGsoBDaPi15bKa+bRHHnnEk1I++LtUkh5DPj3qs+FxQ1W
UIk2X3wAcRASpUACf9X8J83qEbPwOpYYYF84IXWmMJ+hKfD7UyKoBF94P+2oJEAx3bhZJNQuaa/R
CEJ7ZEe+3Dwas/OAEQQiht0TryqTkUiAC9y0MbTZsAga7MUCXAWhXJUzCR0jyDoGLLgRhDAjTLIP
cRqzqZjjKyfGE5q7xfszTSw2bRg0hDrzJHcOYwgvXzM+aKyPs9QBbpGnD08RKbYywhuhCKesmVSa
zt/zEchl3BQQqOpYge2qlxJsGanDCc5hBpoDNTzgkzKcjovbqeVFe0ZddNOpQb0is2kSa7fd22CH
Cz4vd9AS3BXOds8/5Vsl+AOgkPDnjb73ngGCAkDlhhcqanxUK6w/xiyjA+FbqMsFoQ+NpKgtFnyJ
TIofHc2bwLWbrnrXGJ5aDmOQwwYfTgGo3F1s3Omk3hwVhXKv3DN31ckMRDgbCYc3k1PvXA+wV3XC
5fsAu0QOXAJneHywFkmyWRhfmFxU7eEGfDS8RRpNS4gz4ugvRFlT1Ws7OhjBIrnyLs8iajHMrZV2
kf9B138I583BZHt8FAx4wgAQFMpPMXxITzZ+x2W43d49qDLmhXqwyNfuyaHsgUra5AD63zM8QDbC
vAvVKNAFEwFWSWH5keKOYbh3DMWPJvLJ7g0IUzFrOAxtB65iJNz+sIuU5A/QEMPTHUwZVIa4yQdu
DCN8KeRgQQlUW6p9ChWHcFpb380oua8uBTB79hSPU6nTpxd3K80lNICsYaMUAO0WiCWudOMjDbE4
Vu0irrQrlkKJQgXNz4+A+G8d28dyHjUakSY7XWxxgtddXuSc1b2Sf4tpL83iQgwMNVrTLiDI3hfB
wqFQES+gWGC8KDyMN/+rrdCCXABjXZYimMK5RtvEKrxmR6UxwgOBRlxQxclgt9wK7s7R8hbuTQ6z
OtHUnwTsbttNoVlgunRYxdHp0OAdZJoohyDQNOBUaQvSz4Z1qsZPkubgFTei6MaxR+uixpAmjoDB
KoHeZdGYs3/R0NCZBK+uOIXj4JUL6bgbRMje3WtfNbYOXPTcQ4kjnJvCWxO6Ge4BCyFDHALmW1Jv
Q5QZ6ni4si+mSU9uKDl6GlelAkm7RWvA89tgkL+o6SSDfytNodWXf7TPhonS9HAEMooIW1qGPquN
D3LgejYAvOmNBI6OX5KiZa69OzqgEfL6d2SuVkbEY7RjqjlVRY9JuiTUHQRbMGa5lfeUn61H3BNq
89IJowPOwCxsuxlF89Y75dbx2yey7eCnsOB6TsOR5oxF0q6wxQ4Fy6XrlgqGH/CKFqJESDkEYMXh
NYlAVfkrPhHvL/rtXUgxxvMtQnUsTfVKJrfaKoFp8d/2kjS+/cu4qXnNbQ+5oF3Zft4tRvB+Q0jx
aPbCnlIw+XxP2xPrFVw1ekOzBNh+cwHXfk9xTHfTINtolHMn70LbzXHM9Zg155WCilunQaY392JO
1fy9GMy79NADCJOREBwUSTQMuiRucziZEwOr3RonodM7QpxJsx3QS0UhSpLdM2AK+smQDmfDfbKM
flxPHfRepOmXb0TSRo2jRJOpsh8gETPEFhI8fjG3efB+slkI658ikdrqb7ktCBssnQUwSR7wDJ7X
nGQrV/MbEyJD4w+PH0hYteDJaZysD1IrhfLHv2KZBiREqZna37qa25H+AenmNYnH4Pr6HmWAlE8f
NqygFCm6JYbzwD+wTQJzLYxK0u2DqR2rXoAN+28YLgDLJ4ka896leZMdk28jUijhWiro2gC6pJ+w
b06GIoScs7x3JriUXLwBE6yjdL/rtDNp/+aOSG09jTp3tr2A2KbNF350z7xJAqPs8ZKAAub0SMX6
Eyfx2Ik+a81SZTsTHmayc0HfbtBAiwdrYQJAo80hlMffGGrsXV2uDZYwyHleAMETEelMLOw+MTQl
zbGvNePbiiT1pVUtZiHO0YaZfFbkr+n9ea0zWfu6Jq9K9ytTxpdCTCXLFpdmxQRK5QYAXKNtNNpU
egJtM3DRFPPIWexxMUQRMUJJlPN5M9CostpdFGDUboRjyPTce0WCKo8ZVKFHOYFdAEG4ZInwGfW0
pZhaaVSYWMJbCAc0Rc7GK30XwMCoKuUFv49bixwyO09BTUwe5oap82zI08fhVHFLAr2gu66rwvQc
emM+ATMtk5g6y3itQRqBcbZNZ31Zqpq2P3G96ZAFFgf75ni1xmefFfmZxrj9+7MDd3ufZUVKRBhc
/AOxFn40Z+7xetvmN3PB9qCdwPUK1DWPn/T1ia5h/B/t4dLzZ3OTjwO9SrB1fkgTgPUkAVcg5Wb8
paDGFDZOXivxehPjACJSe8H35mvgUxakzx8lm2AF9rCY3s9ueO6aeEmHc8Af6I3jezwxZSfdV0D2
ZbuRrF0z4k6cb2w6I0+AC8P26zaSN+r6IJzkkZzVWyqwqUJf/6qz9a5gFU71R3oQthAhMNSuDO71
boQ1kjYr4n73c2AscmG4bIdFHryoakypw1txzOPNQPNrmZ3aN4q15SYlTb27jNXUw+de6mS5MwCm
y1DI7liaRMI/wP2XI05aIWaV6/NHNaXqD5OusdlqJ1CjJSKKG9Dhn9MPmcmUe5uctlbaNBF1BaDL
k37TdxHMWZ7W8YXBNdsK++Y+uz6GIxDRaaVnRkKcwaQDqEi6MJRbXRVOwD9V+E4h/903wF1hE8Wd
umAWF8lXekQoMVNVdnrDbwVmHlT7R+2gO8s8xvNwRIIfaOpPwgBvh2uKE3uymWrI/B3/jowlMFli
TZwbSSqtZEohgpyUst9ownjJ2MgdjwMgtz2gjvxNa6R24U2NjE4s6Ud39LP/jEU7rgAq+AAM3Ecl
luLTRAcsDD69tbKXYEMJuR6g8m5IQWCwIyb/E767lz/34xbQLCKf1J+ck0d9s7BF8rJ5n/M7nNQB
ZgU5o7jvEDP4/wG/BTtAyizVquoFC34x319dm1fEf+Dz4OmPrnp1Iy+FQuBtXin2odsh1nT+B/kF
E0jFNjOwmmIczmDJXFQh58/JfX2D5tQ47vOK9V/PqBUJ1O42hUzPt+/UUMkvQBtTfEYPBJ+F50Oi
NZ8Ls3F7dP3rBVDliedJHQLI5o29/grRkCdvLlr1B8wVHPS9E2/07K3VzPsqkUvhQGIPW5tJru5I
VzdD500BSDeMV9UeP3IpgN2K7+gKXh6GoJL9oN1FF3nE9h+D5hWgDEbeFONsfCPYftmObAL0jGX5
xJSJbh+ady2DZkZwoesZ+qyxJc6oqGSkyjNBQP1bvZLMzQ84a0euAq8f09Ah0fIMxfHLBKZ/61jJ
yMrwNefis0iOR6nHkNnnHVi49nwr1Wbww5KW9Q+yX3n1yl7+esl9MtXE1ozH4HLtLD/wYfwHZWdC
DtxY+u7sMHDH+3jRWSnJ7WQGiYDkg5zPZxLTZRHtl6yTMfaXj2cw5ljqddmvTKNEGEeuVvAMgSIh
ZwQFWCWw29hnE0T92U8igNvgzPOQJx0SLWofu/aZOt4vTirj/HZrmtf6s5VSF7qiWZ1NKg1JGeTv
ZlZWoyJULUGHI4oEazsxBSNbsfXCGgmoEK1rSkyhSw7f+MVov2JS7aXd/1SLTp/yuOVxpT55gDcA
mv2WXzMWvB8WDE+1ac9WRYUA/R9ecX830/08NMbVZg/q/HCwBj53/5rIr1MqblZQqrg5rut07THx
HXILEhCRj3ZEChfERlV+XNRCHlg5hW7/lozrIiniHmke59UA3vQqfnrlmO+st+z+/bMmqLwMDxAe
kBoVw2F3nWVsuHiOgNICnxZk7tHaB4s++szShvt1U6RdLkPqopeJnzMGoUY9dnHbMahXXmy7n8a4
IgqV+T0uzHm9PR7LasqQ8K83Oe9CZUY8L+6acLxsKkDuSS15qzhJIpij6vAnSkulDwsT3fnyqp2V
LnqVyVlZwgFFh+vrUM6mCbAovKn09Sd1iRxGKzJ0dMuwitWi2VfJPBItEChm3KVO904CtZ2hsYYg
m3k9rqM1QVfkhIwefxCj+V0dbasNV7Mn1bNHDoVMjl5ofOohbewcEnqRkcmzOMhiCgeBJouiDisN
csCkK0g8mWgaCUMomIlpTDuGLrifLMTxSiG/wxa/0XFLFWXJunqV+7paZ5es8s4VEzZYamA3uLIP
x9IDwPGCF8JD/Pf6eQ7Pl0bTpQs1LKX0XFdKrHXp8CwP7GEp/pJOodu2dSv9iiAcRJtnT5xMNrtJ
3kgqwEnlJo4UGNXNWohgVOEgI5ZE8Z/x3ZfGSF35bkeiiO9wrEvSm48Y02NoJkiQRqRXhmaF1RcK
xITCRgBvE0d2ZVxE8vop8P5s4abqQ91p4bMyHZHFOavFjJ8i5onbCOzRssYwsxvM0CJX/ZITClHL
Sca3GbRt2ojEydFT+LDd6ldmlhS6i4s0a9W+x7CSBs2wbYJJuoaGuq7N2wunMknoZKLPA/DennIO
sP1izX1tNlQbw8X5cC4xRz16Tsw5wPyNTYGv4vPschpzBBucvlvjSwqMxvqqLJTK/pqlM1sf+5Qs
fk4fXQWffrV3rL+F+2B5I6OXCxfKNvpLqAXKMO9pXlO5FrhgXTfsZjAnNWAeH1VzXBExYbvWObmx
ej/F2tPZrVlaZbqzNkaAKli25Y+hUctw2YdPQ4PbURR7YVpBMKwLWD8dmLqxQeVr01eln+l6CIyO
OL/QVMQwi1i9JZL7sGGM3QzLsVaGM9hT//Db2KmaCQ4P/U2aabMu5ySgWllnv1xy6EOgkmKZ455+
apaAzpPUirXIQp9oZSv2LVTsYOgsLUrLQ0G6IhUfMjBs8sgbt+3cuTimRHkZCsSyO/u3q492LRml
ohaS+nZF04+aLZCc2p4mD+jxEURsvK46xXiGT3k9yEb0lBYfl54v544e5PD4kZePzLgTUIS3j0zs
5SUOWuXhYJv7+/Fpth3HAF0g5jt69gJ210cCkCzwn+1W9F6gqP5Ms0hIhw/bX0Iy/NQBy4/67sZO
vV82n5cCqz3Gv7s87QwGItyDFm/xEPHXXqpYvXp1ddqRgL1M5+5dedBweQyDZeUIIFiu0tmUIhdE
2ngUp/5cXyhUNwMKAV+2Qpjc7HfhYDgMJk9H2Yv8vNGdmo4euNelDK75t2wElbOYL3sGi9wvAz11
XT6QYoMY2XD/DsHIO/Se4geGYe4PzrvHU33IqSYF6dPXAtOT1ak/3OX6UR1JDhnVRBdcGG8IYSsS
I64GtxgthZIM4mNU4G0st1ZzheAzkrwqYh90rEvl3wzrBWPIuEM/VLR1WXhnp7SxE9lblYeGG5Zm
Y78JC+rm+wWAK9q9fSOqpg9IMWogItq2gPv4Ru3M/OmRXeq5RIwVyWaQ5i7LHAdhxFJZ6etXGlA8
4Q5S0NTX5qbT9baIMtd4eO66AkN60agUybq4tZ/W+0TYCeYqczMYYql2KpgAnmSbLEx/Rb9Yi8cG
MaJ633kJPWI0Sw3uXKCAlemvDcG8Pr8RIEmEeCxtIvbL6t+OFxKB54R+1HRfRKSGteoyi91op0Ue
Keo738zePqeyinVW1i91zb/5ug+z4pQnoSdPXsZATyyfEDBDffOgNm49pCVA4DmmfDOjyNxKqxE2
xq+qLdD/cv9HoY9H5rd6xnCUijodfwIUkNKS02pGPiCzOL1Rycx3Q061b5wZDXB2PE9jm7//9uh9
/PK7v7VxXyYG72o4WQfHI/qh2iX3aPT/fGJt0gRAehD6AeMXun/bm5y8huDKaSABdYE2KOrPJJ92
DhdCd0Zl/phbCm+1n7ABpZVFxY2/DYGVj7kNXWHx6Y12Obctg3YzDzyIbF5pKylGzK5kRO+FCy4V
BHg22eh3TRMATJM2XZwPNhYEyfh0+lxrz5vbsmhMSB6Lac62Hv3oqFaLkTGfhszDOaiqCswMXCNp
2skt7fN5tqKfTr+l97U10wDB8/psSMjrCc/NiygGtMJ7lsxDC09YoqVNa9cnFsXrDOpI8QSAQqcK
3VooBtXy0oRdxGtvHc6+hK/0hOapr+J1Qi5gvV50uqAhp2du7DXnn3Yu1ubawyJdqBKkSBYbZU+L
O/Fqkf8XKI5IdNjXpReC9dEtEb+a3UnEBzw209wI9/AFYWs2Ny6MRNUgHagm46YoWfc4zuaR/C8r
4TU506VxDzCfol+Fl4yH0Qh4z/+1l3JR6Y2a51jkS3wKGQevNYTqBNzLNQ6cOA6a4z5f1uFapAHH
6N4qaEGAsyly7GvpT6r9cMV5q9kmfbvYOKTM8Qon8IBuENttizUEaTs34tqiymaOME2hHY292vuW
REFuZmDMj2x/yfyIQM9ZAApxaOw0r5vC+wlUZOQ+fAHtZ1cUaH24UId31lJoAwnga3FoROqNSd5c
EFAoOBJdLkmpuBnhFuNZ2nC+2+LDglRjjaeG2X7iAcHIMmDW1G/GTQueCDbYVWA8http51dj5Qb3
L+w55dqqMxdzJWPq9jk6u/PIDrp/trh+l92dcxLakCz3bd4ojTVVpT3skm3kUxhFK/PBgVCZZ4+/
KFeZfdcAIWi64HhErAdylnXqFm7n3R9w/LAOvHMktilH6Q5ApNHkHxKcM84lPS6h9B/x8COsPoQ9
Sl8AIoPNzJUFkWrgJjSsiv6dLKf7HNG+Bl1Jrxd+hsmSAa71l7UjlReNgELUXQ29OhjljE4Qx69h
K1qeu+b6i1zZvt8/LHPT799kN/QzVYVSkC1tm6jh3NO8ybsM6YwDADpsPM2NQCut/193M78YM2TD
eN4KHTusOH7f3TZI/uGpMOw+Zl48xifPl8IhAKWLeKUrn0EZlUPK3AEd+T9OJZyYuiG8m7s9RxCG
yAkTToQkV29L4Tg2U7kvyGxdTHj4ZZdAodR+35gMejpIVgOTrFMc8lnoiXZgGzvd27de8HOBuSwz
PJnIT6kJ+x83ASGZrbT5LWPp4Bbyvk5eGRrEn8USgW9LFn53iUYPcObHjiwYLNYTsxYyOeYXteDL
43JZoWkD41sZSEDO1MwqSfV459TCnEQAuBYBvc3+DZIiQkS7nK1gQOWCGVCsu2+MwUIOpfnaygkF
p56kP310glTDbHSXjJyKwHXVlVBKRruky80z5lZ6dowU0G/oHA6mrmhdv+EMiWkeEdIUQg1o6yJl
G8CAUP4UFlD7DvAwNeIS6rUSLAomOeAZ7VOClilL1z93VzYmNv9neTF4YePxttDhq1OpJXlcLQYg
HZstqp2YwXCK6QgzFIBLCEL0koX/hCQgUuhHBB16NWuG7VROoAeD7UNzhTgtY8fagx7nzB1iaFPm
VGwm8moGDmV8TSkYXl1RgN4Fp/VfQtvr/dIWxepDOzcizjENfkjt3jMPBzEv0FsDzcWFt/PCTR/G
4wNdj9qngt/QwkmrbH5wDhGr0HjeEuhe7ZEZIV/3J46WRdwH7P+43vGDt3QT5feKFF/U1Zh0pJjQ
qJradxcePIAnpBPEJbjY4pAK4eWBTOvsxOcibuKaOXGha9LJq3Y3F0WtuyzbCxhEcv01YyEc9tDt
KoluY+RjjozaWH+cm6ZYxWOBTOPS0WCYFC+fGNeBhq63gzwEzuM2LRZX4TKQv+tP/CeBiQNQ+T7o
YNyTOh+kb4QMASztieY6Fl4QJlHlRhgum2dGhVzSdY9CoimJsgYxTEOIWZAuPB4ah9O9uozgd1qe
uoS2ZGJTqkGYC5VwDNcOoX77eQUHbw+s1XmdmHaDeyD3GfYRkE1aZLML2CKKJAXcmn3BDtZJ6STx
YLVCB0/DpXHjj1Dla69WrO6MsFY+9JdEwRPLFCTagI7HZWJz22xVgGRFJ/Z3aZwFqQWZihNb+afY
D73jZYihBo2UPav5F32WjDnKUbD5P+5fwl7w11B6i5XJdUWfGs3dWzVX8wmouZTU3fszdqq7bWMG
YERbDlc0BHAMpG/bbiWSnBsP9VvkwDrjFthh44OVM5WbRGypRSvzzGugr2D6CKcS2bGbVb/2ckBo
HxqaKgb1JWzVRUDE/LK+StBCU2mp0AXNePAsGuXAt0jNaCwWlPhagoL1dAUpfOMdVZ1gaQOek204
BnK87C1Qu3S0FkJbHzcV40s+d2EV/og0gYeRupgBT+zgrltSdmTgvWDHu6VQcBguzZ7jK+aA5Lg3
EoGk/Pck50so2QFYk/r+OXpzVz4can3cwjFZAhH/n7maWXpH7GYFrqKXelyNfGvNdVKZDC9Ubrel
Jdl52ZXDXrX8a2zE/E/QVBu19kvboF/787beXXxD3EKTNhgEfl1KSwyS2IQ6k6TNTWMU2s+hNkYW
7sUPtiuNt6VN246yipyXMm1kazzIqP3kbGzG7dlPSYEbocE8l3EbAnWJ4SAzQSXLgaaxFp04JEZr
9/tlXnjSp7hSl5hB3h9ErhG7cpnqPDU+aEZjSJTh+uNlwXbdQdmFFhAE6exav3OkSGoqUCmwWryY
F/58Klo9JT7reICy5XJtjl38vt/vVeLWYvp+VuuRxlHcQHGbSqCzihtwz/vCCI+nVYf74+wmL8YD
dlGcC/tNHLTGt0NFSZd4bJEt131xwGshDa6fkSKzGM8r3r+1E6ykex195+36i72wRtcQ6Ox5GboE
2R2kfXniMn31nYST+CeWQBS39H/yvkjYaeEED6FNBbSN5b2Ae8MO5MaKOaQ/jvvu09UsEGTYPg9A
WJJf7jRka6Kx41Qvgvto+DIS9RmYFOanfCtu87j10M6QjqFYXV0vHHAx5p5O3mlxcmoE5OqQtFye
iijWqEaZB+AoLBktlOpz+7YmFID2UD+QYNaLCvADTT+0K+Fk3mFzHvso4JZ3cSmPy3ajUkioAPEf
H6TkczeZjhfcpdXEU4pGMWGvzHVQlAEEMAzivVrqdUY7n/z8LVREt5DBJDJYiWqgFDSTh0PXPNtW
+pXVSP1VQKMebJSdsyj8NcVUZ3joeCwedbrexYjzb9+RpQP7iqzOzeNHNH+Pi7GvAP53rupMsZIs
AAY6hSu/zocb2bLYRPdZLTNDViSNAQV40P6DNQ3ZQR09+bNb7byI9eSlE13Kv+s0bKQyaWE0sBBb
9Z0Gwp0hJGwFKWJCstyF0UUusS6K3OQdF7mZ2Y+fZR/jFQXNx7Wrheky4SCaR3ocgLfQOGkf2Fp/
a2XJtlavEfZHDuQ8pDgRik29Lv7UgaB5c9lnCkjQggvilCNfCxN/B2Lb3wNREniBi4P8hwe4Xexx
Jz7rGOUBzT/aHfUKMevpsz9Fnx/mZITOkSKHAj+L6Pecagi7Jm1kYvKo0ivQKgNzcJS9CaEQIKD/
/nibef41/bJV3ntp6OBH/eN1I7pK8o2Nn1Qffptf5zANyWPpHE5d3GH1AGTVVBCeOoqIx6LpIP9x
V5GDqb7YqzYHzi3DFiUX+pML8oVkCTVDB7u9OBRj0el3CIpMeYq8nUqWhEuLh5Nj+yBF4L967pMc
oHYPtv/rxwe8hepfsN+w/LUMzs4LRmxjqYdxn7foCUKRkJyVBPk5omX9HTIxB7KPz+Fvs8W1MylF
nSagJndJBbzkGMi/ODtpZ2XQttBK3E3GTuPfw5wg4vocVKEWmgjUB8J3dhpigRLc9kw6Q8yMigIe
LtY4ToC6p7aukWqRXJDZP/vO6qYeQcJnLzpCxjDaDTvcwCaH0elfU4T8k6cTFSl5vKhuyZRBy550
7bYn+vgXRz0UfzxZEf0YVfCw8RKtA6UZC1S7ZSv3afuulCtaMey8kTD2aKZn6xLcnIyzk64a/r03
wWgGyQqo2vvqhyaDEfT1kjC+QDA9pkCuTsJBWFHCfb6T6s7nl6xDX6ajQ1PXtZzzuH674fQ5vMI5
oYocq6I7jgzQc1eIceUG7rA9ViRB+ajUywSXajju/HE/8yRVE+ihX+LF36kGyvkschqPI8mMucU8
vT5LCY6sAMDFVjiyFqMfmAsAasGzRS2b2gNjYj+PD+GIknqP0KdXh3mSlZdFmhYalaiXft5hpymV
dvI8tiHJCYd9r5uHGY1rZaus6TPNwyhpZ5YGeYXk7h5a5XCx+WtjbhsVfdduzTEL1J9PZCcIbKHH
c0+R7Gsk6QJ1JAATHRUDdmAUIuVIX4qDnMjPNudKIyY4pEP4ExzaL+aj2Wz35KfKyOUdkG2HumtA
V09oSk7jKd7kPhFCEyyOTy5ah710WSWqgkBmQDcD5VuJPG1B4KPVAiYZ6Sajgln1aEja+nW3XaMs
uEo6BZR9rt1PI7EiM8YQfmmD8+0mFRF7DHr0eOkAlVf0DZhphnWafhJxDrFsTsfAyBPhdyZiG+u8
ossL5R3nAZnvruBjli4Bz2V5tqe/WORrmVhx06pZPfuy1JZWqeiFTZKsgLKaPnQhXvhju+Tw2jjN
oWXETAmCNsm+MrWw+4hIOaWZURQTCFQz0a4nU0ynfdshse0n/IAxox0Yl/U4gAEHHjoK7NVO9LQv
kY7Zojbd2BfsAiIvkVcxFYastfHzK9TEow18VXlreJKOJAnDHrh2lIY3hpwYn4Amn+Lm4z/iCL7J
xwl0KdTRrjwY0WLcnhVZQb0j/HkS1rr/yyoPRepQOJ50c7WQa8Bue8hwx/QfHVMDNGDvMXponQKE
ILtFVl59ve2yU8JBsyNihqgYzARYGSKb2tC2N/aOSb0qsOOGNdcK2QjaFeA4pgsCjjGyY0zEoGYi
Z2mILCu9WznLhLsMPVPpJr28dzDkERQSzpOFK/yJpXQKpg6L1wsBTcXVDMouLKTg+t0quDfP+bzH
H/lkTi7g/2g2Lv0ahfrLYO8ir7p/9LLU2xNkOVJb/X07Fzs1mBfsg1xpb8vgkDM4UGdJDFebbXBQ
ZpVNa2/ViGGEJQ3EOIamuSpQaeFXCmt2oZLiTnLghNR9Pnkdzv8II3loisbYQg9uh+/k8+Fpf1vc
RpnvnLAx8SN1ElmTOZ6v+GlXA5Pg7Xp4irbRB6Ldrc93VWBM6mUgnk5Z+QyCgqmAo1N31hgKGd5m
1TANHFaYCL3dZfZmTXT9X7d8qLhSkAqVmCUNANEgA1dPxwEP1Y1XRM+R+4GqEroj4HKxQieFAx3X
H1guH6+dvIttJYF9Qpor5WI70ox+gLJ0azvq3CTQrIPXOz0oKYgUsFoL5CJu99FpJrNEy/XpeF1p
WqKaU9MRfbqcd/NursllbaGGBRsJIox7TnhgF6aAd1TC7DPPSfLStxLU8i2BA22bjegmss9VJDt5
ilN3xzUKSSMfRTL/IVAclFt5gnFoFAoy+/6rxTP6FWmwov87FR+YAtsrl9XrVsU0617i2bsdlC84
pJkB9jQOFjg9PiURPVIo6j0wShESn/+vGedBgHjflBh0qorN3hF7P9LvOgXMCF7SldkwK9oLF8sP
EUUDAlGwRi32prgqLvcHVGfRFe7Rq2F5FuRVPuAsdaisiEIk+C8RGS8CdR8gMuz2a0gesPSxVkKM
HDzJpQ+5xL31qDWRuyEATTMaDSGCZ0M1Ats7gRp6aisVaaIXlh5hRlS/ZlXRJ2AiDSupf+db0s5V
bk2VunW1bEeWv5WBvWs8sMZ9+vruFQlyxoQuEyuP3VKEAIioAXJD4ip2MiiZnW0LPdKZmWvFe6z9
cOBjULsWbZ0nQtG/9mAm1mplPs8kXoS4t25qx66ZN/57MHtLlziku6PDQNCO7BdGgzcGRc8m5lRd
N6Y+oGJOJXIxGNTdoJmraGl8d0iolNWwFQdNtwk61e4kNJv9sIhvEDvW8VL9D3/ofCVZ0lMKMTGh
oEegE+7eKBufGq+UEIXGw9BCJeZ5SBN+uZVcSI/SFOORMt2NETkuFhe6f0mzYwSFixkVbTefBdOh
4WdL/QXtGc4FEZBJ86YRJCgVTG0KH+TKswax5p0HVasWxMOcSdEs6yqsj2kLgFTEPKrdWhXsFR5J
pDSa6BbrEByb2qzLILXMxDPoyzUgvXxPpfVoY5qffniHuR56uI99GvPqOSKoQ8kjtREcUNEcWxIV
nA37/UGMbxOvJL6t2Ztnb7gKB3HUnjbxO/AtWMQDzMGjEFbCdTODv6urHKJE5Clj6NL1+gQKKBk1
hJsTpnItq7UFCvkWiphClgJ4Q7JwJrGBHkvpBI9NcCD0e9yc7IbTgRTTipzg5ouuTvGkfyA0EF1L
WlRc5DThUZ8UUSlxXpzgTcyr3+ECECWWMlPQnvE11E6IcPrWJbJq+vbEbuJ7IP9lWxqnSUqJmGxV
6gy5T/60MWUmjskCd5reTcrgTsCoaikBfRxtrXEjcHgEI5taVS1GFz0A7Xm3/em5ear3e93eXUFs
80av8EYdcZfUBt1D52CRmigNAXtNFjwruHTx3zToVoEVIO2R6XC2IDFRfV61FH23PcSCxJ+j+w+U
4JigMDOou2TPg5oQcNPtJGU+4A2p4ENcO6Hp/8ojS0TgXem9vmWPVPlk0O/x3lyzje2/WDQEwKuP
oUNRdx1JVzagRIYatTBmvDAPUO4agL3Ncsd+PSOdl39Wn9AgAroi7f/GSlID/wXyQhO4kJ8dsAZl
eMp4h9p98tpzVD2fwk7ENlSjT3wgWkhUFVO6zTC2YzLD1bBUPw+7wPQz/PUKMO1EBpTnHXRiIyQf
I/ck64fWCz88HflsUHs3EDDsWXDpvLmuFcgccfM5YOUtHe879lOUyc2JXAeU6IZQrWT/4fBI0q6J
MP/ppe6ktYcM74hF44uMdue4kpuq3NZGpUw+c/uMAzM/f3F5bAy6g8AEXp6iwMYpV9vIb7F5PZGX
XWtNFFjnZqM/RYljqWDd7k7Mr9y6zFZJS5RX0KV88jo0/UfFGghnOfiTCXOgQzIJGa12Dk4en/oN
SIdUatw87DJy7Va1t59LA4KCRj2sPc/Hy63M4wLit4WKEvLCmplPuvrxMRygRyMyrL18oEa3di8D
7hzw3NkiIokyIFePox2H2K9Wm7g9YZI1dnRxHwTwIvfH4q4nQd+hN7Qho08XAnpo+tarKsWKJWyp
A525yubL0108ZixGbeB+kkrCijKjQ+agLkhHFdCz6pFGG34mQkEaoOEvABOVwsFJk5Q6FgCkzrwq
X17vwAHDq8cHVloYKF0BpXEkZVkYMEdJtwM3zjtPn3R+fwFm4pYF1eWTkUiBDVRfwPLvetUuNorJ
hSiGYjiHb428SDLhDACx7g1FJgoFbyP2D8TKWuHIQr0+nzcOWmj2itSbN/W1wQUd18emB+wQ9L5E
XsB3Y79MmmjzCIgWuQcL0+9t9dV2a73Mo3sJFHHp1DHq9DqSNpSAYNCIm1L5dIQg1qSQipCRPziU
UaL9M+jYxuZSye97B+feSemg7o8IcBrkhqVwo78wot8JltKamBTLI9Mtn2CcKQDadAObfl99QEkz
/6iWD8cmg1Mb402vMECRPLilGt9PaRdEKBr9X3i4wunJu+miN+dykJPYZ8zgBMz82vIXTTSZlbHo
ZVThxpAGytcm3SGw5tX7+f9Ga8A09uRmZnPayVhQArOPLY5wVHtJRRiHo2Xc4y5PtmaQhzv11Eh0
3NCtt7JPSeqpHdv0B1kKGeHrJ/yxTOWIWsX0w4XblESY1yddE0AXZy2oCjsr6jl5sUQP2DwuKMHo
1dEWg/PODZPcuI+AudH0MAsFR8sUqflhaqIY04QQH3ZDPB3pKdmTdHaqudSoPXmg1Y0wcsdcQj19
MYZSqA6sDnvbpW0XNHzRxxyEcCZ3oR1H851hgJx3XJWTuBxCHcMZ6H6dKQhbRwn3ywYvTCuL2SRh
/+wGJ6+trQMQOCEOGaaxVCnSXeH94a41xko+QBrsykZbpqR6J1unkIMaBxsljV/RLZ0Hxuoc4K3W
0mTY9172QlKE83WE17W9QKcxj6fEICp1V81aQ++ybkER5ti+Y14U7+2454in3mjVcLZBn9FvLw+d
XqNSWcOSgaGqITa+j6pQon/1NRH7R4WFYFZ3KjcWLvgAKMChffNiaERG7HodV6ifPaQcGsB3teQE
hwO3AeY9dagBFI0v6Fc//jULOPXxugk6D9i2EfOf23rYJxhplw3cPYuk1tCZZjfupN3GhGBzYitO
i5yXaC0CMxwqBf7qgefNpizR+H+ZWNcTBuASnEuRR5hWIMHHrqMybsCzzPrNJg8znxicq5w7OFXK
3hZEBIoGwuM0SQ1QpGXufpMBmy6BPnVRvpdr+xQuYGRL/JfGhOY8B0JP5gJpM5zNRP9VYGGO9MfJ
RtKpEBkLTwdCn7cjSlfe85KTkYWrZyy6oOQD4zk4W1Ni+OzQ1RD667xLqM5Ihd5fHuPUUXubGx5b
qDxWS50lLrKtO6JhaFHz+ngJMb6OgTeNLEH3/FeQHPwzBzgwgS21jr9wB0vBTf08hS1+rxdI3ZhY
gEcHhagFu99SdkAeibNXciC9sM6CVrSRhHzfQRA8rQ6ZjJvMb+qrKC4XtG5CquM7KzZOFiqegP4J
gLW83OuCYZpAMyz7j3+jF8TNqyzJxiQ7D2aqz9mE4NEBPl2ahpi1Oaf38GQkky9RA1eIlFtu7ylx
Kqy0JxCdd5BeHZCFzsHLy92f8AcO2Pjpq9/DBIkPzVzmCvyoQ618WDxs22ELO+l+WGAYrZL4NUMM
b0utPdJOaJ2Vw8aJmG8xccPFWcyKxi0szH7U9IlnTLQUUrxJG/FqG9XuwW5PSCa70pBUftxjlbOM
Wk975+Oe4BMltAjfVgfhp5baXJHSR5fOscrcwUIUm3uVqT3se4wCZQ19Yh2utbuIZiOWAIoEw2yy
IprWoN/Q29TH1texsZElR5/ze/gm9Sz8mYqn59nGb8BXSuoLJHlTC/enAWpqlmKhNU9wfjaSmz+p
Z3pYBHDehHpRNAOAQoLwNQ7dIExYYbJpgd/tycTyK75wjyQ74aBt8onFWZMg6mLvcsPdj5dJK7Si
SH7IrMQNvGSXFdf32CPpx+vdnExOMWRAZhldVSisb8d2+LigqvdeunvHqxGwnTzsgOoGc01weFfG
rBuLstBDVLzrTm+zSW5/RSC8p8a4vSMs4NXpTCgSZn/LWHawCxXuvK/sJs/vYV3D2U90k//vqX88
kV5y9XyukwsSOG6TLw0K6xqwdCFrUyDnmJcD6xFBM/Xvbm7tmTAqel0/b44w72Rgm29cG7w5P7yL
EWA00OlMZt36oyQJ4WMy3goMzLd0SIeD5wD9ufo4Pds9DXw89VF8gBiMbxqJAUALb7oxp0pXCHrK
sUq6Pum1N7HcrpqYX1v6e1a9kgfNVylYdrRzO3I0wgrvfc4RJJRPHoBiSK7R54VcEmcTdRfKHXPf
hQQ0tO6G1A3sFzhHGV25A5TAPczSD+86ZfJIn+mSZPojV9k2i2+GXYhfnxON+zupVlVsHrU2ywmj
zHLRgMpq5xp6oFf+zN1Tfv6UmyZgPt6+AhmdE81+4srb7FHVCdNZmAWWDfv3DvuDTUZXgf2ZxvXR
XJoi7pil+uQNTrlqVXCtkjhzzOghsRR9gtVr0feNmm1O5rlc/dv0mS8M0+x2WsVu5clYwndq5Lbo
uJSaBbBUlgIMT8rjSgh+qeXMM2tXpl1LvnqAVOaLw5Q3B35mUNAc8owW041NV5yl2RYN33dbB9H7
7MuTjfF13A5QEMAUwdcgU6vXI0p3ex/n6xFokrZPWj1iHqLNo2j5n5BhPcDqBMKLi4YLZOJMuMoA
0y3dVuLw332SvHHLuzYztAiI9Hwz/0h9sMSoFKo51noSbd0alVj3/dt6kt+v/GGj1KCE4EBLd2dm
ySeTuHrqlFjlv3ZBNyM5Ur3f4sXyFicJdxhUYBBxYUpCdQOFRMoW6psIzlYYH81fyhpiLhP1JtsI
6h4ksUtFmCcT9/zuB+ktMulisn4+/vnCIjYAYcIqzr+0uRXXJhJN6wzhO89XWozFrgwFalCcgOl2
zKDx5QvuGbm2ehJ46Wdkr6rqXj/GMd6mGonbkTQAGxLu54Gq+B9vqLaeMY0tBP/nGjqpovwrXnKH
y3D6rL7H9ypIU/0d1ZcVFhzOvVWYH3buwacu6Ef7ElSXn4o+uUpA7bS5LIhp7MO9qPP4gmjBcVu8
raDZHVCoMdD7WVWisto2ap4EVI/2bGADfaC9CHe1lq5+t35xeX8R6MMqDSCso5OLhJ2CPuOmV1IF
EZW6qpy2RTV/JjJbW/DQtVuGIN/eyShdIKOyNl+Fj/tkKpcOPJqNbSiuuhRy4m6b/zt76e7UQCCa
N2YUbBFyL/vmN90t74+6P8pwrcCg5lct+h/0MB2o9MRE4KTUTLuYV3/FhuD+WD4K1eQW0/5lAF1e
LrSl6UMUpX8PA3yzlF0yzbFVVsF5inRrMh1rhQaeFlxkwye8Ess1dknp4VSdFJIVHR7Jg8jjRJ0P
f+rp82+HaCFgbcOHa2mABSj5tZCt4Hg/Dijw9vvyypXhtAef3tx3vkU9xt4X8uIuyjjiFPlHVS+W
Ie/qwJlR5x8B9dSKWsHAtqxls/4IhkuqhuwvcZCB8WQaVwNAjfaNJhaFPZOTOXLM97jhaE/qgbTm
hnijbjKF3LmonwlXhnc1vhRxhhmBQQqnpt7MO5RGkXFMAcDnlqb9OUB91NEKst0cPCovibwrnT8k
ZDxACvisz/SnW+oM77bzorrzsedFvjU1SyznO6tIhvJ+Nn6N78+LdNF1itiHnFFTVOCjz/RvpOVX
b5G8jF3w7TGzvr2/I8Ni4FjIjeZ6FZaHBKwSkeXMfEzZ2hCEouX1b1PtrvSoMczBZxqZueS4/4Lf
5QXFVLzFVkb+Io6lKFFrWx3jtraeW37IE0QYjofw0NNxIbadTV7J5556cvUwdfkzHT6GvtFy7smA
Yon0oYctlCGoVgTwUZaVYysaNwT4QEmXDB5RU1CpnwcYsuH5DMse/MvBGH1zVDqsGdD/T+zroLVQ
yPwVUwLoRpu5aItHT1ghALtR731sThYc9gyUMQwpg2BAzSmtnwBHOPaaOxBAzQF2cfUcIBpqb13T
obPAZmHeuR28yWTDh74sKmeEdld+Mx+NzamT8lpTjzqMqeY2KfOwC4d0Hp2XZoxuG6uHPB00Mwna
FaJyq8KjHnY+li7MB2KFkHnKtKvywmxLe9v0TBeiHtl9eYvRGxSzGFMEMjZy4ntyMBJ8gDzn1j7t
qmr2UCVaZC6AcaMOuNXlL3yHZpoSYhXTCpETDuUhE4pjnH+/BRMMePnERfG8A+/1qbcQie+xwJj8
MSf1opI0OemiM8WUCqPC509hDJJHSc5M2hnqBszEtBFpnBxR9YuDZ86Q2WpF1mN8GrhU8KSBizcy
nQJ0IfBP6b82Bmkr1yOMd3PvS9yc/mvnlpPtBfzppMftIto5FI2jTpzGglN4ShGxQ6mGlctihbJh
CsFVMRa1gQJUzXMoE5t5K6hBKNpFtwntBQQoFIW22Rf1qgF5vCbxFodP44KylaNERPZwlmI9Ec5h
GX168zIQtZebSwkeZJTNOekfv/rmOhkpzk+aSr4iVgq5SGx9rV7jehwbzYBfAbb6DTupLfmVkpfC
MLny4EG9YvuhyCQmmaKpjYd8t9Ypd4wWjKGVS1cCWkE7sT5WsopXxjL/u2mkTORdJ3kA/ZEVbIDC
h6dzbnYGr7PCJ3P1T9FHQvWCQkXVMDMrUreYM6KulirBIHJwUOIHwql1GDBQizEJzWSwf1vh4L8v
mjJriqRT6XRucU1MiZfE4zDNWqeA0dnW5XiTEPXe43DEQVmj+GXOFp5QZB8isq4ASLgHPwQfk+On
tlo4GJ6jELI0MIGQgPexZimrPXUpHDaGJmfc014XFCDlbMXUCApwKeEJOeGa9Xt+qiwRJeS8DM/C
k51Sn5SMz1kPtoG49xk0inDDdVTg1k8j+jRjC7GNpavO3NJrYnE0us2q4jQpZVU42C4ojfntUxae
SbPv02CrIlNU2c+J4PfWN0wv4vou9llMBOXy2ZNox79yYn7omahqNy5Os1lxcI6Q1G161/zDW2+m
NRApKCHl9ueDXdGMXEzMAbK061IZnkRpkOBLbu4lIwWU515WwgsgmDnrX8JmFd/PvEHyh15QKt0j
V9x8DRMs0h7B79dTqJZCkAtqLXuMaFK62LKLXwN77n0SOLfwixZ5gyj9h3Tz81SqNXED0O7Ms/yl
9TTb6dv5Vnb/itr00xVRTLw1V9+wsgKhFIYftZRVRTWFndG13ocRWbuCKjn0Ofd8buFPY0bLAxQt
eLufBAmoncjKGTpeCM3OAXrDQsRRo3IjMCaBsDP1Cq7oF33qAar7UUOnO15i0hXxQcKvZvcA6Cty
N6ajcrQMlKzSyhmd1P9/hYRVBMxwlEuNYV2DkEQOqbjERTs3n3CUSt3UadBvuOIqXJx5zg5mjwri
pvBRpxffa8Ywms6+UdgNTLrrED9TvaghpbwRXPiJhkIpzUYrMA5+k8MtAW3hKsP/gyiZJ16D8f93
BQwjNgiXaFbIc0YhfZZ/QoyRQAS5VVRWT/Jo1Nk96gAVAjJCaPM/iP6TZVT6Y0hcaZq0DBP0zt6N
I/7bmAi0Qe8ig3gNYRHGKfT/q9XJaJRUVn61D6EkayYLUtNEtU5d0/I7Z8/32wP0/fEDVtcZWnoY
JGVBUSgxz04KCj4S0jVFBCUx3W1zW8Cgso8khccdfKeZKA+qKdA26pR97E9f7j4ms9Sq+MhF4BVx
vMkNvDzdpxCu0jd/AKBiOK60C45VAAfL7hDl5JaJ6LmIxE3LhTY7alK8cbnWq7Ul6FBT0x/iegDa
2iQx2GkOzDVDCM+caFuTKQADq1Lzts5EqqsrnpcxoFK4/Zd9iJfe1E1Fxrum0Tuv5gp60wfVDzLL
cnuqi7QULCvxCQb0PKkzX/eIqKWAwsUOlhXYWtPtz6xoYy9P0wGHlCfgqmjf4LzkMMVTb1oPXzgL
jNVgLqk7lpyBGYwOK4Feiq7/+d1B5j1gUmzcNmINklNlDYmCpWNYzMDdZ0L/gs3rv/f6ckn/R2L7
lHhrTUWyVrNkMyomuLu8nK8cX8bqUNhR1wyjvXUhKpHbbQBX3nf4104GehsK1ucALqSSAgFjV/yy
UhCglJVm/pjGkMWSnj1oWSx6HDPwCfBIYCJnReWC7IpPn5dTVFBLZ2QLqAp4iOpWfprfo4bk//1k
UutTyNpud4E7dlgUxjuTFdlFCojKVQgpyTJkxV9N+If/aZtXicNkiW0LLvZYcsJWgWHHKXqKgvh6
cZq/oZ65RshH+pHnB5OPgi2my6NKYvWzVauVSFZbwCYsu7sJAnRLnUeGry8rsOd50JB77L672CBG
OyUm1C1GFeXmuvghou1Iwcaxon70Sy9/6jAXQc5cM5lddJxFoK0rH+zc5lC8RxnbiRkB3zObzRPA
Uhpp/GLaGzxbV+rL7WfXEf7NqP4ZLHxc4eRcTE4m6RmchV4PrX0El/9xCMb1Qu9K9gHL7y+RBq1Q
m8iXeLklcdPxCAM7UXRhPTwolyjTDnChIg+Ls+viXomGfRjzt5egirPSwz6R9DM4GbUwksgyxxFn
nuPncPNMM/U6Ojqwakzt+XTMVCyh1IdfX8NVxqSZnxeQjzWG4ae2G9uDjiyq3wN/rp3CuqsyoVnb
YOBOT7zGsQkv0Tq9qKNqMxbM6p2NfcLPUGQGCTwvi2h5fMEe8PppFbyxNoomt9uo7njwdUktWSIQ
+oaaGbQZkHc1+ppCEg1Q/4YaeR39KkjW2o0WwTf0O9TRIqN1xd3DZkqkzMZk3fHUJO8zIo8NSeWu
06hAyCN5SQTw57f/FQEm6plgZkquYgW3NoWocqdpQI7yKTjmxysZykgAQ2Plfo+idNBi24qBXddr
U5hd90JTqe6WsaKY+9s0UJBYRNNaWUw4ewnmzlyT236iwWv57W+74HvsQC5xPPpfyhTVc6xfRfUy
PPCzxQv9k/ggxDeFpPOCyeizcJ5GdQ9ZHiUTD7mdy1E74wE9hf2zFA5MiO9NFGikpM31orrZJtUk
hQvhexS0rNBWSOyInZJ5NkdRUi7NqIDrc5bmRzaG7r/YCfY/KV1p4A3F8EKLqK1svwzA3d1qK4xb
GsDr4RujtzI69xvWRncGyXT1guhD1Zi9SR8Rsd4yXcTsSNqPCsw9St/a5dOq6wd35uOgh1MCDkPD
b08HHUaIkt/5hQ+/nTKUu3i7IPsol0cS6ewWkkxg0vCwWkpdjfQs4+hf7JcrIn1mOru/bh+rintO
Q0eVHjmhLYynAPjasJ7Za7rfAVloD/wV8OrsZ6EhT/YmCkUpbicrO2wuuJRJwBB+XS215Ir16tXD
VcwEITpaNHvQjhrqUsHiH1sDlZb8dawMaSCx6IwJuzQzyPDCBtjeEjlVLcztrjRl2RK3wgh3mqaw
6bdYxy/SiyaQN8FNHDLW+4y+MF2d+GYoRu5aYyG+pFY9p6uRD+Edm4Pcl/sgFBUGqR4XeKF2UPsK
t95KDSYT5F3lDX9bELtjasoPeZAuQ6+yzZ75X2uSvpIUpgtdF0+NHb5yScTCvuyjowehjQ6yfJA3
CKEFqZCnWRCpOjTABimu9GlAQDERzABV1GYiz7OsmJKfSmx/j3dD3H6Yz525fnMhHTrUm+/o6DSk
JK+oBUKaEFeFb8cC3o3qFHaLf+bRH9aaUifeZe09q9QqXaRGKyyo+hOwmnKgEuM4OaHId8cLNvYz
EisowxHji34DlvwEh80yIaUi0zaF5XM+zzxDxyczJwiE3hKD4bbDEpIpjnKKAHW8VGwB0IODOB3e
NUdsWdL/YAyJmCXH8ZhheGebQi5KfD3rVCwI/YEwzKziL+TsI5VwiHe3T41oyCTNy848lCojQrU1
puAeBqh2txIJnWW/DwQGHLY9dLzA5031QuOwZjYIpnNP9TcfkhtR54N+/86/BoZORenUnEmRJQ27
1gs8TkaxV/RDLn8n8hBrGhOTDqpOUIuyWT29+dIiWa+zPbGFC/ox83aPMe2qLdPxeaWkDimqliSn
3AAO2fdzcqKTfuZ8j0YCG6Qleu7mvRpKULcaaX5xZRI/dS3GlGjDf9gLWMERALtO12D+92/hALnD
PeV/MaapXF8tXt98g7PjoW41StfaJzqI/wd3LYfjCG9j9WezEnDA6MM7n1JrrUoNz3eOS2xdpmAo
Oz6sKcUfgbLRxW4at3qDwHdTlDO2zb+j6IRcTeMHcm6gzyAxRafP0NkScxXHoiTqaroHk377b3w/
RMlBV8g81FN/9J3xVgqr3R6uRHRvm6eDByZhGIfHhRtu5ScbZHlSLloAFuqIXVoGyCKruSdpj9Up
0UydZQACXB6RVFn/+J7s/9gVnWQYJdRVaUs9W1R3ANjWYukqkr33/G8jMwf/m5QUOB/zO1b1AoT4
VR6KzGKW6AigHKBg6rBbg95QpWyp4nD3G47DM6o+P0nFsO9f9UG62KRj/iRCm1U0B4RgCbGaAixC
6nRhyrRxgNuKrLiVGtMKGhDnhLnbdrlDakTsOBWp64TUY8IqpQlgE0Q3EYxzeWRq/1kVS5vg8d5d
OyUiIyeTqzJ7JZnNRnuO/dQ3nom8lj1V2ZVIYNRzYuGNZcEGgag/bwfGUTl8kg3Usff3mx5tng5Z
4oukKlqgEJAM9ElzG/WcEDIk5ZjTmxrG+hxGNTDGcf1TLMuO5Q1CCYQIRMtikpREURffJCtQvTQ2
sQkvM4/PGGWXUMvbThwL3R698LvrUS6QwA56IrViWXbyd30yCC8tJlB1LBk4Z3FYKDSlvq8O2/3d
jV/j4mx4U4/YFVMDtB57sACRIxs0fs1htxWhoGxl62x4gZqk5mlMHuoOfw9K2VaQfFxExQy75Etq
MNMX/J47zgwhp+tKeQvNmHkXwnwNGqPuZhJRd06sN9GCP8QCQzc8VpWilyoBQpIC8b3ibm7fCPsc
qzfNiL8yOqIK5V/LJ1uPgsn5sBBZAKjDp4lKUYqe4UTKUXIpFWwt90vIuWjVKv0Y9yILQzdzrLVb
7uTRbb7no3BZrnFOJuii+ydiqVBQOVao1aNsP5G/IhKIFmZ1khXFgIVpKJnjM9rkM9QWCgt//uj8
q0uzmQLbyNX1zRC7Kh/NGB7S7EJlYOK/nF58ATW0/hYpozdiIVSBho5AIv1Fx0kYBwco7ilx+yL7
iBtK9HI9h7zyIDijts1C6+W3X51fl/TYo0wDu/AXpejFjHIdLjeDvdo6/VwMIoSTXzuZf9KpcT08
ubAnY+1RyGpeQH4/Mx9DD3yS6+jMmyDefQG3TVXCy3HawXLAcYcIjeI4w0G3E82kUzbGO3Y6O9za
6yfLW2C4Xzhm44WClQux7Uyf4Rt3wv+t1DPtm1E3dkLcSL3JZdNLcsq4+YGtBpNFoXp9k7OvQ2Ke
gqCgawtXzSqHPSKKAXs9hpTe9+HA8Zczs+mVI5SC6BBoh38iKXTdZB879tukws5ZitQ+XPBpwMPx
ExCm940He32s2hwV3I6thcokti/50R4RIjeSsNF6n6xrAo3fWQfmKJUru4MLVJYlfyY4pjbDXbtd
4k1p8bcFOVDtNNHY6cCQlsoYHT+k3KBD9A8itNmM06mzFoP7ZfheZW39ohiE0nsprZXTzbf84r4G
bDYfAL+jougIcBrfXJgeABiQ7+u5SeZwKFHDvyAq07pGPNuj0c4BH9ucB7NetPCX6Sl45owyWSte
gdVnJe+JBAOvV2fOB0sWm6nXCPz3Pnf6cTNBFCst82YrEA6uEEMhTxAGlI0FqQc4Lct+pnXm/pwk
iOPIQPklNjdRPmNfnX81Oxt/Nuzgl3pP5d1sguoVIntVMqPNEMM/bzLeHzq/k5QnPzJxIFIoAqqH
1vL1uPORgsRdBu3dv0UcRabo17GqikV7RawTgpakcyZZ4tmI6gYWg4DEyisPZoO4jqBq1+FPCTUE
WvplodUvh1QwZTyen4pGJMHR3sn9wWl+E1IN8j472di8BfyaCtqTQUWtfEvRLxim4NhQBWBfkz7K
WyIjDC7A60iDqhdStAzxCO22DoPi4gojs4YzFee7Mx9TzboCI0OAC9lLDjr/C36zdlaysT3s5zK/
AgJaXWftrZDyfDbHWT7wv/tRIUs6hiFQ4XtJj7EUKmLeh9aChyfIVapR7vFtSTiUUaTocPKB1wxJ
LL6oIx5/JR8CkjkFeF8Mod9IUwxHgKZI6JtELHKe2/R6SpEGFifBbTEctaJ1g0TkGMyxpKzNp1/F
mE+Vt07jrhTNrmSz/5WuAvF8kimuTkEyKWXusfmfg4gxkPccCV/LG2/x/8mvpK+fNWQLNgICu+8G
D/JcEzIttMerq7ZNtVpoajPBKWG6CZCimGrcJ7ABV8HTkbT0ULca/ugUglhdQ3hQjDtmiHNFLolz
+IsmOZzH2hVEYhU5ssy8WXQ4tYFvFPubpEebieeYd2EgP1RSphtYV9FX6j6OC/NrkRj5GEdHP35e
aYc0XoFc64CBvDL441B3RVxzxbyIRguZmhC11xtxreI4GkvB750fgMWbWTwxzA56UDDJhTpT40y4
5MIjxP+pLcHUvKecBaCkVKImAf1qSxdMgaT1QsRiXk3tXP+0+WZ2ojSHBpRTrOXBB9yBYOkMSCDY
t+am2va8CCVeV1DFOfswm30uC7tuEXOB2XKOMsRL5s50+PnuM8U/XC4bA4q7OXboN2MEoBhq6VCH
2gRvFGHSHJcfxtnfeAPAoek7+frzaHzLlKWdMAR7Br/MRhn9n9cdJzwUk0FCpOJlpBNJHXF7USZy
mp2ocTYe03u3VXQCEOzzhNQo4u0vSQSXvc83mXrU1NFAhCYW9IE0M5MyzfdE5pIexl62BzpBb8yS
u4M+aMedK5VslAiuk9e/VG0ilZf93LOaxNY9qWV91UUR00b+NQxQ+iYsSFu4qtAoSMBOLmiMZ+5h
gUw25x1nFLCnih9TRGwOmGejm6g0PCQx52idc08QMYOortfXgxJ42LUBikhdU3Ydh7ICwIY+1wTF
oDZvG2geJ8EDrZjqmOf9dhBQbY5G1Mymu0Ij4gSrMT1rCLQb3Bbte5oAGK2wRX9fbGiYDAita8y/
r5y1RTNJXNL4jw63OQNxye6O/LZDPgUBp/3egPKYx8St4eovYjOwFeXripi9Spy/vAwTNY+nWQrh
ABLQimgtM7uzSTYOvB6DYmNHoUUzLm++KTjX+vE+jF4Atj8viy7ihPdCzyvd+ceBdTutiICR64AY
/1kPXfu0PPXpLnNHMTaacJQTDvEJTMerB16avg+5Ri6/3qM6sK8awrl9wESOuA7nDCoVo4Vcpima
59oxiX0b5AcXw/FE3gkqN8ysWu7Co4OvHyE6D5znzE03NXYi5gIgcTz+0ep6/QVdCl5DYOGNOLJY
/z2tQrDOMtvSgSE6aO+ekaxj8jNVBoPJuIIRi/durBiAzg/xnA5w9iwUEZL3yjtlylyICpP/tTNR
VWFYZvHpKkAlpBGCJVqf0ugEH3SuftTMEbh9TDA6PM2wP6/jd/T02rXWHDhPSmKH100ymtkHka86
kOBOsxtzYHnLVWFEBtnXNNd1xIsaxNkm/7k23EyeRYzi3P4NJ3Fj8R2WFomHkvlnV2oKgKcZFSqJ
CDGgRU7fTFqyHIorAsl9w/w5CppDgb8woWLp8qAyvr317DL7GoLK9PU0KlpFSy5M0MxlcKk+3Ui9
6A/pe8D8KYfjhuvFLXmSKonvEnFDkO4G2rddO69rL4QmEkGBV4Gfv/E+rCVdqe5eQCUdEo6qg2ta
9GlOA3WlOBXj3IjE0TGLaffKuOwyV5dhsqmxk2pmwWwumIiTcP15YhSqQhVC82ySuMyruk46XNHp
YoIufn9GFYsIzFExv1S870S3CpJoTfjRY4F7oScdDZtW9nCk43B6OhOOrQZghEUdz9OaWeLsGilb
Rf1WSNugfLUmBSRKi83FYUAN993Bi9NwhsEQFHLOvNS7vukRLCT9ips3Ij0tEiqm1VPTEYjYD6vo
rBDl/aqXXQimBJQEPqHwFVS2m2gKINNKh+oRbEP+bU4TeUVIhxAUIlbCfIQ7bPNjvOKnncrbs6HU
8TPR0y8gqc1yifcsRw0NFDprnvfGRqSqPEG0jmpKjWl3VI2+x41iXPvO+2qli5qyYMKIdHFm5HiV
m3HYhpehPg0YF/zlSdqahatiAKVxV0JruoFxTYgtzM6rkvVogd6z0MLLR7JaJR4YbwdaoF3ybZBB
hwC0IZnzs7sB3g0j0crnqGH0YPN5poV+W34aOaDaHRBYEQ3KKfpca8bWSz3CuIL9VDS5r21xEdKO
ZcxxyIEuRBDTtC1lBpsykVZA2vo0n/oWrKtw9xKE0tMhVpRHF4VlTSCritMUXkiYffkSNqHazEYp
Fnz6c6H7HbObq+Hpg46oRWt5fwDW10ZNszdbXsfekaFqDidZnGDomVryEDTr7S3AqoKfPN3ftzZW
m/uKZFiEZPMhKb4ChNlviMYWjyUqzNfxAZrwqm7nmRLDtayc9moTfL2c41tXU3gZwq/4ZHQAVF+t
MmPPU5TZp9hqe3JpeqviKqUBq4dUtxovOQkuH8Q2VMuU/Y/Td/F007PiYul7aOar6smJRLCgdL7B
hLbk5yCKndYo78C5fguwZNQ5jCJjZOzAVGQNUcR6NdYzaXLSwjjhc7X2jhNtuuE54XmZez1gUoQY
KkdTLW8xRfiTGQA0//rTfVPkW9+yswAkpjHbowS9/RnMplpMrGHnX8eqdHtjqCEDlQu1Bjh7oAn9
rEgAAaGnaVMff9iH01UT9L8NjJQr6Lvw4bM5OD9shektpawsE3qYn5evNoUkvoQ3eQRh75l4cvGP
8D5mqf9nr7zE2KKx2fvMWxPltcvUgVirY5B2+fCXcjx6CVx+8c/YgIWAk8P7SzRIPOm+K7swhq6D
X8+jF+9ELkvK81GuJdFEaaC9lK4bMsc4Jux+Jtejz3gtR9BVP7xJTlhoEfFwYcLgeAfm+8rHLE1M
IHosGc/0pRZIjaK7feq4og2n9dhAGmvMZb8wopmuR4KN97B5ZI5zu/ODrrVs61votM/2jO8caVVT
Gm7358tTOLMUiwV2z03+1IeRZweDOip36tKyvLgGCqde4gNsqVTGIG74Oz7I/Fmpce90c9TQ9P/9
KORf9h5+SHC7gz4YoLNysE7Qc2DBY7c7KS5yfkWZ8Qgmytzn/aMaejngcA7XXkqVv0k2F176eyEu
tfGnxIHTUcZVoYXl/4BVgv8lru4/8VMECFm0ExGdcApxCJm3AKS/d+9GGn7RBDLWNattRpPmBYlL
hVaZE5p0fMPsy4HVXgklH3lToBjtUFEzXkykrwk6aUqeW3zJ34n67KopzTvjCPrUJot03LPCVuxc
OqrrQZt6uZvWQfT9bwAPYlFdVQEdA2zFnER6ye1K+IDrXgfrI+JGxSxJnJYk+5/vc1Fcy5U/A6T1
3NoYfusLlSHy8LjA2RgRW+jkk9kpOcC8QhWePPH/bcEDiC8/6ICvgamTArtx+fFTjM373AQ9aFad
HKh8t13rWHXyi1ZZHdnHjC2Ju3LyrFTHv30NEg5nziOOT8YDf2dvaKRx9QtpFfyUIlmbKKgqB4Do
fTz3V+sykM6URDh1Qh8bKbUmGfQfFvgg4UdcUkVSkVbwA7omzYwuQxZwmvaou2u36HIA2UnBVKYD
t5dvIwP6y930terAmX9b44Ixzqbr+EBcp5e3b0xAQwi3qgtIA17dZ64by0PHrklE9nm71G6ByCf4
+6tctqPNgP4iMt0GnSeKvEjtEsv8eUFJfqy528KUiclJGrYUtd5wIBw3xl3+Fx16TmWfN//z7klt
ooMQH2WvehttUyUq+0FmThT5xDQRwZVJmL63Fi3qkLKoRfOZ5G8xcc4X08+lMMcg+OTN2nC77sVD
vgsl5K14phGUykT4h4APIqEzqmigXU5PTL5U2nj4w9hQ5Ljr8ENCSKwlarUY/jgEtONfQX0c7JRe
IV45I3dsQqkmmaMoocKwG5M5FFXyGmuD+Bvt07RUpLet3ZYJ7r9oCYeSw/d3+gZ2BU4+XZwA0p6D
4e45HpDAZWxsTHqQo/Xi++OecSY4EfFZnuIziGTP47k8PXzzJ7H+7S4Pt/iPGbTgJ/6/L03JIFop
sHDpvX79Lzr2mzHSrewVn458s4ET69wFmU4svdzl46uWYq6LcHSEP9jUiBShhuuZ/2OvpskfzzYn
hsmwGNXF7scU8+k8fktMRdhC6sX1QZtTBsDjHYQqrD6enV9ANtTc+SmlczHgGPZYwHkN1bZTK1Tt
5dxIb2tUHjT/0aER+ps8xCTCp4hwZvsPzo1Aj0IvC6k8UeCFWOCFvttpjHXQXEuGhsoBb4jX5ABo
FqnqshVpLuXYvw+cYRQu4V74eCd2CubDvfqnVE8Tk0zlaji4T78hnlpc/q+QoS/yatzphVdzffdb
VvOX4oAABTUfvcPuWzJzf0ywrWq4XC0cgGlPO6Apub6jpIKFlpTiO+trjaS+iSgCvOwrmexQwHEG
+TGoytOUHjjvr2+Qg0ciy4Ck9fLHTptc4ydMs/z9Yqs0U3ZuN4bLjWyyWOIpVUeO8ZyDg+UY1R9a
MSWLdKACmQBZJ1QPTxT7r7ldK3W6eed7oqVP9mfSP6dLiYN3vw1HwiJyaytHKro2M8amzGUs2AUm
uc22pLJovR2ozwyhsUzIm63k0p0PSiPGkFhywopxExIqkBc0KDGRJuH3la4Q9xyFu6cNwSKgAAU3
eZC4IdgVE6hlks1lTdJAfly8wBHyetSwoqznY1lLT/BDy9ALPVu6o1GpVexLt+idRyMXBbpbzjUB
5enDrny4BDg/3uxCtIWoOdP+T9iULezCm0e45DtlZSUu/YW8dlUjTf6WjMn0L5yZc1DFYjRzXPoN
F3BFpvSftfUJHENCYEHSUaIYDV1SZrm9oz7tdhAGn9vHtokIqGMV+sytuwpMTD0TS+i3xkaLLt8W
U+DqEU3aWjOyjGaKSn29UAWMwn6JhKQ90MGhvq5ZHfaGgeX/6ptqQes8pTJaDEPNtBEt/jOBqsUA
aR/VRycfeiAb+DhYqBBRPIgJKl31hqZZdYuPp8lFdVCRmDegzrWejToXuGSRQMKhNkdoQAfn0NIO
3MRK+baSpk9KraMawnVFm4oF9SMw6sMReF2rgA29c21v1LMBeAL0DtF+XmmXnB4do67zTijVmy2g
tP/Y0VOg6ivh6OHiW4ZiwpaTyuUmWsnUit6gejHA8k2KgMIiPGw/6OxJ3OOOjBfhNsn2WLCh1B8u
6c704UCWPU1iY6kvZlmyjnHJDZk8mW+fQ26fe5CsjpXiijDcCqAwJUPpwLknTRk84DhbHLSMJ/Wy
RIdxeW101smsBnBv7CJFQ+P7P5ul2ChiO48Q0CxSVqHoTMzDSeAcv5WSfj5HcWm23Uud0JG6bfTj
xV0yxbkzAUrc4ocTy1seeg9YRYpC298CdoANcf7+f9VjhUqvqNBDVTCMau8spJSgPLrmGhdU0tzk
T7q974/kpi2ypdtushXozCgviuWCdLBLQClhmNGljZqdIrSGmePWHF8oKtoJBTftwC2Y2XlY8cmq
eUz+FcsyMnph75xDhKt4kog9/1RKrViF34UF0D8KCtWjVpuTqp/hWrM7GSA0K94yTbvZ98/q3KZt
XSSH/cZ+3rzdxrTNq5neqTEcLiYAz+mSjwTj5tw+KiQ8KxYCQLBuKmZGPPSCyC7TfR/AC+3OsaIA
7yX3dOzAkk+2BiaSReUuDy5XpuABXWSQJohikp1ZM8sKnXtlRynTbDk1WmCL04hKIrxR6ew1fcYO
oB/j54CEM6FUYK4KDLqziRrAUlSuduCR0cn3dVMGQVwpMquHV+5q21jWmbP5Qu6QpPhDPcurDjN4
kIvefQ2h/ibOyWwDZMh4YQ+7wjSINFy/5j1xfhA4f56+7EgdCpmtl26DtBBHPOXNsZrUG41V2LDO
irKCb1flK3fPuEmSRGzCV1vo/v64PxWP1Tdr7la7Nh626dHT/K0upf9kq6kuovL1RhEORtjKabOU
IanDo7lpOXFHJ7NkkN0QvP1TFUsu7ExaiNgOhC1KU82oWNpoRZFOrjeJ80MiLcwYO41kaZNd70Aa
jxGwKhUZK/+iLtssK+laNyOLc9uRYYysW9hNmQBzs+jRVykKpdywnpDTrJkUO85zMvpmlQBajyJI
B57Li4rI9y/NXulWcD7adpBLS4C9EqHWMmTOE1Ftdg+7pYkFbh5vsvwlDD95gcKn0LAak7FOZfGW
wkd2omCfk5chKsvT8IgMIj5c2Vrrlv4dANbaPlNzpFXa6OPZQqTMkUV6qV0L5N3f/kT39CoQixQO
o4NvCmAIVbhZ7sAXzY9Vl5J50u7K3UCzv0VLdoTI5ujJ6P/zW+2s1z+oSBD2WWrtQ2S7TM5E4QHc
aw56ZajeEAeplsXIeJcL40ATLosTlLZSc9vLOp8tGCklHFplCRqyYVbngXBqG6WS0uLnVcdS2Ibn
FpPyxnlPNbMoN+fJoWSID+KtAMB5fFSG4RP+/9fgCNF1Hr/kqLMqBoCueHcwi0p/imZhrJRojT8o
gZ+CFU1hnbghDkr9GCEYT7VH0b+4dPCDQA5r4j3++Y/NaiyujDpJXeYbyAb8HlVfhnzTJ2wyeSrb
ziDnrm7q+4VhhGzZbcOfsJTZNv6mpUe7mAMI3R/XwbSj4uRooK1eMC9TeaCMaxkLCQRMQuJLJ72p
fjiwmO49xEZMPP2SsyS8hjNC9fvcQSzL6OXo47/0uHE07GEy01lnfC4jemMPjWkPlyNmj1T1HJ+I
emb6T0pUQI26z4ItYXPBA4ZEg+xSRcpB90OyRaUqeWei8UMzX+8NgktFDzLM6OprLDVHNEU+8EuK
fVbBh/PhIskB13j8JNd11aoJo6J5V7xHCe8Q3GOnTLNQlITVspV2E4KUokfEt3Ed3z5bHUZ1R/j3
ravKaVEN9069DD7cv/tkf0vLNCKDilBeyMOAhB80xTx/W7rd2Z0Whv+xten8fDonb2LF+Bee62To
WaDaJOi4rV41B6Prfe4IIhGpu+6WPHA7RmzxlkHQbRz9RO9kPD94LsFuREA5Qm/4NQHsaXm0x/2q
knqouZ9mj0tRfZbgvBTMLv/3xF2rQLJJ/OQOiNP0evd6qt6UF+tH8gQ800WlS/BnvDpcLTJ4jtcH
S6UT/xxBfYptZU9/zmCrjK8MOzkyMsHKbEzlSZ2PNtEGsUrWLSg5YUTbCyg0bcbb6v+E/HFlBhMC
EOaZ8RuRpevH9BqpL+ens13IIUdNVBkhC05sJVJDLgt2s30HL4WWSZWgaRMxAkB4d5lAdqVMS/Se
pY+z9Qp0t2U6OwiuZuV5f0S2QCadwenQ49IUTgoR8Rnp5c1J2b2sSmRInYCNDk9m8QewusH4qeVr
pdUkrAKdVLJfl43/uxgT3p/eaHASvA0Gd5D3R0KlzBViyUgLJQOADDF/+sALvpaSZqzr6831V7eM
sKt404av2ZUBfs2E375gRy3NE5wthQeJ2dl8v3zqRuOGwjKs02EpKls30c4V16PnZri5T9uyS3xj
xgKv2nUBqILbuccgwqNoqKFNhk/0LTgfj/y233FKVjHpltJM544gWo5A/GHIstVlNXdhH1PYgEV+
oZJLusV8oHkrFJE+bsuWCJ11f9WIgXb2x9SszPqRP9aYTuG2nKSHb6X2BN3lCEqFh0uMnXCYE1Mc
aBSeodvevooirixjiTXBi3SMZtUpstEUVN+Objd80mQplAb54BVOSTpbWtPVvmOfc5Q8mbxaniiZ
Ei2Mihqvu4YBwKFGjzihQyIWqNrNHICzSw+v64a2Hi7Ou0yl6z3sZPQ5FGdksJpconZoXrH12SBG
A0iHULLIifTgfozpKnsojIk+illWLcYdvxKq4Owr3WEnzrU3K0YhINQ9gbHCU/tmWNVxyjWGM99H
mLwlacXP3xzk4OGuKMib7u3ZtnCkwtRtOWO+69O0rvypxXuEFwwbcnDJxSDiroZE+VxYsJEMELaE
9+bomfYBZiOnQXv3QWns6RO/wzfpgnNmSIw7Tg34mOGNNVD/IlCRfKG3yjuZ+jm3791umS7m1zct
wzHJFozTeTGke0sY0yH652NXSmj7hWiHJqJ6yDzki+reTd9XH6n6zUtA+MOBpWrd6aYn2kZURJCq
OKdKIpD5rsqTUmPV/mfd4TpnQGXU2OEGLZoLQ6xyrmXWWRZ/Y5juoWbdEG7Rv9hOVUhT0AYXR9uv
wFxSs5fvPf2uWowGJmo+Uex3HiXLLP1tINtdvCEnCb7b+eNazADkMFRJdoxIWRpZh7R5YAUWc/Nk
A1wtV5Bzr+ssQfbGJ72X4xrGx0iMYacwGQ+eZaXgWF5EIboQFjNpQrVp83kKF/9DmC428gC3Ylp/
3U+uXq1HTaxkwpmO2ObynGB2zW2BtccUv0i+5gu3LiNUNEwU14SqStxVSdS0TEpeDCeIp5ddfdwx
8SQZkoTKOxgcI96WlvG7s/1mPLoM87Wy3zLE6wrWcYV4Q5CNBj4O0tsMjasiweMKzDJhm9txyj6k
YfPT2bT4FGOIILYssw4lCZa9RCM4iW7iBjuv42317NpZ+LpVzq0KWhQr4egRvF4htoX/g7QriviG
RK/MvYFmiJWvA+AEKZXqiuaAk6cfoqFnRzm5goKdm+Trsl5CfytINd7pfrAITZeq/TKyxiwqZRWx
S0H0IKxJlODF5AgbfHhjuZVYRUzutlnbq8Bu0FnJhCloToT8jC0TGA4Tfwro2n4BPUGLl+cssi5C
nwZwsnJbzr6UtgRbcgQBipuJ5JNSeog3ohgy09oy71xcvF288o3XdV0yWjiBaTQsJL2JgTzjsMsF
nnnYzR1jNakjPmvFRvcfEOVY8/c6br0DtZJajQuJo8EQUXvpQY1Y9KAIUdSAxv2pdxzTyH7OFogY
WkhgQLMVlo+5yfuHZURMwj/eGwEtwi9tfftqA7vVw6ZAK6SYIqTuVMKhPaYaRmuZc0xy0JTfhjfD
d1lsNaIGnyLHlZIl0CuzMP0hCNmEiMjFIhFWpzW8JGktJb5cSKEMlHYyilwG/AMCG9YOQDnyR8NF
/7VoiKK1IEL1ynDIkhNSXUDhciSPKGR6OHHCk3vhlnFB1R6Ocl2Aw9hFFDNr6BIf3I4L6jBuB2XF
J8CEMf9uTQ6PniaGM2MD/y7xRYqK465opy9XW64GCN7SOIFZreD+CZfAchiANZ3seot/pd7o4dTI
h0c71ZTulj6owCBTB8Ln/OLLhPJKVfcTTDn0CHhdkZZD+/LiMOOH4cQakCiRX3Bnle+Yd6jXoGOA
NCSV7/uxtbymlC79X9+UGX4e/6Yg/WFAYBS6oAs5LQvSM2DW+hQrNFQMapz/bhcJY10yc8AQ1Qiv
W3qgOM/stbzQCQRe49pSxLPDNp0oI01amfU7UnwL7xYNLvQrj3abDdFm37Y3+YRPu5RC6UiVSf9J
LXjmQB4oGpxFdiGOjJGAcp5jXASlry67w+tp/srNyE62IMKJJIBr6SMovpzMB5KiIvpr3AIcmptP
ouNQlrvAXCiI5tuOFNkQJD9Rp+k5YjlpcX8QHWQs6ld4s86MZBLDFSgKq8dmbb8xaA0Yp7i6URnM
FoAgVTtqsY+3a6JQInQKpZhhMrkCPxxlVC8aA+IqFLEQ72CxJh1/Oh9/5XHWuELfCTdtJ2W4r5OJ
usvUaL4aBIUVidEFrvOCJTs9o2aawlH+OrVLARK/JZf1arUCGtwT2X5wleP9jZPgnFx7VbidA+fd
U99MyadCD2jqKVqBRA5WU41cwqBnJAKpSTBF6x8NvPrRwy3eByX3W3PeyHc4zqc6Gvrx37FxvDnw
2AP5LCh/30RA9unnV0NCTRtv6A1GvMHMx6jm0EknXct2WGd7xdNwCtHypaEpsfQ3sl45+ta6/jVu
Y7l4qRfVwF5JCB0eQZjJag3CiS1Qi4fEqkefAekVbevLY5W/FPrOw0Ik5EhJef7Nd6fmnP0RnwbD
6vzJa2t/gbA61CXHJ6LuUusYenWlydq4DCroxZkwPIpGKQDH9qve4KmTUz9vbsloNYPp5d4jn193
XvKKhPFAAhjto/Lh/ftcqzGQC5oYlblf6iom35R3K7GqUeezZciR3szoCWDLpxnEQkDH8Rfyh51l
9ylbNxCASOv7rqUNlrCR4xRleD3iI8pde9q9Pd1qlfUix0fccl0oUOgT5Ukobp5D8xvnOH86jifI
oPSbBeWAo2Bjjn5QV2tCtNOfgZzqk+Mkj2mdiNk9auN14hfgFlUOh/5LsDSKbD45SrZhPJgJyDYr
kOr7AX0Iml/Ng0dv5rBrcryy38SFy4Xj9Z6z7SXc4UVPoWVhaMjau4levBCPclRRkFkEhYXBdsV3
oILu3ZC4fVfpC5icxJLMZa0d7kA1X654dKwR9jalDoRaI9vBfTgpJtgzBNq7E/PDh4PZPrz6jkQN
bqXhplp7exxgIpieLve/HvdSSWQz/JZuzO1Pr06dk7T/maaC75ms9jQjwaRtMseT5/mm2xz70NeU
0A5xAqJv/w55ENQlcJpzsrcX3qGYhRmcxAuHd2Zc4PVgj+3FQojwH2yZ091VjgnkoSuUyV5Qq3Ji
XYhRVmcl7xeUI1VQLyBRt9okg7VnudVYOlhG7ocmj6ryKBipL+f4UY1Mo5Zpvg93bPnoM9edig+L
5o/VGH7TdH4X7dUPVET0SDN1wA7s5HlDinRioBoXhETzDjxtMnAJOpbGHQC78Npd3mpwtvaTAA5Y
HlDMDL0JhprRBOgkJOgcGEd5uP3TndbqBMym8+2y/82Ai87dTeh8kcLgvlGxIk8u135HO4Dh4hX4
ORG/c45u4ixl+XjJ4L3Wgw2GoBlulolwKBG1nv16tVI4fdNW5vLsJvDPXcg6pwsFtHRBqTqtK7Rn
Qn7iRV/596mJ4SQ1Kg9nEflm8Z2FY9ICOjM2mT9RM+WtI290YTX1Ad5sVExZA1skAwd0HVpK2KZ4
eXlZbZs0InZi/gmCEAAD576rltljeObJ4nSPVxJCxVNhm0Vp9o3oe1+T/sF0Ir2BGAiMNiUWZCaf
Pu+Aj4EsZ89xREDifvEhUQrPKzH0XwBmfkidJuKyFq96wQcEE5iZfaZyH+4G2Ss0v8HOhohfzXum
OznNPbqqE446/rWf4SFCDqEez6ZkWit99bQyFTTHB9qs8CO0a0StON4bKjVEF3bA5O8va6D8r5Pt
RtqCaffR5fVy8w2CnTPeopnQ9V0AsI/Z83mlALr5kDGYNmHn0MOtuUiaF0ywcQCn/Scahi5GzL0v
OJi3FC6On21UhOcTio2h7RYLBvrJSUaMVfyyhhnG3t4FvSkUqg5q27byK8DWRT3VjGHTFr1W9uN/
Qf46zKlQFvIo08chuR0Oqg6zsRfr6z04aPrDj6fN+MoQEo3HyuNquZwSy+nPYqM/g3MnQiElMS7C
ST751SAbGiMwCp6jWzG5V2Pp6gXpZ4tkKoza2H7DSanzIUbfdDnTKPpeZubpdLaog8NQRZIxMx34
ONyl+9ia4pfsP75GFhy0ejtxR+1lla1w4x0JJWZomS9TJQiwEnmVB41JDcbx8dMpiZvj6V/n5Ir5
Td2Q/0ZQBrIvhFzd0uksiB6lnc9CzS/W36cEDchxFgSviXNi9SimqCAxGqikBU7fePpJGLL+aL8D
SMsdfwQGiy8DL9VqH9KjlJF4wOqnglqGEpaWa5DO6bM3JiW/LdMdBDaKucf0ki+O1c0jgvFbEcY1
JZiiql7U82X9w9FJnhqGs9k7PMTvul4mg5BC+d8n48WdUrb1chiWpLPEB5EcE5AxUTUsl6eeab1w
1gxw5MmRadYVt/pVHMpr/f0wlMhekFqAZ4D6IxP6DWprkzRO0YhU7vfhJmHbhKDxVL/juFlEfIWC
OT7zalwavhu1XS2lechgffoDQVtICAFPVNY8/Y5+QjEZKxYoyn0bH925pjTQTOWP4upFyFnCVdHL
wmxIzGO0ESDVsVMpTlFypvv7y+VTTwOLmbIRXrTNjmy4ro1Gi5Nv/FFNmdhu1Tv+h/6LufikcF4Z
i16HqvTbLDg9X8wDAxi8tvFFFsMSKJo0Na7wF+vTf4NFye8bjgk8N0PrUua1x27ZtStLz3qx3ScI
EFFxzLXDTK/WMSRv0ok/LWVWVkDJE1Ss7RIqQfcoRecWb0u/I9JaJ2tdIv+wWW0satjOEoDD4MA1
zaeYjs55reG7txcRZ3ocnZO7CLDOYZ8qxu2xS1wHFnCW99UDNYatujn6YafKw9QZ88WiGCnvKUls
uX1N/ieTdrOgfDULo6c7e+grH252WlDqKAhFoRiWc8BvRZxTKnjCtJ0f1aNffIhD7surldDPxHOF
F4bfy2GXecJa5BHfqMLvWrHkRVTGGFefx3227YCyY0SXSGk8zwyzZWgN58NuCuTjL1LsKFvINoxF
tLRx22I7tesTDY4NFMud7+91QsV8ACtSV0+aYbHwxpxwcv3AuMKpvJvI3zLj5aHFRAN2uyrDZ1RS
C4QI8vGLRJgISKX2K6pqrdpFZoZUp7J91l6HPZyti5AaBGzvliY2EJihQXiN00GO9Q8UVZEack3r
HMKZ5cw4blax73IS6riHwNqyKwtNMg3JgdHyqNTXLRiragh47mcSYLoMt8P7/rOuRueE1XER8PCB
bjgiCnilkOSGHBuyc+1P9U8uTKbRvVbj95VmEstuB8DLPiNwMXvkFejOPYCMSnPY1lv9FZUT2ze9
ym6gfw0a4tm5FoYLMRjwR14Cbc6OIQBI9Y/WFTFqGeDaMhltE2m8x0/xdagKWKhcmBm93yBTPFIV
XmbAOfClWlGWVykEf9QtRgt9PzOEl1Z9ccx56VT6sXgVteZ1FvIPOu1qP82oCCwlw5DU8L5fDwMv
aBeVgVGyyFZqTh5kGaqWjK7OvQg8lUyssDm6fq8Ry7kNfo3vOrs037qHzza0Ntbm1o1AvpFOlDAn
hj95vJMhrEpHwIJNarcHKFODMsoR/5yzV0XIj1socpoyesCMa1AfzRTzktfg9LLE5EwAiu8Faz68
edR7JDXsc9RlbolY9a4u9MMyVytszoP6SKH4spYf2b6+4Q+XPvfZ3xbHEWhQNRsfMwctViuEMBAX
SJkXcM9i1oMKCrPgjbC6OvpkAQ66DfhYo0fayquCwSST2u8wBO8IEBqTk6QGQ92oAt9BTF0GOyhL
LMh/gjndErSZ0CWbc09bwL+ZFm0qtHidRzF2xqEFtaGCVX8I9uurY/1WiePpfsYgjMoraVnb/d5T
JsZFZVPu/LYVsVprIqnu5GVw/rZLfG78HR0WMkL2PgVT8uKcjilBio+pHYFOSthDrBiOzpQt5PSu
iqYBWp++NZbe6+dIEoD0BEf2YfszYsHRA4HIGmg3WVWlEunASE+nUqRxz1IA5ni7NW3Fldq8KdVw
PBLlhPWWzYwyfSkERatsY21BF2k0poZ3hd1ryyQbDJJJmB6k0RZIA2ghAeVFOrPXl+igxF/xiAtW
BTpVkiL82UE+tYcXNMh5svao4W4sLKUmkg7WZA3oOTonAFlu6aFTjm0T5Jgk2qZoastOTofMysrN
41BV/GJsk1jcYXnECV4oY2OE3H8gNwYRjBxVH5fou5BRMvObtqQ4h2SCZeWkHdXrfrZX8ij+sIcZ
uyh/aj+hFRxQIQam1rFZZ7AAI49l5aYQLTHbNacdn5DO6qDYCNjOMtMI/yL6fTPPGdqEOGSJ4JF+
/6rTcyGUBitQwcbPei6Uzql7XvOTCYhJ7IDDEoNjs4+of5I6tYpD6OjBcsyLIvtzMV9wOT2M7e+J
5LIX/BXyadeYcylEWfAjhnvtcOBmvMaeAMv64S1Lv79JwH/BCg53fCfsFOgz5yc4Tkd/m+51AIrT
KqpBITDb/Hk/YB6Mi3weQw4v27jLIX3VyH/EyIXcazifrkC96nx8GE77YNDhYBFNPmxnRwgnhE9o
K0cmUzHfoucdnxdDTR8zVls5Dg6DrvPCZHMvdAVjbA3Wt/x8HFbFoIP5eyGF5gQeYzsJcepk21St
S/zlvCUzZQbRHdH3wDbPFWSSAUh1e7ooqr0S+akJJ5ZD1I/KMzSRKq7j4S0B9paMZNLTAtz7urUa
YasnZAOau1QYJrJ5vMQ1oVn3Yn9uwgEA6eSnZ42J7i0AXngUmdapBHhsRi4xDRwVj14zpm5kf2IB
/CJ0YWejBwQSnxD6JGRQmfyMuB7RUPFODdZ/xvNyzR4IevK963bQp3RiKlhNAQ8z4cPFLLGGexsg
IRTb5yA8tHdHgOsVXdyZ5pzmp9rH7V8I2AW3CAU3qTXYUiXuLZkAY/uBZRZdm8TvfX2ZYP1TS0zK
2IqJuLLojy0060A3ig+s/Yss1sIW685aoTpJsYPkpNnSs33dLBWsISXd277Rs8ACXUvtLtfjyZAV
EdA/3wja/a5cHNoFVyqbGqZsNs6uAgAogAF32F2A9JrNpQj6h8NgIFTphahcQndOndoIRrkQgYgx
nUWsadXYHfH10AhukqeRnUWDyKdmQEDC7Xx4+jG7cGeAfzsDKcxWos8i2uEmkLWqdnDZTYBR1q2g
559oaxCCNkNN9wogKD3IgxkdFaAdJeRc9fRn50QJj4gRca6BKk8lazAhfjLSrgWqFAMMSikkyn0u
cnfwtZpc7KlzRTrRCLgyDNi5k3atj6o1KN3H9D2JoyufCj7KLiXsOz3XtQ6WfrIg/hZjlasRXpju
/JFxz85r1MZVcEgIIwd6jWCWG4AYQ7eTOpAPmEhBp71BjzfvTOTFtHWv7fjUt2eUre06MBT16z5k
TYvaRhcDzuSyepJ1gwCLTcMnqfJTxeXMgDHeZksCmkCzaoAWooAyNLUKbqf8P554s/mDp4BUNxlz
dJG6ZSeUsKyJWogxr4+ACg28lEDXmTG/FAytjR3ct9Fr/Ds/gweYHkvBTSN6pJgAUa8p6h8pZgkN
1iiicFuyeD4uA8k57tC3Pz1Q23ZK336n1qT7mcegvBr6jGrzeFhVkm0+/ZaHmHZD2nHiVcZz0chv
j8mt3VGw6tNzDzmFLJF7Q9Ar4xBmm3JXhNPXuwGKc13c/cYRZJ79UazHINN065fCFA6ep2EvkKAL
d6pmtRIPBSwmhy46O5elggd/D96Vkn/a+VyJUBz/1BjOa9Mg6tYExI9gOEfQ3a6A2jwT1w9ynBk0
8kDXhp34HpBtWo/cDUbelqIlBlQvsD+zS8aJGoMDEIfkvK9mV+QOWvJLBKgLx2JRu9K3oSBb6ZBG
KWQCAMutAap0pQqE20R3llcWtJMLyndvMO0RHefk+H8UVTy8h8HVGmVJFYKp9rwO1SXPdLZBwerl
DPo+0CsimZu2UVWXIEdc1ySXPM1tvhqJKKhds6f5AE7ZbmYULB5AZfF+6k8SCGJX3RceOXrYdGqL
xtXtFWfkVtEcp3PzsjtpNiZTtI3wBMNDa80FEGPFQTjtSWQ5uhNt/+75Dq0JEBfMd4usfv6tQ53I
OQhH0nlIBC3VZA2/u/wYr/HLi6BBJUQFeGN+9FoG+If+q2ujIAYXYXvp9YacmbOpmGn4dyAsFYUn
fozoim43ePeUpPxM2IjuPD92bkh0PEu7ru1Ry7zbbDugkf75cDM4qe5R5XEw5FUfV6UpcgIXxS2O
HlGBms1eTQfYCHSaRlYBJ6Vypifxg+aOytImrfDrnHbD4GIAwgC/OLY6wC0WHHTO3VZJ+8A2pzQw
aF1dQhypdCyPyFnG57pMc86XdbG/NYfI+OzKKtE4FPp0rcD51p9lwoGWbGW//wKI6MQbuSSLJAkx
p0ewzOzBhcaGAFWeZ5DuvTEgxzTnKVNwcmRvfl7U7lZ/r4D4T0/Gx89iOd3rTfAcRWYgsvMbpeTL
pGXDqO4pB1XDsX116HH8oZd0ZTGrLX6PRuLGKw+qJhiUQmFKGAblOiJbMYyB2iIoxojPXhDWGACT
k+cItmfQgdqDN3LDs++heDw3eBti74PBBLlqJBBr4nKYMA94wuK3euWUKmH/RjpCbi7y/jNXi0wF
cu3hULZfflzZOcHAjWTbhziFBCjie7+3wWnpk/nATn0QmdxKKyj4n2EC1ZeiuNZklyMK5WCWYU8S
sAXcHH8vyA6CzLXbf2nqdPv0wEmRBoSgw4NN1kdL95saqxcr6XOd7IHzDVDXnNXbaE/0gGmF5BRf
2PRf/u2ud5Y2UA3TzrfjTiHjdiJyV58D/8hVGXCmEptQhdZP6MQ8epD+yYgR8svWtX9ip9/3LIpt
xXQZg5TKGnOW68sMXwM++D4ZS18qX3vY2rJhA9g00eUciik0qXY+Ge3Uq83CaQ9u2G2nl8cf7rzy
k5vvO8MWar8dQHBrr4myUYJrztMLvfR1f0iX9swIErwxIIqOgoEMG/iqbVCqn13CCHriZuHCdiO8
90MnjmULr6qE1jYcrE/viCD+e09XMs3JLUVwK0K+MTIlBIM5FuAzZtDlIJQgh4bko4090YqmVXM7
9udPb2rAcDN0OeWiMujwBgWkIAED/c3SweKZXxPs0PvhN6+vezMmOz6LyyPrSNxzOgPzMrEAflv4
Y/v6EflMic+hnYgdES84I+hkC6I1f+Ki0dH9oeU66FdE54cPiNnXilThtnOlcIq7MNkb+wuJYGOf
LGyf+vONSR6kuwK5OKbkW770zYgkKFCR6u4V62hRCE0YPIysf/GyaG9j4AGKqpAOF8Nq2ZTxA2pb
PNQj2chsMniho/zic95IVcnesrMKmwWL+g5W1hj5BXAhTcjzGG8GEeI/NH0bYed89PrGK6Yf4maQ
J97Y41l+kE1Mchg+NQOXwUj3PBZ8HmBOs9CYaBysmRnnJ+WDLDNB9vkf2z3wbt+ycqYH44btGmt4
nkodHi1PLehzNf3kRMmRD87smxNx7xR8tNRag1pTmiPDJyypClYtyQvNNiG56BvBF07mHtU2LhLS
CnCQ+W7qteSshn4O3VlB0AGGY0sQdYwZXiWKiDGFw0iUR57fQzsUQy4tC7GRCpgGqEa4bTUpl7h0
2yLlBLmsYHAUkMXJJLAR+X02vlg4DdO1pU8OE0LNMoIMm8GZdmsqqfnhe74lq+VkSsl4xoZfhJWx
FxpdmpSphhXeqC2NUZp/FrdOPzTBGaTGIEGiWDdSMGG43zTxp0joQzA+rvcTXNvU9dlUgJznn+Om
NNncqYPEFtUCrvS5v9qXu7VJ/jfAX+NlOisM4xGuveol8gk8XpJuRmn8+7lpUlX41VncMp3KaLzZ
7LbLd57ydi2xjqd+i2t/S1CnZv/GhfqarQXd5p+0WytuwvX+ouEEcv7R36KNjeOlpMkIUFPpSyBX
q8LTjLb0NvCycPdmiOCLpa5quko1ek9PPzYfgsD0C4JUiCM9jDV5k+zuukzNhTJEYYZ6YNi9Riij
Ks79BL0r+LYiJdW9xZ3u56Xp9boPAj48GZo3V93WPa7YTW+EW4sWHGDBn8asxmdDAK7g4rAyjPO0
wlIPXNtbmdtyfRsWRyrmqD1MtX4ml9Fa568C8H1o7mez705uBy7PhbCWCcyxCdvBQ2BTt8RSUUgl
w7iGgb8UXZuqGKc37ThcoCE2kGeE0/UVutER4eNUM3+47SDE3F1USAZa+CHHqkpMPEjVUa8J0fOs
dewv1eUA2E5E39d6OEyG+yEcFd0RGoN0JBOm7Sk+2Gh0791374sR8YGmAKAcz8MEcbLy3ZLcqPqB
Oi2tDm/q1Ze8Z+UdkN8K5JipnohJyUXRgeDc+8W68GxgPS2g23YuUQTDh+s+4jU7n8Uw2yAFklJ1
pb0SlgWB0tbS11+QhpeCMG0dksXla9t72zti2QVp/vQ9+Xjp1FaP/S5BGgQvpdviofOrQ1vBHyTW
Wt0yvacQDzKHgzD29LH5EnmCGpjxtKgQ8OwnxSl3iVtqDsoBalAFZC0abwDwG6wM1SXPTMPrAU5e
aOZ2ADDx55jfYij7OXHdJ0GyRQHeNUFeBxXEdaYp7grpjkaNSw8T+YVRznLVTqgGgv5tHxSyLopN
rESiqSSre9KdQTkhcqhzz3+nZkDOhdWDcH3cWR52SufMbC24eWJl6Jw6H37n0XmDnBU5CDBm6UpJ
Ipo+xCdcK/VstRxEG0Uhdh+zzdD/2LwQKsyh4J5GnNGpZ90tbuh7KaEjpn6ZVNoPOAMiMZCgHy+x
ivv1TsZBpLQEGRQszhTYPvCCVOwLUTaR2CuQD04m6oS8ZLHy2MFZoOoR9cBi1vSvojWFSlzWQsBR
zH7aE86r8ycdDMYUGVnLj0eF2F0miQZPGBQb0FEDeAN1u0qVZpV1WRFp8ZLs9kbW6cXbYH4oyNM6
MeOsXaBimBiM4qdFwLvfpWTziebgryAlJNDG4YSsZwu+4iCvonhkvbcCzcW8oof2iRmZOAWnld/U
2tfe4v7kxuGEmX/jgwN0NWNjYvIn4G2pqTyP7oLouGFsf8yR4+y76B0TdOpGZTjTvmZsBaRQHmNT
XEKmG5s8i28HzZtf6jsSZYVNwdTvXvK7C6rd+9a7Fb0Y8+BnxZHWL0A/707nw4109z5W2ksRi/KZ
niqkPaG0jl0AvkJ2tXXp8NIppzhb5iwCY4sQ0lbdS+7mnTn+kd2N/F7msN6iKg3WBO8u4sjTw3RD
F2DotBR/8LM3wsyxlK23QMBcNWFobfCmikR2SA2huC+WzlWm70El2OhwrlsN9d36TZYv5MOEY24F
ru/L1R4oTVFTV3DdZIqNPHe4GRyprFx+er7swMqbkGk/84JvX/QtmRhHTtn8a5Glc28jIb3biz0C
89b2LbYnl9pIdUTtG8yBy5S/5eEoCmBvaLCtEmTKsl4Nrko1RStTZMgIaYrJKQQd9qkbo2jMjiRL
boDI4WnIKoUW0ts7pQC5qJpisPP+8s8YvsSvFWHbA8iapg7Hiqp5wRF44yNym5EZ9jA8Cn2V1qIE
yRQLu/SfaXOSiwfEExD4ewtoSCgDxDqrhdOTGr4EEREVcriCr5PHMLVdegZlAjV2P+jJnwomxJW8
1sA25H/4hUgBKYQ6E8BVkKbx0WHK3DcSpB1az488Mrcb4JaAwHtdVeMD54XyxWt63Xxat6ctN3U0
wem7tKhzhd2hjL+4R0oW5Qq9SsFZUrHljeOjF/lXmdPdZjG1iqxV9JXN5JSQKsWAfLNxHWet34Bx
dqH5DG93weVR2stQ9eHrxekD0pJnbVIPY6zNsnF6KQgOpo1PORAw+JBx6e5xR26hRnGCeOryAJdW
/hLuq+XfU/JtmYnNqTVK5B2KVQIWDWjS26Vsqbj87msV48Dv6+b1piYnxOOH4yKqypcSlpbirL56
mEoXFlTpDVLlvkxkYunx28oIchQrY8A7P7YE2O+N1l3+Z2Q0ByMlvdTngt9Xi7ORZ+b84GM7RwPs
SX3kcd+OxXYfvvEUoK1TdbHRi4XYN7kprsPRq09IVN7Rs9ffGgwKOJ/zQdUiZCZ3vukAxQt+CyAb
8v79wfQJjafBA4nxmmFBAgf0rsbUhwoxpF+0nmCDygHq6jEbk0aKLWSBdwMcIGS63MaN1GYS8Wks
l2Rl3wxPkpBNNxgGAS9DY0J6o99tlLR3iCFWVMkngY8mFfWt9qnszArAGjnIhoNRwvzHTdPrcuxH
hZr1Dpv+nvBw9aeXcLjHatAW1ziB7vTE73WA6NUj/Q9HnEtGh0uMk8hd5ci6UQ5scF9/9Z6kAC10
+14sBetKRAJkIn7q2vHSWFeYhrSCJ9EN3SiyB2+8yqOqcC7e8io7mQtGS8O+IObW0otyQVdtOfBy
F6ECotJOo5/8e4JJtnfrN1q3Hga1WbVEtqfGyHVJaDGz4BbIZUrW5K8urpSSwekFpAKe2j74lbxo
xxkAHSyRpnHTi3hUkrt7ZOMIXxi6tEsW0f6O8fZOrSFSg1J3f2BQBU1SVBNNQQv1CNoN0k3lF9r7
6XkIm1I07toZb/cakq7mT+Ai0eKH/SV6m1FmBJFMTzqtc0VyT9NpO9lm09J5SteeyWK50xmR30ye
O8Uq21Gw6W0k28MlF8fMXviLeI6IEs6r4W/A3o4ai17bUWeI9qFcQRX1d1uwIjFXPgATmKEIC+gk
QmeQEBHEGc+WLblRgxjdgEr1tqI6bhmrsTvA+bRtSR4P6X6EZxuxvhEeVid0FUcGIvkza4BVl3LR
1onX6pLNyZiMfDypI9Q7IIXBNA0EN962rXEsm9hS3b2NmFOwALJ1epZTd2HJlgCoFLoBCtuPFvmZ
xucJkUoITwxU/bykd2In7mLCeIG0zStUvcvDxlnk1sOudajY0XZfd3nfg7Wq8zPNeex842rv3KHa
kXa5nctb8ZrfhvRXPaVj1BdF4eWhmBoEUxAPd//pKVmbprMN92U55uVSo93TF7hRjasKxJsQVOXu
ZAhXpMEnWpI0E0bHsaKucvN+3aTGH8iBcjoOnaTzI1PEKedR+xLYcFaQ/lnk3HHHxoyupV8fknnc
TWED9KIgupboEnElBCbX82RamTeiKzK9tazKthNlbdlhBORekkpBzcHTW8OJe+Vv/An6AK47kG9v
uYMcaxjGL5a33BWGx5VSoQ+ZkHdvJR0hIKhqH6suLp0ptmzi/ZCwQqsCb6TLmLQiQa7qV7YoB2Y7
njNzLNMsFlV6oge/S0OQu8sz1npYO2fGRHf5SFmM6O79oLCasGrX6z7rmqdca9sCo+Vpa1W27pgf
+U62feXRQA1bRyQUtTRh77cxGdw/CFgQzzlitLSBngAT/ed+kzMlGeC9+wPNmjivwtCJtH1CoVHU
7HULiXuAGBlzBgEndr0Qw6ukfBRK0TRibHgEvyJry1uObC04emYwoDa619h+IIhNgcSCS12vjx6T
K7NUn6Bax4VzsDSp/byQlZG8nq8w+NB+RtorD3WzqwM+vQQGVSHvaIiPzSzLRuM2fv1fGWUUf+Sq
STtMJ+rkIM2UuXMgn5FjR67ifuY2Xl1RIBTTPz2x6hXed8FN7S3E0UmDEFGbN5REfwBHzECmOy2D
vzVs734GRz06oieJrREXHYDCDcFBDRULxjN4bkMx0I2Dhn+by+fu29tRxKk4PpYXbTohVvMHje5y
enC0Ef0wKfXxpUkUkoHHhPb/VwHEOkQutwNv9OJyNzz5RV4Rh9Cg2lXHUMHDq+Zt3wxByYO8qVM4
gHiCQ7J4vWcGzUH09I7Yml5/+RSC0Efn3C2+gzl+t82z+INWTScxSH5VWx9ggDSpb588x8yMMn9D
7DYFW4Ns41qj8apwgmZaMIFNy4fASEUDRmyRAGyUor1Ujb6K7DzG+Q0RbhhnHvzGB1YskWjVKO8l
r/bEwLRlHiJi0eN6u757W2GDwgN2qZ+WkYlI5zPEOGKiD5l8DfKk69pxFa71yd1RNKKgxtH5bNx1
i2DacZycoQ7XZrDjm58VD4D8IWZ6MV0SvItzDaYd8Y+0RSsKFdv4L8t/jhi4qKwo0lMRlOnEbRv/
JiYN6TGk58rVGMgWfbZcyAQ84HIrWahvcwmBvtl9scBKGs1NuPQx8FQ+lVvbSIejro+DZ7w5Qo78
qfWlMDSL1pJf2SEIqbn+ZDlZ+28d5rUZpOMiYcZjeDR4NkqUqDYNbvDeiOCPcPHh2XWolUaR9puQ
KUC6vqxFBwPvsADW/5Vraaq8WuknfKjJuaH8BY3k1IwqV+j36kSD8itJJ37AWWXdtEaJTUnPWhVu
vzit27Pv0oxOzs6gEq102Dyws9GsPicOxs9agbMd08riY1WseqvYaPTudv/9PzlFXXDDmw+DBkvg
jP0/CZHnBq+0o9bZbj8g6JX9svO56Kpr2gudm+3pXcgl2M1yA2uBlJMXKBs4gFApa2OIlxvtDeYQ
EaR3kw2V/+ccZ746KkfIK4sMtPT7tOKwWuwWDH/HyRglomMRliK8uzDKlJEswmkBMTYHBspOi3+0
rjVY3FQkGIUP9/xZOW1BM0cXDMQssAwCRZSSI8RwLppWSHQ1+PAQsdlYIC3u2gaNewBzcbSa/Z6e
f/eEqAEnB0ama1oVXT7WtKFS2FN0MNukmf7HQInKJoIMaQDvS0xhURdek4yZwmYnsWD1zHxkZqt1
yuNqVpyKPA2COV2Aod9yeUvcgs7b6NHqpqPcsSgA+Ja4ZYisEjwz11L3QIuQR+6UVHzfewBRp32o
DZ5JdRwFKmi4E8fzv+cIAbDtALDHWwFkRoXbsOf175kI8IS3hq0yo1z1DaYwjZAqVYeYHzgVWHL9
/3aG4ogRRSfpIdd7NXLO33q6y3aTQRCUQ6nZOBmB8E7M9/FskRLhW4R55zCRlw+kU0p4bbViS1R9
JYcYahBIcT+NA2DlhlNosG70/4cvxF+iL4xt/+Iy52VEOYYdEdLuFYNDMTaUuLM4GQE6lyAJmqyH
LG+VkdS3CI+++6QCExaX5o7uY22gUEkMCjAp3u4AQ+QN6RlvEEyzGXMhBmFICX8wBGVT5ELg/qMo
VHiq47C7u4i7XzAxoUzkKf72X68HEW7rRseMWIz2GhKfPMMxp2bszEQOwMH1nQ4jgke/SIkv/hnz
bqZCQ76do8l282+3Nc0980e0cQoCEuNq4QORDcPm9KJ2FyVjGtzy2uDLN1F+KQJPHK1XP1Q3KubS
l9Ul7Ahns8S4eE6pNkRzLkaT5CoYY4hV0VItDJBqm3H6CKDhSwWpYtMcV0M5RDGlWtUbTJfszFa8
n0EGnTfsYZyZCN8a1IEqZXQTzQEePzEXD6W/P77NOx9gboyztg2Y19e9E7ThrD11ZZwZwDUYmsXC
bFDUpR7Rom1JQS1Ec9WgomRy8GC13dg2AWbQB2gNOw4pR1YrjOYZDzVDVwGIeZP3Slq6xBo/E9nJ
8S4rz8XYnI9wG/b6lXIAP1QHG9HRDlKKpyTgiRs6wqubKMLNR8HfCHXfVSxgl06d/sH7Pg5j1XgH
PKGz2aXKtvy1xSeipS6qHsXOjcE7aRfnVxLl0uT2PyfxCQdeQTWpVtlPrJ1BJz0JbN4hRrArZ9Pn
O2j4J00LSgKb/syZpnfZV4Xt6449HD2kkKc6Xioj3Rhm53xg4FcP9DUudDKBVlEaCNVN+luWB8eM
W80cXs0g+GfX6B2piCHdmA9VdHNIwwwom1ja3y6aCoQneH0SF7HtEfgwE8lGKww1SoIg0+iJZfRY
epwYLklEG7PkM4ApBVEsWL2ODyMcGfR7ggGkz0blO1GInD1KGq9DxECPAgokMtkUQAev9ZNbXlze
mA/zpTlGdkCD6zHwJIjfYEzIdCT6dpYDa5FJ4Au5XNvb052sum4S3gabzodkTtHWglbCT6RPizGm
togte8fkgtywZ0ZXgoeepNY2iBxt0uz3gLy4Oi390FIjMJiIh330Mdqwc2aa0E8+3rc5ZB7OAvxl
hsSVAKhBj4gLGkUF/YkyWRdc3hJ7RXEGKLY/kJzb9bQ5T8s7BURlq0cuhjNABgzg+dpPZrFgXcTc
Jr4cxM5bU/uTz57G07ZPbkbefTF/xZeeGx602piHDvg6477OTStQNBKEiTfReDAX4vZJTAmhtpUX
c9w/3ST/bX53xDmusGKJG2anZMcxpFlF1LbJu9eJMe7fJJmEWiD5hDU17BE25Osy2KTpDa9kvykw
+7Ao4hfE0sJJ2/pB0EqBCXwUy5bwCALjinVZmB++myFtIcsEQFIH+0SoRP3kX24oV5S+4Cev+8Jl
wDBSllSCxLk50MJKbx84K4rMznyRebZltcy6iwQmIpOoCgHVsIuPesoK/gFbktYah1SxvOzebd8C
r2+inq8djY+DUiBF5UP+3wRYly9vnMccoNspIaSFtMTszZRILf8ZEDyhXrgNjQC6AhCS17BKutIb
o0pPZqWFWlQQy78qpZ3gFl/+J1wSTpanDaywwenFZD0I1V3HTr97SHI4/PMFH8JOsjWzcYmHwhl3
NC4HDXVAdUnPU9tS5nVpz1PzVRUmnzgLt9jBLERE54w/mmZfpa9XECum9r5eUisYRszWuOOnYVEb
os4zE8rhDymPahEtfG/ZtIeLnxmW210r8iVElYa/sgIhKeWeDlXsERQT2p3bSeKLXxwXxZewDdzZ
OhAj8GF5zs2QU0LvavEjhxMvbTzcG01D32afwWp0gj4o+5dNZIy3k1gGvu8pbGYnG+ONzFiNb75Z
id4VHN1fWX9q64vgU9q4lBVvtVn17vOlfk/uAvbL8Ei25S6ZIUU+U0xh8Jk5WBSxa3iBBkYiyyOC
JvcY6SzROHw9i+fv/Q9acAGYcN+0RtBlIU5usfdSW1+jLqUZCDnRys0qcLF0foWGWVdzPXuXxiM4
1nErtd7LktRO8Y++F88btbprb+zK0iY+f01UxuAEJw4hhiSBcLKoKEhBNXpDVAMZUIifowCGE2SO
+b+8pJwWIJpX64q3smxqF5/Ox70xoF7xXqtR7FCsNLTDcGS+6cIN8R80qzBgbTImxngAoBebrxGn
chcCEfu+Xsdn5jTVLNUrwaoKtKlIY+sRTMRYzi2iwKDmfxY9Y0rGDga/1aZvPdIWKrwG1hrj9WjW
q1o9cxrT0g7f6QiHKy+xRIV4GZ6FrctPiRIwLwX9idYHRrIerjkYBrcNho3rIJIzFWXXipaQPW/H
H8tY1ZCyg1yRcfc/9/vbeEkfSNoy33DnT2lNTd6b4oFtaNnyWgT9PE85A087JTSe/oVBIyiYIy1o
Ncq7ftuaaOWwqXr760RyCzXCQoKjABxHEqqvHnswbFHZfAQrjPPX+mllY8Uavx+pqXoBmASt/ujP
Xlo5qPN9Q/R+4SpGdnA5/V8iQy6rwv+av9mimbRzsDBJzcrTMaLW2qxJwI2qrtD71R4Ms51hf7vl
qD9adTUMkMQDiHzGW76s/Mw7prDbNk7LnnzoweQ9+jUPCjkBUDM2rrREz1JP2mSRpJBP9r7ERiHZ
sPykLtK2ct89d51HdFUiRiTmEP8zshj9hNVg5hR3pN/rrSRSs+NZqmjGCMW4bwZbU555K4bR4Krk
j7XNS92g5Z1c9XY8oEZ5qCyWnKbY+1idyB7qPwh3kCvkNT7ivSBWs4nQfEM1hQ/OHM97XmiRcoNY
/2G/V7eesheaz3Ro+0gXwEcz/5JWveU/N0IfrtRedh18qpf6LfRLFZR1jQLVGb6/uGpmvuj2ZO/e
6VhbAizOankRKBBhVWdHvI3a8fXxj3cpF724VwlLDhuTe+7cpqjX3H1BGOWOl20+shyfWTydRKwo
ah0UQfQzkF5KHDmQ3n4G0ELKQUWxfbFX/nc8AOrvbihzyM4WajX5PJ9RAwxGstUWBbxNITDo67cg
2lW1Dh7JZmybtj1d13y0AEisSMmdMV2KLjo5PVjelW6wIy0hT4HBocTzv2Lx/5iXsOZubgdF6m6/
7R5ydsjGMpf8BnyUG8IcMg6kyby9tCsexHCO7nMf70lf5quvKdHIBUG+mSkz3u4i5EmeP1VNHj89
gszpmuvuOET0tbPkcoaGh55keUR83QP1FNlgjN7Evsdf8wO5O8hyuCixsz5pSTazQFRvGFU4W7VG
kpSMI5A3bEgW7I6nxVkdpzP+uk3NNvvWoeLZpHg56If0a34P2mtpbeqQBpYrvZwZUs6GsVRyz4Ke
QuZpX7PcBKMkHwNEcvrEdQtRfcAxb4jM4fD/KSX5U37aiYkYI04739Bq6XeTszR+VUpyUNewBCZi
vKenQ2oUNW2EkaAnO1WIdeoCQV4Ilac6vBMx4Rx6/q3+ekLbu57goY541GTRB09UTXZ03XDyyRkS
UXZg8Z9LYmtuEDx6pP1rdmN9lsPo+GRAEXX5V6YHjTFBA/q6ECGn/kftqWsqcNZZTGboBgZ2UM0p
PojXwRK4WxqRTizfGPkqMrz32UiDkbHMp990GOZBjlxOQSmrSB00xTmlcm0ThU6XyIuKJR17a9Wq
EfOFH7Rn3B4Vh0DKcD+FCktxU7rFtpRpg5o+ep6FA9NzSU1KaBOkV5mjuUEdd4/nWXFZXQj5zD36
dB9YLgHfWshdvPcqu6SWvUUqfhBeOn1E8wND4HAUbHKVycVxcHZNoYRJ7d7tURNGvDCfrTY+ZyzA
WmC23QJVK6xeUDReieqRWFnKrDRikRsz0IRB6a4Q/KxJrXVUbcwPnUM/5AJ9I4N7LmpKIRGSsqNh
0xo+9Sa121ojItku0cS9fjWK1DLhYP04cQgug4bB9eBgAba4yRvtVtTNRrSi02YS0WmZG82C0VUy
o+ZKaW1p4acIoZxqR+5e9K0vLVkDezRGjMoJvjIAiSK6R7BPlFbQHNmY2WZCwos/+muCkd9vR1WH
HRU2CPgQb0CPmlTu1WlIvjEjWnG6z+HGCycf06vIm0tvI7/bErx8RIMbGfMWPvB5DzJ4ZgKazbjD
HEWFpGUmsHtQVtuWhmgRqHpndj8xPphLcM5ki+4PbdzktksWR+AsE2qNLLE5lXHwWoGYdzh8BPLA
vc5vSqEuTQW4VfLq6T3Osm8e9LyKXFAvW/tOnke/jzgeUz/XmG5n7rVUj+knKEWXNX9tC2moBtcq
Z8nBobOHkxMQYoAFiEi5oqZtn3J228zDLPETtCiFavVY98McwWCu8SSJhVVs15SGHltzBNoUSmDQ
ihdujN4AeZEJCB8eUOOUWJBxGUmQtOP0TldauGtgN1TTolb5aq2WmZCXIRqddDX8g2B3qst3wOm6
ZE0OR5LqXgqk7SePbvByR5o+xCIhtroXbpxMTBTX8RBopo0qX5PpR8Lj8T0DzzMeSP2zLZf8WipG
lRicHhdDpsM/qyqZp8+Sn7/Ai6wo63/yu/CZJwjbbpSyE8gjwmLGjij7S55BNOetVkC6p9BqEm83
xmSAi7wWZ/7F1YLqxMhJexFMCA5J6CtFaOv0iSCFSnj/++S0Oi3KSa8uUZMgupytfDkqk1iKLkiF
hSksDW8njgodbSLSqeftbncJBL8eaH9HLYJmS15wrJPV2PlSjWX5zbhsPoBCM+OQ4DyhSHQZIY9z
6X8u+waZR4dmxLX+l1vkl+5vCC0SkVmHrl4Mp4CHV4rMYc4THSZtsA4AVQl8UEx6WvVpYp5Kwo+A
Gh22GKiBuqHO7voJASaV2raVeIj7T/h4eDGk8CDtaMdg9dLaVgZy4Qaqu5yyEXtLLg/oZZJ2gdp1
7MpnZstF6StnxXinPcgIJHbcZ3HxT+HLPI8SIibgtoIgPK7deQCflclfiyTshpeUWInPxlz41U1M
milDa6kyvIHd04pINo+WBeOEJi65RZh9c1vppWe1uNKGUGwJspnnga8DNEKLj0sl8R3OqNR5Rihn
Cau077w0ONxEauTnZFiEKhfEmiJ9zdxRDlxnONVM3PVronePE+a2qWomhCyIvOs63X1NvI+wnGB7
QE9ZByQgJs/hdIhlUwP468zbAzIkbPHmZ0sNSj2hpmQrGymJ3o+M+nH+NaCyKDWDptj9jryEC1Oo
PihPBiOv+7KJX+Pje138Rxa2VoHTbpXj15aiqCGeVHLdETge26sKvr/+ToPkVBLcdBZ3OHCOsTrL
iAJG1ZcyJ+oe9gEAaC+YkSIJDEBuRCnX8IMvcPgKDOH0H8DSQtfzTwhfdp8klhwxKBmuOYpoC7yw
JC0X8QiCIc4J8w8PcZlvD11paHNluyUJN5MLqp4k8jLOpcVHgV81pPI7l9LtUc72Se26KA/Nb4+O
A3gRWL2KKg+2K850VGdAAb3KeBvnFTU1ZmsoxQMxtxa5Ur+utw818mKyVVwJgKMxBpg1XnbSujqW
7N3wteZpO/QRlGKcv4wsGogzQXYMDJBbX4xgWKQkgewaWMaEuLLSDMBwwOitgv702usDhKcH/QU4
ph5eC6aOji1FGibgZj/sQRHq0lce+3Lv0xSrjAFQn/HB1WUhmIDhw4QSrET9nUToB/KY6HcHMW1F
nxJjNkg3c1ND1zChBU67O127sfvkfmWlCQN33qnePQgrlmrCtyImC6JIxbOIrJUsBs9pWN0p5Y3Y
Z6TnsDk13/R4VO0bHvy3J8mSBwmf1P4PPIRaqi8KEE5vXsR3MKUC81n7RWDxE/GKEC4s19/GurGo
dgH1x0Y7+BIiylCLMDA9OuDu9hG8SBdcb/FJw+Aqy6MsjS+ya7VVrpikkYzHhR5mvS0m071ZQ8VU
3ZKULIaPOeSXjBkq7tHVW58KMj7o/SPx4Kl8zpB5YXO9vYYiqEbFXJaIOr09qZwCHGetVcyyDZEH
EaW9Miduuob0gds9Jd12audDGcqZwF0wooVukiPMy4AoPP5QdU6Aa6ar/IsViqwlB4EttV9TImIK
61eUGLgh45BfKM7ktihdKDdkghZ/gUF3cx2c7BRaGMDv5BiYlqtzePEczKpIAkNSK8dMbnaO81gp
+vEL9QGmTepBvePGayGqcYdgH1tauwKbI+JKrYKqhbMpVLUfV5FUrGyD8CQToXA8OjQPYJiEAi02
ylPjva0irSrvwPvBuBz9izlOMvSeaDinI8Hq0mKoWa4+RGcyfwmhO8x1l3yGklD1KMbZQucVXH7W
ipl3qTXtAmLbQ3TLK4rMrS3y/CbAJyKQP74Dlp6zfuPDq89ZapIjJKdpvGrVVR1rirYTVv+ROsi2
96K2E0EerjKG0qtjfJ3xS62OM4NPYWWHM8df0ef8Wovt7Uf/BajdcDQOTe7e9tJiqIBnr9gOt/LN
2hYQRtf2bWQL7xVYWY/lnPNi9T2NyolyFjmHRjkudKEHmFnwWq00dF2a3SrsQVk44FGmT5vuVGP6
8D5SfnIs3g56NrGiisTSxlCbbliI2yPYQ6gtWHbuQvgY8d/RS1tr8ImB+iSUYvZEj1SYUUokcUSc
3cLYFROTHkVetPZAVXI6mwqxrnNw0q2emylZeGVuEmGphGOcPzytHcVJNuliMlnqIf/qcfuDN54V
aSahILgEiGepCNJC7GMW5svdLKNa0y0lxtNjQPfPJ/C0n0RTIef2DiBbtt1pr6En0LCAAdaskbUH
D+1BkhCpz4+y3BJ+HYlBGeQfuwDMOO39x2eNYbz9oT0/55Le9nC0oa3ssW5/DMULNheEm+bKHDfU
YdA68Ueul4Clnh/iwGcNQ1X6BtUdrlJGDwmIb+eFgCIPcoal781iCK2HrE1c+hwCfsPx8O2OdmBt
mFcEvD9C9QKNeAA1Zh4oMPk5Hy0VO1HQcVpbUKaLUddqz40sVbP4yynOjgG1SpcMGB8llcpbXlr1
d2cXNPmUS4cVnjSkdKH4aSa0FjnCdB8G8zGkl2bhhzW6PtP8/NetHthWATt8TicO1cBbpz2I1laL
4Sz8M6OPHjMP5dGyvSns3kUm15/o9WXTj5YcrKewk9Bx0qGfNb7Vzqa9oX+UCS8fy+nRC6yewW7t
R/xTb+IE3YiK9gyiMBJoaKQPdTAdYvY1pBFAzGjhX5/tyusQUF3Jvfda60O2AgFu+AT+TiWD70tt
AMWdgn+Ny5FZ8xXsg3wN+e7U+ELorhfLaUaXEjETMSuGUt2Vmoe2m4xHbjnwJfp0UlKeNe1L+pS6
CWTLVnYy4XOC+PAkV09xc2RFdNnrcQs3HI0aLA4AfwIbsq365qIeZKW7wEZg8nDbE3+TdkLdsRts
/HPZ4vnN5rr0NE83YMKVP+D7kxu74/V50+5NcmIjazR1ovfWNkPq9hUQkfTBNsRyHvVSGHP59g/t
nAlYY1hZv15Xv0jc6pt6bgYAIAfmQGiU9GkDocQTlOyc3bHsYa6VaJ+fcLZDfOrSGtJ1abs7J+h5
WyLxQC7KxIpFhajJiMLmD18AaHlZhoOOgzOPYVdTBypMHKRyccoxw75CW6+gC/GaysYwdFDH3VNo
ThpW0f5dDJTx9YuXghl/gZ2gPVMG51Yyh1DaoVEA2gXH6/q+vxq2UJByMFW3nfGHcRj7Td3opEaA
wRbJrg8A2HhqfIDMlTfXsTZzBDkMfDPcWFmV4Rc3PyeMFS70GTaT/X0XuynFF+zY3PCOqwO2yMWD
Taqi1imqCKkzA57ENuqG/TQ3Gd62vmbcFNKm37cjGccRpTmAh0uMlIh8HvYTXRmKULkhPljjLgnW
gbldF9FLBToERu2HftdmkrlmDzt9+uHiunvRYnDI2aHuczuGMIE65rrXLcvnD/jmmrz/EuD88oqC
B/4OLnblOdZEI/E/kTeXvCisIu4wkjUepqabVZdVP9spU+0CsUDkT5aIbOL3pA9BFZ7sGaEGa4Bz
5rb6pasYTApSrp+lwzWkpt3stkmjRfniSurW8jIKWLtot4zg9E8MuHBDZCpMix4KqlkHoe9+VfBp
RKrcPSjSAEM20TqPjkVcy/GKqAHSFvByb8MspYT4LWQLLmRWLfqNqJeN4KfKG7wisPxx941oxciY
pMQEwcSgzamUOvhsuZvKbm0fGbVAf6D+uS/Fr4BF8e8IOB9EYPH/CSH+Wkw5Cvop0ryqef6nF009
cCL7cJoNV8/8gMuil+UPOm0qK3WamnEMj7Q1rTRK5LxhxGq3T4cUDsjfz45yo2debwMZ+bSRebxg
Q0IQCzsHBb/PusrITlR3PyqOIjWSHAbGkj75YQ9bLLFxkWrwcF6i/7TMML0tMJX1LHDAVBnE0+EO
nxWrhyIYnVOPNXD57c714Y+/L9pFJLaYWFoEdoY2fxWcgtdBzPG0mocF0ihQfUyZDgoPuJfouYgy
HS5aG2EHRNzXqt9TquyT4t7qSx8a7lJVgRmBdnfwv2001AxfsZVE71xSLrAN8Rw4x/+yKYFTjRVX
CijVAD6VdN9JJ22GjzDTb5m+o+NgsB4NzPd9OohhDtyYSGk0lkr0OgDSBkJjZYdnBYZG++1nQgWR
u+M5yIqljdcHFdCDKFrYi//AYovfvrhXttCTZpCHkNKPIfWy85u+cojPxDJjs5SexXjfWqByAeRB
vOY8bGlNn7NSlJMLdPidTQ5mXnuXZBUhq9yzr/zSGYl5eCwN1PUlmd/1AuZhrpF87QCcjWXYKfh3
vLYgJi1PsGUUFIX7Ag4mfCu0HRLq+Mhhigrip6Q4YdtUATj4oB2aYtlEoKXWGrowZDrOrHzVl9pz
JVDLtn7Ih7MclWXdl54ZJdHsLICMU0vg+Ne0EQJMQJUVMWwoTqRd67Od00Pu2DWMrj0oOpjFmvak
91e6ggTbKY6EWyzRQGzSiT9dKMhjthv8sMezOZy0f1ngqxGDrBNCk48cxuCLAIVnQ/uJLl6oH6Qe
xGgqK9sRMn3dwEz4Klcts6AxS2UW5/pVTIzjE0rdD8QqnibBoefCDgVEFtfyNK3/ZM61x8mzMBeL
HpvI32bLw1OB9gvcbqIyqMUlwmFWA+KZwBIuXZ8W+IWBPlDwKhO6pxT0OO1hvWggSAEZ4NDYNH5f
3Y3jB1pqeEK9oJxwnc1SVzg/jlfGiVPVlLEHrCs+mD48xK9WEVvSj3dyQ9HyGh3lPhK/DRdfvI8u
U5SWFQjCrYVTq5pSvxzRVmai9QHsZ6ZWerHnPwRS9A75lQsa9MrQ1tZ8PO/h7HoFapE6BOptTlZk
FcACNhIxXjtiXqvxZMtil5KNxH3xyVcfWYkwUbthbsmjQgonzBgO9tsvHxMGF+FX7NMyaxvShnMz
/sVHku2vTUboD1ClJ2Qe19FGLg8n6iqggkClARBxKxeo3aZDGhwGf/oKJTN79iJe/agwSNZ483Xp
u7mbmfjS7YxsIA2UEH8qmnfp3mbVn5ljXJOW6gS8T3/eEkceBsHw27rpj65kada6bFHCK5C+hi+G
dNqfR2SNPDZBpCxQPLVuW2t7UsTPfCQjr/aSktIh/dqQRuxcHpoKZ+hmVU9SD6ZPeyb5Gs2wPIzN
WnBeqv1GQtF7q9BqCQtBf3UKhYfcSdWOvll+nkzHDqkB8f9jZiGphjIAGwslY/aOZbwHbcFA4KBk
AzzhNYjkxbG1Z5Mqn1oNBwXmLdhP3SI5seW9AIn7dlEHnUsSwkUa2KUS++bnBQ3hSdMzV4XEM3bc
rBUtezZW2ydpwgNGq+dbTeQV8tispLDlOFGuR2UhJeQqvxc27Cfx2KeOyeDvdhG9Qc+FEaskzQhY
020ax5JLpyVVcQ7fR3Eamms8ZU3ZaPmqgufFjdEgTD5FKWNR17jRaeND90WDzTaGXUOGcK0G9X8J
A1+9hgHUChU9+82jrCM4WSK/SEYqQ8FIWMqN+zSsE58Y8KPU2C1AhK9sgz0KVyBZbaLtGyz2EO0A
VcwFM80YWF3mtVytnb4u/FsJLDd8t6Etbc2q711VhqvZEZ/qmBJIqRF3ocHNPl8YTI1zO79ufF07
FecsI+41fDYw8dEI5+taqDk2KnAeabuwXbcbhK1F+r5738myR2AauW1J/8Ou7c3Yh92+UNEZBgZ9
UKAsHXPD94Y+vei/pLV7fg/p2YYOUGEJKFVdF2Tz/5VwNQ070CT57OSIFdb6z7o+4cQS8DvX5ZQI
cIM+Jgx9nmb5UFL/hz72bqxFXX7pwGo4R/1213C/ULfAaQjPkTvktzQJQ/pzuDUIAeXoPDEKcjUx
ZQkeSoc1tb6jO4Dgsf9gr71QCj6Y7XLplt6UPqezGYbHwHgXMenKZyAc7Lgi+/dsZStjBRlxzdHX
6brBYdBRPVHf1aqNp2JfgwUsQ+fxBZLkyEIIzz8tERTnlbR6IdCC2zYJbCJJ9gc6T4VVUnwPeAk2
gj312lK1drwe1xjRK4tlJF81YkKpG70+mF3JZQv1M8sO5JZeIGnMxtNg+1H6Gu1huaBpS3GQSKqV
TzjSWCPqSnlsxlxY/YGmOvc191u+RRbhu9IvVhR2zvigTy84T4uVi7FtUUv+AzA/uxpyMujJ+X/I
+4ZhfvWlQi5H85BADPzbJ7b4w6qP1Ks3wLon9FS8E8Xyyyj7fn44eAV+eqJSAElJyk55YcS0DxET
rNnBhp5Z67hNCcq78/7CVe3GkZFbISxMQReHgp4PPz+KwM5TrRP1JcFI97AAgWNYieBjZyZPp8ex
b+uYksVCcZJftO76j4fMumJuanEW8cfu9pMDP8FmTPdsJZLAZrKSLoXMARDMx/gB8dZiywsGtJNm
nfhipGqFPu0/rvgoQeDgqfVtA297wudjLc8LPI91YZD4XGGHOec5NcLmW/9P8D1kh/Quet5L1sNA
jmRjyUfnxMCST6kqR3AH6eHUpIUn566hIyiLWomxEw/omihTlyUMJqhJSIhY6WDueqEMuprcGQoJ
fq0pRs/nWWP1jH3Sat1kpCni6ruOBlEzQUSCplS2adF31fU+j05vbTWPlPA78v/sP/9y1w+BVRy2
NI3HoB0YR9YtmO0J1sY7fudYC76fs3gd5611j1OLi25pNs7YoF4CfQM9/mMo8QZeYNsrfFixQOJi
LofjTUK+LlnaPA5ltxXsszUDUaTN47Q6SADY4YkR/x07Vwoc3yglRsvKqm8xyVFQ1vI5qhk3hmMB
Oz9A+GBkneLv78qZlJ9AQBn+pyRgE14Bni1a7u/hKQ8W/PwO4Sk5Y7UZTt1tZuep1jpNLovjTuki
donV8os8r+nulYYnmlW+z5pXQ/1RQttK4whWDYNvOCpmXbrat6F7Fu/Bsrwhz7297ak+qHtCdeSN
dSlgjfbIkCYrVUyRxkzFVfMPHxMGJfjysEg/OqCK+bH4XFRz/Gr2f7vsuBlSpaQm3tOlHZGfbE54
cmOp5Kv83PTroZqdzr6T7E4TFqTPB0WLxP09Hpz5N/d1aDCOm7s6lBDhJbKVzMq8uozlvZBCssax
uwK7mEmglLypurW9JW2RY3b1a7LOHCdk/MGU9QW4JysVDTzV+Yw/KIxGINLNQ+ZCQFuzyXnkKtYn
Fpr445a/PBNRj2Xxer7IjfV0vUZUrTRtc2Q526Wh9WiB3P5AQupT9OTn9iIrlK5jTmqMQ9T4EtFZ
AiZAl3Esd12dywBSYCKKKy4DpnaYB7k+UECrF+OjrdUgP4jfaTxDPxJWRqpWPBWjlqT31wuCXTu9
Fe/hgaItsDhsCUzGFK77DjhpP3RnYPXIm8LI0c7Y4PCUww7Zwybd50GkrJ7Mp2Aa6v3utJci88SI
tzg/XLvPQGIaIyi08nGaJILmiRcY4NviZhhGj/bRiHlSTmF2jZTBv9QBlvl/ty7yv8zfyXoUNLVY
OaKpNHL7aChsoLgUd5pXAPCUBu/g22RxLjvsvAxRm2kTwH3gH76ghuXpAaN+AOpSF9hI9rPQK1Ie
WQSAzlj1H6Bi9Ow4ZSvP36gWTjAcU5kb5UADjNH49FB5hyhqgH7NdPyhotd1ewTBSgE6TWyBAAKB
sh8M/nz6N30KzGAuLo+2+sb5W5CiLhQ3pksXBee58etQeF0hFRtgRnjBnEeuuLWeRgh8tBUm7n9q
TzzWWcT76vyw5ejZ+g/Nx6wr1qp5SOjCx5BPEmktMQVhTyhEsKabYVz1l/qbSvZWVafHgKhfBEtj
BUDwGbAqGeew9RBL8rPKK8bH+10tXMcRHsMAD4oU+NwttxpUurDvXqO2KVK0yALhP0uAmQCFeIvZ
XFBnXdQnyRSIyQhYWRMTt4E0X8QvUkYMldp/MaAA2lAYNmYkb01K5GflFZz1aWAq3oSlMBfCIujv
oH0SsccpFacFXvW6vfAalqCzzhx81iLozLDdIAlFToDkrLWS7nuxo9MXnLIdV5gAtYCMNriSu7vU
0W9ONCczltXXzXAQHVchPHzlsRbtCglyP8CqLzKF2ZMWUZPToZyWKBTnrR1ocQTYtddaDWHuy8nN
Ty+IclyYY2R3CQQtUdIrbrCm802V3bORxO1mVXHkPMbGLrjmpcqi/Jx+LCcDC8VMMWQyYnkzewda
kbVqS8hjUR+ZRDxDq9mGETFrtavhDc4j1tlBeue7C7oM9pe5tcUPahsP0FenNbXS2dSbsOaZ7sBk
5Ejl+r4IKBbEZbSPUirjh/NWsIaRCiuQrLg4G0wwH4gVGhViNrHl42n7YWUYrcKxJ3+Na6qX8Y9r
Ux6RkBs0RS/kCDmpBnZEC+G1LwpXnDuRsn0eB3QMcOAgYQBWt38eR6rWhP74Zgj0y5GaWif1tiu+
CiyvUREZ3M/bwU05mPdbSog2wRfqQJus34o+IJa58qTi4o68PDTzWwXd4jtygh4smSEnKYhoa100
oiUK11vf9FN1jiR1zAWACF58Ilc1ui7wNb6mVrpqSdYviTFz5/0da7LCJ3NXCaOZNSBRsVAw/h3s
ZTwbl36N5QsUqwBMwS39ZCFquitKVkuYRh3uNoCyQ5QeHYR5Sx7FzKgr+lwO/QD6KtSBi1ulYhac
9KA9B4xXAte+rUYnPriy0obTe7pgtg6nd4KTy0x8zLQvGSWb1tUVIE6uMB5Ioe1VWvCFqPBAjr5s
+F5u07YINdnqHc6qwXmmjkGIn8PIu+ItODciPJ5FeVZUczAOUMKDrThwSVNex6SJli3fVLg9r/2V
Gcok3pLsMF4uyXQWsPxnUMQECIEUkZpbXaifq4Q44VGwOVIuKuXpCasTLauZda+NJPWpoRnXX8Qc
vzqPSU0A7pGTskq1oKJRjotRchaGaJ/eEIyZ3yhzqkw/8asw5ntBw3bCn1QmLdQAEdXWWTC8hP/E
oLG9tijAn31UbDzQK9iJ0uX6Jk2GrOVNHfRjCdN6LrxvVpOG14ltmBXMKJN8jHOMHeuwiJ3cejPz
KV27RhIaNl8mDmp7H6zGAUZVXdnKva5oshna4vf4Qm4rr+eS8bPa5XrAEOIfJpY2IgG2NCAeF+DS
JFlZ+xIhCs2gCh8OsJLJ2KI0wfuxe9u9d/PkUfmmxDF2s2j636lrGSMPZFgmH9ZgpfTHwQjm3e6C
WFTGcO6AeQck4MzOxwqxCuVQQgftfNNJikr8BlVN9Bm7QFZh2L+cOCJPVQjtWbOltjntsc/8PA1U
UOPHISwZQK1t727L3c/LpCrWnwSzWzy+ATEiyE2Nqxz7j6NeH4/PbLM4cr9CTbBLUI/FIlqKIy/W
N4CsdLuc1Ehu2ztOIZtWVqXVhbeUHMHgMOJeEGhgCFsDg2evYOyqnkEUAnhSIFNvv8hs5jmkMJCD
lnjl0SlCHZ6bCAH+m1e4wrGCKMhvyGD5Q/p1/CJWLSJJS0I2j3Tqq2c8fsTn9JdqiWjvSd9PyuEK
Udu5rwehqfDkNxeVh1i51uhe6cjuQZRner4e1eSwBX6B5I+D9YR7FkX8fI3HL+DK9hr/fk0hMJEf
27B3WJvOfujBxA/VVN6oaCbLJKdsxGciVQhOcjhaOW1PEcZtsj+dJqe7hk+B/GYJSPl1PUjV4fPT
TZ02Vfzwq7nkZVWM98sXLsZz3+1QBuEPUiJvyOX8KFF6S1nW9dFL9gVVRA6CRmW4r4UAQNmk1cHy
4f+ONJgF90nJjSCw9098m0WdXRwSdKsm2O/HZsnFv26r9IGtRZwUrZ3IR9+vPXAlP+wyxiUbZCpI
6jIDH/K5puPTC7ZCSlGDC92n0A6vJQVl6nptnlM5aq8AUlCmqXy2O5aqSf19NzuYUqb7njXIc0xR
A1shoKO3xqGp0Y13gctkrv5HM0drgneFi7XWc6TK3aAxobXoj9/6Rkkeuq4+APfBBPUkhlZiseWc
fi3q6TgXEyVMV7HR8I3u443yBVB7BfpcfyJjpQlkX82blwqVmExKqPBcdiKdJoR3dEPqAznbj9CK
CfSqw5Ukm9/qpE9yJHSPCH0+bMQ46tlTNOKPwQ5a8WjhTIr9KxFAtFweWoeR+E4w1+lZB8bDvUhX
DuKvSnGZFdQl56KaF1dlxHydP16BIIiDRtARoJ5FUjED0sqOqaIy/sxei7rPhAu+S73mvubGPzm+
q6hhdy8RZfnoQhpIZNtvQEJ6QPtVU7UDKy76d+8H/MrPOjWo2nyBKDNCh9Cb9GGg6UqUYaCLPIwU
RqXGYn7gcbnamxWvnX7wxJz895lzq54rN+GgjA4db5DL1TSeWKEYdTpe065p5013RLV2FrdncaKB
qxVHCOzRxJLIBY8MuDYiuL1lCeLQatlpvs/NwLO+YDNaTK5RI2F1CKTl7nU3tULhxRJ/E1nNRsBq
RosINWANsaWaUX+/tgE41NY8nLdre4Y/aDfkdN23l2ZdHiaqxjgLyLL/Mo9KMMJ433EigfVvFHi7
ydmF0m6K29WZJXI0GZ9eqhAvuiUt12lhBaRtse2avpyMN9d9OJ9IpVI8TF8HF9hgyRXNX1xn+0ZG
+c03lq7EuMQGLTh4m2WDLSTMT25IXo48psiYN1JbwXp2qRhj7iDI1+4lElcHg0PovyPtSVYKorFZ
F1+DfZsva9uWYT/E6CqRz7CyDWIMyGpcY0/t6EikkWT+hsPYlEax8c5319TCP9fbeWtA5VLZj9P7
oCrhd8ajQT/AKzK1iGqAgixAe5/es+Bjy3R3C+YYr+/r0lHbFtLTjpfrapv1QQNTqF/cAi/0kbAI
ZsxkCPH64n7nGGlBzhZpJ1oCmms62bS++yRLs+p7Qy9lP4G2+h2RVgYHKz9gdMqXw5pg8N17zl/a
a9R6lnrfl11YGhXJGKxETP/E5gK+EIim0G51bkSEMvLIb6+7aUlcGImbrATmnTVKPzAKPTtScNSb
PprGsPsrRRaqZA45k5EVc2tb1FzG9PjMfsj0ngUDEGcmv8X3XmEUkvcYPa+QrYfRLKcyEWYF+GRV
DPl2T+fwOOKCQdmY9vrVMEeHvxqojmhXAt5yBMsGbBavPpZy4xUp051WIIcECDIIvbM6ObJsHPU+
yUCR8xzgUldeE/Ze997gDgd8JqMQAcpa2Xa688iEBxpEWCe2IyXoVSLa2D5OiFpgQ4XQXzXRe2AE
cIHTWV/+qOCoy4HYExc7/XVk+GaDH2ixM8G/AcQuZilbSGDBD5J8VEOSchqQIUrpX5N+Cv63/S15
xpEbvBzkNVtwJe7hkcdBFV/HOn1Gca0XElTOBlK2ZpNfc2PmtEfqdTEdlxGG8xjPcVvFSJcDE0Kv
OeRWtKcGUH+jXD1s6sKkqqJxTOYQtlu47D/fPDAh8FHeLBk85NSXehVPyAWyaFoCjezVa7qh76OS
TIbohGb5gGgNPSdWlyLAokLSbp8ScEZJFDIcMPb5enND5+yHchG2qJhPYeTqljenbkwzbnN+dilk
unTsWkmZDmvqAL8cMqO71/b8xZQ54fNvkTL5x0UB9jLKC7KdV8CW3YRIfFra/sqjUbG/X4HdOEpF
l8ix9U//SppuQ4cxmQg4bHORu5k3S5ImbIOU9ctbIU+PCrvgPnqftm889yHxTI2m7QJ3mvawuBsP
wuj4QtNlypfFkg0yQTA+somiQWruIMV0I8K+sIAFrYYcMVFgL7VxOr3wqvVQxVBblrC7oX7SYwzh
3seVYPHwc5R8+TB8AFGetirn4reP3UuSs3YeP2VseHrS6pIZzU7mHacDpNs620ioe7LxLCUpWuhL
oVGexeEN8WiQfT3T6CFOeIsFEQmw36Ipa1KorTtxbkpnse42S6Q2fAiyZPJmpm2CYJg8o0rGf+Rq
irBLlPao6RQ+mRG0l7hODDwG1y12v0mGNvOU9UKXEPytvlXYfpRhnsfGL2Om0klL+vO04yG4aJJz
7DfabLqiSHVTtpk7mhUYp14KeNennMFMI7TLfBtWfb6t39cyRlJJBYdErX1/KOiJ2W/pk0jz6v+f
CuY4ejYw56H9/HvKpBGSO02IrWDMdk1PX8SqQxbSprV/4FuZV3ZEsoCgpOHF8RnBy3FzPIhTgrbD
4QZmEbKIaLDyqEEmPRTHRQazptzOQ9HdBBEl3xjT+hREv6/t0BNQZ66DLW4VkNOwZgma1DOG5sTI
ppbnf1SGcBQEPV/pnoahiaE8sDfn9lSWoL+4ZSvLMF8IIg0RyIzacWkOMoYdFPHE30UWnV5IRXZq
ubUKhbgVBABJu1a/OBGmsKRw7bldZe/PxoOC/J1iBTjRm3m/2hKiTYoc4kgW3US5UatiBnCfRYkE
0AWCvUMUXNZ6Sj6tPwwLlDrEkqw3OCBawAIdU7Dq6BG99GsWMe0w5555QJVcjKQsyQMeTb2hw4Hl
IZprkGWrZR2igXQ62SDcJJezi9wrRP7aX8ZDPYzu1p7y28jPATVbI+KpncFFUmI7mCBsv+/bRQRM
dsLiTUz+DxXzX3wfI4z4LaVev6hlZ4v06PoIq0+ZZ3Nz6u5gtuNQM0ZKL8y3yQkmAoRnJcNia4nU
cHp0oj1KpociJ5k7UsYwD4AIaLcOIEgf/7N2cWbbfL8LcahPSFleHu7pGDR90/Ovt9ryM0ax4Raw
Q/tNr9Lt+vq5RrgS028uCeitVeWli1mzuxsPkyrfR5GlPFQ39Aysiwaeu/bFodu/WpAaUjCA7/TR
+3lS269t1kDaic0fzVXYx3KPOR+1DcDEeggs1EuwpbwKKWHmDL6kODgzK3k8Il2vTeOwPVvnnFSg
yDnTIuZ/pA4fVmZ2XZxEQSHb3o/QMmdkyLmvshzdVu/KHXdiDA6r8qQlSojz4KZcFQ9+UaqIaupV
ZQvBNLxg06sZ/CS7ZMkZkI/xc0SIvLvOxGN9o4PkSl3jbG/HiSt/Oem5Jarne89MO0uBbq/uKudg
4VgsxwaYu3YHmx1QZwsLsxRNLCL48BMr2igjeC1wOIB6pu4HuYAyH4bLc5+scObDvjcVGYMDv/iE
88XGaJYB/cN7k3avjaqdPoDh6CSV3QUR0jrlxd11ai5t23znTIU2bSRbGCH1dS9zj7eebJtVOzo5
vZ+5rvWZsK2fMWfLi09HtwPrz4vVzfyTH4PO748+PKVPSr17ifCmLrTcEmFcO5bogLOWLyU3SESs
4m7+12aq8T1aFxp+nCnDtlmc5+uCUR9V1gOgEhSi8wZE/niHCOABqXMkCu5eY12BPgV1DkHZdgPz
lUo3ZdhPosKQlxRis0WEDSiBj2ndBtYckylQlvF2wRVVBd5fcpqScrKU893YPitNyx5wAbHCjUFm
zq7wcXcPqF/j03JRh7yiGJugxBGVP9izULqPyPT57rAIevHW7gzhKVfdrMDNqHvR1/TUK5zrVrf8
fvXIny+RKovWmBFlvhVfyXTpxdIczQPkimcRXj4E91G+lQl1wETL5Vdwri0w/c/UZ4m424YT+2vA
GtBEqKVOIrPfPfy1MfobYgVd6NBaCOnqHqbOnMEJ+TFlJbhMxfqdTPZlGlMyXEOX/yOkdrgmW2H/
gZxjCWkcYNevd95q7V8RphCOSiKTL1cO/UtoU0fXImj4hP7rhRkm23fX36J4RvVhdXQaQ4HKknuC
cblfXj6EQmJ4rBc1IAcMfi0tMWWb3XVse3FuQVzyqDxZPKGP4CVEzqtkoKUyK99DyCI0kUDm6K2n
YCAnRnxbyELHIGpULXgo3Oc395amBlOYefT3XJ84lketpRCvPOHxBJ0LgyUlRtY54RhYjiJYXm1t
rLy3+bmq/ugkvCCAxlZ6es4nyCILg4qATZTX77CHP/Af/gDwvdO7EY3Hns7K3st5MSwzDTbMKiqd
udgDJJsJF9ghTrbCSEgLY6xz5CrKAzx7TuTVR0/Qco+7ViTFH8ZuyGM4OzvkGVHPZt3wUePEOBcN
ugEUiyhho61tE47IsrfCmCJjLoi3KdvFOiSnWgo1OY16pllaJ3rr/4Xr9vSncj8f88vK4YCW9bvY
YPS/7ZqmN6t/+GBmqeV/O49xS7sCGnEa3kg8+nNamRtUQdAuIYTWhe6A0BHaEG6Om6pWoxJLVaOl
grjo7UTr/GAq1DxzGjUeXUP7UNs42sy0QdgJ//zYO8lnnfHQratCd1J0eFLAyBEEZcv5iY2UXcnD
r2MdMSFmipQm8kGPsaookwiefaIVrwlAWgDkp4xQnv0Y4/aPy/9+dlcCcMRTdXh1HuqHeGmU/HnE
PE8YmRvGelShfJkRPRlerP5Ueu5//IzhFLiOz271ubVLw7X73J9crc9l0sx5REfUcakXChthjem7
ulcmV12CrgeLPmSbUZmbkl7KYZIensnXoZzFNgOGmiJUNr2yitRqLY31bZ41KRIuR6HkIPaW/WzN
QRpAUy0ImFEarV3oslEcsPtHWA/3OWsmuazs9I/XrZVChhYn3+68aq24UYrkBGaPS+wqDyQ+B8CP
te0Kg/bhyrv/1FwYGkdJQ+NBXZMYXy/T4ok4BWVonY1ZEhxhw8w69oQ4U1T/GopC+OLGy/cL5Yp1
OQ+45FC2ROBcgyVjmzumbDmkFG2+JtXl2KZ8Q154lkUlB5fyK1/XS6wIK7+nUSxvFSYmTdmeLbrG
KdeItbSOD9LuQ3+3D+L8FAVA4cP8j9BjrjltgsuN6p7Q+0cqBkZx9UFdeItT4sFqUbxBu8JNv6du
/T4wlSB/qV4rNyU8xsXDu6+B7MBGLH0o6g9WMUQtbvDaRx06Rv46GlBBcI9fkX2Iipgt41kpEK8a
nqG/T5siC9PHSstOdgfhNNcNLfcnfwRQPFMTwDCV7AAJqtLm28dCthLMJJwHCyontDkt0Pz5qy0a
ByFbwSfxBVPiXuf06pSiLuDS75YQZIpVPizISFnwbPeLSP0k5ysO2G4ZG9p1SnV2dlL5op6/sERZ
2kNfVSkKZ6dfSziSX/GAlBj3e+kdoXQMaPL9KwuO03Uk+Vu6x/KI+mhIj5UqtD2l7q0+uEVfz17q
diFM0KoSR/+jVIAxIv6weGbrOBAJbIVrej4rAwf01tXV8UMx7Zv6iBcOu2kMEFRgAhm0RIyfYW7x
blUt6Bc2svM74fyA+jY15LTIgP5UNN4VEju9RHFTdO4yxKQFaZ0tf6iizefUoHH5MAJ7qd6Z9pU3
6D0bxuILZTJzHRkQSiO24Ksy4PQHh/4STxAxlXMP9KiHo6zi4tfWnEWrITfqlpMD3cyWseJ79mX0
qxratsFrbghAkhuLAws09gNwr5iQ4x+ySh81zdN84HdCofVRY/2HEwSQzsm9meJOse9uWzrkdGti
Ov66Wf1bcTWPBhJgNFdW6BlRhzXqllPyGpfAiqGMU2UvLDqm2Fvodrq/KuJI/2/55qAX9iA0xWyA
LKTLMvpwfBqGENdExTAPj+OIKz9VoN9bmgsN1OZXktzNIrKtq6mlGN+7Wfk4e8oe/txB+/ac2llk
9dgN790gWfoIVM//luh+QQNRNA0gZ+n/ReA4RUor7tm7arrOGpReN1SLvcc68fP6vBBiedNU+u/O
hAIg8TX6lJqHOwJN+EiypjE3/u7w5e5wZ6cUEAkm+i4VqOWgG6L6W5B3Ggjz95StlMq58/FtmgHj
NisDcqmOzo9ItRA7ydmX8G0AhDVmTF4dUJ7ZNCR6IN30P99keou5hg361EuLIohGqfcV/WC3J6fg
D1amsVGz5iBoZ5ksVDVBPdrlVfp0QUxc4H5BhZGJTKbKyxc8/HpBMw5DPadiMHon0edHa8jwzXz9
4IliNrL0l9d4aIa5yGqbgFlUhXhFYS/8kSXmgXGsK9YSc1zeRhd4Pc0UYqV5s8RN6Go8e+Ei8F6g
zUaFbnUh/uQsfNC8yRVRMYeaHMcf1NvGrWcIFV2x4YzUcErENLmiUAE+8uV1goDxoHxGqxuWYHo5
QCAjj6+1CSdTqCKJNTpiKVrIN63MgyjaewIqjND6okieAOs4DRXENiHgL/3Mgp1FTLlLalJsB9IC
VIpXxxXfvaDFQKNSPHLJQzYBMrQSySzWRXJoxk/kH38LQ1Dnsn9CKWhGNP2r8wmEdiiMjPzp+alI
Sc1mAIPc52/xzDoRdgLrnxAaOsCl4ytrhif8WjD0Xwz5HbGwTTV7rVcPZxVNEkcxv1EAQvM2vU0j
nAOEvDlez2lXFRyBYv04ASxNx0sXX9M7TF5777cA+X7dMjnDG0dZOeYewI+FXgBgbFtiJ55SK68O
2+HhHvoDg1ourCED0m+sLN+/BsK8vHir/L8Z7s5Vqn4KjOyPVJsXZUYY+v7f0qnAFqFVbz/k3I5F
eFDlTg0m2+tPxW0j34XoCD3OXjS2VQkl8sTTHA+bGx87bLICykbWvOVnZPc2h7NIAVMQDMwIOVsz
AYjKL8azf5xvsHQYckaIbjyyEtL5gs9UfGG9T0sXjQY9d0QykBwBg3zYYMwCydj2TV+NWhPebg31
Id5+6m0RQU5SuQcDPxEYdwJdNuibouW8kqUQ2XBk8N+2/Z3x3g9yPUTt6I6ry/FwZegcftoDqY2b
96pKsAV56+hfPpF7EKQ+wxJNz/1f1RwisjaZGOV+YUwLqegBmoIAGR6VMN3ufKNWHhQ3aVTrCmUB
9OKexXzitR8/GpaBp4J/9ONOwTFDIg6cowwe0mVq0gzuBWtOgHsbxiLeiRDXSh9qBXN7zszZ40yh
RuFgITuPRQLKor74TEhz3nnCgm9Yb1hOWAOQ40/okASVFdmY0RbH8p3e9+zQI09l4RVgcdI5ad6A
gSdfRZlMwYZJ3G2JLScHcQMQ2VIQcfOdKvwuwb0u3G6Y8rR+z2vj/EaPxwX2s/qPNu5Gy4BnIsNB
3i6avi/wzif1StSIG0spL6y3/jZaR8v+Htumf16nHEPLaxjqYv37wuMXLfjTzzSmElvYhDK3rnmb
b2miBYWY0JmLxksJCVVjdqHnN/UioXsuu46ZJuAT9nus0PkHEoNBQeZkFB/8jW18I169AbDeKMwe
wra7KfLNr+kow9ajxu8Bww7gaW37Lpk+rmQIa/F8oQTdwHPNz3breMTtZa53Co+RCnLgRrC8lAwj
Q5/njqCQVa4hU9umSVY3a6AvdlZa+Rj6/TOCejLvPAEu1txxUKM04IecMEqxmqoBAFPLUUS0pGMw
9vkrb4yeqrpCXO+E34e9VikGdJfsIZwq6lGOINJYnc5DEa/EDzom6/JCZDCniqD79+pEQsUT/Rm/
1gHk5WuwhNJzsEjlyOnQtPngl5wx2qeLQ0GNv0VH41CaE+/Khh5DGAWDArH2dd5P6bo7/Slbnliw
H/E3j+5b6x6SrNFQsvxZLMuvMDA1H/ip10W0r/SYFSt4ROEtRdBFTVGz11TE5ybtlBBCL2vXkA6w
wER9eMrQHCm+SAF0YVIjbPpAjN4E+Xqv4raz4eaSILfs/pnDd1hYG2dKQJNX/xfTODzMrEJBHPmK
18uOaDKDovhpsvA9x21utLGQpmwLoWcGTtrZ+GY3UPRVVvJSdy4yKbPndfozcNSSwx2erNErODGF
yhHpbDtGFoxCjl7bEfool7aeF8BnHS30ujNZ3ngdwZZRk17RKaHhSAIgis6zIjJ54yOyC6W2qnOf
FiHMcTR4HarY1HxgmVLXjeZaokqxNBfrVeHwrX5rDs4rp8bqxE2AsS5DgE8ozslGXkoAc32Gvfsc
BQkLmJVH04pBmHrY58h7W/0ojo7Tmu3BGjfwNUMOEoc1/ETeWYKdnD7ySo54GILaF1JIVdl2bVhx
acNQoP0Ql9mtnP6vNTCD0k8nZSAEETvWhp/jFlN6JXoCZq4fTmwvpyJN1B3fDRIyMHVQO5CRG+zm
/YlNfA5THZWge11Di2dq73F3L4gUkaXnSjQWNOTH0EfwSc3Dl4WBVfHTsf3mw2qn898cXZvWCs+X
PPq2FfgjPkcG+LpfXywJm53rjEVBv8W3cJiatsBd7Gz+7BAZL7tCsysmDVAdoYWaIFahLKOqVZHE
BQIqJie+NmKXYTSJ6CLRk7hyiuK79ZSAwQ3ODOaQk3u/mbZdBksDG0PEmPapao+ywZYEM7SUDWC9
2eL5+3mn4ssllbb6OaDMBeUzkwP+91pDb1+t0iJqQXqqQMj9kmogyOGKe1uULmkWvf+hzyuC5lnX
DIohA9uJ3DgVDuoOcEDTaIj7IX43ZYNtikVfmsNNAFfJKhFT2WVMEH533AzCWvLcoUV4LaqcI9yg
oY+wxLfnxM95jDghOiIZyVqhQBGdygwhTstomiU86kZDJdad0S2/1CG762fJF9jPAgRnChn11GK3
xwrXsFazF60O+hkacAMlpo1yZ1M//qI7jfD598CGy/l7g8/+iUVv4PkvI3fQqjgtAfAIukqzWL5T
yFQ9mGRheZ2nydx1YM7y+aMbaLdq2SWzqe9pdQLq1A945RW6fny4FsAM4X8wrnq5iorsqwynFeCc
FaPaxake3DWOzzyDNlrAbVJhFPxOuIe9oc4+TtmuMMJQhmRZl6rXi8JNsbLoERfU55CHRKLPu31S
gUHTy7XL+eTEZyj4D16/ByNRXy+6b/1Xt+Vv3BdVzKDDARkcBRUx/ntwazQRlvbdFoiNWv2uMikT
7j2HBqEBmEOM0CbIn+2KI3mSpUfIAHqBDGiTzf8Inh4RNl+1xgd2VI2dhO2v9saEll0KcmjItePb
scH4IswX9G+cxr6JuG559AvbDo1BX4Vp11RKGSlysBwYBhCzEgLbNgF9pOG2CCnV6G4lzaWIOzcM
+wCADR0zYg8gafLT9ii06MiyZag39eercpbPj6GDXtsGUbAep65+z8vRmp0TJY7tZ8uITjaXIxM4
Wc1YcO31i7qLePeHdAk1f5UVwU83oY38wu510n9nXq6XHIR3p/aRueKfZb4cS4WpNU1DYXbFytVq
wqrHjDvNCAUeFnNt7iPZLdOg2BcL1iNeNXFvekNCqlwJoB09nzwRY2kamE4fOz86Omma79VZ1Dr8
E/dYvUZK3rYZZsQO6FRs5QkgIFE47tT9F0TnDuZR5Q59+Q6Jx12cWL6zE16tc37Om/r+ZAoDRvJp
LTNdkjnKOMoHsx5EbWmZViquTtkNE+pyBWf7M7smp5xrPAh+zuiqXvt22T7PlY0hz2baPmdWPrI9
CkKhxiGFZkgRDwM1ggTPw1LZy2hQLt2PfAg6nwHhOZzkmxK/y+e+iLyS040VO+1DuRcDk1lFYDxB
tJdHREWevnEoUlofue55x34HDZ6i2qVYiMZblhvh0L8Nni+s3A1J5QUSqxlLl3W1B/YPebLUM9al
49GEXZ3wgJUSAmlLsRLvfiLSGurRtmNPaDw260gNXBn/I1d8UBvlYadXM9XdLZOr3oNHFhXqRtSG
rN98L2NziWO3FBwmwf6vqCp+Zov2idrdhDFl3owNgFbT8coQJdLWvaIcVAcuFzYsn8XAU3oA2j+9
mI+/D3IW6g4alJROIoVIIfYLzx70r1W8Ldm3D++mOQVH2UjLzuQyyidha40HPjKWdMbTfLTU39gE
tDNgfE/R1Fsdb1wtcO7ZMwGfIr4CM5Apqyuvp7thLPeQY2skGCOOkcGHYuXZ6sImXLynneRsK6sO
mCXZ+hPX4q5kSIUmaoBAz0HoHejfyJ7L8SQm5MTX6xiNkroXnO+u7dbaqo0RxG8dU+ODTzGakdxk
DgxZ/s8qQxbE29UkQ1ge99KM60skeRyAv9VfnxloKrxK2vX77Ir9kSFufRaGMD0wrtGZNR6Trtow
bFnrBYeRWHIzyvpvDE8gxqwFGUqa6moZX5uyfNRlmIQ9IeYer+NRowSd9fomGfIEdEzxdeUroi9G
6U0r7kbWFvflDVJcQ48r6EajC2U/me8+zfSj2KzOOL7jY/Y1AjPMhFCgRF/tVNnaE71PjgpcqAr6
fLPOTv5DyjLZEHlig1hMyzilIOjjpR75S9X3j31apU7QUn9JpmvQwutcr735yz+z84nPeEGkhavL
75ClLrbyxkubDVhtg/mpJih3qu1NbCHcUqXyyjwpVTXn5HbUaOOKUlPEUhnZANZN01STWjpdKY3D
npsGjrqzDQE2QmUgSAl3MOCQjgetMzkOG5cWKHat2mM6egGPluXRE3BMaxhZhJdTR78cCF9KPrPI
Bu4CUjen2unCFGVLh3x75wE/hhSF6BzFca55PkoKuVI7vsc5JbC7H44UX72kajJuyzy4YwQTZ2ha
sPgZqHxXi8kIEKoWPi9S/0bD2yqfPfa77RP9IpuUxVOYf+wHx9D21GK+WxjyW9toTcyoKIGuKAF1
QMXZ+uFh0S8xW10RKtCKqR/VDgIVSHy0ts1EQsP5N38EHROsi768sKVFc64uAmSC1QRYIZRH3HT4
/QlAc2e/Lbf/3q7c0wUgAF5+nCDMvsmWGWYvLZbtjF3LfESxpaRkMhdHRstS6oxV3KwoDSzmrc3F
mydAdV+bx4vnSkK9oJeyLlM5/bLJA2wjl7+9w6t7eF7KZqOiLeU0al3U/mf4yXMSzqmVvTxqktdP
73oYCXBAVpmqH+sr7emY6Vg7qbLa11cvASZgzJhoHpMt+uHMaeznVNrck6+OI/Ab2WRIMTIhLQZk
Xl3ANgYe/Mt153hHfkX41TdOcy6PAagHEQb+EEGo95pjbDAw8dd3kkfHKxgHH0PjPeqsvaFY5blU
95X9JYJJfmb1X3y6CtE5cAmC0kKS0H+ZIfyMtrmA4Hxsj4ddi9WwxmibxBe1hlgjXMo2pSjx8EGG
acFb8wzZRBxe3rGRbtcNRfhqVq66al7X9rlr1YqeuV/dKTY0FissjxwWSHzaqVryOLqHVwqiXOOt
apd7L72UiL0mFX5lXwUxRIac663Lh7t30sR2NbePx1S9j3E5F484/6gmBUCs16ruXHZcwVrAGdWW
SJKbjqTqKJcs06bEuWY4Bi257xLg5oBV22qUUeHuN4KdXyiJfvxaPuZX1jFNPXg5vamgHl70N++u
SAVnfm6GiTNYU1qIhD43WRbMwPGK5m+eQxGjaxxLshg0yC8HqknkQR0KokFezHBfdIjK5Ip2QUa5
bROnrkqiIVCC4zsECH9C7pjRD8ayFHxtxrvMJwf59cY8uT7hB+51YxGqhMp5d6eVggX4XaJRg8Pk
ZU+UE7HN7DPWiUxCqB7RfvCC7bEHHJhBIET47BNuxMFSGroWBcCjuDa0MwS0LO9a8u0O4pgdqCyC
axMSvxmGDBWXAZWbdMXrRTnC5+S1RKME9eOCM8LKvyYb6ZzYZ50XX6yt+X6XHmeVLOkJ0WjloQwt
VI7fpZCxqxt01UMRnD9KcVcs07fblACvJ060XK7LqIXdIuEnj5GIxU5ENRwxfiYsRn4+qpTGdPgX
PRkmmgNyb2yLVRwwO1jbeSuTGvW6qfw4ZSYEtILBI9BbySlIr3eGxNCkYdEA/W9xCwplQ29iyGOC
dcgwTRMjIrutyYhyNOTVq+aYjL+6m16MmbhtyKsDtcRDBmxq2nbc9rt/BqBRbR1K/3CkoAyWkVIo
CxIKsMEYLT2y0l1Q2sSIDSxsCMuxXLAWAhNGTb7/6r2nATbAbA3rabRHKgnfQcxVrc/Kckb+EY5F
n590N+/QcCpAasHzCohjPpDYjhT4Yjhvm3PXY+Xx86TMxFrE4S1k03efIfYy6W0Xi5guxu02OaBU
SeWxiXBeiqAQUXeFihYcU5UKgAHjD8dVq7bPbIwqqMyrq5oFMJRbsdyLrQhvxI5o5kJmNo4OPY9K
DLAUlPZgX0CPg0DJeZGht/rGtei471iy2mSZ1rjqlVdna8lN5P9k6j5lnH6572S8aKqDyntc8Hxe
07pBnkRjFnrMnEhZCOIkH+duf4xHgkUqjRApreDYrrM2FFrJqAmkcraL234T9WorhEDFi2RYr3pE
SBElYgfCkpPM3YlTKYAjBymOllQNu+BdTg/VJBSjhVKrADEG39X0uHjju2d4H/wHu4Z7JyqGAb5A
i2bOOheE4RR9Vpy0mIszYr6SGaHxvRbJrSzsvOzigIv/3k6LUeQCkTUOP6ilBVVSryrkQiW7APLN
1muFPJd3dItElXUlUEUqHW7dFCXWtnMHaA5mH6LpUT/CwJtZTIaQyV2SbdbDbVZNFXWwfaw4j//l
pECQmRi0ddWxI8y04/Xw3zS7oy0lCKMHV4nDgAWeWZRrDuUlMK8lDS6W8WuEbZqqFcq9zZquRx5I
I2t9tXv1nEOxdgUFeMXXP43CGdcQ4NsfHQT4HIFfQXLQwy6Cit2bf1ocprmc/2mvJ8F9XtLg71N1
df/wuS8tnhb5f5XMj4f6jdj3QgaSP2XBei0k8/BVurJTNUlTgALEca054zVgMkXyhzeZqFdM1d5e
qKNN7nvGNBgmRset9uq8xWZAAXsp24sNfBLg5cKr5cNUryzjLTihsX/PczzqmVf3SdlhmmKricQP
XsjPXVQWMb1fEdPqgWCyzvyaI3j9FqqxlmaibwFXau6t3I3PoOGtkwdkPB5Jd5tp9Mqqu2VASsa2
IY+l/eUHBqy+kNDbe4IJpJMPQc++CslYJRexKE2caVJQgusTUFLyfupA8HnWs1Or5pdO/Jl7Cxmm
L46v1dR+Kw63BaV2oEnBcLnpaC3XchG76LBrxYcODz+Qbeo3MC5Nln8bVLYkOTf9wb9dVF8Z2UV9
IaSnfswWQIMfiwg5n57D6Fmw6S9CWqkZlji8HzZQS8cSJeVv96mRYcTsfPkWASEy25Ochej4sjuX
vxicKwktd8qPbgNrkh9DyOE38Y/FfYL98FsnbjUVL/GoGUS8KWCt5D4meC7WIa0/zuiksJCYZISh
EO46NpzC2wx3u7uG/28UZv7Bc6STtIAvAnjiZA08M20PN3AdWw6ogUCe0DZqD/cv7Heosk9xhaGT
VmW+t4O8coeQbRA30SDZCGIagMjBIvzd45VTAqmNEhrPnI6/O5OCCpj1PDy4TmyqX/V3OcmSZHfY
uGs/6Xr9xDsKAFqv8NEkjYxxLEP2jilk753WN8BMh68VR/ByFS+awLgLkJ3qKCBrRHLbm6iRR/DR
bCfHr9ZIAtOYmh39X3OrgFjJg40ci00FiuvhWoVff2jyoLho29PFDOezbwBZFPmdX1ai7+NuK5lW
9qG/4S+VWgG9pT3jc4tudzBM17i7Y6cZlcvQepmDBYdokMrqUnpu+rT0B6iY5VSNX1i1iLVfMuY0
3Rj3RuvAGAremj8JmqfRJbOnAEyx10GDHaKf5MGecR2hkFdvgt62uWMB9gV5QyGdLuI9eg0/rr0/
fj6ty4+eiRN/OWyN7v8iMAda/o40FhbVwyZXa6LV8Jwcy3jM5WB8GYjRRTeJmbRJhMR5Ns8cSYi7
T2L26IjvEBcKj3mo36ivmvj5WLr7FjRshtvCU4aP/Vo+sGc8/n31kbLJa0KAM8rwTgaNdBgTJBsy
32zYLsTOHJfRBLq3m2wyWSE02LQOENEKKEkxE077jZOlDiJ6wWE+lCgZcwgRyENMUwr2+Ou7Z68W
UGjI2MZrXxohJjc7yVC0eAGweh/C7VJPP8nIKLYtziaubP+CQf6A6R4qjsUvtNIyf6HtdTy9GeCu
6faOW2BpnQNOYzOf1OId6t5PQuPp2eEKBItbf1YjBtAWLnyI3b7WsbBXLakQ//LnP0EqBw9e4aVi
WaFRAzLKVDm7QdC0kbsY2YbGBj7ie3nGdcEuhJ5nnAkpDFZXpfcPDgGB/CMJCMLN/AVc6jxq68Kp
RoyWuqomZA0ow7sC88Ce0Nz60tovdJ+iPLtHZdbOHxs1+RTxBrIdEsDioJ1yzpFX1Mzjxu8lJSTG
Hkp6gNyEJ7N8XjmrIe7GmZbsQQl5+yv40YGbItU13pHbWQWVeR90EbnxU2RJ//jDYoLAJF4Yrd2k
313ROHRlmdLyQ8va51TsrFbtYUKZ1JGWcOfrVTdCJtqfFv10IZEI3wnB0UBBVj3ON5ISNIl8h+/I
A1+RPeM4Sc3lwl+oiny1v+ZI+qiMIBGcGYNMAKeZnblsDuMf98ZMFJrtje9gqwgUhGBVKnV1jg3a
TMwJLE9fet8c9J+MYuwxaIfihlwvAq3lsXaoT+9h6K1SXkZN7wHFEx+Vx/S4xGLUBjgNoqFtJUyx
JYUbIJCSWROsZ4UobEHfJjafSXKg2PK0F5VV61nkNU4k4sSiJsTmAuSKCh6WODOzQNPAjL8wfH80
9/vSeKkTKreR4ilEIsgFPJWSAO65/G0qOhazOMqSHL9WA1NkzY3+EDC3T4y0akpV7RPcc2ZuomiI
Kdo8AJtiaJnueaDRwzwa6y+IX04wb5CsJenIAu3uXuzmVKnfvrRaUWWprGwQ7FFqUm3MGQKqzBrL
B36+K1GeQekNveMhXRCOLqFbIpSOsXsl2C7WvAiWPIpkF+JbW63RAQ5qB9O1+zH08YrM7uarzLzO
TtmjKnXt2TF44auVBAN/lXxJ/OJFgaFjTGE5AKgFKDEwuUdrlhJI2AQeqbCFummcuyHGOLy9qEjo
URHZEye74k/n6LsfaN8nkB5lXHo356+hq9rX8lzlvw604BSv5te9o+boQmZg2PudBz53x48Pu3aj
zpGp9pX0o5I+Qq2KvX7A2JAGgGwS8BKWWXKKjJdzrXDjzM8v1GmWyraB8ReVbBZv2S8hii7wHdBq
+i+bkMxeHDpBMtvvtM4YVL0gLiLvdtEIQiiL1Z29QgdaSvvJLmzgRUfEQKLh1U1k41+OEr8Fq8A+
1g00BCW7aPOWX3jdNutbwTX+62N3CWHPD6ZWdcYmXh+tPYMBK9JIh1iS8MabFV+MzQ6d6PUXG7aV
k1kdsH8H0xClEMgFbIHU9mEVlX9uC5gl/mf2epG7jsqr8IQ5lE9m+E6cODr44IYxuRlhF0ceAuo/
xoJ0mLDiU5ykZ2gzFL8TGebDKlnAiBHZoBnLvfEoMuODDsTSlJwOu2qHSdpFPc3xMEUiSiWKghtt
t5raxxnWa0LqVe+vQxIJrzk69///NAoM0jmifmh5dTzg81C2mflXIGMUPHwxQNJ2RrWyfWSEPrnh
RRA/AxB458Y1M/v0bqxtJh3RNqwqN62P6cnC9PTFeEXQpprv9CAtH7Zc12iRofx2Z5qydK9OQyQ7
mLWdJK4agGBzCh4S7qFq5KOjNXQUVoily23aBqwZFSe2vjPnuVSu49CcZhDm/kPz7DKWHeoGM8LI
XwS8swkd6kbwr65SnPfL+HhVS7DDbRYohmaULp8rEY79hDeJYSg/eIzl3p+o6xD/dtQtKlJiqgDU
gaggECG2TqErsVx69Dtyt3n6S7rt0EHp/tx6jyvFXSawKHSZZdTb//psIbRCnQj4GEXoOVh/Cf71
xHRiOie0JpGqsLWA2HHCXYZWw/QRhNWIxPu5+0w0W+lJdGzo0L0LV+eXjvPp/Ea6UX1ywQGLkIP+
PUU3JgMK9aYafg2dmalRLPJL+M2lBWic9bKT6s2xwSPPzoA/lEy0d12RAAqZ8qBBLuq6mcfKsq1p
i6XKaZw7ji+Vm+BNC8sxW/pQfNWT1aBAx0LJVshjK3ERzF1NXk2pJW7aJ26QDgqX3wL5enhdbSZs
uJDq0yeTZOmr9hjT+it4z6JvLDhTkcvnvXZaBxfyjt8ZCAXQBIBxC7OO4rs59O+j5PkdFeNUX/by
pzxH32p/LWr2/j87MxF6cVYWWIYD3u1DSqpqCmAGJ7fTsO7LpuEoNZJld38pq/0BGZmB5XtcdSZi
bqXoTuhVEdLMSWTMqfIpQEtSH2r8uqqFaoKKRxJ74CDXtwljRCPjqFEpd0Y/2poUJXG4E39I8YBB
Vk0KzdxHKvUBSUJJoeSJT1XDPyWgClnmL2FajariAm8cffXClLjO4W+KktkWS8W4g+haTiJI83Az
gB2xJkJY/qW1h0o18xz/4Vj2AOO9Frhuc807HA6BUVb34bcrg/PxpYVh7FxZb7iaDMNV8QL3VlGW
pqLd/Fq4EA5cq+lEVBYGswM8k1bMaPSu7YC/ERvBEILa8xBFyBTbwenT2FpaJgB+DoXwx9FmbTs+
XrnPGiA9J7vuqcr5XsRDy3FF3BEw0OLfvhSp07UvTm1LO0uV0v8F677Grn5EsIlYuPCA6M8kPa/A
D2D5rpROMKoyMKp7Eb017vNWep46SlSjt/ckKJisdnjIZ8nyWfiI+OkoDq7pAMBth4RZY9hwRPlD
JbnpW3e/ucsFts5qpal7bwfc/PYywOl426sWIFdAMG7giaGuYteDTNHNNumzAq9kMiVv2Glp8r8i
KMH4uu0zus/J/GFLBNjMfH7kXXc5ZbYGmOSum8Qxn/iSGEfu+QnItwFNVho7Ialzg6k+AAxKvmDa
Bd1h/b2u3a9E8SQt0vShFxAIeJNXWubvUtmMb+xlKhl64C41M4YxIekllnLIyBYi5c/8cY8CxqAZ
1WGUIuiUqtB/QHagsQLmbuikWRDbbhdV2IKMq7ktL9ZDd1/0yPWOInzuH/tRzWPD0kcGnTdeD+qF
j2uhat1EMjhzKzjgwXU4eObHlRgFdxPrTLpVRqCg0lsnFU3TrvV+XtnVJAfXEloYh02y/TQVoQPv
0opesxci4z//3NyUIl9BmDdxMyU0uvr0iX36C3LVhlThTEKVAtBSTUCCF9Oh1ohSqMk0P4gXzECT
06aXPCQ7Ufpmp4cjcT5BAJ/zKlwhk0dj2m5QbEkCsvSbsRzuti2fJDiGwjHLs080mOo288+V33D1
PUE8a6a8BVHlpdF5M+JNqeEdqEcZ3ApYzSzp99GMrKijO0xqkdKMTn7O3Bqe+ziAcJC1VMyEVjNt
zs7eNxzzck6NFziqDBwuSVnfWzij6yW8XG1EiPC6I1xEKubi6bL5q+CYIIKYIuuBdMb/Br2LiFnM
Vd0vZXaLz0/GPEwgVRtajJIgEBurXZohQITBijvxJcSay1sqI05xDcXKx3EfCNtmTDwW3jH3zhl4
S9B/EYoTAwdtOO4AGKHN/+w35VZR0WYDdde7NORINLyWleNE+ODN9VJJ2dquVO8LNItvbCi1KLOD
JJ61eRyH922kCgrwbA0ef2GQYxTMWDt4YlEXeWDEjkEqkXnfy6U1pz1HGC3MtNmoqbVl1eKqwq5l
lcVRgO7m/J6eir1I+1czfCcVk+7xhPwO6SoIgGw5EyV2BFluVZQs73GKxYL6QXYjwHQOMwactlh6
yUhb5GTjCH/V2ScwrCfMM495veWSy2LQVhsytfLeQxXHNL22aB+VH02wHdHbqD7ApZRCd67h2Yl6
8rr3l6NIMwcoPUY/WcW+nxOVgOLnwbLuDf34JkPL1jeVpPLTKon7dX+F18p7fVBV4F0pWUXp8Qs2
EJcF8sPPGuV+EJ6gtZEw5opCXbu9OEJxxDjWovFoNjFVQMzHhvVHL7aDHXP9uxG2h14D3kGUrZMp
7woClfmRbOEsx2avOB0wW6NX3JD5bqWEXQa8BYoFfzrKltzn/wxzSSAM3VdT66IKA2YgVGkM8zgy
gQGwGEKF/ZT8UrMQD9AaGaizOZX6OOicgeOSlr2jau9b1vlF+2U0bFOBlh+n5zpTe/qGj8kMWBo8
gqCEWQGF+1Fk13d2x5wv8qw0WvACp96sE1TZC1Ya1LzTUIPy2O9rxLOdjjGhZvrtimQ80PXt6F+f
UPp93SFmqF/v7A7jZmSZOZUF0/+lBrFtuDZP57+y/jr/Purzuyewxv8wTxyJ4Asc8V1rt9e7Xggu
zc9v+xdQkBe8fo9N9LaaNfqLyJyw9/6Y8QLWZ0mry88dMe4kvTrgozqLZr7AhFVjndQStUCz1q2+
rcHEkMrrv4zLwkcLkfddNbPXDoaSrozPYpwiwbykn3CMNB+9C7TLPirXTEx3ki2EErcKE/zn4qT8
pWTXAL2htXzk0yGMc9eO+4HmoPmVMwSP5TaXcc+j/FE4FfdQR5i/Iky47u5M+8IevDTdxe0Nc8ep
OQGzkiMOp6Fl7LECLgPwMbGh0m8HEkTiQUSUYYDpSidTD2lITP7f8tTqTYzMyzTa6XnLMaIs4W3G
QPKB3ejmp5jgDhL1KnAx77v79PlF4lLEdNyeHRpE+ezB4UWLe8viLiCr38WCaQkVfpcZVfzWyfgC
0+ENBuDWC8bnOOx6a5L+EBPD/pWmHuk8iNO4DrbpH5G6zas7Xmniw0sMRSsQUE5Kvm3WIgoHo9of
RiO/FZuQmRvMM3lweU9VEB0EDyViiXR0H8HTQ2yZvaOjRvd6fIevbZPcHIKznfv2vedAXd6v+L3H
dQbyOMZ4tqpYLGnvg2xK00bM3UvDCXtR+2wLnFquM9UM7qxefUJCZy2K1SxgSTet0GG+2PqIJOCK
MCiajZKxfnNoud2FjUMVXpNM6Z+/ZMamQm5G1fH6p5xSVvGd4vR/rxUxtI0P5BskBE/THIY2oagu
4BnzZvLP4OnFS0F0KllPdE0HThPXZXYKQRy20fgfLgsBkMRBTj9RvQHKs2l2GwGsA4/Zg32U0458
THSPcpL5Grow8a1ON0vLhEOUU2XRuOO6wRcjssgDjqNrsIcUuBhN2Ad6+ivLhB0y9lBKKJIfINBW
7fTUxEOVbCW/I06mFUu4DZOR6OTaPFu1CE3MZCyqeDqHuUTXc2Iio0xB/HfsQBo7OVXGvuCpq8ob
BfladOprG2H/POpiB2pKad03AP3syoWO4Mkbp1bjqhzQF5k8opB9ToxERrk0U6JgA9YlDwhUx8Lq
7Qx4+Efa/Ny9EELuqZzQe8lqeu9V56t6UpZaFNRIM3i1iHGliZpbN1zwg+ExSQebWaD3KaTYfsEw
5SvMPClHycazfBzupHnVk7n2gq4oH8AlncK4TPM6sBJTRsfUscQrxcYAp5FjiI9lvRF/WpuY/pOU
nO4IjmQZCfnh5UyJ4UtdE+jaVTV/s1Pr0DwWTd+1cFhym8LflCt/ssLUr4Mi9ebghTMTsixvibzC
VxWZFGyp9VWo2ZlcgQrH/7ikKJzVl20Wl9sZtZzPRDFkQHLUyXrivJa5R2mXwk6/x+uR5FRNT422
3bcIx0nsUkITn4QzRi2NFsxQDjiBQkDz10yCre/NfDhNq0M1U2koNl1vyiq8hmsT8AYad5oM9cmr
smksmoAXmD6+l5g5jwhI0nApIUZ57wbeanKR/Bwo9vQHVX9BReZ4GMxdTW6lkf0HAFDIwtZAkGrj
hAWGyoGlDKNbbvlkyU+NoRf7tqcV+Isl4z80UJvdPGZLUrKigVIVEcYznQBm/0cLfndh8xqOFIoQ
DTfIw1poiFnTk0rdGktNtoXPu1/LqF5RW6qwyUXgnxC5r6igFxl/77VQ6o1/dStXxTW3wb12MN/V
CgMDmzRf+R6/Gbj7ZA5JexHIASk0XGJ0x1Ydz/bJ1UT4ef2pmx+qHiynSriZdepJ5VjI5NP5g0BU
GfCar40qSWzi4lt+8lBtj1FDD/pRmUwiLRip5/mp2EH5nGv2yy85b0lFhQO8LQfx5v/j22PkbU+O
OzYScaSSDIqYgU7lkNK2phQQhwXi7sEgc47DKiZB3e0yL3sgjPPTxH1I3O+VnENJLlM3cAEyEWk2
YKHERyT+H3bTZjxfofbepmnyxM3Hn4rfv6i0BvqBzzfhw5fvtRUmQW2411AcyV8UCa0JXqi+SFtd
gpd/s83M9zyWKhcUep8PHZw/367P9V0Xa6CSOXJguv+rooLx9kZq3EeJKv88BELzb64aW4h+RNhL
sQ7OVWsx6UQfd6KMDNcmNkBAHGSsSl7f5SLGycTHNE/9oCp/B3NojC1JSkrFPFPJevYtBlKx5BkY
KBHv1NfMEtBdcIxjyLjeVRWVsw6E+nKM4YHBQVzB7w1AgaxaB9/OA6cl4Iaq6SO1ge/men+Wp0cx
HXZpG9xOBlPzfaQG882ouuB9vpdrfDI3iSYCNsBVQAA/SvgXU7DZugCqTbPBCuv8eH+yiVF3jrA6
5ezkjUo3KYJ3bzCndhFTMJb18lJMq+ijrjfTNMtMX/gFydeRtWpb4LXM5VXwMZ+CFVqpjUcCasdD
g3v33yTYNLzpleXOHKNp+71AQZWdSsG83J9tuo4GSedAi8dkuEYISeldaCfngnUAgSwfh/ozGi7H
GR0Hbogw8rIZX16SWoSkhN/kTWr1G56iAcZ9sAjq9oWUAL4KREA6/UZ2GkKOyAfxBEVDoeIIIshz
ymijKQmz96At8VOrDr2O9EKH7/hNTg2RchQRKzWp+fRuB1AgJG2Fo4UlmYLdsvZfwey7aoobiBT/
S8A9/PaLGfug5tFhjlyWVOp6dackbtS70WMTAvQSyqfucV6piAQejyyLRsspKFQ/iu5SW+CfPJs3
cYC0osbMU1nSE8kMX+DkMQMTpdwKNStfAmvT8uoVKjdwaLVF/UsczLjT+u3dWzWrI8tRQJ46Ky3X
gwOFs94Hma1x51qlwkgS1UGeyNWzEMEvDBPYqBFrt1rvkvzGXXbzpU+Nz5VCncfRO328R3C5vTwb
Vp4xOLkmEpwV7RX1qMpGZ4HEhtNrsV1TSrAXYyY/UY7OnzRzGyxvajFsnAnoumMzjmm1o9q6dbwR
7JYdOqytsENT85IqdBboerPUpJYVU/4hAzgSIR/8BIxr0+Bb65VEdrHqktafXBr4c2fU9tFR8f3G
aUE+c9DlAWyBO2+/VQbUrOQSPPQN4rTqMsvQcExGyobfgMhY8uiAYc2uGU9CHLw2yUQNpqIgrnkt
LYa0td5F3t+kKVJmJvYpeQwBZP4o0J3wVCkPlOGEYitmOufNKW92opjY/7NkuebxbJveohVNd1ws
1qBWFUPSU1/M3rPs/bJRoTq8liDhKiR6H/CgtNzhpdubzrTJRUGbR+md5IbxZx0GTQq2ujLtNl7P
KVASOO0auycildwo4BaHqg4IRRsWnoItYCJ44HumZEaGqGDkiQKNuQahf+USY6cQAdu7VQgA2yqP
rZqoc7BeneyibTBFLkJH7up7CfZN31Oum6J03tQ5a90I2EMXo1znvMTsewVfnYhATvyUB5lJLU/l
gYd/o7QAsaREbKZiutkUMNsTnMrlqgchu7BcRCRXmFIKMdwtiKFDUEUhkXT4ORtX4Yf2J8yrYOsg
ErY1//BUVKO9lhdWeu7yAdeGf5ec6NWzvlJS9S7wtQuawmm+iA8RIy4Rrbl1xamGVKVqD7HchkPP
C4CRsfMazZQeRsb4kG0oI0ZWkgrmbe+WdLydGF8i3zQa2A7XLMRbKt5+kzO2TaDEtDC0dtF0hoCi
QZ0cSWfG/Q8B9qiUBMFCJshByWHz8UNzRID/vyGvLr5NEh0huPP20Mz6XCp26d9WAilrQGIUm3cy
ItVXrRFhuXyBR3mnkEH94oFcbN2gUllvcB70aXJOYzf07yVUZaHIMNiXxBsnV/AFOWLjBfEI5avJ
CBhWeoBt5shfNHUTn0avd8ypO3vh4c/3IQZTqIi5R0L8sjO4dkvW+ow+k20wtiXNyfTiW5wWeV6o
hV9qh3+8DUEWtiZrKAPR/9ujv9jtQMfSTGDqEEvtoj+qb+y+8w6TAH4Tsp8U40NgCnVPPzUSRWxW
MsB/NVY4iL32m6bPVmyWbvwcB6Y4ooelSZIjjqNbirrHvCwSOPFetquDTKV/i+jPTYGe5a+M6jpH
sAx6HGg1tkur1dfsWxxps/be5zHpEnjJ48JTfjY23PLiaRGnF6Kvz340C/H+IMQcRgqZaNVpOIov
HIA+tieRhNO9fVNEWc4HVPu9BAluhf+7j0UIV7rPlQA6h2hSAU8IqlJtUg6HS89kbhgwjwKv4exb
72np+9o8mu5AZMcRhUD64bPqRrU5askeNOy5dPo4d8ThOVeL716xWHyzNsyzbAQIJRr7xDfXrJPO
/ALU9THZKWdhzN75s7zSGKVJJ5NhWuHOMNCaCjV12zgwkqSsYDu3B/jEhnXln/9pStLK/TSRes1Z
U5nWXrtRwwIBtXw3TZjfu56Y+//pBYoQ4DTnsyCdTWzKaUfNwLZ/XR8TR0qq9d8Co71yJfmFvwnA
SBPAQo/cuNtfqR418cqYaGV8LPP478co/qjUbkqm0g5867+rZfLDifDAmKDOSwW1SUsMmupknmBt
783r/S4foG6Ex3Nccr/TZ5/RW6rfBPzL0YX6MdnHSrPMup8h/RegKzIi78OMu1AoqZD5avF43qZ1
ql017jgIlcQhu6wSPTxUkfbgpuAhgip44K+Ekfh1qemM8IMsk5l+eXmhYj99ptY01hB4OgQN+ImA
NZYLk/h09L0lXPIwKMrUTITzy2jrgLPXdjvEnTEU5mDrBzFtM0pvX5rOZqHG63hGW1WV+cxkYXxl
MW0zQT57pomdaM6kOkonzg6KgcN2ig9PvSWDyutB2w3LlmngBNrUils8HeOq2ZSOQNHOLy0zB/Jx
DuQNumU4re9aKzBHKSyqP9idMjVuX228acsFeIGvcIABSUYaE3oEn4F06NfoMZafuGqyRTe18LC2
Nb4nGT1pol1rGUPi4zwJeXV0pRx9Mb3c7UFHpoK2+ilorhZkz3KkYifs1eWntyCLGN1xUXtYQ/q5
jcP5LnCdnuPitQk6gZC1c1MfPV274qjTIf9C8iA6KefiFw7coSg12XymkKyNPaxr2Ef2h13eF6Op
VFyfzhB8YVQdR7Owjqbb5nzaHHwDg2mekozhCvUW/jnnmR+YmdsVZCGBDUSdgfclWPqJs3RH2vqO
lFVxTm56NxHcNywbFQITYDYYVxcI+WPT10y4tD2NiFP/g64wwohk1TS4CYxdrVlEMc2pPaeoX5kU
yTlkpuL1HO1x1azAphtOisIAsvRCVGtSqGHK8IJPpN+9GpoJvjdocnwWf/y3YXN0Q8mzh10QKuw0
OIR4iWgLLxtZWj/ad6jJHtXs+tR9xljIPOffHEkiwQ9dCvVHMO61VAtHeRJcVVhv+kKPalGbAw8u
60fEoENZxwf+pX0Bmlz3UybfOfXJb4e/gHHtYEnBCGcYgiGXY34o1yHIPMfokRCM64ImC2FyF1La
YgfusWUseEAlSSqJd8PjA1V3Ym/SmqZghLW9VuLfAEY+uzGcXuqVBkn7GY0H7KsKW1jYAkKHQ41b
0NLoMZFwNHFAg9lOEp/DTewJVT2umwlWHDGmUSjMQPbFXE9jH2erL5GniZ4YXAkllF4Jtw/5ARZY
iNgVqeq7R3+xDe6nrEL5rhiupWi8elsxwQhabS89jz80kRqvO8EarZgXHYrD4g6Ao1/FD1+vF+bG
4iLnvdjDi+n09MAPxNVaZMydYFNKLrYykZSFaAHQmR6XPcf1tXQ9UwelD1GlSTFxCg79ZbSxgDig
nw9QtYn7OaqFLjWehSca2a80HSrxzZZw0s9GFHtnsjq8NaZpfKjUkvWWnqVf2uJ2nLH6mteCrlw3
ahhHbZ5KByp8azpu+KhyBZ9FzpKgr7m2W94NPoMkCYoMQeRu34jHUZNLVuMAY0Pi5zx/p5HFqAQs
gwQ0TMOKZyirPkYtBn0DrIRhrMYVjttDt8OscnrR0mWL7FENKdZJ+ELbt5FWQs0z3mI6nznnrl49
9jkqx9rPbRJaP7lHAicDsDRD7nP+gELx9HBNV9dYn9g3+iDgFTqHiI6e5xkWaxv8OXeQ8WcBq4+b
92c8QVTgz1yrP5rXJZRCISP7rd1InKIHiEYP6gMBD0ttQpnsZL/133sEftrB2hOeSRk0rInFBDGi
oCQMqVp53mziSXn3QgpTBQ8s+wu3snLPlPiFYvUKmPgFLVkJadH9x0nddYFzPUc0mlxGmylSqjfr
V/KJTzS+6I/2KKVhYP8vZaFz+i8AAlkBwqp2+fkW/eOTFPeH5tnONFVcMc5G13KhZpp+7itZl5XA
1oOrRNHjH0p3YjW6FRUL4UpW2tO0co0yo3SDyLE8wKLOOZoR9XmA+AivnPyXKA3To+s0klAKa6Yl
CklYsx1/dLDA4MmY0y7LNM9BM5Wlll539UWjMGV+79WbR9t8F1m1rgVf+Cs7yoka38vl+ieUdSnV
4K5rxcyCEp+FcQ8WSl+mVwZ/451CjdlbMuGaIKWbs+OIgH7dM12kGR68bXHG0KZjttR1cECMb3S/
/5RCt8G4SAaMV+S+k6uq5i80iO2rdhhj1p+2I49yhSE5cjt4R8TA1mB3vhEWUA7g9qCUZdcMzEq8
bHhY4TQiWAipsrLUVwLxSN8hBelN5w2ERwSrSl1SgYSyOsh+UP3/qfMuYQzwsmuy4DaNvljyE4yg
CJsL/cDFw5Z4L7N6YEAxRFxFbg0tFl1SarFirj8OWLfzB6dLR4R0noa5saF7KXWcGFCJeAlQ7WEI
CAiz1RUFosqeBedUXm3UYBYyKQE6Qgjun0Lx/ufVt9F3FePbJ9Kct/c3Vit3B2a/1H6LxwF5f8D2
lPjSh/RyZq4fovRJGIukBaTtCjYQjp9rghc5pnWV3ydd8+l0djPb7yNz8HnMWyfLMTIyY34Lxj8h
6hQW3k0m1e2RqbC2aUqMjQUrROiHWfq9dmFmVDjFU3mWlNRYe28mXmfKQSwliSN3YPuhe1VSYjgu
/xQY2kBUc3h4Vy7PuqQqiZbYqaC6ZYAVczxPyOd9+eSlcYaeCusclREGiO4+O42/vC9B1W5G3RDf
f939/GXWB+W0Wyq0CIuMK4hzlsEtPzAw6zD9A5uX60fSmWu5EafM0jq57LWIykauOB8SqpKESzlt
r+wQfDLvupx51FuWtRACjyOLNckGNsttZMQigv3hkbIPuvSPHbflM09HY3mO28Cn9vbiGQPgz7Qe
tMWlOdz9nxkYNIi29QxUipdArty94tBn2KmeWtTqvarVxkhWbdgnhjyvxgKxcYz/REHxqMie/Kv8
2YPfvxQU+yryYmcb96963+oNvAwT8gxoEAKyrVMxpLSe56aqD+dx3TlIHD+AH0NqsAFz72pwHP6c
koJHwD9Y2lMD6dgZjMQE3zHY0LzKjJbgCT6r7OdCI1tVVed2JI+INZwTw6mtYXOAvEt14zarTysN
0W8G5nFXsvTllMCPLXfgiZjv8T64BqBRZEl2K+gAmg0vlvroBhgdgh3SJvOJU5OFE5xkbN6GS4VV
fbbaWFboEcTK9Y69ruHxRLwQYwBDEhp2E36ORRm+i/thXrVxX+vm4xVsTfJufOwaHGeetZttqwyW
Cmwz1/CKVifrXuLEIyMQTnFVVaPAP3ldJyXW+dXbbc7oEZ4vNvDis0EXszdDCof9GYmJ9+sBAYgC
EZwT9EBd4VJdw2wjVNVl9Mc0l2ze9NamV3VFOR4rw8SBDS6Exy3gmWrrCyI8EHcLvM9sHLjl8dkO
BcvZZkjxr7ZB86vZnyVcU+JEY9W8hT4zdO+3TluIBJaZN2EJ11Rg0nmo2HKuuZFDjfwJBUKxrmUK
pcYkHO7/PQst872EQC2ANahvQcKZ7M+UcN6Sm5XTZkyhBiZbPPZqOWElnWzNtqdA5qtVaxQ/wgym
BfYVtF0qwYmDPoXWh3IQ7x11mknO1QO2ltdbzI/iMVn4zi//8bSjKClzQk08XB0GIHVYRJOYtzTc
KDpgKGtHJRos1dn8YMoemVYMoVgDGBv0e+q6gYYVI2Uq6GdG8myDevxMt0JeA08BvjWvlNCtxQ3G
A/0hOo+WkqLStTH2j79dNKMaRJAZermD89t78EfAo41wLUmz3y7JOkpa+ChZF2TcHUi/z3MFbHCG
OIb/nFgam6mZSRAUHw/Uwx+75GXmuPJQfKiqgdp5cdiY9YWERoKfnaytDfkfyPGeYRk3MWFRycnL
/xoko6BUKAKOtA+nbLbJKj1xhOfrqPmByCWNl86WCo/jKBfV8eiU4ihRuSVXOj46lPgbmKPhkW+I
J7BdaXvxtaeL70okAQtOZAF3GpwiP1uEDIojksgCg1yDSES1JggBPLMRAiyRrJYaZm8UAeegOU0B
E32uA0wNpdc6Opa3rd6CNST6VCfB0UTe6UhG1nhN7oMlvrP+hX89Ebh7mKdbVIKfit0pD9hufARH
UC7lE/tBNRCWSqUy3JRc8d9wYqKJo+QQ4yDHEg+Mbw0WAx78hi5dllpBEU6OvIa4cnMAoFSLBy8n
7nMcb+c832O1goebCqKCROZuqCX/6oKSRUvBn2qWA2LhYuNxNvJeBW5ySN2gPNn4ADPUmTxzFBvp
8y7vGivFMYSu8Gnn9u1R1ds1/HwOAEOCWDgp7svvw/XBaYzsLBpgoSI7fFsdX1hYWiEIacryBYGm
mtcojsrJroAfgwEihHOQ2fXNQI1qCqiodbpMSnVC+6LUub7Xx8bVhS621TrCa6SAxgKKxxkg4EEc
K90uW614fuaqtp5grDUe4PeAMUS2d0x6pFxQhB8x7+qogjlgdt9WEbyCHrX90QvmSpbCilj6ojSJ
y2ygRhojdqpQ3uPvieyveZ2TVK9omIx6uLqgylUpOxfbJxrV6KWy6dm1NTAxaNUcjFcX4eMkv4aA
/Tbyz0RYl4UslqAYVWioGC/zKJ/v6/EgoBfU73VOEjOJo7Y12kt204t9V4okFpMW6xNsQvm9SSxo
B2r8OUDMl9zOdSYC9H0hPjY9IHPpY6xwdFlnQTkrdi85ovfGCtEddUpxzsr2qLlx7OVZX/z846Pk
GsUy/31r1vpddDe6gjfIzjEMDDB1VU71V72GC0fuhxLlOxy4bksTWqt+24QmKIoLVuWdRyp9PuGZ
NCxEDwQgohzJ92r0VsDAVxV5rgT8EFXefXWeLlu0IEN8UKAzdr4/C5+vopM1gp9fZWNqrm8pEtRn
eYk7Gj+MI5EiUJAlx7ynwA1VSbDJ7Dk8Z8+zO2fjHsYxIyyHHVcdjQm8ZLyBHOMliBNWS8kqdZWQ
vNuORafHq1b4+ViY0HONgGcsfCSGZwXuaCouG1qxZKZ4o0fHA9Npo2JG3UIHJM8cAMz4igau1suW
/ZvF/nFXvEdevvqz1eKCFPxo6VtRPZsscpvVz0UYIvkDCIGOIaOivj4vs18nXIWefcUSAURYip7O
GTRe1H7JiLx60JH+EHfTN/TVxHxLoiI087+3egEeiznLgiJpOGc5kf2g2e5EMad/0CrxP6qDS2XB
vrMemoPmf7FkcOBMj/BFJme8Hwc7hhWDvnSL90uHyikqpg9MToEmcx9SpgvuqOnm9U+q7bUesN89
3RF1FCu33JIKko4mksBYLv5vUaddiP+ZKeyuu4FgQA1ehq0b6wrtkQEHoJDFgpdnaJP02WB+y0kE
t31LBcyFRwzNGiC+gS81v+XwG2JQM/Rm8Y2cQsiC1aKZbOyaEaVRRGWuUUqbpgw7mD0+U2a+Xy3D
eNmYEJvUz9G6lsCAcPqFFe3JDcXDWAh2qK7XmOZDh/JivvlisAvhdm5nI/WrFc0F/JIP3BPC1hBi
7P03/q2iuudZr2JGG0T1NYyIpiY54RvoDXyUGfsdYiqYNZdISZttIx5d4zWBiyCf5acyaYF+MW8/
vS0x4IbEGG8sAYQ7GNxOJ+2/3Qw/W/NjBNgGGgjNhmG+Sos03UEvUMFqiJs8H6XxtcULfSpjBXzV
RQ90ONsn1zBTJ3ELxUM1dORS4eQuDnSjRWAf9BPSSFkSe1TDqwL39XBZQ+sFx1L7DYytx25FqeEA
ztt4gqvf9z/wj3hAUpLG//C6tQgl2oGTHErdcjjsDvrO60yaqqkYH6VrZutxJKENA+m5w1ZJ+3gK
H0D9T2rbT8auES5asODLFGVveBdmST/nel6M4jSNBlUGXCYlwQmzJd2LhfFm1QPAmDX8bVOphodd
GhsnlDp8Hqn12+Ppzb8IAglGfadkOgde/F2dbmas0Hbqszl+0DgEfsHeDjRyrW3vw5m1zzz7/vy5
fJUA/1iWNdFUFXITZEZ+lwxhZorcqmjwJH8seY6EsIJyWPckzqGVSBEzmbZaI/ytXaH0V+KoeWkb
hrusoHAwD5T8a/PPb7+QrCe6cdDlGS6Ln7oOivwXbr0C1AomTZGaxKpAQ/gTFMm2iaw86V9Kw2PB
EOif1MxNnB/2R+Yv23r05jCdjYGm6aovq9DDRL1YwDE3mq8gT1VgEXUuNE74hu0y21xkpaSNCfDp
1Jo1SVtSztTi9csbRRT2SvmAhmiVBV5+O8hkpwy8yo8KNaA/0L4YSLrke22t5kKDfAGTSZFd791u
k818fWPitBOZ96DyPbEGrX/oSYcR50qgtyUtOUW1dap3m9U0qwkbQRg3Bc5BszF/fPNYKjQQK0Gd
f65GNZzsiMF2FP3FZrwcl7WVpeYOGXqL4x9t5Rk2UnLIaGAZZgyi/ON9WKdbhVOTe5UQMpLxyprU
8Yn0MIda/cZIPgriQR+Bbt1Q0Gw2BWhWY+4WSvrjF+bywYbZaBoQmhc0IKVsklvkCP9HmE7SP3l9
QlbkuDni8K38c26MWIMSJGqjHO4WZdEG+MgGAiaMBatM5BIUx5HF+pG4VvvbxJpM+ZEgm117Y7hI
Hz/gXvH/iv2rEAafdr2QRUAwrMZpXCu6bQOq4cJG4jiWFYWGQyfXUwMZ7CVnQkRI2Ye+MUaiXsdd
VsreANbtXKs/uRrW0sNduXOBl5RCovjdyipf7yVnJQwWQgFnMoJFSnHMkBJvJqhtpI9PUDOGFybz
3L79XRmvSBB7WRWO3wMfMcFzVMGKjcQ0tDirTsCyCNMSUfFDQrVTqXWEDZ/5qQfO3Gfv7Q0qfyH5
pwn0BJES7sd9kNYyfzl/o/y3XkS3CRNftyWhQES8IKSuv+seJW/v9SPV29r7qgyy7PTEgJH3xuve
nHFad6DyRcYwmIa+ot/GnnY24maAkt/kHB3upYhTgIgSNSZYqAtWKh2Dl+QN/+Z51jWHKNfWeNA6
wDWvrMoyanDYtn8qu404X/yBYLcVEwZxFiIXr++f0lzyiErpGHYB3woMS6DXtU/R3tvzJr7bg9zb
IQ511loFucGldWsyCUOCo98upRTWnmwgkllmtTsj2UkNejPCVCPb/jSA0K+JigAT/6BCQ4va9EVM
3+qhSEef/iEwFlwjdLIyax0fwmF+Q/Qp3We4a4JCviGFqm4uFkow7/+9rtidH3NTyn6OHQbH43uV
y2QRBuObtfEgvJ71TVVkmwHl9CylgzRLXYo3sCeTcREnR5emvltf0kvkgx2dIZr4DL8f9XkYA0ir
lDGM5Pf4zXhfdQc1laQ2pVfRJfZRc6gh8RIEVSlCsD2zwRikFBtRXLs8rpfKjMIOTAoeyNPnxREH
CSjl0BX6i8G0q40ZzlvuN5TYrH+bU5FYNx6v2ZIZ46zkx7qAa9Vxmv3TF7GcbZFaZMb2gnrtBIAS
teKmZOxUy4C/1hvBWPmqdVlFvzFnopv7Oy+Bp7iY7Dinmw+zg/BeVKCOWNVM0AxkkFgQ2tAHYgDx
32ucE+VDtAczzcDsG7PNdjG6dZzn9gEle01Xj69yRl59BtxAa5exz1nvcI2vAlMaGMqY+u0uYXfS
N2KV03ZWeMU8V37Ar6YlDupT8QxsRuT9pLH7EvnXlM1cOIi+ZBTR+gmdSR0XVlHyTy+OnP7jvqKH
HdsviXYohnA8xagapGYO9Jx/v4B7jv/UCvZUGwRtGK5ZtQeYMRA4L0Iuykl0JAbOfxtbcTRK7KJP
enm06EjDN3eJYKBL4oFO13ohT6R4qxTD2fPu+dKV3CWkuZ2kh6aR6tQg+ehbJgF0P1I4sRRHJ3kl
CJ8tWjIX0TnG9X8sIwfuStyp4PQ0J8mmLn8QraWLOHfZEThyM34qQBx/ZitTcwP0B50lg1WKbj4q
/a2IiPSLl0VTFTMKLAflorxQfPhTkecXaWkXrWNUBqM2YKbOL6GRsb9Un2/FNkdnRp9RERCrnjaX
UqAJisoyLqcQl0r1nhIpidb7mWJfpHe7vCV1CiPwGyQKA2E/PC4JUnTbyiN00rhmZt1N5Hi7sN1c
3uWVR64T2IRlonq7ZPzuhoWTYVwUC6kiuOBAj5By2qEAvOsfgwjBGeFgWev6P3n4qRYh6BVROTAn
ZlqmDUku5eTunePMmWsrnLCLly704zW9ngizfgRK+m+G0Q2/qhW4/HX02r/60fStBxYprl+/QFPG
ft9WqLELNlmy5HD2hL6ihqCq8hWikQKCcE7DcWjzr1hktrH4lbIV/LHNhbki4XgywixOTP2N5VuT
TLdhgvJXfIBk99y+pwDVapa/UZLKnAXkTadIztPXFRh3tOUJBT5XrdS6EpqqPLK8NC+FvYzSkKBr
c9IRa8qcDxu8qaHZQWnp/Tw68Me6tEGtPWCgsKguXjKqJvf71V32GAUCHKUiU9xkoh7v/r2l921p
QdfxtbXcxbROZ3xB5dtkw96Kxy2VYwu8MZQEqhO3lb92dWfW5CsPm52+Yg2FyQHHipc6Qri6LmpV
L435VFTIg8n53Z/p3V8LorCrUNpu0RwzXV9JEuwJGFq6r3nBiuySL9cZQnCBMak4OVk6k4ARDNVU
pBPeVzD0KeuTR2eQL+C9QvWo0CHyvd2/uhO/u6mPSozT93QeDGLobIaFYansxPt5rztK6ppe+3dB
Np0xqUKROMBvlMPAachgC8zvmUsZClmWn0NjjkY7eWzh32I+LN0qa3NEfcXzOYkf3joI2URTqSwO
cboNoNOsNkWNUxlgzfns99f5aAMLl7PGnj/XKCXX0pAM0B5yw3O3iC6d4a8XMPQ9SpG/1BwFmCa4
WO92OUWLCsfQTrH83/kyqywba/uJKNc5yGLbsDGK0Gy87EJOfPa/e2N+/2XWsZfEQp74JohEd0Ou
amgS8KjnUyUtuATMxEBcvHnRN1i2JxgEuBa1ySDo8Fn5BaSQazrIO641lQcwhxAeFAI92V5SQUFi
udF8IeSssfmoDvn8wI2Dcv5d1QBcqrhmdJW9C997hQfmGAq96vq5nTpuI46deyhIAk6Kuk5kt7pb
ghyQ30LYFmL9kroaQ74hCPbbj853Dn77eW1U0ct53nB15UAqpGxowkdseqvr5lIETTfXxKQYJKOj
wRzpGz+CY1WueqQUhDLPgrhLUMr61g2z4+dPGVet5i2mzRChOeiDM0OS+v+Q75THQ+R/MVnCcDkP
H2Ss18TB8n8BYIcAExougK7UI8MmSo8u67SbGcqxC+3tkZajozR0/x50DtBvlGaQ9F1s86mbdjxE
0Ja+sFMeZOdx57pGEaMOH9vJQpZnBhSM3i7Ti3gCPts9MnkzhlUEst+ehTzLnoApQ5wv9Yv/rUIk
RjKDC4kCglA8YKoh+O7EiJyCcz+6VM4eufOCIq/07Q9ebqqeJwRmUWU/YkKZXZaTEi8t0ox3NJjc
8ILPEbic5/Oivv/Yg7d7NmiU31MdzJaXeWzA3zDH4ruCzIT0JUCW7e6l6F3z40HqVmn6u5zVScBu
ThoKMAd5Ps/yyRaA/kNBjk7qJ1blsJ31pOuEeHApVdupy4+efRT+8HuEghA6aHHVBnmHgJ5Oq826
iM4dbivkt8JL8tHbPbk+uUymkLeFYouNWxZ+2dkRXrPOdiyGqoweF3auyUvgt0Amjbs5ThjmXg6+
+EnOiqmnvntEs7DlI9e3lJLCG6NpsWUHbM0SBg+J9hJbBjcsvBp2n9qjFt9Um61JP6BJTAJV2CX8
VFhuEYANFoWYgVjEzdNie5YDeoApLMDuNYP0Nr8IhYZkckW7FWnEG1+77PWwuLR6oZcUsHid5ZYP
Wgpyi4jvJuwwJfMm+x3ioaRfhy+P0VPwxxHjs8ZSHlw0ThRCMiNhQncRWwe7vxQ9GR7WOLXDIEDN
11nSjo682V3mkh/4wQkWRyyrAW3Kfm0zns19jWAlglmYcOw5RNYWHsnnidkMv5uXzv27bpSYqusi
pXd7GLBXBouTyMN+LkyJGqjJqFrmCn7zYDBvVMIzJ3P9NnDUhS7zxtQIVDkfOHuSdj3mFfSen5Fi
G5P7TP2lbJYhxRvta5/ftbbwtZKZwtoB4400sNFcg+gez/BWL9ZCgw+b12XaS/2h4C+9vyTon6v6
4EJt5LCdCU3xbmR7yEs7lv34fIpkoqBcm8t/D5xtIM+hN3+Bj87aqyusHYSH/7KJxAT2SLAw4XWP
1Pg2e5R3iZZWsq0xA+6o10etItTtDo7U9qci/3R6pUTkfoORgrj0NEWuP+l+oE6jrikFpNLaNCrR
oHgf9FpQjsPdjWwbVs1kPLyTs087h5X42/lrZWOHjSn7C0fB/g8Bc5uDncLBf2pWAcK7PV4m+fLj
pspwidN35cAGJfi369LYa2tZXPXPhwGHJzrfHiFfDJWfp2snEGLGSVLkEfqMP9QWSH7AETzlRiOt
Z2xxiCyy16RMACZlPjH3vUHqGhjrtRgUByJkDkRT+tLlSLfOREEJqYrkUc/OYGO7gQkp6ulDdQOT
/bmKTm6tGc7BborNwyqy9qHT7/E/+5wgwGg1Qbi6RVpw2FEqjW5vgz5E7JPBPl7axdfTaoDxoLnN
UY/FvwWSZRfQ/YYWP7VCVSR5uC9qq8AoaamKdAxAh4G2kddcSPkKdErqiak8AWXo+SReW81vlmUY
YajZIHXZfKOMSfU8lYsCBvQ9vx0JTob0Aa6NQLacB0mFFuKjudFP6re0Uf6HdNO5vTAPQ1V38qH7
R8S8Kb9xEItAsFlSiCxzfsPnNvGSZVtdFUt5TR8iK0e+jEPDSNgxzCxTmd9RJ/7HJlDHGJdp6WzX
lxhatTkmn60VwQjBH1pI7N7NV9HncWaOu2EH0P7KCzqcGzj/RxW+YH0vw2zGPuk019MPOp9qciHN
bTYwqnRd4xqKnUg9+CcRmbgHpZKk0dhiu2hL195ZA0IfMuBAI8KXq4uK3iFgy+x4h4t1Rbb6NKyr
7wIn7RqYAkISxCrQiPcBM7/a1joogOjIqXO5yB4kPGcA0C7oqV92McMtoHD/sL5+qrePB2Y9DbsC
ZF2+w/BbpLy0ZvfxtlFOB1jMhFU/UtK1Cn+QYt3fulMFxNTOFTinUUoiWnHTpZcB7FJ3PntBIyXq
bzkvHaAhZHBHR2Ncjc71EaJhfdquxTDbW1F0LVxOwoHgk33VOVbd3LHHgUocxWTadTasbBTyiwxb
TTGyeKhoGkkigrHlThwhrn9YLnXpaBlu98S2md81IQcuyKBANE9vARRZQVIOEfutJzwfShq+DZ62
v5LgsB+PJ/8UHIwRMfOa4N9WRuFtaKdc2WK8HyXj9aQHP13ReEcDyyjc2iXxWVF0OiezsCq5jXoo
784sGtQSnQUn4vO6JlpT0vFjfYJdwx/VvpQ5Zmo4qJ79OB5891IeyzjmBUCv+7dMxO6pcCGEMIZ+
Knr4tmIPgXHATaYTO7U0CP2mqIMq55U2Ckly/V4Hk/gsZo8zTPmjruwKUv7OR83TKyLq7Pz9MGKR
KJTm2Bj/MzqMVAfasttzHScCXJLgxX5OhR3H1rrGopA/lGFmZO+eoYb4gWA14Trtzlo1VRfQmPgC
UgZexaGljcvXlLcDliwHM12yk9zyN9bS2oVj3zC/6wMXAHrke9fMO9YOrD9PIaHF8tYLLkc6Yn5l
OPfYfmfNUUOnyEoLLX+JCYxw56nkheo04aUHuoVOgNezAGdA/FzkhI0mNtwJ2ksVdVVzCvlpsgCF
P6cOzZC6kE5ZzBGbGIXlv3QBiaGx/M333cR0wQsAzhZ1xCUg9w1aNT0DW5RAmyQmyQhCe/EvRNIU
amwJqUMACbZQPGt7seEJeXcIms4GejkOpb/OOHGQH+IuC2vdXvYmLk2QGsTYLqkOJv7JaNjT6nZF
p8QpkqzzLktqLEtU8tWDq8dzGc/ddx/MeFlTDtBOq+TkX0EAAHQ3udx5mycNVHk3U9Fbhov42OBm
FTGYhJLlu+iYcOmh603aEaL0l2gimbfyDKlLrBxU8Uky6SqITdq+xll5PFcl/VFLNkWR807qP1qA
bq/zEyBa5oW717bU7MdgSgb0pguD+cSqqemzXen0pfDsiCZeFT/ZtvremcDcT8i5qNx6IGWc6bHH
1FQI8IZvJZYqriMtx9wtsbOEyNkGzNk2kbGyJr7DQoHCvA6rdGkSJq4S7b/cMQTdtNL/zdcXuMfN
1TER6zvWX41xZQadRI9P1/k0tit4OHBVZPqOmpvfDIhTvu7R3xVjlzRc2Oz5H+DR8QPXI7BOrt2q
NjI9+p3KKClHILbquSmt7drcSPbOCdz/Ce/7TNopDM5qx9FrOnn5IDjdjBUfA+ynMJJgt0qY0XCe
P9gco00qA2TOiTQLXJUcyOEZs1CJ8sijq83bzD9psmAV+D8UD2Zj+RY3yaOVNYWj9xOOC5xLrz5y
j1HcQmNNSA4oMj7rcILDHoPOYak5+5/3L3AINvTG2xUyeM0jOL9lm5ut6xO0vC5A3L2ZQom0qj7f
imPK8fEUB2Dqf+SVbyuUiEvi4rbhBMAT/voV09U8j1kH2vB2nBwtBvsC5dnhMDVI/lFN7+txE91G
zd6oXt6JARBFq2lLySJM08gKntL6e1GJX3NE20fKY4EQYI6iwnbA++NJqjqS/Gkb/JAY3WRPAbPA
MOSBUNcZ6eiuw84MUChbRhH6oTCCDMCJjInKHkh4tJ8zl8Krb5WfGPNPnRB4cxdyD0e+YMbcWlvi
FUQ9Zq6GrVWJuFxv5PBndblXiMuvq1sZEtYu5RExkdhpGLjUxuEzRMPIphlYgZn9bx/mcxxaFZbb
NamiYE/WgVFFqPJ+dsga4S9MC3mK1AY4Oumq0qGIJmObDyGWzisdjJJo+xdxTZ9/YaMT6fJCtLXI
05UY/fTwQm13Xu9MAsjrw7xgBwMss8J5Q6Wiynf4cCiiotaclQDhe4OfRmXNYpBvdiW4VhhvpzDh
NczCVXgO8JlDNaGNqmfopCd4HxyZtN0uT7TwuE0WT8wT0uf8mTj9dvX4kS5Fe8WVlQpa8/QdAq2N
bDwdo5WQWUch5FPTXjXMHrZd4VuTajpD2w+cax4q0s2XbPNlZtgbr7Lqhckv6YFkSai5SVS40YbR
Z7wQH7U9+Wg7HYjtqSeN/I4MI3tJDd91Xc746sb0bPH1bOqAA0EWoRq1R0fWBR3G0xTIM4fGiBg1
A1DdG6mDnpFJ9svuTOcbSKyjISaKQ9EYPx5l7NJsvSppyYrV1e+MQJDBRAimdQAVBGRrrXm4xYMO
ep7xbEJPUW/ftDMuQLWbn82gdAQpYicqaSMthczeMw2iRZIaGGjgv7kXgTnz3lNcg9la6JlDBktH
5Q/3dVDGrotec7xh59jr7m5o3jMC7g/eLKubfZZbeB2krwSBRV29LX1Xx1Y+BPpuc8nBFSr83nlP
XpJwv5gVf72iygszjJ+tL9w6MyKDWU9zVZ0FhLX9iBcvVM9DwpYndGpDKaAFVNXZOHDqGkqHtucN
YBbbPUSOLqLhIOF7BuWGgQ/7N1diHw0wVtkSAhrlKZKTRxqtV0LxDSL6YgXnqqlloN1CUI2N+BdT
eAJMEj0a6r2DZB4GCIJmI5ZIiqOXgUTnWjmXCkp48/wthzA3m5N04Ig2aPFInnlu8sOtIEkw+azi
mD2a9BhD4PXoHpXcsz8k+7RapjyhkDEIOy6iwrJuhkZxCj+3EXG4rqXLGiiova9MKly8rce1qWdy
pRRN5EKsgcm7kzIuCnTC0wkxjm4grI3KDNdMMLMOnW1JTBln3W1Ox1MBOOHUwCLg+lbWfab+ExU2
B26cbOeFUJ6ZlaXLcBVsmU7WHcJGhuxEFvbgC4t/Y33CPRPR/Hmb1ehRECdQVRyFdkB0gfXnVTSz
MR8Ql6MTEoECLZCslGJb2SDQpz23ZmzUusT3wOjWENoy+XDrjnwmRIigaH27hf0QSBn1UNCpiO8W
zx2RC+TZlrsimmTdtz0Le9whsqkOnPXCfRENCuBEDiVGmoKlKUDGRArvf0LK5giBstiKAiO0/eBC
RYRdO8TgX0+jxGzN26kOVocbFv59M8+ZFwwVPHut48ldIVD2wDc7ymRCjY/vLRKrIRtMFhdL3GC1
roS5/Z36KcwgHoCC0cPjiZ1mGpAk8FkQ9ks1dT9T2LWJP/VQ5WknvpYb1AXltmKpVMBLlq/mScLh
tCf8vomId97mxM70zK66mqbXURqWM6rvZsu5ZCf5a4194gLSnbSIy4Qt5gaJ+zCJ1Hzlwwd7tEPw
jJ8b5hkG8ZRqEY56lgjj3THCwQXhaeVN/OhVxGz5n79BE30sH33Q5gi7jQFAh3o+TsenikGdeQFX
gw9g6F5ZFPLt3IOh2Ra8V2rZ7LQBZXsYXAb1fZSwO++NA/I1F6yLYyqBHD3ePrIamIQzTNhKoQnR
fSB3vQQzMkwh1cobiXQZBVJkmpUgDko7KGiAymBW+keAyRSFeb7UMmriZfnSwsx9YaAzJ0sADTZF
ukEevQOF+fJCwtMPGTUNoOJyC3UUwKL53k2Ib4CHLzYFV47Z0WacVqFarR8+Fm84+wBAmzvWg7v7
chyGSGh/LA4EkSa1NCaO6aPCPpUbag2gekZn/Cnr4Cy7+Y392Izx95ihXuqoHOsfhm/6vlALlrS9
EbVzTjiDozg/N237q32+yzDgeCbOayXXdYp8auFVz06VzvgQgM7YyBBPIpCp8GIsX62ksQpQ9BYx
4yrLc8lTAx9tqGUmvne0VEfNw4eQIp4ayTfIltRasJpjWtfgOaawq0QV5OrtPZRm7AzXX4Uo+dPM
8jlax0C0XOF71anDeugw4m141xmZhRsOQ9wMr9TJHJh97SRgDSZ7jnr1be5husasYfrwa4pKehNu
jmZDAxud7M4ZF2MCvYwf7LAzEeSDH3UJ0wB4N/lt06HNGWB3PytBi+B/nL6C648b3n+n7j8GhAVn
3sS6zO1cADnZSVgxLzqhMTioH9kqJpvKk+PA0ZGZnL8oC+hU0swQhbq2CYpBtcO3yJaWNTFLtQu3
JxjFlUztzmK8ZbqG88VfMy+oN3kDLqUoyFA6L+0BKtUBvECPQgcER0jUZ9I0hnXnHK9BHqCZ4cj9
4fR1M9KJAr6ucGL7uPCmRfR5UqiRPnkWUr+lGTlA21MdA7eHFSsTdlWW5BJJAaV4rys12tE4Jfp0
+qUDs0lmPHB6Kq8pim+Kv+RWV8OJrr/WuoJqVv+dMzwwtuaEhhtc7qsBC8nKqWhcpX4PjDHvWRln
+bBjr11JbFpaxiHkvEzJec+hojG5NDcO0hvr3b8fk3aCQsfUhMSfqR3tpBO6vSZDdXDY6F435vd3
w7kkp3JRe6WggOhuzZZ0ZMV984BvdnF3inHxFohVCscoKwc2n1b3QcZ/FpvqQH10F6VojHq+0+JM
WBDniVGsUnMJWUkKNFJmlxb7qyQLh0MbdXvQtvvcs8sry/5YL/FhKA6VLES3WKC0KKJlFPKxChGr
bu50drwm8RR316he/uN2LgFfHKS2/E5+BDgdzAp5+KtaWIY+TL4wKYHdmOx/WDqeDW99HiIUybq+
pJeP1q7qBTT01vLuOC8W8+J6rFumsDFNQDykbGgvyG4tqvfVVfL2SKFayMNGnArEF0NxcZGGZQP5
Y63+RyqyQxSQBfAHeTusl5rYNxwPfyBUyUwlNphb4I8Aj3A6xBb0qiN5ovfK6QavUsY0y8UKRRHi
2zHDFFusCfS2E0qqmhiby8Nqy0VfCsstqN/snF3ls1YMIedI71KOwER5IkzGtDeUaquDmkTFsbCk
AePjU3FPEQgvJkzJ2aST3g/Rha1ten5TusxsL7fH9ZmoTyTGEhCFDcEq/Dy2gARPCkg6Ih+dofWK
DMCmE1TtVJ9vVBBmOad7EtmnRPUP6IF78HdVbOzGhNPDk9IJ8EZFra3HrjcWh1T2AG/Je7ypTh3f
ampEnRN0ivTI1PnKhNIkvHlqkOGB24GC4lFszO2jOA2WLZ4tJJ9cZgW+PiOkr83zw8mOrVyWgsaf
4bJsQhdiEPZpumloHLR2GlJyLpPndctlXjP4TtQ8ZqsLlO84rW3vZoRaSGRdiIq/0IIdO6GB2kVC
abiqibv3rzCv3R//jPkEQ+2HcqwDFAmSfPwY6o0P9YAPU6dgsOuwcml9fPgbt6nH1a9WpVwgOlVz
A07yHkHYjbc7mz4JXJTb9Km4p5EoJXHxQdA5z0Oi+b4+zYY42zhScfs+BOLKkwMdVOZky1a+oaHL
d1fVw+9wH/Ej2yPKZ6hLvEJGcUYHcMDRQ13CAcBnz9l/Xe5FrvkGn64vt1Dq2wXCEhduHu1N9tog
9Vhf025a2lGgDElZnR1od8hu4sCqxV+T9uiW60+HEk0+/vY3rsuYpqQkzIXhsMz2I2S09AFO4cqD
92nRsw6UUgHrgW47Jy3jHLCzP/LING1BTRYivKi46WvWOk93Obwm+HXmsmzGtkVQ/APVnVGx/4Z4
5lKaI/7IphXOBGPWxIJPzrOjL+UmiZdIzakw+KggFMDrRy+mFSKHhMeIzorviDF6en+HIiNgRidY
2sXQ47/3eVrdezDgt9VNl9k3qX4ZXx4Z1mwTipF6rAGP+I8DY+cVcOfMF2mYTcnnITii8WjtaNdr
Yam+UaA3+fxjqvsUFfQ8+5FFPL7UusqokqdnitrrOnPXHtd2a1c2/gfHDIgzCokA2cVu7V3v1qNY
+V7avZXPB8cDS3LApZiomLl9xZ1e/RzN+55sT0CP18ke6PHq7Ii7/89pwXotsViNhpDCqtzDq2pl
9khDWmOhIYwPID50O5Pe2MtYzhxcL+y6XcovzIp/Y5foMjpICmjUio2sw7NTr1hdjklH2/Qy7YGP
+XRE5OiDXTCATD4vLIZ1s7DS4kV4ZBLJ/s5GUYcEZx3sq5jiuFB+qyKE0O43BOD3wGR/WvkkIdox
4BlSCrcCnVudMZDRM7gfHR+wDqKp/H3oUOkIf0qAluxSRPQ7PzL0eTgbVafft3X9BHgA0Lv68C1B
r71ILs1Cm+ft8M/ANvoqudPozcD0U+9KpGYgX5pYeB3FAb+bXUVgDo7NRWFlGYOgKJtIU1+9CB6j
u/hY/ageJ1eVI+zm4FC0nWSlNnTYP2mvL8xPJaplcErzfdl6QKvf17WJ5eECJbo6n9m8Yz5piX2D
uKal4xNx0h4JgGwAqhvgHeQRiRCNig3CKcO4aECrkCn7PJLt6UGEPgwY1oeGs58EnPXCrK8cMBcs
re2IAdaju+Xa8LR/zc7JZGcKjst1TWOLXuBNIOH4k0l6j/TBH0B2KWnnnHCcgmSng8Ik+vsKIEap
G3byA1f5lyyDaQxG77/Jr3+JRLFlqmLNRcsDy+jIA8tTBlLgjOmtie/N09jHsZRaiWuF7HtLZGuk
rrjvsLfosdYTTcARMa/3YQpThzn4rJf3PntJc9jvIj3evZzdPiZkd94Rr8wUSuvC0s3S+p+y94kY
YQVitzdiws1V4DOUtyFtCO86susz1nHYclzOJ/iejQyBAHtky6sdCMGkFuM0ZyoIWppxnTa3aTUc
iS1peVc5PmZYykDLAXsbKz5smoFtEYJBZbc1FolpdalECcPBeUpbQPYaSGxcZYAlLtNOBt9BX/3x
EYcy5MVjwJ9IbR/J46BWw6s/VW6GBh4zWf6Ndp8sosPDeorzKNmd7eWNSeygKDjyxxzYCn2m5yrF
aBleEGd8e9AckqGObeM8aKmKtkMaI2SBxLwL1/cTgTZuaE9zJ3+uPjnupFwItdsoOU511NyHhwMO
c0CROgOaN6jwUICQy+34Zvzn/87pTyK+XozEsOyVN1FPG78Ks2HE7ubBrKCLL2hYBi9M6RSVWoey
YOjwrMKuJv7iNgQzrl8K9VUxL8hRStfTqHVsg331PFQgc5KQJLz7KcO+hNeYXnzs4+/EBePqqAXL
TKZ7JBVVog7ebIzdKdwTMDn+dM0I4+Esc7HRPFDZEHWLoYnEItPtAX5a1vSRPUzthpvCHX972fxN
5Lq8dHxGYTwTdn10ELj44pueuwBxe1LXAhbE7VNbKpjT0W45oi6vl+w6nJZn+nx2PGVi1ZZgf/Ip
an2+4bxtpC8IoGh+rV4I72C8OFoOByG40VNb7mB6lnrJWK5XkWsehJuyS4hPnOFHp30cotGoD6KM
4VrJK6i9infVrYxXh9CE9Bd//H+da9krHf1PYkSQUeJ8rHOid4Os1/Hwpbm+3p2kh08zqGo03rOh
HFmlaUVZ3Fj0dkK8o9GDMkarmrg9Ga1/O1u5oqn9nJMkKwcfkiDgykbxxtU4BDzlghAw2FvIqI8M
4cZoMA2bVkEWt7dr1vJ/WgC8p+og1eEMqqcQYzhsdjmhTUbL2xCgX6w5hBKmcUGE2MnGHv1sEFRU
2AZ9dPxN2MbphG9con3KlA56D78AAYu3Apsr8Cu9YdXYdqJMp17DiaODRoqjsCgRL0/G0/+P52iC
M06Un1HD06ruWWdwgFdGg4bRevgZUXgMUVWdorw+VACWkKA9uQWOq1r86NHgEybwUaoKys2+HL2D
r56NE09z4yNRYWLvT6KNjR0qR9on8EzcwUm6OUpD4paXCOkKKFPcuyijj3Yz4ewNLx43Ma8vQWqu
7KnSU8KBmgQdFZ9T6Id1L6ELm7gDLU0kLVQ6wdjKx2wtEbo4BvlzVP8U95tlZlciRKUprBAS1tl0
9vUo/YdAFXXsKwHk3BTcf0PUusg1H7pNEF+bMVI1TBZmzsIJvbASi9FGWpfiz8S5Wjwt6tpov0nq
dczLqfaKiJZbOMt1h8IBGS+PbVzVQM09m0FBXbOxh3ezIDg952+bs5rsPwzYKefwjfaCNLN5H1D/
1AOgY8KbVk0X/94kx9zubm49UYnpC+Jl/jxA7n9iVxJj4AfPGhreUOaUy6Kr84eGInrIozoFSStD
cc6FdpQ/kIeanbZe1Wfdw86oXMW/DgS7pV917Wtv/X37nrMpJOMMuH1cVQTm9wElfyO1BIWLXU0J
N+oYG/5rPH0uM4u62ghoyMBBqW5Tg9FZH8FJr90MlN3Z3a9ff+J+7c0ZpcX0FaPbH6qVFFWrqLCc
hZCIDrP2Q3CKv8nUWz/k0z96E41JT1Bysulow7VhgJj8SnMQD4pIhJY0mgnLWR2YywWA1TMu9Rcw
irSM4vim9688uEXWUdVrr1mLm+urrmGAvW+X/C5deX+8DEGpPrkuDIvNPv6fC93gDrZB6X3g7n2Q
Xe9EklZYpRk0DDN1T2fpLWzs1WRNxmXZhbtJBiKmv1BNpbC+vXNnSRQqHCIgjJaQ3G0JbNSvOD6c
Uzr7wZhurw04AG223wA+nZtIgXdqMeg3ZqsjNn9fdL81dVfD6dN3ZCjpmkMH3nvE6iKKzpIpZu1C
motQduTLtI07KwwPLx7eqsJgSEMLR1ufgVdCkKuKIfxWVpzPSpqrj4oIrpp69RNP+qqtWFQnVfc3
xXuJsy/Ch73BLhmn6aBUkrfTY6mL/5CC9IhOdy4LTI2R9thljaQFzHpb3es3Rj3WeBIJBk7ZhWF5
MWQvtKP166xpsj66jJqCmi9RKmU+GCUlpIVvJopxyLFNS5GuvlDKMmGsFZpUN4lKb75oHHiU039L
QviI9j2HOPaBzVpbPGg3AKm7IkH/ua/MYosVePmbY0sjlEmk1MC6ogn3ZomB15lS7k6VoAilE5Bn
srCbZkb5JgN7/zzYMS9eqr9yxj9zWv91RNG3Eih6IRdtn4DTkXPokOZsR8UbuHAPG19X56065TBl
KqGDofuF1I+tMTIlYY7+xFqBuaNp+7Zr9aPa5gNckrjPF5v7b+ONCTL4qgtNOpbc6nG9tFM7plso
XJZlu1pQh6ewy5KnXq6mTHew7eUgyM11PFb1CG7dCp9zkLubXEb8M4NYfPwlgI7JPIKfxtyXSY7A
ZLWPzi95tUtzjIY3PDyj2NPVjNEs5N5UDK2iZmIeWmGG/4N896qypOBLcbBsMiXv3SFpU1gd71AU
glYTzWmnrhZE2zuMjW226BpSLuG6FDJZ7kfaJByZYDNVexn6afhvacgNzAIQW/XYxQ9ebKdZSy0M
PISCLobgHvhL1p88Si2QXcuTamnl4BBzgUODadRLED9X8vJm3X8/KDVuiheI6byfECiOqSuZVNa9
gsk5GI8crL21PSfuILmj9Qnp+icRRXdaW2zawAIWQpT6cW4+venGwoO4ngizClze0nt0aPsAiOmZ
L4PfOktoJ222Zx164mz9tdOQr0QWM5ogtE1zJIeMDtyOzr8zLbJIX6btjR5VAAv/plP9NzbVaQra
aWc1aRJBKaf8jxpCz7l7YV+Apn8TxLoZVx4oz5MTk0iUOLfXILKQIqxkinBm5wkbbbPuKTkRr7n4
xkp3nuzZ6E9OKgdIlbz4SrGhi0olDYO9wSqiisou46HfE3W447/cJG5Q+D4DAE8LIxFl2VJeyh1j
zBvjMqPsGd4eVnEcZ/GLKea9MOZvCho+vWaekltVP0Hd3UUlqYWCR0dBiuq3oVHRW45akUb+csdj
UPE/QPzaav4r8zKtsRGCfYGQO0dAiHyyh4oKEk8hlR/SHqygVspmOLXnTzWi+7UU+Jf2urIRhIUp
/mR6/4i6ne4cGp4nS+KoAhUBHaEE3feqo8uYKbDAWwLoJLCeBlcQCymOeWjBUV3kSrxN6NyWnRAD
0mI597d5BbdERVVyBFSKWpmgztB/U/Os9leioJqLTUcO0uDuDzFz+JgNMfVFVzAb1ViySON1VK/Q
DHc5G3NwGeTBB59gIMO909XdDp/qhmMEz5/Tx78VedLZ3jdHh36s/NVPBjuU0Ux9gDYfgO0aBVLA
CqP/Awwv387AA6SBbW0vbD2Whc1DERI4Mjo6VWVvN7lBV1Yl96+0LASsTGB1i/D5w1n593f9AFCn
iyNOR9+2hUiZtw88ZvWrZJXDEEPYkGcXPmK3pFTI6HHlAcNiCuTC6MmVRT9VcUHhudROJdqeWscp
ddYlHJhFPutT947hzqoNj/EgAqUcH8QzDPdUJnGAYc7cnAzBCLvrSt4rXaBibpcelxaBPtclnwS6
nYk3IgQfKsdEBsBpdmyhv5PQPDy0Pb7/LQtkqXUU0AtCYfE2nKa9OLpI8iOEJc1rvE2BtYmZq+qK
W8S5nHmYlxOtdKVPyLjns9wyUkbddyJizRIKXRs36d0akSM5NS2e654zvMzvPg/tHddJMg2qhdV+
Y38niu34nQNnlNb7zGwTNqts8N/+bbAAPRLh5hNbx3Hcr3sCUwbvWS1vt+OCGArtL3wt9Tm2+L78
XSGkAIzU83U6FVBtMoH8iDdaYUX2bxzw216keYa+iGgK/8HHfwnd5QM7BPXx4zB7Thw8k3ZFT1v8
QuGlrf9K434sdqhXvkecAuAncxhRwz4QxQ8fENbHgx1TmqhpdIACbQ/cLIeckP/BXNh+RPuXBmVG
vIhttdZAMqA4rlf47EssJrCdjXXuJhqz/prA95YgN4rQHDlnVAp3j+lUkBV5n5opY1aQvrE1HFuL
7semdGjTqwrZirtwWN2lVjPLHJSpNrtxAtAcJMxqWPlCmxVIw3euUsg0lrNEtbfIccHapPKX2eQM
e0YO/1DcV0JTRVDjQ7xZQm3P+FGgFHtfTqqwKQIbeJgIR8ijl0W/o6wrPVly+58tMqkIcDwoQHlR
ueeRnZyqThfUL0GABjNaLkYV99gWkPenNL3JDl1/qJHva2jpqPk93MRWsY7r2wChtaZiZc8iVat+
JvpoPtTuquzyxBSlTa1T2ufCfhfzr+xx2jxRjM6+ametUL/LExAIHspEtRf1dwKA/4GDXferBoEQ
kvvXgvdQfHDuwxxVoPo6s2KdabZuRlOw5Er+EeBYNJicAGWlSd571BzDVz9OKYnspx/o7OufKvLt
r02I2wVxNZv8zXWG2szwr34u7udjenaZfH4ug+ePUxoL//c4loGsA2LNG4Oq8kFluJ46G0ZNsYPR
q5okAIu8xjaKxjyABY2sZaZfNbFYe04BDU8v4Vn1+k8w93/ba6PzTdF6eEwRxbzyU2KbhnrqQBV7
q7D3hCd4ucFFaq5xzUYwz8zlLRcxAKzKdhHAqiieLMf1sgHUf71QgEL5ioXKGMTbS/2/fqo+dw7J
J3GV/rRlMnK8LND9PFW0CXYGwx5DD7Yv1yVPYEV6XS+AET6mzp+mlK2Mtl8H4XlHkv036f5p0nPm
ttcce4DGmRMfLvrE41cFFSRtoSS4Hg6/vlJeJbnn6lRLV+luSSPX6SUwJH9KfBMlZ97VMWovQMnj
mNqSZeQlmXRMh6LLDjXiwxZGZSrXjc+rdHlv8FB+Kx7K6/IsU88r9M4k4UiPs5xc7eOOQE5OSoTu
DUKPXNTA/F8RQDPUARQyMC/OUii7RYc8dKXu3jMjVVM2XfRD4Qi3O46rbst/k0TKJ20wDNLyZRH4
X4RlB00xa2H35GG29YCCMx1nckQBCFaXCHAlLxR0lD8JFJpIiT/6Zpc/NVw4iLtWCCDY367V/nJq
SnuEoI80zhZD87Mb4iOTFsstQK4UK6O4W7InFzA7Shp+Tms/wzSGHhWI8f/c1egYtBxsJxDrimnI
QsLuo4JWRacoKIfanqxaRbfGZNgCN9QBSjEciY3utJv1b1qiIhW9MfTKZHK+P0VVlSEpf/7H0N1z
cW21m5w2pGIFdtGi60Bmu285kpS5I6d8c3TLFvdWJisydYhRgUVhBpkxlou5eRNII82t0mPUyiOj
XkNYqJRop1r7751+H9Wd6Y17CiyHnNDnKDicdgGPCJxsavc20XUN5sn/CZYjmQl4mSj0SDGbTxBT
aYcElmKRGPnrSt+mQ0IiVTsYNByroj5dqfcDulW6HUMlwj2bArHRPfLF5brRS2HpiS0O4T2tuJ+X
DTOXopDv/17l8jUVNxye5caFl2VWWl2yFN6jSZWl9FdSLV9vNIMvjPXVIuosJrBdx7JGiZ2GZDgT
/XCMDvQMwFN4LKV2n6z4JOmF35K2GK1OIu9LCvCd9WQQJtS4ehT+teve/IGJ9Hrh0xggyJTgB7Ld
8aSNuZiD7U6oQetOCYLpj3RpBHnuCSTXzsCc7Uz0JarwvH3HQ4KOSLkj+puGsP3oCBxn2n2AfxrT
vXVQOtKj1W5Yu3cXpvFaaOpxFkHec/34KkjKHhrAEV/skjGJvNmPnalCxTn6qldyu2LWThU167AO
TftkEObjZaCvnL/WWjSSzoZsKlhjVXVwIqo7J2my8u1lpdX1mkcjwkfrHaQUh0vmoVuYATwTek9N
FtLFaelCckjhg0hPZIpK7D4e436F2HATl5Zvj3boxSPlwlHu+2jxDVVT2HEaCSsEqqezZGv9iUQw
k9aCfCh77f+VxHwfalpuV27gJhXtt7nilzyJNM7tEIztcqyTCDZFgmbnkbMroDj2PlaYynK82YHQ
7XR2cQLjUfRB7fljIjAJ42llFtfylcht4d2u34enR4+LrynW71LagYIKSSyPhpq/G8i8jey/YJH3
tPVi4OoevOLbfKhsxZah3H1QDDCQBnyO9V3mryfHntKuxUkgrT5vzlkp7ewpMj/nr4fhFFFmnh4j
dHmoz32DZaCuJtY8Z+rdiZ5wnR8FWgWsCPZPrMqVIGAix+BWi24s5VzescuLOzqMLfgDkVl9R9BK
GVrOcXOGZvjf4l1kDS4SwROCN2dmYe6JJUycJFZymLxuPiiYKux8R6hrJmImila088M75B1j1cw6
M4h4toYq1e1RvANwfSI8gMCEEx0WPSOVOc2qVGcldn7lbnSb69WWT3gOvYvnMc4UkpLBnaTj1b/0
GREHXXJ6ZH4Gua+en7G1FvsJKYcxlVFSjPLa/ou/mv9O6IAjE0/1j1pGTgPhUBYu0kD6cTlUhwFi
Woq6dyEmqKC3C4B5N4LKZZT4e4lodZ+MqE+7e3UL+Oop1LcBC7+YKEK2Js3ZtTjpR4vgk5Fomnug
kKmeyKDupeC5+0mKclHCczmXMmxZmXK3fti6OuWkf0SVUM+vpPAvE7itN6y5cUinnyt+XpHpwome
U2DAKtQC5mESg5L+bu+v+fD8oUyo0lcAl1fBDl6xrPQuim3H1s5VKMh/sdz06eBJqiamKFnbUZXz
Ve9fq37z84ODe/HYoASW4MKv77PDXD6anhCcFuWpfRKco2ks8Rd790XIx60Hd1wWQ2GNJLUbLgqa
SS0tq+M/2lEH2Wj9CK8Dnn46kJj9aHKydl1sjHFpd0oCTDn18by+eOGlQzagQYuNWR/SBPiFX3YW
FdZ7LKi/Uon1Br4bp8u/qArZgTj/vp6hMkeHBB2FXERedcgk+8AQS4F5qic8Ogo73LziA7rYf56d
OU/8Qyh+TWd2icm3haZ/yKUVhZMyKJ2KJQLqjP15yo4uZ/r51p9OlLgFbYtzMYmhBDHsCLD3BoeH
EiO/ipbSzkUBLlXERtM8zis+XF/Om3WN+YsX73ZlkzughQGofFNIS5/pxVGuJd7xKorl3XwNUJl7
PEXCnOHsuiaTei7yCFN32/seT/5/RfW06ZHmUMkNM3ExohpfHj/LP61XdzC5x0SWigI9EDyqjqTw
KuwyoNFSVd2MBfpj/taBIMdZ/AqNEEJrE2MwW2JHyzlOvFHZ3bV4C6t1m2PdQWTRwK9HlBVUJZtp
grg99XOuU7oXeLJn1EDD/kJNgFLDodCV438AG8v3HJ/FjshLkOm/fzY2ojWQYwQSFeFp0Rrm+Br+
x09N98+qZI/LZSMW0o96Sw3V50pSZPgyPxjsSP6lYu5RQFNKM1wnGAEMwyzqCgSQEeKrTBGmapV9
Q37L6Oq9bnZw1XvYTl+xDmMokaA7wBXgHOLxTs7rkCJdQWzEEc2JqoxbyscojXLKAd01f/KmkgEL
H7SbflkFiclFimqFoesZkLrmdPBYNJaon0DnE0NcnMepsbko2IbDBr8rm0At5VLT+m/f0OrcXu2V
q11Ibo+taF4GSq12e9fnkTbHR54pFz1e4Vvd5lU5JboLCI6Ml9vSbuyYJMwHGXPfZTVqxhH94nB3
x+xjDBzMAKWmQo801OEEkOwNb3ItYT7Mzt2R/zbn0WMpCO6+BsD9DVz9ER+ekK0QKbXiz1L/MfbA
K/5h20n4qr5UsCzp/R+wPXLiCtCYXFnRlyhen3lq7U62z8Li1p/4F6zryzU9C1oA91HpGLjJ4zhw
rRbs4DSQQ9gj6TCZmKwKlmlvv2Cp3xxYoypWzzLf69uG0xpPMxZFmXW7EBKueX3Bc2TMbgv1GMRf
LUQqlDPngf4kYZxKzQaQonGhQIJkRhzuxjASTBBULhAKgpjL3BMSDluFqRRYHLKqZhuiQLzG9FIP
4+0IQvsQ7V6bJN8PvejT8vZp5wIvSiz1hK3si+DWlVFOmiNljQtMnGdXIYp74D6OhAFp+xT2V5FM
i5wvHiYGBXiTcrePEL+GbrIyQNltcRNtdPpJW/qEiRk67QHkYXSYP2WNf77O/5z/YzAMqSgx7izO
Srik+Y13zvVqB27l6qiDe9oNLYkIPrBMpLPnhbtotTzelIoO4qEcAIYLOO9i3BKHDgqUYXE1Yjxr
CiR3kfWu2AT7lMl6arrJrJfFtftmJuoDfJxVHGB30VTrrVMGVuiz8XVSN3SfQlYBK37eNwco1joB
Lw+r2f/Rfji1zLOcEuEiQSzyLIttQjmBCQZYz6um1DYnTkxWFkiFIFRH3qU7DAxbNk4tAgwOkJ+Y
G2WtQqbMIrwRCTX+mEAO0yGB3s34O3hG+YOERlp+O/s0TcuGGw6IUTht2Ys4o5Qe5OFicL9GDFw+
QPDPfg3Si/h4ZN+MxXhtWInC991mFOJ+fhY1Y0iZifb5c6a3x3FnVb/FVuTR6SDRSqslIjEReO4d
K0aOIzKjoDROMqK3Nhkz3dmk4MNqgTVScjolaryI2vXvkYZeG7VAtElqrHjozq5h7Bzl3JqZZ5tE
1iZJG0szN56laqqsQS3ubnOcSqJQm3/+6C0R1rNN9K0Rd5O9F3fTQcvkBxJcasmMWvrKQFEju3ml
V4ZvrOMMHWyX7NtnU7B4ayUHHmXPUgp5DK94ImYoymHweO6nyIk6MuTetEJKDM8DaFHx1RPU8/Yv
FNHRhO3Fmep8CdzMqfXH9FbZXB/gPiVOH771JEL63EouFTJbS+U9kMu1FVcdC0WYNisoMckmu7lI
hKo006ZyOtOKFbpAfJAZ6gY/mM7+fq1nttvqsloblo8KIytSZy02467bjKY2wlomkGiRoV1JykQV
rqt1SnuRyb06PCRM2BixzKEz7oAJ/qdEyIc9WwyUkg3d9Vu/RkS7DwyU4x5Aq4DJ4eQ80ByNMvmo
GAXaKLNryTHPgtvY+teaKDdjFkKALXwZIz00sP2QvLboZKigjBeRExkxoqmqmafOF+sTVCia3lts
q3bu73umWh5JJ6r2pRJ3ir60LJlzo/wYt29tk/05MkU5hOGuOBUveYbRbuWaQlTlwFfGv8wE3KKy
qghq9TeU3caoV2BUdPhHRj30F1OCUfuWrXGBSK4Oe7eF7b9oA5s0LP5DX5R2KQl9KQBiKN14A+J1
27YdW/Lk3bbG9XkeE77sVueG1lLfn+90auu511Zhv2M6tV0uXGYfgZ9Q4WTCM9A7nWxJH2/cyDNN
fHzFbm+4k2Gtewppy30DuOAs78o9evW5tkrxwo20TrXMbpKjN3f50Wfy1+wEBdeYv81TmlP0EUai
FM+QP6K2njgMMlvBgdzgw1vIGBHI6g6pAf8fWg0zy/XiGnIy9TrYHjvVBJBH35nGMZutYllgJRgd
nKCDy2RNXDj2TB/TTUczl93cOnzzjEZePDP1Vpll99dZGKX99JPI7yPE004HFvBMSPiEx/YV3+dw
mn2GSvhPfp5q72mShQm7Y687yPkO+dgm5QVj/1tJvlIulCY+k2WmUG6gHE5xEckkgAmGRPaLSiek
6s+m3D5LfGzf6DPCku8+nu/wc+XoxICbNKxZtnGHY/4Jkz+cAerOvDVi5Q77MtGRqLMCmd5zzNXx
QsjhxVfkraBj1g37IefQhJnnJR4JP8EzX2PUKny01HaIYiU7oZt/yG1uXJQp6giUGfst5rABsZSu
/LiqYQlDNNmkLjQyi6IgclMBmPC9nPMEPnIHvPpFGhU7+LLfltnfliAFkgYp6m7mgY5pafWzAGmx
G5Ba0Cs0mED17HLX19hqvDxL8Jh4q3yTZbS8k/RCtobehh5K1lQaV+GGU5qWJnAMiCZWazpvBxUl
ivea4fr0WT6/E8aMv9Fs1jfRj2yUsT61C63boOnKv3AtxJ6d6t9prdS2qtwivqgN+au7Y/ZM3mYu
9w4XZ501cbTQjImW21RGNyXsZkhH4etTfrvnRgnslriKtI0uE8qx1PQVK0R6m8v/fp8nuDJsRBqO
CP0XJq7WabAKljakMKGEIVbjNS/32EQeaGVLII/IWy9yos3N9NiBA0k2Y3qz2EPWmL8IfqbYeW2D
WQE9ZkN9Rhrpcw1Kv6x2SlhUXnLxeQvKosb9kyt+eHZZInEiVK56k2RNOe6GUz1kDiNLMR6VBszp
XfII82Kq4PG8kEA1yKpWmzRC7movCMp0U3ngIRKVgg2L6/yKKBxdoeQfUILyqBsrpLTDtm4r7lF4
fCpcfpebiNzUMe6KQozpqUr6fFLj3ufhU4XogW83GZe9k/z3vRzipFscC+YXaKSASkeY3zjOvfkr
53nO/4Yi+oDIhEciFcj/pUZ4nx/dF0pDx2rkMwAp0yy2XbAiJny3Tkqr6fY9a5UTTEir7L5ibLpX
kAwhruVITB/PwaSOjytjx/yz+yF5/d/qx/oejFHNoWa8lTMAvPzqeauhEA48DHn5KUt3sf1y71kU
2Trk7+kCvAlvVA7hZxm++2zvkgWDP/QDmeYksluOuKhR5xXjSFzVvxXQDxItfWWBjW9mNqFFC0JR
Rke+j+05+wEfVURiJ7PfF+jEjcyLy70RCJ/i/YskSSKLUh1Tq2CyQ1KGFB/ZRXhwMnpVgkNsdhza
6aZrNpPuKxFN6XbwxF9PCLNSUHHMdbGEmSVlNxuR8vJkNNSWc1iK5/60ZXT+dypc17AUVkUN2EcB
lte8ic54IoJBURl2qXovLhC5K1XkUNnwDW1MXNrllTYVLdadilZucA0fizILxN5unY7f2KcYpywW
lee+pnPAJe4FfsurhARtrrvVpS27nDqiAystzSlMPcBhASetU+JRSFGaluBG7G+pFjhjDlvJBKiY
MwIfKrDrvr5rfWui+Crgh0RXyRf3IfrxeShWUpZmNeMP6iZLw+07BZjcgiAdmHA/99lrCWjv2ERo
cc3KiMixAzZwE9uPQ6Y1k+72Drt/cFKn4GUQI1+lKTXoL/PyUL5LSqadFqI+NpZFKFhVolgc6QJA
yrmeS+DzmtoY/iPYmedlD5uelqA4cFwYFNdfKchk55m8SNjF08IaNqrCZQQS+MYUcwhXiesD8Vt4
uxwX7rsljUR50YVVQSyyhbEsdEb20NcyzKrfUw/JRcKV9SFO0VVCCLQE4pqgBsLnfIUX09KrbmUX
lUYylR86YaTu6nHlnCv4qoA9RfTQm8g4wjHjCKfkdBSVGe0dwmQ28RVFMQB9Au/MlgfjpVANsjYF
sTirAMvbcmfrx5rsw9yxKxO3enO6hMp7U7v7pApFGwPN3NSVYFCT3GuIt91WO0K9yNjo9V5zvT2Q
5fXpgpuC0fmnxhpQPRUkPia5uecVOWN44UZD5tLbJ1uCS6HAhD/ORqTsg4uDpKXxW76Ejg5mAhYl
EWbyU20RbSPD4ezGvsC7seDME0L1JpWz/fxm9Fgv8+qDaQEIBv07ss+CfFWjE2QyQ1xqfon1FG3f
VmgVurBuL9KHUZvjAfy0vVrNVjDCQl6Px1A9+LopH0sNHk8YTALWM+84TelayPHeNq0x0v5/+SpJ
CWmUNjDXV1XtZv/cbYAXpYhNzKh1Gxqgm2uJT1fnrO4WQ+0tf6LCym0DFtI9FPO2BUMaENzco/5o
AyCBa+nesZzFbltEu2CUGIeC7i6q+O/p7qu7h6+fsYPcBMIY83G32WDLLuTPYyiZpgCotQBLJprV
aP+vhQkCBGNBQvWOwn/6Tx/2QxLttb5kok3pA02GdiOEbXaS1Mm29eWoSqWRq9xhVKLTwEGr1bmg
bUreGIxC8lktbfdzmzIbBdxEqGsB1IM9U9ipd6PSLD9mbSGppazXQH3pZ9RsHY4CfeLCeOjPDzP1
iM88Y+qXEOUJkzYtrtkwu5CW/8KPeivZF8APmyQIR+XeZT2idWNt6Ic6qdZ+fd/mNHfoa/AI84K9
Kxv8ckX1LRf0kfvNj+GjsJ23dxEIKjXitHGmWPVRJmN7Mbw2//o82rdYGwo8QL521gGAh7Ep1tiD
iDPVDQ9cVdgxiHRQdI1XzwwlCkOducMbUbtjcF+qsMSJe24L96osO50tdcj0Y1S2PrgyzdyBjd6c
n+6lZkLUIpMcrvAC7DbxhYbgNO7zadWTe8ldac7iII8joaBJqxWBGNbxbiTaFB0N7Nd7qjRodIiG
65+6b8AWzyQacQuVMBnSm4KRBysKctwxQlWM0F+IEfbnKogOXZBjawRTey9Ieju2+lAJSQ6pPfbA
JR+b/QDl0OYqFOY0/+wrR+ROwvg+xhmiJ2l0UzAnb3B7OT3jCSPVgGGNfIxC8bCeFQZA/aA11huR
A/oJBP69AZUG+0sLlI+BpIS6yrHRS4be9Bl1p3o9Cr93rBLnngFY6pEPAEH5+snHvJI/DyctWZMc
9NyeatIrK8QpSuBqIG5jlIXqz6dPoPzr5uQGlfoDdS41ZQud/dsgvEB6NdiHxPwLrvn/qPDEN+rU
m/XMfDZMic4ujQQAgGIs6sANw0ZXHfCEASxNmU8EuoqTc5FQvjVN4QNGZS07g3ZB21D7EnX8rFUu
7+7V5xcYcpom9H0pTG+CNmHKIjkXK7VMI/UFWIx3KwlOtoDbpamn7jy094GypPIob/OxXP5pSWW2
yg1UvvEWuO91rMA5n+jWmSmVF5o3efRBzwU5snEiv2AguPzWRM3OvHKytujzldrspHHFEQ8QwdZD
Gk14saEeEbaacvT9qGd86BmjHgj+5ubyB94d/5y+JH4obrzQ9hUyEKGwpdXu5iLo2Q7opPE6i5Ac
xi/7tWQXXl/MQhc7TL42diIsmsE+3QpN2qGCR/T1qqk4UbCGpbYwpIa4nULO0iBPzFjj0WiJyj91
8EMvdgV+G6+4/4U0AKfcPGLQCWcQf1HcSYyMDtCnR343iD5KOXKTCxy7tbkgzoaLBXo7kfVLfMGc
bdrjAGbt/Si/tzQ3tueSLKCiCZw6+DgLoE/elJ/5SkvNrktF2JT/2K8geWe43qPjQPbaUsdmEbH9
/i6YrzB+2lpnJRrxj8SYCtkNZm6ELZwZ7pHd7b01bQMDdKsVd6gGbTcKd6nJMe/rbFst1ER6eEmk
HESE4f7Rx6HRvVbpZwyOknQpxlZl1ega8PxNp58NJAy1qH0n7+6SveDiiU0iA7n0/GEES+bIfxwF
uShRAN0B0czt9Wrbpj8PyO6wPYDuAY/Wl8wNR1pCxIJH8iylvGwEwtAhvckSX3x2wq4eIUtRaIrN
keke2Dh7hNnXgtP0anIouKQOCHqtXWyiRuNiJTGE28T1F8HVmGHQ+MKiL059LytDBOfWHtmZ+Gf4
nlt0Q277fMvF0c2Jtbr9LemDrHGwc0TJbG16HcYFHOz7PmO2oiepNWCdSyUSb08am8udloysqLpL
CdUfbPP6GOkhM2ZXvZWyRqYJvahMQh3vXvg4KLUAK0eDftuK+NWAeexkRPU70uBUgpSKlmz3Tmsn
CvybB9jwWjx9KTSt2dfgKcsiVs1BSU3i50LtD44u/hbWiKP4wkUqLneTy8wL2Z1iXyyv4yvEwOj+
h9wBrM1PAPss1xUB9xLZQKJxppFVp6ms2rhA9TQrCt8/N+SjVopH/H80Kimm3YvPi662XyQuoQjW
Q29VJjNtYD60SyqJ19sr0a94JCJjWPYQHoONZHmtzfGW4ZmGaYI78cKiOeK8q3+NmB566d8Z/abo
TvXXSCRkDjOzx+BpKWdg9zIwwYDoG4/kYWWUjINeEXD4F2r51IhK3dczRMw/c/MmWkpFopu+L4n+
RxGfTGzZgzFyyKUGkgwu5RhSqSalCzdjB9L6ulCQY7H9MP8PWzms3wl1ILJnkK0PIWJkNQDErS13
zSPWgc/fwFCwFMsOWCnAbrHlBoNzMHUlEJ308MSqElmJ9vQqKEnS+czt/x4K3SfmJdGVWct21bVz
MoQmOyWFR/sXgCetL692tsL/nWMBhr+yFFqJa/qL7APCketnyid6gZax1o8OwtACesysp1hjzPNe
TxOS27wNrsH7xnQI/7sL0SurGKa/CdM5zubuss7wL3tTx9WzCHYXHSKYmFQy9OJL2Hqenk7Gs4Aw
Q/ghH4J6bAk+OGfam16J7r+WjxfkOv7gnzkWEwydN5E+zGJ2sgExToxsM40aT6YRvWG5jeQGDnkG
i5f4S+q8IU/ukIlb4gskw0WKRJ9d/9k/eSfWnHHB7819XegtRw3uF0HZfBeohQdeuT0f0gFIWFdz
xDEwDx5v1KnXyo2PuLLGdzOOuvLcNlpCZMazG7ARNI0ktr+8Pro1x1Mgs6B8xy7nkommj59wKRqW
Dz+YT030PZXTYn4oIbZHRWFTpoDCThAc/2e/HWMQidlpyl2lUIFQOFeNS3NfAHONZ0brBkKuhIQM
BKqmxkygLz9NurgfI7xvJ6UOHGFP3L3zKpiANdtTW8cSJwInuZIe43ZOwti7r9KgWBmucElTpecx
MXOmiSJC5fRMrijIHNrrkbAE3UHQCB2Scd5PAnWsdhoGbGw1pYPbWPryhkGj3qv/dIhYpc6jN2Vw
jSBWTsKLuITUiJk8G0cd9a5piA6M7x3MuOEhAnlE2rGt6LzwDjAN/2X6od0BetArMlDE+PXfR7b9
gbL/V1VlQp3lbx7qlXBnfaPD/JWjNRpWDd55d5UCwdQVFY9dmxgo0OVtwHn2DLVysYiKAh3NK1MR
xvRJoVNFsU9yuLLkxfr0iwO/DKht9tmRaWADOjbGE4l+pG59GkWAoTYDSSdQbowXA1RM0QCFR9/a
75+saxGz7oWsW6UhUa1VJmPj/LRHvteZmLo9bESqKhoKDLWxSw6ptasD3nBWJ6zolaV96srZBOly
nGBXy4V3GcOSWy0rfMXW//HShEl1U5Z1vyzOYUB2Bi25dYdNJPN7wAQaibgwJEDRrqHy9szLj21s
eI/RyA1TFw3CAKkm66YVpIBCfkLPReSpJRWVRehNY0m4xIlkjYOZ/IMODeq+BWdS1sb4OwdmxH9f
OhcBSh+qEXzJUmkhbKLnNSLzxoc2/kgHsPSNk1PChuv3TJ/SayXuIpPipOq5Ddw/RjVO/xjCTcew
YmYXcnH1zZFy6tprwdmDWxz4p5335WpxbVyWWDRHj+EppS6H4dKXo73LQV3lQlkjP0P/UDv1KZGG
uuksCv7N7k2TyCw3LZkSRG3/Q28f2kEVAfRqC7R0ass6C/xc3hV6nqvMR2HFoKm+kUgDX8ndE6TS
GKT/wS0MzNGNAgR68WOiDg+cT3IDLLaXVn+vdsOGV/xbvt7oRaB0Z07yaeZQ0K/hxEnkGRRQJUPY
0E+xQZCtAHfl7xfNCSu7kj9GZ96gKkdBpePgYEar3yU87t89R//jl4uX16zYhsb2ZGg8jdamWK98
wF77+5YZc7RexwwkWrOCqnJ1o+Jh7NcLqj034ENezhPMLozY7M+NcP/zubfAqMEfxPmjrDMysQdM
7jeIpEkwqhdgStNr5mbnFfLQFZ7fYHRoFY5AKxWP0wL2guQNlzhOWwIg4Z9+WrQ+rHQR8n0bgw47
1bM70V3uj6SZ+vmKTryy1Ebz0xfjp7mlFJYthdI5QJV+Hzp6TNye8byzPUlznU8uApByN7xOWAC4
G0TMod/aI9uuwq6Jn3B2NBk9SCI3TqANuyaZ6wy69C7TpqJzI+JvGOUOIcv8TvPLdJ0hCiyMSiaE
u8e+0iL4+dKou9OQA32fZZMBjukBTAtfJQhurQNuwQst1Fit94Lz1xcAyk71gZ6Stni7YVphgmRX
e4B3Z01gZeU6rFntuMHImho6pd5nVlMQp3ZXycG9JB1WRHhyBepIwMQAlpsJKI4O6BIT/qS+0KOv
B+47z5F1cz/ekT2GgljwG0QmxxRFajZOznzCZUZGib3EqvsiaN1P1e+0T+hVwj6sZcf1Rbp6bF2U
Ui+Ugm5hTjLdMvmCCCaoP5KVCssYXNo7keQv2SW+fzATEpBFaRCNpupu9YhvbrCQca715VXKi5vX
yr3tJryLjDC4OjHPAjbH31S16JFbX/PfVFEISiMMr5qs2LqrDzKWeqml7Us/HMsRpmZCUdIIzZBk
z6B6nedzzVipQDBmRyS5p/4+9+PGaEjXEAoEnRzh2M4mnjYmZlZ7KOtyE39D3qB9AAsOUS3oJRpT
UZRiUQi8vRHrWQWtWGbzWxLvSjnCvzHcF3Mjx/bT+EOjKyPhppIFUbMs4rZtJRZuDIlBVg1nAiJp
jP6Voq224FdJNCeNdFNUjxWJ9RNVZ6LeO9/YlOyzMXtXYVgQEG3+T7o2p5dP+A7bXe1GAkZGur7d
JK4QiT5fJ4QB4CASojDJicj1SsrfiG+zx6ehXs6Na59Kr66nQYqISlp9nm+4Tg3fnDbsqUx0XloI
i11BpiMKYK4FRmHZy4vW24Rz1BMsK0xDxLnDxigOSLP21NMgtGDQXGwadZMEVxrnrYS7AlpCE4YR
+uvuCxy4ToebElFIr5fpSkiyKmiK/Yxcl0raF9TP4hQ6CT5L/hPFExBdTN8tflQZt0Pjkl2rhnT1
C8W0bjdAVohun7/7A/TB/5KG74LjTRGY1uftrn8UjTqYextTskSZ9GsYchHO7IBTB5W4bKcAnQ0A
eP5aJ26vDh9kGJSX4ZanS5VDev01fJTpwMEPQoUEEOVXW+RysbbT/cYGqdEgHDXcI18kNZ0bZthx
iKkWpbnDddTnrLQE0jtSPY2c5SSlNGXKi16PSLOdMbwdhYyfMEK9SobAa1X1rpKg1cdnj97aShsC
sB1F+MnP4UA0qOD+Gt0S8O05v9rxaUfDXYLeZxQK7lyX/M/6wJGlUEfFatXww8tlqP3aBGXUFAA2
jI2K9qHi82STzLFq/1zz9QIvCJgM7Jy5IURrp/5IMTwiDdlH3fQl67RQf3jjT3xyPLYldRaOXGs+
SRK3SYJQgc3NifdUC/vBTkjw5RYYSxBAUkzi8WhK/L1YkAysoMmVgnjbUM7t/zabV1k+fMfzm9fk
f4iYlRYGUPAqDf5pPvJdjE5ySpBZY/Qrs05ux6aX6s8VJr41f+35dZ1fXHTNelBwVJ/BA3bJl9Bs
kKtzDV2ONo1nbe5h4GCBeVyX79Iim+MFc4ZSpTTcy+egUriYnnMKAB190pJANDy8yCkgaNUn2zXr
xPtD1j60N4ykNX//0ywUTgl5JDKagLIvcVsfAAGAERfOoQs/0ZPiVY03g2NcpMyEjxBiHfUyKesK
Z3Sc1TLy6q6y7a7UOjF0WiusvowRDmISChzSIyKHGBF0/OMiN7vLMyIh3SrMwFdS/sdedPl/BvFS
WQqP0n9YbtIJkxVj/vs3t7sib2fozRRI+kXF+MOFjzwq03gtvo1DY+2fRxSz6M0FnOoPKPV5xfoy
kYZBSTm9Tya8Qd5jUUa9G1TMCJBt9hN6a8PB1u6PBUZ1AIrUNFkCtWfXWM30aR46VaRbt/84QHcv
F9u+WpaTlwWnUVsEj+UqPcSVyM9IrTHonNIe/Jf7Bu2oCPGsGP3NpyxcPUMKfg8vZW22I+92/gXj
wpb5rZK/b1N/pkjQOIi7JAS+68pNF9cWXGpy2/EIgcts0Y95yfeP7Dbch1cBpfYHbJ5QsJby5nW9
9Q2DjkXV0ef9B97p5DovD9kYyk5iEv+nigtm5wcbdp3rb/H1TMSv8Nkv5ZZvpslYOT0ONbDykDOM
ajxW6OshrxhTBFXM16bRJWChIAM74xKXYk/cakf4z+/uFf9t0nJUzEipM2hZsCyxF6n/SVBu5Bop
Vs+fQ/8hMqECkCxCJmjvqOokj8jl1RTbkOK8od6OVpBHwcNH4nmRBhNOWHH2IWmimlq50j6Bd7CU
3SQTDYx+XrZg150o5MvbHA54sJ/OQZn6PXE2KbqvtxfZNaNtAWTrjiiMbMaalyAL3FMsxdlcLYpr
aAvJNTdp515nnfTZrKXj4+fFvEYA+rUvRuWlqs21aH+BQ4AOl3fqGNQitg7R9Q7M9FQ9Vdi9xAXs
+Era4WEYaQK0nMOYdJ55TzeZoOlV9mo3FhHiAFf31z9yPMkqEwhhlCDZdi3eN+RhPOYb4COVh+a7
sRRdEbLyJjAzYEsgV9MBbTwbgKkZ2o1VQaymQnIqetbK3LSMDKzyEVKrnkv8Tv136frZo7wljE83
8167PjkNy76pKZfpWDgrfrEvr6fodC9Bn00iW0TM4sQ3v46G8BymlLJ6ba1YRxG4SJksZU8D8yUA
IRergSEY2WOXZ/bVfz3LdqhQEqaEXvhWgfoC3unbDA1xPLiWFuKuM07rN7mWc979Kqtl46cBPK/J
LQvNJ0bXKyFKPjdBLk6txl9dUrbH9Sh63fwTvlnjy92fAfXx5Pn/FBpOE3mzt/A8ihZa3LlMMC+/
5DFgdr/S2RSheMbioVg1aHWFpOWMzRfZHHp1Q25WaytlftCP4BgPKDiRzW3h6qZapDlLJP5UnFy4
MeK6aMdQ1Kjlnw/Q2+6EIm6mYouUszPOO0C2EJq3Ycbi3LxrnjU6URS07aL0CwNeHfZZzaRvKzPM
0S2VOoTCV+1hrsXxPtApue3n249B2BhwYZzpeTISekyyHvEH6CGCWL46G4393XL9nUPP6ZyY2Oxj
I0L0QRj9OqgxRXJumYe696989Eyzq8g6WQZJGgfTvdEfxafqCOoD73JhJRuOYYGKomCYLMux7yER
HTXF9VsxcgpKXY8a6q6l7FGkvGd2mAXSMoo1jEWkboL0a5lgbauazSN++iX5lK8yWTn/cge1ft4K
o9TxJKOMZOfKS/98XFvnBPF9rOTFmsVc8wNiMrmiRul5pOTLYBnIR0Pr+J4Kjc2baJqHC/Apokju
BLE1Rx59GdX4fbubT3EXoF9QC3YV+L2BjFUcD7Lgr2AeZsmoXp7FVsqF749Q4Sv2GkdPrhXaqOvK
/l5FmjnzphixpmLxYBYEYCkz1u3d+IQZPbDbly9tsdtEwiJC85hGRKwWW77ZPNXfVq4SmMmOI+hW
lC3ymHfWkU06WF5XgkMrV6Gt/gjG0Wr1vf+BBOHHz3jqggF9i+r9bgR9kfj2I6taozsS6XlD/zIt
WtIBp8Sg9I6NvFv1vj1Dm6r+H9cSm8riCVjHPRHixJj9BCz2SjDXNJJvwliacKr5rlF7JGBuaVpL
Y4FJptb3mDcdsRa3TvPgala7ejlLT4vjl3hFDcoQHaDNfmQ66Vl+H5GMOgudXb/l3bo+pCDlGOgt
uOxQGTtnVXMB6xT4phqhzThgbNjR4Xz6sHO4zFlYwZYKxPTwilx17GdzoVnie7bkW9XvZwX/9S0D
AjAVqQ/EpV4GfqKr03HMVXH9Pv/8WqRp3nrV3JPXbkcNBz1FizQhI8f8wC31A+KkcKNo+bYDyg78
7mX/t9A0RlK6WsQGOlB4JJCPE8NYXl23X8dcEU9RDjzW2LbkyYLje4sGN7yfpKM8Yzn6jDu/5uUe
fzukk/OdJ5KnHvKSzk+cNRl1RVEjHVAlaZojoDbQQDQyFIaqt/Pk3eeO/W7Uduz/eN+BMpnMTq9H
LeQ5K1Bd6YfILbPnD6mNl5xf9XFYWiWvPGEYATFVu3aOWAGaGGEP4jS1FSC4ES9KyhNou/tUerCl
i93uZYm1MGX/uVNca4C5QUk8dh9fEg64sPD1e92KkLpCt36WKrzLF1Z6z7Fl3XfMyjDFQpaVTNiA
yclRZYLeqMWeo4RqOZEKMMplJVrUzVWvgr8eRjmxTu2Vj1CwhaEY28dEQhpN+ra0DQXnXp68C3n3
6cKUzabPPk/H3qLerupu9o2QHNS8oOXvhmMIa0pGDCqEYK0H6wIJNQMxuXvLe5bCwHUF2K/d3/6c
aSqKlH+52ChWg6+0H/+sM/T146BfiYgR2X4pweiq7/fVhGGm5jH7QWySHOQw91Ui8c1wZRsk3mJl
yARB9lYJtqd+maWdHvlkHQTa9cUyV7WdIVQ8u/zXCTDv5P3H4ERyPBLbHboFGd0hUsl5nlBDCDd3
JLRMzLWHZhxaSwArCHLHRzucRQSpAk4Pbfqn53uJ83U6ZOEYY1uxSqKC5dcpqrZ1usOXCpaWwxTw
05Hfvg0tSPQCEGdsQ12NpI0K7saj7XAsEFUorWB/jVNAfB9cJnZDObVFJkfIcUX51e42UaWnl81p
HCp4TUJ8/VDgWbq+qG0Y8GASh+LJBClxLNZW5J0LHy3mb/+lUzR1bR6+fmqTsIUp7ZN4YK/GqaZm
M/MLI+EHFn1WuexYaya+pBJtjFLfhvtTPv9lTeeV212U7W0yEh2ZpOaUxGQ/d/6/mahogc6A6nzw
x7DZ1dzl3xva5KMdZ1EmPY+ThjG1RLxe7N8IKOzSf2sCZ9jaFekLgShtGzwPl9xDDXvFrKY7iNCc
AAG66Re8U7P5xCOoK+mV1NDqkIaQyfhYQiHC6LKTyNoa340iBw10+SX9uzEKUWrOCvJiW8Dhks+M
AdAgmc6hAzGYJD+L073JG1RWv1V8IBqg4JJlybx9LV/OANJMpUyjuDEuJm8KtKsrVUMrrfss94rd
2G66MlMUv6jIYhHYKOtHqIL2IDRFrdCvhVd8gsGmzK9p5RM3lrfBx79y4/IxP953LD5ZsYdH7b0e
ab/yHia6I8bpIeE7rBOeAyxXFXZ4//QKo3wPLPzoHEsSjMplomuDTmlZD5itPgTwIT4vimxTU9xr
77AlQ/3a4p8TMVR1XyTv1/JzVVwXfe1MFPd0kUtNz2Iap47zCat11Et17JWMKZjqOj1K3lyl7gT/
sAyQyn645PmIKOc3lzxdr8/gmtRipLLSxUMXV/3VmSzdvSyhrURr+bX6LJv2HZj1cs3Zkb//Bz2P
rHCh0/r8fIQ3Q24R95Ms11uONz7J8x8t+NQbgMiHJB6eZEHac8CXXc1zUbuQycFljKqn1/B8YvC8
G2qoSPm5Qh/sCOdkL5gyaZN46iycHHaB5EQotZDPvn41R6D9BaPsjR+gw7ErqD7eTbtL/i3YuEjz
4n4MK7C+iZCX/tuDIdtzCI7PF03+FQ/pIC2Bwe58LJzqBtKbL0tAcvIWqnrYED1y03jrPc2AEb1/
Xd7uJC/AozWxD2EPMo5q1vshi5hiDulrHwgJWB6Bqhuiixu3JvsDucs6C3lneh/Lfij/lOd6kiUe
kVmmjfWbv+MnEYRblg2AJF85xPtKqfV8KC2hslfEnTruA+fN3bb94ATyOyQ62zguNqZjds/RZAJ/
qG8nv+OqaZxttdgPkjnuVFJEeobtay53X0D5kexxiD45trtZmi2VpwXiovV4xID/vd9K6QH/bQD1
1b2PHk18PXwdG2Bah/RsxJIogxhzqjmN45RDFI8RihPPv2pmAQvSU60V3pOQJ9mvRKooMb5ngywt
RYwr/FB/keyr/RnwM1yO/DgK751BShPymml8LDaJ6T1tthrVTZMr7RlUoN9AULh9BDm8bBR0Ao51
AzwHtue94uyjUgJFqNo6/NJhFgav3kkot1BkUcD2XHj0BQ7H31lTxAJKR1FnttWnAkXu/OpOmbPY
f/WuKwuVt1DpsmDOOKNCaypUTFyaI18XQuUlEAeCV/jJryS4MFfItDRtDenucks4fzLnXYQWunOu
j9sdpcGN0a7sQWHNXmAGjwnP/J6kmejBma969KuObS8pMaZP/lVmaIa3+QciSqO3K8oGxHHwpq1T
h/UycBaGellr0tHb7ZYuoC/QzvpyZqwBG69T/87kI+1Sy7lNcQKvG9T1BoAenrVgg8vYKq4TdXJr
0sck9uqjitUalkH+RnlU+Y9VTTGCHg8Vu5Cil0OCt8a7oMLJs2zvhWzNuDoTmTRlwNAu2+iwPglo
nERCL/r+ceV3ewwjRKqHDw/OwAxs1YTkou9V+Yx0t9vZfSF159l+jOE4YVa37MIIJshN3fuie2uu
ZN0yqXBsPiVxrp/NPxYCCbeUuy1pSe4VserU3mcbsHQekslZgCYaWTge6eBFh3tzycOlwvGrIfyw
oejupWZFHHJRf0VLtpYuBUKJds9DCxkyEVTcQ2Rt7Dqf9iJab7RyUD4TniC0ZvA2LpugeEMciOPN
8L19c5uJOYzt5ny4HK8sWa7z/lUptUOsfRNdxgwZd17fBHkGVaJ4uIuEO/Hus46wzrdVoCswhkDd
qAzoeZ7S9IMhAL7SlhgXCjGpd2KhOQvGmTFsWpcsPooiTPU5lVXEF7O39HSKVa8rrScd2wW1/wV0
6UQov+7nxTg1zs/DQaAEcUWL7VyWiee+jtyzNOKKpdkPn1+GJlN/0ZWP5FZKn5SNmFyoyCPbWboF
jCVS26lTva3GcClKSpMQktVLSF6T7TcjR6VdS+IUP2sfLfME3Ao/L9y+LXV4ONxc/4qvfCnNimV2
34v6F4BfbYJ0+TXViBipjrDXc0YOCCmXsjRCZRPoUrzr1WJtFX603PYneIX8ipG1XPb8XqZT7TMe
D3UWnzEzalDbDkMajx5Q2Gaud8yqy7tcG8C6vicS/jZe8Oj2fjf/wWrtiHVbzZ/jd8mFFgNiuo/R
rQMOTyYRWkPM/EA9Hdx5f+tynq0B0ca5lDGE5V18qGJGExMW+9t5j1rCDhlgDJ9cIYsl4dqrPgZI
M8FE8TlIp4ZBwQA7MEGak0u/2EIWRtYeos4G3oeb30Ms6zM1BHNKbF4jZdzjhpswFGJDnQOQQLhH
Rkmwg8GVItD5JLgl/ykdmU6USz61066GVRZzPsI2mDMUyS0etv0K5fCl/OizEsx/ccLTKmU2NowX
cLqjZu3jcCld15MKpAL2isGCxva1kP/i7bBmuc7iqq1CLN7RelwCwvzEHvVz7IJl6WRmJo6n7fIR
Z7giliPJOWWWXmmiEWOBpP9P651DDlFgeyweL8o+Ur4q6z/XmoUhQwog+3DRmqIaEuZbF1Y93MQJ
BMyyNV39ozQ6x2IqqM4iQjpqULMojC8pX2eY1qr2uqtCUXOd336o13qsqLixiYRPprUcBgRWfaBo
GG8sUxbst2TWIfnr4wHdNQftHrXRFa8vGNV5QdI9v34T68e5/M0iGYP/pyVSBDGiXUN1ej5GFGVF
DB/evOQGHDCdvYD715FDk6mslJIgzbDKq2ea/uXxr3Px+80UAYUN8ryIO9j/FNzSJBlED8/S+cKu
vVN0+6i1I3SUrmhvQ3RIePUp5G2KKxpGtxEdFD2ksFmdK959dBPzXwtHJUSN4bhAOISIh36MA7p/
+e9O8+NRljCBuYd37kweJ3s6maYiRc7IgQw4RBh5zusGaqNQ3ID8v7beyIx7WhIQrhvmFnCU210C
hyhkhJxmvceZg1IlcKyO7OeWKX+3jT2yvBsLhs5NRnNCLy7eURHDFimXny5ssaxE8dNE6bCvRGpq
KoaptvhJWJW8AHelKm2VeRvRHbbDc/bmALMJNDO9jH/N5vmvINYKgKrQfX9vshRT+IC3B85AYG8i
nMcwqrLY+rC2dRFgpieZRzukn7ZOONL2I6aayyrevl4/LnXOJddmaIws6XhVNq2sDmj9FfCn/YLm
WA+7GN3XXP1ocnxq82NRMV/a+ieIzgMQOUQDYN109fEyowG6D8CzBk+niyIhabQntT+lIRJTDgqW
wIQq4PgUbhM+OjPr/yZYjJUGEmxA1QL4zmrkl9017Wpm77Fw+3rqKECJfoE9ddWUZJh+mA2WCyQs
dcMK4cPrFt+LxOwpSn3Bf5i/Gr4dOuQFokioOgApml/KDXxqf01IH7CU2E9YUisjVPN0lAIe52O6
7jq3ngDYGVyWcsBKH8pWjsD3sNJptOzQ+JsNaQp71s6JSpDH++H2BjfVZsHxoNfxQ4oTFBAUJZps
vsbC98nfHqKChgbN7BGcn07/E2cpQnbXlqgaUCPX/PwC3kFjjbXvKZSmmWM4OWmsSxjsnyTxwuJX
y1X1RyxXse75LEAaDFaRSboAn7Xq7fzptlmSXXeqag7RKmFLGz0MXpgYo97o0Lsu1iQC/c4CZMCn
vebFvh7WCa6XgS+Ggsh1bC5AYM2ZH4FmhuG7hPw8torJLVnxR6EqFloYK8yvTUdgg9U4Rvm3gIrK
u6xO43LEcg3s1ygajcuAN8EEYUlUeQeLLm7DxWTgThGWPipZ6Tjjn/AKlZ6taeUpZVVd3g6BDzOG
qcqHZs2mzSHWPszBofk/h+utz1Ad+LA3fooUgU8bTqc+y7TY0YBqZxRqKzIBCqvOFuJ8wZhMDXgD
zw+SAtYsj/1Lp5qryECXE34T1beEcuwrsxweaSlDc0m1srVrfuK4HeqE3Sht6LTUCM9b4sG/acVg
+l8pNWrX/Eoky7zsRQq3WR60SpbPVLZ+ZXUDpgR+0NFAF5QX32Qu+c4VF0aAkKM3PMbuHGtMgZOx
Ywj4mdWu7bNzo+ig9+qvRS5ALtgi5Qc1VxL4XVNBq8ueiHW5f//fryTv1v3nn12jPHL+pE0xR9RE
TRYLcrd/iTiQELm8owrsUvAfa7SzD2pRCVFhiwt5MJIowNtwt/o5gEw5WdCNHIWq/JZpVJWj3P8T
JMWxV3tPXfZyTs0AYe8YY1zYOE4OGwrYwpH9W0pA3leZMb1opqp+UeSBiZxLUMhkLFgvkK7KpPyG
8IKGp3riXXKli3Q3SPiz08DKNdvHW5MljEWb0QxXaxx+2RcYeBdIW0lmn2PBrfBePhpZPfHF0eMK
iQI/ClE2TWBxenL7jyiwZ0VlO3AtnAE83Il+7cEHZ8Qgb7LmJPaHiCJXS+AuvffprJWlcoojOSls
R3uxDUlIKSGN+pLrzXDsfO28bLPnESrdyyfTqIfP04MmCPdcKfsZXxSqGn9sPGD7QtkI9AO2bqEs
KFTf+kRld5SDEANe2pEbaccbBjZl55DZ2/5VgrCQVcBiguZ0pTqgbzvRcYCoqYVlgp8xKFtSb5QW
SYVm23wa9EaaFlxanUIJxKeNZz18HZOc4zyZEW4fE5hS1XrYVPb/vcqUY6G6DX+9y3BI4YtHIrab
JFOAI+fWGrKCYr45JMkLVhGKoUv5oIqVTLFVIrmzlXMcOr9YPQeKtQZA/mNB/g53aIZMnLQYsCuP
nvPRzqGT6HE87vyydTwzYJ8NSa2QvR9mM0ZfuQ1atzqdIhsdJI2KlXZaOvmb9i7A7E52xn3bNiIo
HPVhkX7WCs5EY69+Yy9OSG88JmQkRxxjUYHXBSww2KYEZWQ1YNw4G0kRBhaJ2Gz+znnMbPkIWTwZ
PKXLyVgj/pVEMHrjerbLFuuWN4nFieHkAOwV3L5oMom0ENcRM0Z4vEoAXcgYmPUR/AFIZP+6CcHd
0X1TZ83akMPz8J6M4faWtefgOMNS62Km+5ep8egWI5Q799m1EZpKCDAmv1L01MDhEd308W8ly6NL
hmDM6+IRiOf5iCPf93NDTC2od6ukrnsxxeFuk+J6T8L2bUtz2MJMruuBHSiGBsTr2IYlZSiuavBJ
YuXKQh+Ra9LOJ9JjafkslHulM6gRoz2zhcq7ICkmguH+avQwZXKHKP0hxorkos1TZqIeZcAXgtQP
3hpzPSjVgbY1+m9j2dVT5QaTvdfnREVfb/c9b06hxTIZ2hfE2n37G/kFzXHFoUOmCgFnpdsDAijA
Kp09zLv0B1iMb1fRpyGJp+szpAb6onoSMlY8kKgFh3AU3dnO05ScvZyudZxcbhbzuFa8yI1ILdBK
ABUJw1qKFX8j+GA5zvCpyeCLX+O5VCOi8KQTz/SESEdXUiWeKq+WWkswwjJuqcdpatakapetvYAF
xgle8DpFw6C7PDsOPwWqQY8y05vMNch2qF6w6YIaKfB1hYkY7jVkTECVBURG0oD7an5EjZc5gPxM
Mw3iC3Sd+mnkS9p+yhWXHK4Qqx2VpO9agGFZf1MNtjhUjqwgrDdT3vJi84KBh5RFbCCd/EzgcQyS
iyCwkkbkBRqgysy3JR6hc6HWGgRbKOf5D89HujZzZwFzDfVoAKScezD62EXrzS/72g8xeEi1xK17
2sUWFgbTzFIGufcX18BTICumTqPB63G4KdlDYIajj7h0kZRKvSbQLincNGrdq/+LmbgS3tyz/2j0
q9yOhddZtMFE2plAfXGiGVvezjhx4fPa0bAKtsBDRRzI5aGRBO0zV8KrRgVIXrJcsHKASdTKkHEh
/BWthmrojHvBdOqyHYPfr5t+Po25rXlNzybQIcZU6Bw/Mevg7SXvWp7E+JRutS4bUn2y/BkNQefR
HBlQwMo8rjdnnO29y9hv5++knq2SGNMoaDhilZSU1534obgc+XgKKskrSX5qLspYSmvnc1qOnhob
ykvrP3yNKGiWKfcGq/ZvWF8olcIuIpSIOBHiGwDS5YyQvsfj6ORgckPZrrc75WZBjHULOcSnIqX1
49fw+tQ4ksfdmRUMYoNfetQv7iwxwL3D51oKjMtZfl20QhsbawdMqwDjMUnIYZi0obKFpxBfj/DH
L9esOhx7jFuqWDsdp/fOyZOlNVic/23nvCMCbNxnOLTwkj/qsUUCMPAuuxIpqiEAyouwMOTE1Oax
xhQRu8fgUQVxWH6wTr/pha3AQyYh6pAJp8rjLMNMWWfpq4yMj3PvOP1KX6/3YQ4beGdT2zwL71IF
LQAuA6WAWjjhr4uwFmpD08kN1ioWt6O8ag1VRExlQKMqqiiSFb/KOjm/zJLH1sRHCBEXATNxUkT6
RnJh7cPkV3mFHhqBq/EhMC2gncMacVIa/R4ap9Qa2LU3nR17UPaN4sFKnRhphw3U3P5wnRuSTz0q
wkYdEuKIRnw8vNKFMYFG5qjQY+gQHj+fKbdLH06VK9nEFNQmr2wvdtvnVEEF/Ftlkwwe3O9svuWM
uaGh0RKBR5RBZwRtdLy5/qtquhmvfmSxajHou/yvJrG8XQLUUFGj4xXsMPtcCrHHOJJbwQuJeWp3
QbMTWqQXMOnDz/Z4TQmE3DHifFR/upYZftpFMYrZJ1gVUwcdwQ7lQA/veZMDX7v1NX5qioQ/Jynf
vTMzrVEWJYPErM5MFwe9BGuIGBMjljXP0S+bVgoLAEbjSS/zZviouwH8ACtf9ZVMbY+1z+WBAVgF
6R2U8PPIEuFpQbzjgGVbeJ1bikXusMIeOCm73mNYDD7JxHEpeca+1LMir+u2n97RG7r6SYeYD2Ql
oIbUxo3mDUshe660kWG93tTVasan9NH0FQnrvUYL8fTuHtkWOOVXXYCgasB80jWcGKJ7fz6QBeSJ
MWUresFOjBmufH1EqObc9z4CdDVYp+kL39/kgmQn9Ve/d/OCQBQ6UwkLcs/hEcvPbpTj+ZzHHTN3
93T93V9n688/ibeifjeoH4sI2jMGGkqAoQkOqvR+NNFeoCOW6dHcOmeo7+jTL4sYyM4GYGNHgUK8
imyh8ieTFRCP+sB85etXwZ3WZLMfyZx011d9s4MY3kTHvF08ec4ZtTGpMbGsCWK0yrvhenSNh/Bj
PexzuTpLAVko3TIb1mRCNwGhnUiCv4zGH4U/ADdRdh6LRybsKGvlQ7l/JlT6tkggz/wcNJ9lMV/L
lYew9eJhTeaFYgHqCMfMOnIGlBmUBuEbph/OXWC85jxIX1QMCYkEbwppfMMMGSj6V5YNnDmZqLb+
WHy3XvThHt1bTLxIBWpq1eeZcXAwZ2iotEau/c2BHlUcNFR6lzo8mgXekP07QKgZffoSLnasubII
uvvSgV8OXxHPFObPDM5k9+IQdlwopVnBJdtyzTNh2kmuCdA3n4fOaNDPHzxg126Zp1RULQf75CrY
8hz2tJ6X8C0gGPJH4xlmAFr4bJQrWMhM355QsdLRzDiE998GMZajT3/hvp5wqe7o5s3zhbrbh607
3O0i7Ok2EtkTvaGasi5xWyzfnx3yFeLV4na2tPIBXYp/ODRhqN0JS1it8V1bMUExl/wTKDPzDOpr
Hw9iJQI1UyfLWjH26szJSo/awtpM+NCEkC5VptogPiNEgQ5hu8oS55JvqZgGfqaBif/ZUM+YZ4yr
gFYTOIs34ESGQB9jzU3kxJx9LNSRwavuQ+rKV6ku01DXHOhP4HBiZfsNfK1LZhIb5L9/w4EiUq3A
kxjYKvaji5hdvKfpQvCoxm3d/AzJWNoCxfCBmIhOiOY697GLFNfUNaeY8AMaUGSK7LXoHWD4/K55
faO4oHLEghY9uUlfXIGoAspAyBqZ64RjHwXYrOQDTll6jOT8HQVzE+S4WgNf4B8NYmAsqwV14B5F
evy3b4pti6P4XUA7PyoAsBTFWrvqaLcxDZnVhwL14spo6//0S7teRjGvDEc/p56yi3/frd1dBHFm
mSi2ZiS6I8bgoEmP9Irs0MuTEaI6IcyJ5rXYFcji+91dUsPrFePvFg65Is0LdZs9dwCNZtb3QP32
uBe2vByVMY10wSF6DvfuVETqTNtQXelb9IZo7fmqDTRO4ov/t37EZCjTq4Bix60BxGqDTnlTzoRH
ybBcFbiSsZyuy7YqhT0rOK6VLmV2/6ouK3Qk/boCSJc0kxrvLTNxiIJmWC31Dta3STCvjB+bCQ+n
xKTV7JjUncKycUs0mnm9GsewFxVMsy76L132nw4LRKSTmCHgIK5Nf6q0OgaPW7VcejgFGtejD9Ol
fPZPgiKo/VbcS+IgfbobwZ/sbhOFh/1wcHha+NBuDWOTJjccKD62AjkX2f5F98+/bipV4CfzAZHz
oUC8/Ns++MsJPgpTDbsz88ZYw6c6yRmhefNgnKXwQKZaJiy2HPRESQ67fOR0raO5RTvllk+BW3qY
zrqIpAmx6+z3aX2uTts9dpeRQRSZrd9zQHFDzaDWkrnEUjQgEJSXvOEZn5LsLg/jagHkAKjIhQZx
RMdRm5/6pvR7B49TMUrFyVmC5FHXoiT7uNXhbcec75XRsiSfgxy8REsZxO0pOsRLhZ4y7udG9xYT
OonQRvd2ybhgTZNMBPFokDUJGRt7Gj6vE0j1CDkwBVZNcSR82MZFg+kJxV409EkjUCXW+hS7wUY9
qJRvrCdS31CjywyxGkulKr8+t4CUGbYirzWtBRwjYO17eQpA5ItVTmVK5hJT5K7SJKF3Iiryo+C7
mRy08INaWEAHhoY1/F28wlrZC7BF7xnjK5raCPE3QVG4rocTFAlVcKVk9icjqF3klzy706Q3vrY5
v+GoZnw4xl10ZnsS1jqqm5CVtH2yGtVAU3pFV7bshtmJVi2BtTuZhnNXQvEl0KXUWZrYKZ1BEL0b
KjsgkfW8HIzAChvRy16zeDSwsOwvaAfciOD1Lgm5u1ahgJ5c4WS8G/GMKvJGkaa5QkPxzBxy7OU3
PV1whvsey8Al8+qsrSzpEpKLodvw/3uB01ehuNkx9+6O1krL3b34w/2SlJPufHP2iguPHsteVHCq
6h7rXTd+k1Ze5WJ/50v+Ob+DmQYWnYvsXpf16wfIXbdB76x6zwpSHgKH48xj3fear3/YuTu8/nwh
zI3qhrFyYQ34PH7y2VNbuvR7UtqqawLWfkWSia3dIK1r5J8I+4l8yzcyhkoRql1nJhjYuMV72iKt
P/UTzwWPATSa3tZffzl3F7vls40AVJxDXRVoov/pVIgDNi3ZtNSVTu4mErrTZENqy633H6Rcmkmc
Sl9NM9bUUY8UV07SJHnuFgo++FMUUmldOZLFxJ7qWsV8d/+d0CpjCX9r+Ln/l6kHsy2QyE9yACm6
YsN6PC9nbPRvA0nzCNxsqMt5uG6YKr72s+fJg0/2L7wP6ojOzcHF5jNGvPtYbyuV0+fEYeXrun8m
ool6ZG1h79fvewfWuQT7YPUnlAYuLjj4ys4JXTPGDoCp7mRJhQ1WoBS1r/drTEvEocEzEo5OdvKu
dCzRzMnJYZEPZCBHbmaf6oNKuOYbMUFyNrtH/gfSOqfW3qyEWFTI9aGeirR2GUSsWXuiTIxr5Vn7
DG+rF4AMj1xjppdYabxZ9IZ9KUK7BDuMlt96uE1qoVd1HMC7pi8IL7Hy+1J8/gN6g8JjRtBFHiA5
KMpl86L4FwZgzZxi8V2kiqpAMiodpCbXz/skQlQ3YgF7SOH3BRfVz9nF/RlH9g2o3Qi4SwMPrlDS
lykeAkz/pLO29v5oqoozSwl1Itn5DMLFx30+E564Twwlvmcoi3oDjrJgWWFRIqS+117HeL1hBLG5
PSibRwvDMVPNMmGM0uNuQ1R/J2sQ7/oHidJnhwmXzarVKayYscarPF3TCVecdgXf+Qr2pja4rUuU
OlRQDjyMxllrf6VHdcu1CLE/gX4VaiFIHZ5xwi5cgva6gzEgn3Y7w/g/yhg0x6hMmQ7T6Lyk8wQV
Vr2r9qvgWsI/HhPnMaeZEUs/VdgEcvW+Q4fXPFRrZ4V6/bYrSATaHt7yPQf1ogbZg18S2pH5flvF
cB+Dbza+Hg7Lc8knr5A0AJ2obzaiECxdizzoDHHrPgC8Ayys8WyTfueXe7c6NND+FzeT00eCiq0K
d9Yh+4o1WSeKYExc9oB53IQnU/pY/WBcPQ44f826DYH86w9tczYkJrKSggV/iCabYfSqYyXLS8xf
dAeMioRLFE/EJYdE0EU4E6u1Qv1GnJ4pJ8/khfSJPmwxuECNjcUe+7lnkav3RiUKgQVjRDtU1sDk
nsX85gQ40Eq183ANxfN+MwoBpgpX+2npFVhNM/X+0e4ODMVbwjOTcogy20qGbcxLO5lyn6kQQPyf
O4pgTGCcPYQW2j05DprDK+7Kxdw9U2oy/uoQhb8zW76X9jNtaZ/5DPfBy7GZbKzZsIpdPuRc4bMQ
sg3LUabWfPRKWDXc8l+masBKhua1Pm3hShfzyMlvHMzs7WwSCMw7j1md/y/e4btwHRfAgnpTba0Q
Lgfa1vaBXFJ01wwcA0x0m0PljQrfvZEWlqYI2OpnV5I7MrCGawObQChAPH8zD4JlwGiNX6ssIdtX
H+P+6cwiD+AxiwWwV8IOP448DLdY3g5Aft7TXnKyWcV9ZDpX+R1qUPye0NBVBAj8RyCDXnr9c3hD
GLkgxzHJVjYvZ2b7xVQMif+JVJZ3EISuPzAElUaG/EAzu8gx176ptHTdwxubCtIxDD+5sgTVNtDa
P9DFRBNZmkuIIkfCS9x80c+aikum80EjvlC1qXTQbk4RThz2Sb5awdioRKzv6yKF3dnMhsejr0bZ
z92/UiIh79TLk9B3NMuwIDyO7rEi+529PTzbHwsGn6jszQqaECZQy8bsFZgu6VKBKyiEiw+cYDAn
ew37Xs8HNOqr2ROp19RlQUHuBhQHJAkOiSed19mV+tszQy8Z3M/ZCNewt5QdRt4hYaC2gfvOjZi1
Ow50UgaPvjYRqMV8zSxnvfzc5ShgXKIZL9+FLc77CNSxs1oVUYfLDbUIWWqRT+YKyBnC73dJKaR2
jo+5hjKIpQY5bIUDrF/foXJyOfpB4q1kuY9MyzFxqCZNWcHJ4v6KDJVfNrDqukKwmSDqO7gHjj8p
taE3Yh9YkdkwdbvhMGobIs+fTuC848lyG7z4aq3Hx8QVELhl8IR5370m5HGaTCYLf/GUZjWRmbfr
X1rfMBAGmaVv0pcChQBsmx9ibxrCvBTJt0GaRQWxiVY1Hx0KRGMybqTCierNZOknUPlGWfzwa+aQ
qbwI6UllT+G30AC/f/LX/jDt06bmRmLUXbIO0MBKLwkDdC0/BrC3bsahZ6yK/36I2aZ/o4WfbMu1
jJOAj+DwtDBz49UaajTRegNXP+fBdY0wOIz9eulNEsVR475WAUcB78Nh1t63ZK0YuE8PYPDshpSF
L5s6GHw7FXg4LUKqp5uGHCpYrog5rzQdib8rMkL+dWlfaGebw4vbcPKwSsNxvNwo5cQVkckiB3Jy
xCmUHsM4cJSaPUk/d8qEsqlufn/3JW19k4Y3u0AUqgEDagrc5mwvqZNKQNOpu4lmjCKGlqRwu8lH
H/Khw7QRtLRAzQcAFbp19vbHQhG8FqOw+W/GRZ60JaBWp4PIdGQjccSn26vzdiYodAkKxcCSDpKl
5lcgj08y9bZ6Y7Nr5quq0ED60x79IzxdNJj9AApt1mlur/P2WgpP70VmJaW/xBBvyLZftaTemviu
DbX/4l4OPIHSA9FmB0Nr3miTl0p7uVR0/9KA28fM4LesvfI5UPj0OAKtzfkAcTxDzjEfLmfyITV0
i287StuB4FjQhXJm+/ME8UJwbqmkS267Dy+FXQwtCB/5HO6N/2xju8123GyazvlDKZqQx3JEvQVS
d5WUWS0LTeHXffU+vfeqmLc//i6Vog3gWbXkHwWJ8RyZK+7WTg5tReTy3Sfrq0If8ap6gX9L0llR
aMLECMHHDl4oscm6s/NvAZb1+3zAKmYL24uFQQjxdKl8p9q2ac08TiufuBnq1Ez7XG1rjUJLHwNt
9TpB4IdN5Do0qvA9YPeYVJujPCqc+XMT1rQW6HGDEF6KIEbAH7BfmkU98qPpMz7dZSQGJP341C+d
Fp4KTYlglwAjH2Jatnamz5DmD6a9lk/cvzGEaZ8nbw0yWnUWIHBgvGqE7/o81YCJbIc3ZSwd9u04
guBsmv2Emvpx3jQra9gocTC68pU34CfkbRvqxYHhRxse5YhCRjG0Z5GI71PpLEmYn5GTw6CvcKZ7
TumhiUD9Ce11Mi010YWjhot7N3Sx5J+Y4VXR5vqr+qwTiF4f2v53RYdDdjHiOgqxSuXBrBKOqGxP
Dl/gWj2Zyq47xg64RAOuwsgDOuaKIrulHBXanfN6gDfJ0hok0WhDOixejG5kw7Xe01saVY8uMuco
gk6B4yn/18D/jTrwqlKz9Yx6Dtu5xNmVy3OUPiF16z7lTTc5TObM+AyAvLsrjaQBSmSu5YV3zQ77
oxoH5UtorRJ9eKQasKciSbHI0LDg2gVKdIkx/JSrwd8lGILEdG9mcuyvnMP0sL2WTKDY+AgwhP6Y
Ohgxjp+k6yjAr/sHBrwOZ3A7XQ4dvR8l1n7KU91mBX8YS+zXoG0d5nTWmt+D+Hrb2pXY16vhQwun
AHjgQ+q3wigXklc5NVnC7SrmpkcXEuqxJ0fUTWIJjWcN6eNI2a95k1BP1A1TWog7sp1OlpqfISGc
0vujdmH3PPDYpJAp17ROTVL22fAdXXH9lRKMCJCKtBSNkoNCMy0Q4p/8SnzWIHvrqOgSeyRJLGzY
Lx/zXdAKHK4Krb5ODwLN/UfKlzfjEw5i03V3XuxY/A8gu1ASNgwLeTKMfv2w2MgNSR4oegr5v1RP
VYYxkZLdu1EcPXqNmcHSsW5JLxkDfNv8GRZ9ZX/JODMka4uwxYhxA4mT+arrZLotZlAwpbiCp1qT
jxFkx4NeyAqJp6i5T6kIpJKnePFOKj/mcx4oaLDY9MhKugRGtshRRs0FoE0IKB63f5+CtloagzvZ
1KZKjsn6kXIczBKm9eTmVTCwEF7Z3XnfA1XkbEqINOoFTUqkerfNnZ9ePp7eCYMcfB9f4H1dDQ0T
vB7pA2ExZk2gqO8bqiWBfKZc+KKGyU/oudMDWhnbMMVV/21fp+dh8CEH6AgoA2t4O6WQW9mPIpMY
mV0Em0NQtQapv/11qychZCyb+Mj994FUYovHEWv0aSql7GPBANCDKIIvJYnYz98MsUdz44q4SK32
XKFpxICnA/kwNFCIq5kgudIlGLb0mlrccC/R/syIEQFw65K5SjYMXyEo5+Xt0VpdNehjl9vrC9qi
OLSmZwJgdqnXsrD7VLEy09rVaOUblrqtMYY1W4mUOpjFd+OD2nFf749Z/t3t0v78PsZ0tD+Wgc15
QH69Zpr/VIl3RJ3619TevRR4CiNCd8g2ch4OaEYcFQrHuNtS8PcCIJVnSThFSb5Fhpa3nl+ttgzT
Y68Tf28nqXQV4lgq2uRQt8pTGu80+3nhzUQycyGL6KbSUl1MbDAdcEV8kZjaF7WPuGYKIYPKBkma
SUeqnBXQTKDikuu7Krgz81OByeOV7Bp6rj/nc1cKIflJGZpoRQVUXA38LTYWKK3ZsvACL4xYthSN
gSrfGd+Y9FoHFqy6ES+aO/JNKQabBnBI2O3PYBXFng0LuJtBb5vcBxo1j+fyArKc/KUptP8fZ0BT
E8xTIHeFvJQTsPAJZq3zhaIx+us9yLQznVuO6EUVLjnZv6jVxz8ksuMqAl1PESCyfp9QxBhKZCR0
RekGlYjxYY787aNokuWKpTg9/iwI6Oyvqb2uw0RPiXSsRnpDjwm+vCXWdibxXjEUS3/cWbS4SqaV
aXmWiuV/dIQj3bRkDhfPmZoXNWryn/KsW77eboI8lB9Lo0dLq4iM19ggCugbRLbGCBvA9cUomhJj
x0KRISHEhvYA2Zo3joa28KyD8veGXrTi0BcHuaCZ5BDIFgW29zT5ZpO7k7p/RbYcgA+AuSkTPAMn
E+OpDYTwldc3zwWWjPNZBT0LoK93YdOAa8MD0gaBg9/IgqIJCgtHgMlkOFLCarLIitPv2e5VettA
fkPX+bIlfkJhpdpedm5QLcr2DN2cEV8kaZIik+Lac3T18ljViebaSSKd8agS709gmBS9ff+ji8R3
J8VkcV6yi+USbAFKBshgfPKR8aumRRoV0kjMk0t4GHohXZkS1fLIQshn2eQ2b56ggFzjYmnY1hWL
znvJzpqfRd4xX5lDNz2grNWzvCiXwZMco0BRFdQjjHgcNbfloYAqD13IghtXvbBwfpolHp4kVIng
wKK2c2FgETpKpKSupJ6M8LS8x2o3nZgkPwdtGnxC/iVlkkhPn0UQBYUCDctIr/qZOBdiRu/hNRbg
fTJtXP/DEzDj1qmi2myVQKIn4VYAzwbkCYMRwqx1hfbuVFqm5beB4fku0aG5U35s8QDq34lOws1W
TOJoDUj8xrtE4XYfBPC1VPxR8UstXULSrD6z147io4fZ/x1hJo9k/Jo+Ab87QOTR3VM8A7gWhtwc
CqD7JqJLGhgu9d5SBJUR2bIDAxWTnX197xCVsuKzEdcJEjFbzLU2Vrv1+SGK94sHLpKQui2lINjE
QFkxacts4R9bQo+YIhcK4qBTvvVyQIPL+5rZKym6QUyXD+ArmVan1HTrjzYXWu49IiIDurSqZ52I
QLdxe50Qsus9sQqUV0b8fLiLema8dkKWk8yxJwZSim8HvwRcrf8y5Mugjl41LD8i/L47ImOWy7cc
65dO+PXsq+ehLb96ilUCF9pBCeFT+QrwzLy1jD+CTp0qQ9rXF1hzbjP2VnEfCIor8tSeNrC9TQqD
xuRAMpkBBB5ymi7GFI6gObB4KCODpNbI9RG5Tx/YNQEKD0HZPnpCMvqWrLgISoj/bV33i2UzjMx3
dffDcmVChWcT1p32ebrktRy2qdaIa4FNZmWgHjcGDhjQ07NxHVahBTbHijlf6UZiRn3l33+ASlB/
+bDBN1Aqr4yBe81RYcSeS6FaYwHFb/qnIvdUMsjBvEYlfGT2hHbpu/RmP/VdZsVftDiZhRAgcfm/
7XY59CJ1uAyv53/t/rKLg8ongxr7w8+2KJ00bTqJ/yu5qA3s7oNHnyzBLwwdIYOg9eQa5RrRavgP
LuptiI1Wwkg0hoaLnxcSW3hlUkdUnthv3OEon2NLFKPH7pGLwgpL0T1CLVATbPIbEc50t9H9OKBn
7sChi1ZuY4wYmq+H/XFtAlW6iUnKwoNyky0C6mti+KV5lEuwZdFNK0QdZO9RuIBt3QcL8gDoETxJ
v3MdW65Rdsmd2OxF9B/Gn0NmMG54TCvLJfaBSaTgarJiZWpry/Bsa1iHT5Cb9xcFy13YLB0oQkNx
CpRBf6ioAjhZZncmjC9FZTjeTc+t9NQcT6pTuSaFYG+b9rWRwJF1T7iy+MHBYya8QH+AZMA5U0t5
K5iV8O/Tke5ngq5xh5LXHzyvWM9VsUtVu8aR4Nq8VyDF3RrZBuhHZqmjXWxV5PPoQjxzFuswcshS
UNDXTmPB7NRHvp5klReERsfY9Jo5OYHhbK8YxpSCN8CBXPSuWFYZREde9kjoes41AqJV/HMNfI7X
PwQxE3eROT46JW2DPjWyDrYfhQ9utuw48wMeCTrUqORD8+7y3A7zhok50CQSBKobStn7ZHP9oi6N
HQcGIsKhG5dRL90Ve3uCf2uPckwTjfpz5Uxlf2gAXsbeCsBOSh4ENEuNPdcPlF3lMzOy0JqpWtkO
lTCkLj0dfn2t+9gaya1Os3Lgs4ZDatDcLnooSdApjYAkO9p5q4AKtFLu15olmhI83VQmWYCtg1iA
RmhYk3tMnoDMmmNrmQMmarz8To01edoqiGuiU4O8wygJm9gPU7we+Nn/2zECKt1VGQfpaOy0FUfl
+yGt0M+YkbhBfZDESXJ2aYtv79rVy/Tf4NgnR9WZ0nGW9aAvL7Zh7S3rmtlAyfIPr6X5+m8TJ7hY
HLJvIxd+w2bwZsVRSEshF0S+5uMranct5G4y+rGL2xyrijsIgUDG00XZ8gbH4qxEb2GJpq5Ri8Da
kSzWLsnF6gxca07ZSpaYaqRmQsYpS4ACmtS0KxlLI5s3ek/QvKRWY3lMxUIaVw/RuZHpkhwpUKeH
oxKk4I19fWbRHYayJQXDoGbgZawjoMWbf2KInS7DKmcU3JWKiudIowceb13g7k1/6+8F1QeRlytV
JyiUh37ivnOpkxMHmuKAeiWCduqy2HqD/SiF/B+NwQsGdTDi6T51v2sX1xHBEJXbPURg/k4GaiQo
swRzV0FLJQZXCN3Q/mQxD2E6J6jV6W2lqCx6KJWeFnFmZaS2e2/IlF6isLyRXLUireBpTH5XjXU7
cf7LZAs2rdifV0gATiNUmYd/bkp1ofnS9rzvq6Wa1MDYcqVhXoD4qi0dm8iT+bbkrjh7jyp+fycP
JV7+yLnM8E4bYWqxH89vMd5TAFU+ursT+dFIDg/yzFidiaONug8oeziSmL7ERXL8bhOfhVJU6rAF
oeGCz9KruR5sCxzcHa72vYN4oWKLuU1d4j263c1ckpxSu6BuvTSPfLBf1w0AQ1l6v2PU/nKbZvEM
317FlZ8LDovXN8qnv2j/yEHnntZfFi0WOnXYDt4wN590uCCo4IlgHeduqNLZo80crOo7L9uGtH12
HbPuDJm+UgVF66uCxmtZ9nXrnhRnkmmTnIpM2s7fnmhv+nlAmUZZu6nzpltYp7W9rQBDrQJEZxAl
pBw2rlBgX4ZXetNb8FbLnTsYO3nCWhRF7B8LfNuJYAb444jZUqsrI+awtl2dbYfPTIvBJ8E1G1rw
DtHtW3LRohAPFK+ODjzxmeRCFWRkY7196smV9lx4hTaEZ7DGsaBHr/bPjKb6/qpVf2snS/0P42Ij
+zAjZ+xbSTXj2T3vq9KkfySUHS+iCQVljpDTwOqIriKiZ5OJSFcA28/lk1lVffaNTe11C+9QCTIf
6Ng0IAL0b2CN019VBoUtCoJLI6ek3EA5RWWeE0pxLgqp3Ms79LRsID6u6uBsofIo+yRiPXaiRXWx
fLkr0yRTD/sOCDC48aPdLjDncRJOwVc3tdmIO/kTLJeish86auc3GJazuX+fCXKwtsVd+P5W1yMB
r9w+RxS1CSinkPtrd6f3fEo7GRCpaBz9Ibzf399Cj/Kx4OvfQB+KqGOeMOwNmM5TN1gYoFzQYjjZ
FvhTwwe76Au17WivvPpm+4AUwYbI51IUUuJgodDes5R5q13EhR0LXrYuxRFifdCEDjpg4c0IAUfe
xmC0Qj8hNb7UXNgz/A/QWa0Ps/Mk5UCkbM/jSIFKvgJPWFa3oOnJ/q5a+Yc/gM3MdGNf7qiUszqf
2N3Wyn6Xkv90di6HogxJglJ0uN5m0y2oyT8eUTgYSBnYvWYW2SRHqpGhDHUVZynklerUOZsIjTwD
AENcZFu3o8tSQDlk2z6RXnJI2+DWvUIpoSMo7MN1VKqIG5a0G2CMlYSI8hpjCXx4UMHaErJdLOBC
lqw5+OS+D8y1/TCw0xeHr8jVDEzkVN5pGdGuJsbKV/ttKlNnVkXpObUZcM5IVD/N0IPD/vHhjK8p
740TtDT8/Bp3i8IYLRPLclF5fLHXFVFOnN+tzzzJgs/eeUGj1H7/I5UODjERiNeZqF3e+HbqlAZY
3MoP0CwO4dQy3HjnLV5Y+VroGfb4FhkINhuvvDpaJBppz2BJBvBqeX8IX1ELGH2T896otlX6f9T2
wwyrkDrcu+kDfRygN2T2/tiZ5Fl5bQqsqJDA9lBjacUomxzpa2HP1IoH8T6pVkEM4R5IfeAV58h8
yXJ9U81B0B1xMof9Sf4g8lCEvp7TNBUOzKgq5Yn4u4OBIJy2/fORxG6JDK6shaGfRuRhDoBj+8aF
4yyGDpKhWCufLSkjE7SOCp2OsWjkrojv4S6ukmPmWKGyq0/FmKfkxdg+oR2o7Q8/47W8l9Av0lRa
hLRGF8M7z7pWqfqawf9IKBt3yXlaZUL/+z9kLzGcAiBEppH41FTzEzCPwz05ZmN1fanOratZA+n1
sLp+MSa+ReZ+R+e5Voni7oocIjnve7BtT8j5+g3fiHsgrVchPiJO1hqFC5pZCfgmCq7uEDNrrYyB
1yQotgsIIpsmnjxQZYEjq4VrRR1M5mLb4KkQaJpDyZHQWXA0ePIlzhfrUrvsOxTqfl3vaBs/mPbh
yM9icWcUMA7ElfSxbpyMKDLIhaCCyZ38ioZxLbZjSdceeK39rHKNr5FBGWert78Ra4dGtoGGMps4
6eARzLKYa/Ov3zwch6ZzClWLzxSJvrF2Fbl3Lc9JaoBDDmH+aqKla16Pv+bk1LYGL4alBzf34Tfw
ztgREqGo0QQR7kviTv9cgCRjP568aHxrpGf7/I97o9/sl0L5hfuFoJcgTMM/8SwxZDchZLl1FoNV
D2eGfNV4TeOwxaU6GYFvnAV/JhDWNlOgUQVLtxhprdq7Wysc+lyeV1/fjMvf3vlYpQSHTWKr5Lu8
+mUKHAot6PdsTaOpV8vw27OczizwuG0teELOYU5WpXWyPRcVqY9dlfRdgQZcLRoj/JmO5za2FQCT
HA36dn7PnaFSvP+6ZLyk/LJilEPOSLi6YzXa67rF5tCChVACU0bGNYij/usD+jxecHXr3WQFhha8
JqqZbgQy/fftzSqFaLqVji1DvTLTjhfP4/n8B64BTjkCT/g9bmysHnhMa+K9kVYeZ2Qa0H5GeOUM
H0DorBqeZ6QIZerU7o3jhfBrSzRmwxN0elEqGXcervbGIYDMbRRDy9k47UN4IfmsYlqWTGUwHgl9
Buz/iQSfe1Gp6NgT5Qtt0Xw+JRHOXWAZIyrLdfaPCkytFh0IIyn8O7PAF7zJmbX65qkz2dT62F6n
2In2BZXcJvkLLMkhKraNhR6tzOLfl3uuB4CaPj+TmKXdqSTv9FYldgvTDJ+UEbYrZhgFf2k1UrlH
jP6Ha8fcyLqncxWVCvXf2nSc3zAgX4d/l9Nayr7LSyDciUq4f3P5ZMcrY1YnnIEYXEOuhz90A2JD
XtiQl3dGhzyLo2ZvrvHwlbH17JLFxikAN6nKApwk5gNv/2iTHTF20oPLwY0GsDK6fAnPYrf3UIDy
0CzrYrdSkz3VswWWa7WofveljEKEHPnGlp6lMz177IFMycwoyAtH+t8qesTV7y5uotPUofW6Iv9r
M1B8cpE/W++a5yT8mhltOgTp7dvJVRWd99TPBRZW4tsXb0ReawxFVGmNZVPRd1McXOBkxCrgzji4
eKwkONahWlD8AT0oLFnT5OCpGTVhr1xb9DnWmICCn898pB/64L8KR1lj0JX+aomtMEZy71flM9IC
GONPz8lsknEhtjbWyVTn5oJIxfz5E2RArCy1H2VMeMpfthvE8p00J51+46ulkA4t31Dbzi96vcA9
l9KV3p3YkbOjGK5cEAPJyMSxtBt36I9UKGvxGAEtzy3DOQPSeA8H9eQgGqiF8uKWDuFjiidRXhiv
D5fw7v9TQzhe0L9TmyxZFnu2DNBO8n88Hyqz8cj9E51EpemsTwa6nK3VA/MzyD1HxMHNx30exjCN
KekIj5dzIOJeNp+YcjP56syTfVJ2MLeBH8HvjYXwrxGZQD8UybZCi2gHfFl3Gx0uEvrxuk1PHrsI
Y4rkvAnhnw5f+HNlXQz6oY6WJ78sqEM2i5GOGreV0gquIXLeTns0Q5d4MaWJHCXV9thQfFTpYi7j
Wq1U0tU5kRjCVnKzdEVVkTQrfYr2HVUehWUtL2NORK8Km1vf2AYdB5cy7uLEk5HFQQrgc3nwYI4Y
o3wk/NzqcFVupA9kOFs/CXKacY0vcehro+/CYS8l3WrK+4+9WxxdUhkFLM1gcuQcQEMrNJTYI6T8
bAwQwnH98hI3PV27IZSq9cjVoPpCLqPNA8V0+DaOjTiOEa/3iea2OfUHCmUWo0AnCc8RzlCuXYJh
znE0mBMzaJvZ7aIyEOFqTH5v9WF6ADw+namc2k/0ShzxATHcOwZmNO5fpARNLCYlr6oJsBKQdkAq
QygU06RyB5r294gyPiQDVaPAi455oahL3h5KkdCwS7yV4foyTnVWSeUQsF/0retWDltHEKSQJOpx
gQxqhkz29Fht6f1KFJBSFAcFNqtkqiqviHq0kPx14rXblkc65LbezkwTvZsQSz8wFiMgvf25iwwc
Pnl0UQzRAcHJwr2nLV3rqC4PsaoZ0UOt0X2pKTuZYixpKlIYUhnTFXM7xKDmoGvbZhFel1pFX3Z+
YZpYZq4PAz4BGBnH2tId2vWWNX9mIVqA/Y9BQTlNqOqDxMK3plp7Kr72Sv4DTAEcsy3Tq2AnDlBU
04NnYIvtoCUkGU9Mk1qM+y+irssOYbhEhVbU4zt12cXL2u7ZUKqTaECD6CPzrfyl9xYp/koStSxw
UVHpHKOUf5xUfYkO5Hx+MNi72kZGtjkkd9F3ViuS+YRbnAs6usACyk8jKjT7ogKUGRtkLLNCsuMQ
xsk6PuX18n1jwBq728dNwiZoQNm7BI88MZdWLQogQHfdByNJF9aQcY/Oms0yVP14kfMeDt4ZAmX2
4r3sgP2w58FK1VCO62PcOT1A/VYvgZhFmv19/7KofRgHs669R6pFQtd8C3m8sd5CrXAeRiuySTrk
fvOzhaDWrwbpXiuo76Zb1P0kFtelNfqCd+5Jla9u7Ol++UqROE5Bvm4XTxODAIFacAdFFqqqBqO/
sQ3udgpk2vIoOzZsX3O+0I/4CWPXiOq2A/nr5JVymMIDwzZ0XUxa1naDGPswFm+nQeuwIeD7jCsS
cE1ms5xq1dRUSctkV3pg+OZItPhVQ2975Z9eyt74Y9LfvxEungyzkGAvjItGh6MVT3Vf8zG2GXBV
r01ce066z5XeyZgyqiGFqm12OAnbmrXx4PwfnN6kUXK22Aga4dJkjzsR+tZCls+D3vVqxWFkcIYc
943g9r1V1ndVqcp9hiaGEMfwb+5NPCAmihRws0nfozzFjBMBqnm5vdq1nMQtp+w/j3pk1A/OZ6ss
xD1tE2B97NEv2+KGavI6nH9tekWmgchpIqXksChi0gGHVF0aSAE0JQeGo9K0YIeu5LdQ2voJnbJa
/8ISMVLDMnQc6U096IyliUtaseCI6s90nxiECixUNdGvJ5mwAENmcCgyFQPNMBe+2DymDGwnIu+C
g/x8o/5+IYekH8Jml8ya2CjcqzNjcUUtJ4ReFp09kO9J2t0MFjTPipayDlv/J/sMn8n92Q1TdvsJ
knYehp3iAoAxkOlWWLOheRL+Tws6beCEERtjnXiHHHP80Mi609T/sNp/Za6xfgZiD9SNE5AmO4O/
sdRr8BrWE7zF7p7XHyji7hfMBuvvguoz1eLgiUwAhBhLr1+/tCsCzlkshOpFlwiK6u1ajiG4Ic9a
AvSVQDbsz3A25RYT68EZDc6EXqRDcb1trHJtp7xyxMUpUv/Le0wQTJctHL43Osaw5tpgo1e57J3E
A5stmVt99eeRBS9EwU2vBMU75iy9yO8OTcnQFuFZuexiXDcMi6nDRjS31jHRWBdNHxDgdo97A3yE
bjmKGkAaMJjUXeONR7Ltd/ukU2qOYj+Poa8G2kBc5KS0GKNpQ61+zGuubsfvDsAnK0eVv2uYVYse
bnOIK+sIg8ozgXzcpB21v5EGZWRB4cdTfkvFofGWYrCFYGEhbduIMvZ1C2zz/LAt3qiBLmBz49WP
8paeI3SfW8pbyap6nFHHTYTIu4Hlt0vt7+nTd4nlQPhES58UERTnP10kg/eHvF/E/CHypTKW6CKj
7iJ3XvHIJJEOe1yxZpeclBRBXpnH4n0Zd9KWnvjnZXcIpNbLc4+fpWHOlRn+V/SrKOAZ3u7P7kg6
qdZ7yQZeo5VVh+EIVhj9NCT8v3I7HLAciBX8Q2MVVqfwv2MBjuCC8BOzhoBgRco17hOgDkrfkrYt
v7OUnXM9jVqIUZkl2BV6eKSYJs+pqzZHC3nFzWFIFBYaVighvDBoKbgD3vBuLJz39rH3gRvRRrYT
f2jjRYT5zbtJBiGDVqQVHJsjgj1ecfn2+XfTiTZx/VrbAwSCVFxnHxwknXRTVGkTonrNHUJ1GM/k
dr5KBpST9maNABpFsEfVvYzw8m0qBJ2uadu0lIAd0uSL+v8BT6+zXrGN/2ui0GHaagxlukhB5/5T
c16L6mMuOh26Or6GcWUrlslmLH4mp5Adz1NGo/YjJQqyfSjNpYg3wqK5SWEpEjuP8ULc2fxJrS2D
QS0HtmuZL8cc2L97I2AbWjOF51BV32WgKrXh83sbud8qZ0ZkOgtjq24AsuAlQVrLMf3PkPzvetwH
Zu2z7SGO9sHdcQppmm7oUrP/wWXFuK9Vyrf4ymLc6YmANRzxZDLn6J+NJKUF/H5RHtYkIfMDjs5y
6Q3atyGPSuPMBEtzBC1wRgYznN3+IT7jsgGG2C781pnRmsrpYNfdG9OfwnFHTKAnN7tsc+hGxuQ0
NY0RPqEb/cjaviyqbcTyxYjH1h2wMKtu9nhiRRJXknX+sRm3tiCTRsE4ADCpZdTDHcYbCTDHQZVb
URETULE+xlT7wx8kjV6jFk39aT2F8P4L9LHXXlZwiiZmkz8jB9Jyv5aqw2s2mk+JPvhDn95er9tG
ml2nuYU57Ui2C0nn5AXZ0e72CiK+0AwVRjrS9CqPOq1sMFsTKkdWpYZzNwsbIutiL1LfeviPQT+i
R3O2dYsgQWeFl/VPuHvl0YN5mzxl0fU3K721CWD88W/7bQzs/J7BherMxHLXM7yBKYO/3U3SNux5
KPKWD48hcY2Zl4f+Zabj4y9KsC0DVNbnInTfU6nxqhNjb457FR7+MdPDhJ1BQbdF2N0CzKDb1Pyu
kYNsEsfSIyM/pyuLEOtvLIzYiI3xNM9Zte32MPk5kdUSbrulcjc1BJPUK78/BnHE2Ifp4BkAr9dm
+dJbi3MW2DI/5L2reB/otuCxYvdgxY6KfijGuNyZpDWFKSrCSi2sUFslH4MMUzDUm9oVWCKdcBvJ
rbtTUNDFmc0ONzAaTtDQXoa4e3DKC+XRxBeuTOmJdwbKR3Ak/LuyKCW1HHESdCKZgy3YWLc6EWUP
rqsPJVX+pCr3o0xsVCrak41HUUFl4rmgKTFunVL2Dy+DYjSsS5p5gSa//T3zN3yZe8UBjTuPRcm3
cqKGcDbxbNw8zxamo2HohQmlP9DOB6F6L1YBUc+MK9radBfZe3DjeFQMX+05FCJpeTCkLL6jj0k8
4F2K/q0aEouMj0Lq0iAW1dH9hTKQz4yb+S3ETtEE33TrfqQ6zcDwCVpQ1G/OJ7ESmFfaFA51yccs
V0u+76lLWIZg5p12zSn1B8CTVWBevkNiAL2bo6mrPAmlSVmd5lugCJEEj9i8FSb8EsvlnbLr2IFe
iKwil2K8hr7FsgDAoSOxR7wkq0XXSUd3jDf1onJYtQuIrpXgD0AgEotL/NwtPUTFB58aoyKXrwz/
UtyNCEuFTKAq2xrOe/Oyagk4LdXuwf0mj0TCefTMkfjrjXUtm0iU2uYW4XXDYjD8FjpGvmPR3Mn6
4PvYyZ7rE6kCQnJfYtcZz2WTctPTBW56B0aFgNsDYVQj5UoIz7x/z9I7kY9Tr6DtX6ny87+okYpw
qpPtiisdvRUWQuwqA8DB8ifnwylzTBz/O7z5/JZhSgYoEUBJ3FPufQdl7E+9gmVLuRYqdwrUAayv
97VCo9HxsuI2pR8xcMxm+0orXQDczRaMNlC4jtBukLLtechcdAkx3Na6Sx9L/kkBuhEv5HynPPTC
Gw+5Rz2lzo2sm/NTA7kzsQt2kgkpdNDOgA0VGxrGNp9U3rQ4S4piIl4O1vzRXtks2yhs+7DW3H4X
E0M1Ih2CQkiP2N2H3ujEKgvHSZbKbH7jvyj7lcypI+1F7oJlYEx8QRWYi76CbI9JdbK+mL5fxWzP
amxhtF2XISxWQD1hHVb69yQJ3n+UywZcaK3HNKMncF/rnXDi0mYyUKgTiyuB/Yq9Zcb7g4WTuyuG
WlYn6lRnvZ9iF0RQCMbznFQPUfIrz9+2DNwJbMwGe4kwD6rMaxr21HtUldlzSvQj7II8gHqJ9ipu
DEMobm/6uAJ3TFRibs/eJ0Wz6tqKRmWau166onFlTfAg1rbC5uGc75zldxCFjF0/hraU0ZW+kcVd
u3dqHAPqlhJ/VkXCxjLRaFcL+bG1wo8CuGOOIbpaU5L+3SSfHvnbOrTRykqcBNwLDkslZcyK8Hsd
DRTTDiwNc45FygD+tV1K7cDJfLtOqOqTsvAgzeIZUT6spme93YMlVN7Gwzr0qumfPjKwZOtf+rYo
yAULjMyyXCotM0sMI6uMFRiTKd5mmwzZlP9qdjMm0RI69nsbrzj5F3UGTnFhROnx+NH0cTbZfCK6
k2tvprTOfmDm/Hpn0HeqrYUEcRu063uLmTm0SLUz5L2+EkAOqHUzscMoFYUdiIbcjEjja/9rkamo
AyfmGomON5XK3aRjFMQsCcy2NtM2Yo0kx5stDZunDvq4IOhkng7Lq0KqoKslZHkjpsLRhb28Cy7s
OwwjkFVPrR+ye1g/4uYHGX4SPmGUU2jMpY4leKsMECUAg6AQxGFOTJsX7rGk2v4eeQZ4rhvoSkhS
M2KeLfU9V+XjQ2WqscRULVW3PmAhNccN+ivje7NazwcmKTVWtR62/w0ggcff4U7XaZ8/dK+lqQ4C
HLlqnvFA6p3c8x5r7rf2YXniHnhkpvYQ/Df85UzzcMrm6bBDllDAM9+0UxhfRs1PyhYKysbEF4ed
fb+/aY5b8JpHo+ruL02DeEBC0xltVBEg0DshlHWFfNABh3GE/C2i+JvCEPA4Jts6bS/5Ayd6KX7n
JJVrf6+XSTShtvP5vrFeY/QDHo8wWOfbYZn+4Ox8zlTaxo6Ys9ckM8BYmZT0yXIh8czPzozDF7jA
XhzE+SqC9jKj9Q7OKghZYFmbwFTHVwi1gWZYg4pRYhHRV0MLGXouaAZWjKLW7OMtPukdOI57Mpc0
lrDJe+490YaBeADhtu20BlSMFQr7Qh7mnIKux4heHkT6yzjl3ha4rUdtPYmklXaY/c7YGiBvZrKu
QVEMRZ+i619/7/38cMSW12/9DUcMD8Y8Bc1zeF0UCbaqK3f3G2iQCLzLNhWVAFjSAQ8Uj0bs4yYd
RYIGHtTQAh8+g5Vs0XiTQV8g6DbS8QzQdq+tUaaKQ3sVfBOv7yUhoZT6r01PoxVldDssXIfFCt+B
AGX66Es6tZX4QOmByQJxbJAZ92pe3JjIbkn3qnBKyzL9c4+inMX2tqrJCgGyXEipoiW6ZzJo2PRm
PyQe6ZOwgC4lp3i0CQN7A/lrRNM128V3tXToa1WtKImShBjjjxmss1BWYAAPL4exslImWxrboHT5
FrUzsk2GlGj8eOvVd7Pcwy4lEK3STlI92AQ1xJXTz5XPkfNX0iSLBOTZWxF5cokywJGrNX37tdJk
GYzgH0l4QtcRrevxX0u1W1tOZs1XfgixbmJl64kUhpdaLigMKwydfcktg/WiGSRA8CWm9/NrwmzK
eUXPyNJtL6vusUKbhWZISJOQtwq8oH54HQiiZMhiAL35ufehBjnd18d+VsiM1K0wAswQ0dSrASf6
BNo5T3vLoTsu9AWiP0htuOUkRkNBSgxKjFNRUJCb6aELX+KZIgx/c+NYipb5Qyq+2od6jMZgSoaR
qYblwzPWLzz8I083I363fB1irKbQlATM67qeUtnRphJu0G/m9q9I1Z9tZ0No83cTVJHkvtaJF0QA
l0TWSJK/J5MJSeICHRk0vT+l+37OKxjy/G1z4LLlUklA8JGtvpCY7d5bh/KZeBOGrQOunA1TiB2q
tJNNZvhC7wtl4Jpma4ggEoYj8wsrG5sO67BhSpEgsbWUf9jziLvL2D8kGl8Dh3RAAuvl6IDZauDI
UZ6HQ6Zk1497sY9PqvxC1LUKE3o17YtFaR9wAAttqW5B/ltf/WRrf/BgwXqnPANWjc79WdA4ywDs
pADxcjU2FPvWWVjnDHZZRvKFp5clVub9acqq3aIClB/HRJh6wVsCOWZmdph2OG0wE7cP33Uy6K3l
d4Xfqwxqihfag9ygqqnPOpx27YzOseOUPfN3WUOfR4TY4ERTUF1PshHwWz+HB7dwr0UP8F9DZ9J0
LKRPvr+8AXJZkhxLw96Nv4bBX1UNHIdIWmos1GLezvrR6EzHRMp+54bRRtssmUCV1D4DBoARPZhT
vH2rk0lTBAPEOE80t5fVRLmGRzVu2htw1kUZAPcKsie0NWBODQlF+V7K0AdgipdZgRXBf65NEcil
KcIhYf0Ye86aRq7zW42cKXsRk5Hh4Pd7uoHkNpz+Bg9IVtZo0fuA8bTpqPSfEnLkjwGmh9JXiJRz
r5RGYdM+VrrNpBlmyXxZGHCtL8LChb8IKRw3waALwA2FtwjAkauHkETWOTkvfiynCkoUZH2Vg0Qn
dZ/BDo6KHH3ipbEj0Aw1ytPTcgjRyWdbk8kdSB8m7L3m6/wDkD5acCWIVCUpqaLZmdd55rm82CUi
rWIbud2RqQ2EwRcbjoi9IPsqPNY/zvnKScc9v2EoquRfb/08+Lm5JzvVV53xTxGMp1sRd7G9+VY7
DRg907E53VhJuBZVoMRZIP4uoOg4XRFESM2WlFwWf/8pyZlJm8tD8hk+m5E9XBRrVeeGNGep6fXd
u2g9L2g0tiJ9ezSMYfaNa8UFskR1ebKmIz0VzQ7vtTIqdE/cmWkKIGpCrILO8S+JdWvo0auDEXKu
5whdUC/3RRvItwmBvDxtBqloAQBKFT9uyEdpJRMNgKe8NAHOWzyHs1iGPUu0PqmOHXK617UemSMI
84Lbr9+xhcPWkaWsrcbDVUKPqUyGN2Hzz/d5oaJAxZfgFKinj77/8lPtALv7t+4sYRYNSeFTK6tD
9zGaTlMEiqj00BayuaD/TCboOnhZwc7g0vsuMbTIQEffbRYeltKQTNB9gWyIICFN4UCyRyctF1wa
eReLoV3ugcCmyXLNsx66nE8W8s/O/11xMGh06sR/+UbfdHpue+5vBDwkdFWLpsQMNqrQ537DqEKY
86GJi+DZbXoaLknYZtFgr+GDohd/IRlSWfpKrYzklvSlpyccbn7mwbYDBF5ls0CvXTvOOqJ/+5iT
ghI9HdTVNeUcuBxkUh+wBg5GNPILqsKQLN9LbgGj8a+NNLpyrXLMluuCwc/TUcuMfZBbe1LfvZLV
Qb9qlp1oNJd/SdE8jW4dF+F7ZYgkmhDtAAdtd8lunY3dyLtUmqzoq/9qPUp9/dGddQIZC4sg7nfw
v2/qv4hDprzKzXFD2Df+WqvKMnRhrHnkds6/9EkBcWvZ7wxkqZBqxPPYod1dU1sBTFIDRmBxG+vG
yDni05FFdmBIC18GvIJpr/6cefQEYisS3EQedtENdB1PGMT1/WV06SS3Rn25bCkoCLps42dtHH2R
QsC/kQrq9Jr6PRPyGGv6Y/7TJBXDq67mLx+mo6sc7/cVpySjNTZEQe+vFyYmUcxjhRF+JHUmUgm0
DHGXiu0c3pf9H830V+Hwfmz45AigoLOWVbuz2xQMSH2zIJp9ihuPOmSxdxYgQppuO/0UCV+RGp8G
I6FLl+zsDuwtJVucO+1L5kL8736Z+ynkH2vi9k8J2JHQ/KIthkFdtoW6mllh0+eYL5DlFrZ2Yi47
jPkevqVQQ2U3m7eDwCV2VYuXCsX2Kg+Jz/TudzLIS2lSML7wosF5rGT7p1sqlqYgyIzXp+nrwl5e
E4opjmVJEAcvShl6wTbGRAW+GlH3A+fm7L0nj8Z9+s3+jA9+TpJyIeqpNkO5zsutnW5/WkYHyjd6
HWX4F1UioAgoHueUNL75VWRTWclG4cSx7a5by0+viIfQdhikXLKOM40/B68rqn6rWeToGEjSkX1u
bIsW//yfgL4f5hPbIauQZImz6lkPlzHnVLnbkWQTmXLVdpaH+tb3bEfyxjWqocEVJtyVBYbk60K0
e8QGDdVU7+vVy7fRfOC5AH4HU1iUWrb/zVy8n44UoblWNGLMxR8puZWMIfDCea6Kv1eo4DiRDzbQ
ycL4UqRr4bl7nnme/wyGSfrQefs8zjGZapGOyjo5HVnEzXi1h5r02VdC+OQtu9BkIln8PRlTc1T+
h7MsN2Xc4MCGXDYJx4WChMLSx/7yE6LC8wXS/xmce32/enXj4Ech9Wjv3KgS8EcPMXSRQoMKOhdi
hda+WbzZNHh0V+cymCn2uR5vcUX1pHx+FI2dEL+iWV7sk2FkUL5tBSByKhDvqth9csBJa/t1cXeA
RKj040MhefUbOPfgfLgZjGYSDREgVDrRPeH2AdQbcongODdyAlnDQA4iQ8LZixbSIvazpDto6UfP
/+ThzgaX8UYgVU3uv0IBg3lnuYdMAtSooQ481ChGm1OkohC4puvYj+v6bkSWA3olZMtHVYrgAk0q
MZi28pj+HeI38z6IEiZeg4LPuoJvoSSbanH32VQlUcqePqf3PUJFyB/ww6unvbwRo+2pQCIQfyX1
ngRt0c4kUwBrXdrC4HB4mu7q/FrjvXevBBWv6nz7aUOwVmZlbmOIkcpL1kJA3mkDJLA5dP1hrzjH
92C2LTdzmIYmPWblxhxOdf+7z5mm5XvjwpzX2cF7wgInWYzZLJLgWAwNAfTfOmiJ2ySJaWrSfP+J
m/F1v+Dl+OZiQTIv/4v4jsRThbV+i0vwwgDrZIC2mBa0+lPJ7Vd7MsMsdhoa5HZ4C9zz0o00WnH4
vmGpMQs03pxtB1OwG7Sy/Hqd1103TcqaRtnQo8FisU7ZS25aAxAM8XYNctEUpoHBiDM+GxryzJYR
d3h9hPll6hCZIjt+bgFNJcEtG43FMZhnBYlWKzMHYO8DbjtFWSGhnE/rq20xGAIX/5YOlNbo7ylH
8tpO77Gzoog4z8xDp2X0LO+5Nzc8DJB6sJUl2O/QmiWirG6b/hOKD9+84pqQykN+uYXG6fnjCjn3
tlGUjiudG29mVQEqHsznymTKmY8TRWOEWLMWU8KNWUbkpZakeQL5iS3BqGKIug+42/iC77kMxH4g
cidD3f3/AiH0Iaa89MPRIf/RMMP0MJ2I3CL4lgXj0eIB0j4vqSfgP7m3xgCMX4R2d3rcpaLpkkw/
4o4lO62ytZhYIZw1la1YtzS9ZAVyv5s/wtwUhOfPR8cYrPFdrTchJ6t7SJbwpOW1jPFhQhXYLfr4
1mozTkL+/Lf8l/juxEZnuGzGb+V0SkI2Gfh6xE4Yv0L2aL7Gb+cQTY7WI4DYQ8oDt40y/DEr/VFR
npS+K9A1lMSLTcgr43Z0YPkKwkgu0MT1ec6LIyb+sahr2A8kHVjPKxX0ewsTcpV8JAmjBYr2DTR8
gT8WY8nhRcLduUVWvusih0LzerIaXFzB4OToM4pg0D9DIrN6/Q12LQvzbAts7yf1tPIz+bt7l0gb
7YyRql7xukwQOGJxfRW18bI1+SQTi1IMLofN8y+HYfHV+v30tb6WXKkJy4QD5QMy5ncwH6QiWkQp
TO+9eZ1h5W9+BKb5tnvvHt8du7j3G15eStZZNo+OcFrLgCiT2tHof/uGxgBvLz/uRFDzej94tsNF
ek6Upwkjji4sXUu0CusspBuCeH9LEm+hzeKiPKjz4yuovmu+bezwrKqmCpSH3zPHq5F06/hcqsCr
h1zFTiX7jqDeIloQb76DbedLxmrJjANHp0rxicsZnAvmB8LeACYkf5jykO5/hXxy6Qzlc6zkphUk
BLnIar7NgIUxJfc1QCQC2ieos0vDXUp3H9jlekbum8hWTys3BtTsZLbEvIiu546zvQj3xfHJOIor
Y+zLWDN2sx3N0KCtvZ4nHJEkNj/VyTMknJtKPtbN8cCFuSskwEYfHkGl4vzLD2kzQn9jxEFU0dow
KlF6KuG0H9oSgNBcbdNski2BQv1zPo5JtFOlcvjccPbNLVJ2e0wcYXyktmhCTDI9aPKTodgnXeLl
+UbAOZImW7gr5mWanx3j13UEelBFdzGfz36jvY2j8+rIZRRdqhnVlrYyUIsTVn1q4oTy9bP3rAPg
wcKxgYnzvVkQG/E26Pg97RRBeFjDNhr4DDJG/DJqu88+znQu9l6g3RuGoEKcgU3svt5cdlUP44L4
rT7x6MZbKt78m737ptbfWy3ew/kivX5RNWuXnSEuuRpjFii9T7qT0RPIzN3yO691tz4rBvl53C3u
v/CCd+mtdvFnCjPort//PAW1A3XFI0ICFjYwIYZnBZ4vDy28GNdK5CTLIDbNE9ou8BVJst/ha/oq
a+CNumDyLWSMMzQEEhnwxSkiACOIzlZUx3HJnUciLvEiucrmy7yqt+0YKpJDkasTspYqtlSK24Tn
1+ZGXhxdBS9zZabRU1nGsa3va1l9ls3sF+vSBU7V/sSGbnHFlPjAZi8MVNPlB92WTrbb1sCHOpu8
5EiixyuYjRiHJaY0/J904mGMsii4WxhA8d2W9ceBboB1AQAAn5qP/NG88Kv/GlINn9is28kpVdFO
ESO5Na01LgKpvTbxfyYc264jgAn4E4nKomcMRcVQo32n0IY6ho23/8BvBS4bW2t6drW1U4iQqAv7
gms5VUfxkc/S4+Zfdsa3GanMDtrtQKbNvaFNnRWstkaZ5xW2NocuQwahlg6gaFQH9CECkq8xsEqs
p5Wtq+FGc4klpUYdLb0JCXUzXRtdwOnmAXHYdHk1PLjf/jmaav8rnbhS4/q5Nhtx9mjMRFQLm8G1
7O2bnDkvSLAwyAr1Y5nOWOeVdx0CXCya5iHU7D6mmIrv7l/BcYE/fJKJVxxvmwvKE3NN53j48sJC
UOunI9QdjWsV9xR8v4zed5Ji1uAYbNfzKTcQOHxlIA2k7k+x9FtDahT6w0h6HOe5lC5uu3TVX264
V8sOfF9N0U7zDHCE+FbfbwEfxhiPDF0b+tCyqviZH3hvF1mEkQhUMNBKtGdhfteVqHU12/w/QuAh
aRXrnQ/pVBCEMJO7CBqi+mOwyMXOGtmV3kuyot924lZ2P2DB4AIfQUwwTj8QPPM0/gcgmiuVC5ka
5GZGJJ3twbAXICU2dOCDzoGoQ9tyGZnybYjv93hEUj1cxGAX/Lup6wxcY07WkdQtTj+etyXOjB+/
OSaYdtGIemBEL6M39bN7/MPV2ebPJD5qUU2+r5PxiSrUYAe7Mh93iZGoQrbhMSKd9FmVgmUmpoyk
9tPau5jnKOm9byvFpoY0DlzERqXphWGsp8ZBZUTHvy8P6or+sjSc/3lEBPpg4aPOZ9LjEMEyPz7w
vrJ9u/KkeOqg4cPW5og+TqyWxFKu22cbcHx3MrOUK/VF6lJuBZPlxahkv5cMWX2ez/dlgON6zBNH
Wo4uqtuiH3RQCOLESQWyR+HeKR0YSb0RiJ3f4kcuIUsry+xBRP0PVEDxqL3Qs8JagakddoW04G99
VNCGnYlRe7OH1NZoK27aRuYbRjF7+2qkG0iEvTCtt+JFOf5TKNn78lJw24h39XjaBLM5kIpGP115
nPBGsE3FfmEJuQVvUlnide1xlCpYUUbK/wAmkBlCNlAu9TI+/i/wNy8Ql4MDBrPGlDzhMmGTy0Sh
D0G8L+QiOBGazLDDnaSQ8FyaWuHtH1oSu0H7MIA3yJNjx9bqrW2WYLsf7wEA/+9Yyf20m9zSy56Z
xz9ML2I9Zuf+paxQhlaDFqeQMvczZzApWHOGafphsklWLxv/n5mgWUmLpxGPIxan9fpNIwA7oLYz
UtyMxvawvPyHMmkHyUcY7IP0ZJZVTGl+utTuLvZqnRLLxaLeaHsnksrclR+6NB+hyJlTfO3Ci7mf
ZVorQdG4MzYpcjH40jwTz+oOsWcJbrGc65Sjwp7Vq2S0TUmv+y04qVy+eaY6Cy9ZSLNzmUPd1BO3
OnAzjLYXd4E3ULOKm2WuN8xCUIj6+OZO/kwdr9hI64sCMYDYMR5GTnEVAMEjzrPTbWW7ZcQudjSJ
4ByZChy9sE0OXQO0ME7wtnAwoRyFvQkOCWt2shlClVBRDKiDyyZop76x7js79TBE/Ti15ayyHAfr
eYQGujN2yX4euuzaDXwj9q+HtYiPfcQmvpYHnic1MYqcenS3fFhvt7vO+sEkgkc14exSyK4Iwl7Z
G6ApNbq97v8w2EDN1Z1QDhPyQGLsiLqssxW3DKOt3BvUicy6WrapSOgP77sV5tLEjp7fRp8xmShA
ZBoSpb3RnSox3mjmhW7NCzVEj18sG/WaYTMAZnHdwC7Z+X7VuYyM6vmz1RSy2zIA3O3lPFPbcQTa
UHOgMkbX6zzMJyVm/RTqElcYIBGGSwApN/6AZ+DwdFvb0zOho71rAXqJ57/P+GgwkU8Ch+Eu+EHo
R78uTvNs4rLCY88e2j+rOg/mXDLNCWFwul4dxtisFk1SmvFmEMttQA+a0Cn3COJV3CCaxI59R7j/
NvIotjomA3R0Lrhi9IeNbCzJaIyJn5VbtHTU/fJLkdcxF8PExKTO6xxTXgBQ0Sbro/0bNEUoHMah
MA+BVyRG5CalqgL7j7OvHIYDHSdv49YiBuHIJW6Fe5Jy1NtHd9JUnH6J8+G1V4mz1oRC1rU/Rluo
Msjhxkk5pmTwpBMgcn1Ustajf5/KCsg79lvFbLdI2SDSZfnTr9pnvmE+jROF0dXOKQYFXroMmkFI
+gaFSwEMZzmdba4dUqfsYdKdImger5nK+1FuDLvimz1t0BM0HBGpcQytxZ1banvk1bguNw1DezQm
DA8WqwPei/ZCXmCfohqWHwIXIcn019ixUV7nPFdL3/xfqpTDr5ujPfP0yW+8d09bnYBkpM+bXTWd
dqFH/BbLs6dM93kG4Ga4UexU4eUr7CLryeN2ZC8N6GxmBUG3h6Ty5eOmzrWbZYhbHA/kBy9QxcJt
WuhX+ccspG/H41MzcKr7/Qn2do9MRBPuM8hk1Zi6Gtp8rSzgoMtPCvxGcftPDGL4mAbkAE6pPZYL
IzDxZA86twSmbsF/oGYOn1c34wtd71sjxFOawn1E4Lh1QFn6FMahv33yBouhYWluGniAu2PK4T9Y
WouKBDjADl7VjVsMfM4neUC4v7B2doc1+gdDA+QlgnRO0+40kaZn4duf6TvXpwiNApZcEiO9AM6p
oWZ1mi0+EAWEyJpjxaCIxTsUq2uoksfYS8ht3BVNUc/f0BbMwUiHTIVHENJmB8IkgvvN502yFF9D
aeHvKalXdDdXqsaF+7RRkoTuwD3VwjxkWERVgiPEQLkIPz0a6PNLgnzcgIlPvStXOAcNT/hZ31UT
AP8iwq0IzInIK8NTG2jBiU2hCMKfX4LI04rcpqz1wru2dwVXlOefurAQG304/mBGNHG9ijCYOKGs
Fj6GbA5Q0GvAgbIToqyCZqyLdqEVq8XasOz7bTdMDxj7cp0koh2Z5rNsex/ikbJlbWEjBYSKk3TH
uYnb/h9QInFednB+n8ejnfC1K9gM9e0jvrxJQb0OfrHkmUvxMB7k2l255/nvT3pHjnv8pnPWTZKf
y1/8ZF6uBbC4G9UzY/G0QMjeAWbXoPZkP/P42/Q4zRf4ey6OYsG3C0WAhWPY8sgGYTCx+QwIVTxh
b9Pi7UMEYoESQUWtVXrDFvm0mDIz6XW0kX5JVj9/v/sg5YCpN1q+7g4+rRjJrgNY4u1gkBeUb5TM
VJFukuoFWrKt19GvSZjmCdBB4vogFKEmeWrN8XBM7rrtgXMgkyqmWqpq5rHB5vBr4Jtq/rl3DFmE
/m1EdZlFhTXGSUwaOESjSFOXFvkll9kj0I/EiPtgwbbsaYv6/IBNvd2duYbd4yyJlF3HymEhgv1Z
fKi8cQjw933yvaOGClGnMy6daGtOQjU/evw6eSwjBHHVAzg26NkwAbGjMjj9CUKrokavx6gKvKeL
vSlS4mmG4uPG/IENOTvfLy2MKV9MpH4tqGhns/6ABC2p44wNpKEIzkgrWlFSu8qZbvaO4OVbOlKD
2cKBkaAcrMNY9Pd5Umc+v3zs28bdlfSs6NOTYpFSgwd57fTrr+cl16UKsbiZF9bPbr0A++phHDQf
pi72l2lbQHOC1Zh/9R4l57Xhl85zOQgtDlbdgXRXWlQWHLDUxCiBr4tnhdoZUsedi2H/qjuVh+5f
WOHdEg8184KMETZrJ7Q0i1yJOcZX5P+lNHw6sniedXFg6yMEhhN8pNTV3sgtdAWEFSGJMxX+KWAI
137tJK7DFhMkska44iF1IxFliONrj4TQIYD1ruCL6ah8dVzRUE3FH1kOj0AdWSAc3cQ7CKN4KudI
c5Um41nj7AC+qRD+xpMWdcIwIPL8Nl3DUAjtyQugNceg53BgLZX6NNDEB46btW27AykpSMS77N+8
cGVHxHEDKIKh+0LvwLCGSOTRUpzPgeFg3EXjlZdM262a1xYL+MrBWYD9ef/H2tu4dNbPrLNL5N2A
IF3HE/NgmJTkcLkrOaMhuqBTtIyxB28J67odKhFH0Rn8+CxncPo7LedQZFN2tyFVXgaNAYna9Lqj
WfUJH59iXAIC7/xSt4Uk2QvVBAKb+YCz5MpedxEwaBquqOWoY/YIzWj8hpE+FsoTID+85VmExA/F
DhP4TC0smdesc9qoi9FofvqxSZhlFAJjKvq7slIo/eU5QRfmb66gL0BXqfiFyxB2p/YPrdDcn+EB
P4VW8qD6zESjKTU4Sukesl1cuazalTmPCgqnUX3dTtiZDhUHJ/0LCQ6Fi28OFpnhZ67G9TcyqOb0
qW25cVkLN46yUxHRtxp6Zbnz4tu/STtJEGHu2NhLsUQZPeuQp9h9a+tZcmjhOxZOCb/NG3HhjPdl
s9ppN6rp/1DMjZYUJe6PsEB+3fXfcMMnnamw9YcPwoJjkZ9xKlAgu3FhvIrzaTMgTwgFvGMnx9kz
FahqE4SgnJ8lIDaHvjFY3uqVjMSsdGW8V5tLruGH6g1dHRniLl6WE6/QyAIF0VCHtwEnNYufzvZ4
yqatweSuE0jaFvOnab7DjnWopgytxhM7HAwfrhlFLG7glOVpFx2eApQU2xTFQvH5PN9FZK4QKRHQ
FiSZN4ZTsFWvalemAeGyizj2rBa0dGh7zokDb5OvZrtVD9hLE/k4VcfAHBE+Dt2LU9lfiCoAr4We
7TV0rm/fFNuPKRDp3TnrOb7/U/o/+Wcu0Qvo6/cybEv7lJgMm95HoQXbjAT2ShVOAhYOvBjo8PnR
ct5H0nQ4VZ5ajZWkLKL3iItewlh8YFlW2wD35XQbXVV2ddhwR4eHTxl2v0AX1Ssq5HvdeFnK9HJS
bubaNmoZOxN8ew72wINSBMH35HAGQObBI0DU8IU3HXNi1B0HEW7hrvk58z/uLRTpyVoljPUDx8Fh
Y2Bb7Ml/xy/Ot2E2k1IeBsVqjztaADnnSdwdWdHfpog3JlHBfQA17Z3qu/NvXtdw0EQVR5OCm0LX
0whRgniKJgAoQSY/hnB7pEas/T7RQu9Pr5iTOWEKmE2C3xxgodcJ6VzcIbqzoClJiT2LXbpUN1cw
tisz0oCzCacEp6zNOCtx1RAS/6P7v9kf2AmnckGuG8MX9xWNMra+NbBf5ERdbVc537SZdBt0IVEZ
kdzvdoYtsnDk2DsJaLigUDtfZqnywozike3/NB+4XsmqXOIyhWhSdDY4jykhN4mn29HE0gknFVmz
SkMdeIcV9d6EkvYxOgzdm7FJmBSTCRIRCwamGTEMqtKfDQ2/L/0VRnCpM2ZQKpzC5rJS3iMUWkde
fIG+6sQipn1WQgiQqTVzf/QKO4cnB3dfH7ZTFyL8LgCSApuKXnW6FYPZapzOe0U9Qbnkp0xEXWvR
jIBRYkKViblzsM8yQD/6Q0iKs57wjWBcOAYdumeADGodQnGiNFuFpheqABPYXzLTDLawo6XbdhHY
FbcjimL+pcoAYEytIh9pJ7Ve0+9jTPA7lcwxKt1LNdWYZrQYMjusUMdoYt3zAwq7BkyKA+NzbLh7
78QQRFbR/FI9202sLBTq7gEg2xCYJ/RBGpS01xMJQjFqTq5fN3phexUDFToQ3702nV8DvuP2Fbqj
VlZAwtlCmOhOZJh8JPk+O+1ljyQQcoD/uUg41t1bENnDihuc0e81yAvJmOcm1CnoeNt0bgAWEgB7
Oluah5qvHOguZp+XTcDWlWJTeQbPoaHlpWVjB+I5GZ0fBIsaCzGNqwBR3lutVVmFtFUv0m1A0mU7
jXTnYHxw3p5seN9R4RVk0TwDU7OfM00yufWlJcKZsUf72n9VA2yO3llogZV/ZKuIbhjYxh3INdXK
Be8rwFmF7D8Lj9VTY20IWYRgmVYy7v0ETapLlE+LpQLeOAqkLhZxTItlqCRa+m7icrbriC6X3l0N
gfE6lBjhvnAkn7oAL/0eBsw3xNwMlVVrlzh4CtN5u9la097SEf5TEBnJSOlKqbtZmSJfIxjwoNVe
fD7IlcSLEeqvFqe1Tzw6tXegCSDGgAkK7cSn6Ip9CNDP2bbOLd8+6kaS/GfGkxkwK5j+96KyqxVN
IpS8Knjn/+HWMYgqFdZm89kfgFSgmvrE1DPP63vUvLsVYIj90SPRUo/DxKZIr1fGxcHpz1TkO+mm
BlYrBU2etbrRz3ubW1XaHb2Urb5W8GhsM1K6ptoD4W5MqWVsJPPj8T0zILwSyLHa2gpkPyXf3QJN
wWB0/zFCqR/c+mFgPsaqRxRr9qDOmY1aWJTcrwbfghPQGCfaHdfV+aMQVpZ0Yi5vWpz+xSA8dAyQ
ECXPe5fhaTNVyK6gMoh2RFyE1lyOEpAZAFIBSLRNRrphmwKmxUnMT7ZCP8bmLv/cp+ugj+yU+gSV
aEvkBELjDoEqbUOb+KBlT7bv+x+vqs5keE8FsSBGt/E24N5MkEZEXFSPCyYcuWTFd03FPxwmFo3d
zfmL7zvChuuxznapMyWIZL7i8hZIbOKyuic3EpABDcXoFccgbRnlzBbxuWyGBheHZKmQJF5CqJ25
gDzCUtbDg8TwW7nOBxUIb2NTEAUL0HUy7pQsJWVlw5LY/uAU79gZWWhRLzXv3vxSCUo8mlEif+Nx
sEYctT2dML4SG3MpOJTnPiyQiJgwAZmPJFv7D1kAlTK0xU/e/IrcVKD76i8kanWAacpGDo9Ufvg+
wsbSTPgFQsBk1r2vRDCr+jEozebcWVNcHfTrhNV+pCks6b1DvbRPJc5Nubr1F2Sb4otYhlXecZNE
Kp+s2ZN++pwMR2HsbcQcHqLV1ZVf3ZHp2reJdmSkq1Aea2NuYfou9mWZ2cozp9mbE354/FnjddoT
gi34uzWjNXmsm+ckTgZXHi6iUBOyso6svg9D4+lTN64Fhwi8JWAMbfPlwWlWJeqW36ktmOfZLRSa
Y45SqsNQTsyuo92gRo1PyiQL/beNI9oVkssov59bAKFwdx6CenrWWj6Kj2oCtAJTBn9C+8PngTDP
KLPaEX9TAWlyYNTcEiwM9MOeCxuOuspw0pT3TC6nj2DTxU7QuNLolWzgkiwwEN0+T3Eh30iMP7qr
6/OJy43um97zgRe5A01ozhthMImV6RCcpu+1Gr16v7yqNAZ+CK9dCJQZjM2BzMBrU3wxQj3ZIbb8
uGG1o6qLl9Z04YhqtvkVxYCMiCTLFi06n+hmIJ21Ty5TDnPMYt7KBBX7pe0cfs0ITIshkR2b8DDq
414im4A+KH+Vb1T0471mcvi2cqYa5bbCj+pJAjyzMz16GYsT+lIe4d+VtjYChcxygP9EhhamxsCi
Sm6BxXBtehZbqAE8o5xLRpleV9347cPuzvKlPu+d+YruYJd6lhQn1TYBzSn0ywVsovy8sHCpcdyr
f9Pm6tig2e9ZgfnCh2w8QN4J+1QJVlUgDc289cRlUh3ffOa1hLBbZAXyuBZlS3DKpFgQsgdLO5yV
qAAERoaYf23UylGCZvMoIo9tNH8VhhyYd8PA/2VUtEc5+nJI9IKMr6p+U6UbIwK0GDjgNplt5+6I
Y9cZIcXpN2/5QYJiFuvZX5teJ08fOVpz6L8tZH3bB4IK20gGDCsZ+znkmT2TqyOjgdmsyG14bELj
1s9n7FjXcavqFnfFgozew5lPvGfHJOV6JGXYHqGm4JPQb80fjeoerUoz1eVc8xrwndyWM8q3WPfl
iy/SNbz4ZjZUfTBJmH5QNvTDXlpBEYf4fQ0Bi7vWOfhtVmiqwgbDsljOLveDWaLUewPT/fVffT8v
tyWOlwLyBDGpGnplE5OmsnbgmO5+uI+oGsc1ZGJ+FMicdlJk5lSPs2MpAU5UVMxM22nnVhzkYuXm
iPN7w8NOSGiydMV6xly0KhUVatCGchLVxVdm6ELlgLbxSIwgiDvaC1eyuxHSdaQhWQBFD5ZhKg2L
O5vwpdSNyA22l5RuSJMbsu2HZjzLz1Ko5W7E+0j07HAEuhOc+3WtF31BEvAFAwBgp+36dBcr7MPI
vR5pA8b+F1KKsqoUb5KA9uN7pNTF1BxIuLO4DyjHf7xZF+B17HDRAE+wXBP0ih64ajjZHuqcVpaW
nd5P0CgiJTvX19RX6yWD7jNesV0F0+oiMcyrSG7LXKCq0/JnR8vRJtjuhtR5dPnjr8fIkYoM7Dvv
k9WQbkImMIjMEwHkTeGip9tvsPryMewC80Z7o1Wyem5N+0ivAOPj5LXPqYpiSTjq6vu9MI/K8Hle
Tb19JEiFVpNUJvjadPw/BiHCvPx7W9w5YdWxsXVYlfm7m2zI0Eh2fAt/c+RoHg1piBAM/yicpz9Z
eC8p/SbEw8inGACZ/4dz9LIIqZ/n1buKiy42kuIZfQ2VjLmG6yETj2LQs3CDhoD2wY1MllJXX6c0
4GYM5uEXVhzAo0Hew4odIW5ivhengavU1+UBYxGbK5aJNVyoZ/OIziyFOOSnGOWytfpCrRv1x45H
mV5hAnYVeBtGNoQE1YfSamkbFICfUjqJ0ak68wXneGTaTkSCUNQoTukJNTMMR5tFok+KJnJWLEne
1dl1RC4FeqDVyBo1Mei0Zx0/hNFhfCHDVmzhTOeVvHinTy0FOp0MjEqxy9UCkqWLoxpAyvbYtfgX
x9I66sE0QvRJbxLxoyjH/E8BdXISP3pBhxHx5sxEjILqh4PHbPVpiWjoPO4LwveA9SHx6uwBw7NX
EZ+BGGclLm8WhRqzkPQasv8/x+vOWazOGch1fJaOl07/aOedKirW87z4hOQNK6FABfcuds4Aejo0
VYburSi3EMmsC14uRTpXggwCB9s4Z8jABb59nrNU82mQbVtSVAGjpLh77P/2fKPiZ/Zo21zqXzFO
aE1qDFEJ6SA+H2UNAa6yh5BKF54+6tBRwnqBV2a+M1AQckIzqP88ZhnjjrStkyMnqjefxgkgI6g3
eD/eez+ULWp7ppfT59lPP9jaXf7PniFLnGIfZE4lE3hOqnvQ7PxAaUGaC58DXujEaSKIF6IeOzDp
J/rFSlfbwfAnp0S24I5CB1pi5WcRIwzpo2CbEIO3REzrlKZbGOsrKOZigwqJK54TH0C4ikeXCPRI
aIJqXNvmSqre+u6H6xhcg1jkrqvB57j44l3rxziOj+ZrnWs37Z+fTgkE7QV77DWdhyLoaOIyQiq+
1raITnCXPWeQWB/pVDdSE+D78hRVswHJOpMiWfqT1D1Y3j2Pwa/941qpDa3xY05dghimSGNSOIqV
2YlL+tOECTxP9uGVGeqBcGRoX2qnEAa6b6JOcsTMKU7ArLaPeTuRrVPLMzhEg6+CxTmjf8ge57d9
oS6ZvlGWMz1tmjVvYOH1PrAm10jHzWL+xG7iGLNag4r7LLsLdh8p3VjmBInOJ6A4c3RWUyWeb5/J
KLKoYNQ/7BjzdsZCaAzDe01SsWVBhrvmVgY7n7dTPsGBw2WWIC/83mGZRLstuq8MDmx8jpxZGzjK
C3OCJ0sFGpiyyuhrCX5UtrDTksPgA2jh/FyigZyiSv6IrKmDX4ex/h6u1mMfV1zCSropTvTWw3gG
9p8j5X30lQxwj1VUJXt1Zlrc41/pKZCQYCRGYYg0m7jI32deM6xfe3x6Of30DTzEyce83MTSmtaU
bgHZJpSdnH4ex4bFQqZbCr4txmT3Hl2w/hXitEX4DPcPjdBmX9YV8r8X0NUhmMVExsr0/Qsh2fKM
YTHzoV4T485f2XeqNEZo4pe5+oiM8pzjjbdff/OnN3cLQJyz6il+TTzJGQ/OsGuVEUt5x1fIaIAP
RVsfL8ick9FVBEuamNp5mMKgxu0KpAZFoc1UY3h31u+J9q5wTtax32UklN/SOviHlD3qZCXr/t6m
vf0w764iWrpNINRLplhcFRFnz12u2RwTOBQE09gKgMDKM4R1ggXqteZWeaOg+uCqHyaNctW7kQOh
9XrXeMwhbtz9IIVPa5K+XqsljLQb9PBV++poXTusoBaSuJKqGLeOAG1Uv30iTmQ6IR83wNGGktiB
wp6QeUuaGc2FRXXSSazHKDojzOTm6z6r3ZuVsNFII7BoiiPwb74/ZyUi+JzWWljnoVbFilCB/2el
TSjaDkxhV+wpxSD4pJd73FwLscU+6SscwHSPJbOzcA73WniDy3LQTyrHSlkrLDmY3OUB6jvBHHio
YWf5gP3f1P9jls8HO1yA9Xur06FKJUznZUXKjx4+F7URkyCDKIf4V9M3sZ+29kRmf/UOYUaEoKR9
MT0OxF9FCJQuPdNUB3YCAOviThu6U1LAEz47HSKY31nUNHqDIIXT3CyNM5O0evViv6v8YFbiXUdW
zTGHarJm1z1wpS1dprZr/3kvD47+fmFNdQHmJ9D6dIhsiKGATBzphS22lj6/YKBQSoECcYTbSK1r
o94n1ORxoX7HzmT3iqMbrHcIpkYEqlYiHOMPG/0mj04JyJ2f3uLlBICzNiSGhDVGa6WPLAjz+eYP
3eftP3bElWCJOTV+YndSHFb6VJUXLtAx3r3iq+o3/L3HKGQmHSCCWAQJf+w+LjY2diAywVlRZF+9
1dKtIm6xyyYosY7Io2NLrXfa/69YLCn01m0C6oCe6HHG4/RhgiXdbnqyGV9M/xznzGXuccHI8G+r
GYnBiF1r6/gG0qVYsRiJs3GbCmgFsLP7OPBUknvNndEPdvHHu6UPkEcm3I6L2MjMoBPTGK0PeiH9
IaSMgy+tjsNntstqbmHihDalFUNzy26YbvBFAMyZw/WU2UrE+7UE3AGXJB0kU88Dt8n1PvbdJGRf
57gb8z/s58c1oGouEHuffyxrb38yO+hvEPThqntf9idBOi6jyGrVHrlSbA17Sx+FtBy42wIX4q5L
wvG12C3KlGYlFSVf2HPEkDZLmUbhcy8RmS7zvTVPFXWFrA4Iyes62UrEv023+U8Oozr2TMoyO0ij
9/Hps/CtzsA+Qce5DwPP87+drZuAm/BfiwGlSdqzKTQd0PSMluvvJtXcwz51oh6mkR5nNiJXAc33
dmUrQjjNiRUW43yVQ4HobMpEgfDs7Np/TJM5A3PLVwLjJzfFdcEf4cwXtzpf1GYWb735aSfnZY3r
XM13joMszAxM6gDI+EUnc6mnSK9Rn9TxQNS6anGMlfrUdRYCYDtNQLQYLGTcEQ5EO2iDhjG+OD0n
DEkMpmPdP2mtLqX5K4nXUlGtAB8Ml0dqpOcPZJO2zsnPoiEbufW4UjTL1Q0ESiRvPodUGSu4en4m
Re79ewat7JgycpQDJGgJbfIsYMVexHUBgAiGb3d+DqbgqahqVOplh0bqreLPyYRY151+oju7drGZ
B9d/4L//A+Cj5IkDJl55GUAS9utbAslbAaR2zZupQoGcFARK3uzLTIWlKvxELKAIbHoh662ZGhg3
uwzA6F9hceoXid4PG0NXe72dPyCVlfVOLvMzTKAI5o4ojfBa1F6kSizAEz6GsPb4jEEXxP5ujjY1
4MqUbf7QgvnyV9BgMXOO/M/DDMidkl389cT9C1lETK1+uORgQ9bJXJaBtohdS9Q18ar8aFq86qLp
BcDPnM684fvAc5z+6h4pc5/Gkd94SkFLT3uL0fqVwbx6bgVSxQkLgHIOuQvG150hp1ZHSXLZdbky
9BAZjrSag1JuVtviJiCBhGtrwpp1Otl3rOmzafgxnDVXAA980JL0zRNmGtm0mFecGl81SjOcrC33
UPG+OtVku+RicfUbftvRhdhDrG9d5xBAkS/IhU7BHoulJI6WlvsAYCiYCWCHbyReGOXbcVwubkmt
aCR89VvNh/9T7TyZg1Gq6qLuOIwasWk3F/OtojTFYzzFpslEb+2UVluiwHZBS5ucezFdIhKzOWYp
QBY8V/yziZ6uJP0J4gYn6IlapVYKDSb08ALmGcnNtQLvWN+suCOWDWI3QnbRWOc2N9JSiACkDpiO
Xc4lHqUIPOA4u+euJ/Pi7/vumvPIjtaailMiJxvSNRtj5i+5OvcNOITxf8XqrXgAlI+gEGB64bi4
KNN0YtZH3nZbN2mynlLAeDl3T+7o2gFh4uPBwNTyZ6dTzIDESPKhyNcuO+NblFmC0+Lqxj1hV2AY
2xfn56XqEfjyByZaOa2QNrrWk5PAFQcI5yefrXVg1icKPnj9OAvgeQFrNgv4sxhtecdCNkDemRT4
8jmifKhkpGw1AlsyD0vCdZrEKqlpR9alu1uKZdvr+3LAWU+osTlV3/0VRmPmnx2FQU0KifjyldTF
ob32x9Umm5KHWEeBoOKjOXM/fjfSwyFuHj1mnlHzB6PQfHcPNwZW2muQA2q4cgI00Zfym6Nmr/Dx
akFysY6EAJLY/Pwe5yjL6HhFL2aiDNdTDqn0FoukqoH5cqQ1pndVJRMv39xD21BLj3A+AROxP7m5
rdfj/B6qA6uYxo/lKJQx5BYNcUOs/u/psDZXVvGrT7HB55FyjNwD3ZbmmvDzFYalxbm/2JU/Rf9x
qX9BVOZSR8WLK6A06WOaUFfZK/7vecjz/DqN9ogba86X1/6HjPx7DR/Ok+XPYwxZAnQkariCJ/aF
j6sk1ifmsN07OYu1aHGD8+yGCCotbzXZ5O9lCBMpsqIvt3hp/yTvTgie0VcNUEdZGn3PAeLNsKae
jBctDBhC84utHwU2wHATELGuOWedgA9DlqKxaj8HvA6ElVlUKOVROJ9xQh5paP75EILKaxB96QGR
DRQAY329r9OqlRpq72Rwl6RsgaG+w1gbnBMJKWgmnsObgEvniESThW4AlE7QjqrBfzeNFAHN/5/S
gNp6iPX43kiBXW3EANNkxA46Bb+3fRsNz7y6z1ai4gnFyhkJ5lmVr+KFjxvrSWpk0lLX6tWtVOCZ
k/Uk7Jg4cOnTvzIFmQ0iXBY+HFjmJJjwvfNSMWVvfKTr6P+Dp8q4C7v4uh/WRbkA35xp8gEjDwZ1
li7Ohwy/hBu7ukpCQrs94A50USkiBi6Q9TiDGKAe2iBpCwR4lA/tt3RsnCYmDuM+R17If926H+11
VNrN1xDMwGSH3ulOVNa0fZV/bqAZPVLpuN2RQeOKR2M8katrrGnttgTFtw6yp2TEALOKP5YwV3DU
0MfD83K824hePRRnW6A2qfjrhK9FO+NJHJBsGL/Yj97c0hsZbyCRNy1Omtj+zJ7aOylAWucC/hrW
HbSoNkOuztdCJ+SSHfXhgxYFoqVUzkCcMUtlQpGJyKL6I2HnUUU1cT4scLzaio1JisqpM/S4sKZW
+EFNK1iO3gOsVhh2+/t2WULT77Db3zqZqpm7wKXOhOfPgxZ7SUNKIzX4xj7oBgSTR7DaJIFXWyb9
Gc8q4jRiWGVNjokfMfnNmumdZCXKtWFTH1jZ8kpauzO+UF9t4sWLv9osaxalM2L8c8YitL3AzLRR
X8q/H8xUTM1Pi5U2kPPsj5lOzVEFO+xsbLQmHyCjP1nhykso3OIeV11StmbzdO85YGLUIKI08saD
rbUgkUE0btxuNbP9SgDb1C/sLRRvdCCJdiOZhBTnPmy7MQ5SC3iChe91MWBXXLyA3FkhM6Xb/qTx
KWLBn6XaAQXNeWB6L58XYNtIi2hSCa/1LGh2xRIn4NgJ9e+DtoRcAvRJoA6jnXfmg9MfQzB0xwAL
n/dV7GM/wXjX0DXne3+7u0gpodbPq5gmhXQBdbYTt0v1bOr+wHlAm8HJKcUrnkQcnN9d8o0ZPmIq
+zqURIcwHTFDIPciNUzPcfpjcNlGppaD253N5EDbUXCu9rn4e+mPQXzD2rs2c4+/4yt8A58eqNVH
PxFzdxIxytq/NNZ5G97wdh6aZoY7UvZ3k4yT6jk34/tgMYiNhEDS6qNzqM05LH/ch3IoGNiGVf0Q
BYUwHhKxxLn/qb4Nt8y0rxEAd6GKOujB0wcwusddgAtgXuMqwv+TwEJs/5mXiRtRqI29NaUBOcEo
k5YI6Br2pPJb7sF23q9qy+xGlYtYt4DRb5nxXuZ7IMXBKdhblq9ad850zdC3grhhkp0zoWdH4FKS
9VV4CB+C37gZHwVteEx2QhJXjb/mxTT+TZ5B3hJEdtFXy3XsTfrMFTRzKtvVOM16HLLNK/gXLfON
8K1oY4xblsIGJ/r8Lw0DF0y3WLexQQr3Ot9V5jg9F+LqdJkFsPOiX5JVE+2bJzDLCR0sKYZ/Uz8x
anZRTR3WStppZ1qChXxG8uEGyJCNVC2oj7zTNaLMZAWrAsok6i2qqSKfGrnHCJO1DdPofaoj5Vno
3HGRFdab5hD9pyhnlZDL0CcrXDTLk7abu9PXNVt9klLGcPgfQnsx5JnNtoXX3oHanXQD/srxeKPy
kTPpz5qPkI6FyV/TuXoWJqOFvkzRUBX0xMjDnjjGTr+zTcwtvg6hQoVSnc96NwcM7cAue/ajfHlK
hd4XViKLWUAhkq+ZQ3yh8E6slDN79e74FVmllzdx7EKv32wAxoFyJ5a3HVZt9zIkHXcN2/DBJ2/p
bAQhE7MfWNjSCN/WMj8f1kVLshl5a3KTJ8TqQCkujrFdLt40PovFkhabxCiiAExIl5vZqOjZNfQF
3GPEfI8jVAD3W4ULRilzqB5qQK/vWULkn5ZhpkF4+ux3jDLgoRXzabH99J8/aC2Kx86ASqBVIAfa
74Qc4WeUlsMgBEDaNfgfW1A+gHQN9BcQhrIrXVcWPBpFpEpLX3KnrTfe0PTYnjjkLOb+6DpKej9P
AhI0nNf3xC1UKsbAcmoKOohNUZh3GlmH6xjDjvk1IZLWLX9IqmX8ZFgdMnbX2WjomMbdHOgxOQK4
4vqH4OFzEivM8q0XXMpWnUkefoSFj7o1S5zqJxlacK83wxl4+3UV/nV2OS/GH9XvEXAvsOWjgFue
3tZPzXJp55m7+vApeBg0X67/9bP0mhVMLRFHn1PIYfniz/L2bhwMrlBeoFQOeWhxBrZlLEG/wFdU
PEv8wqNdo/sTmVkTR2Ni3mTwse/JUuYMwmrbTvvFq6mEW7OJXCgVTmizcLP/vCpgLq0WcLVzoJKl
sc8Q5DBib6nbz8c0OSeDguDqYrvT8jgStvGZE+FGlimjtzYstpL1TlMow9yNdwNs0heD7bhI41D1
7ppyeNv4sPnJ4vVJOGJFjvkPb/yWKFJ35AfXh53+JwC4cSjfjBCGXh1C2LVEZxXF+4IVWjYGhNdB
MExZknD+kEe63fk7lmLjuYo6kXNvk8DZOL1aDDt4GeNvF1iSUotEus9n+mAASdSk/p+OQsoPcm9B
eGrNU4F9kH9wVJZBl0eyutoMZd7lBgY/mCnQr9g/fq5AvqmFJgrk5ca8DcO373VpKnH47AOJEOeq
i29MSgdtbsLEL9MGsyHLrfgpqJx8IQxDrfRUFcRdDoFLS7uFF6TGrT9uIm6w55eXzTcridAxYmKG
Vj44AK4MEOfL/OeydhwpNK5sqq4wrE0YQb/KVMwR+dhhgsXlhC8JWFGtp9caAvlmN9cVWj0IRPf9
XWmpnmvwxahUXZo5kTvpsexnP12aa01MOY1TbR8BWesqs1XPH1mUZCvbOAxPoqXQlK9UUdPQ8nB2
FZzi38OYUdpmwV1iMcOIxNCLXBprhaaQjEczLZPZoDkXpFOl8UW/bI7mdRDntjjjGvlZjtslwDKW
WM51kOmqFphvg6SjQ/z/161jQJ5toUNVGIZVTpFAHwE1QmsT5MvtDQRZpwEgcuoiOpBwD49MbXtZ
NvYdNXcxdKOJoQZwpy1yEkPcR7jjI3z0urjkFVIYco2ALWlJbqNq83ifjJlJH4dkiFrv9WWW5zEa
LhM286IQLBoujZcMluVxWnyg9X5Ff3jTvUelYYFVskqlluRPdEmxi7WPgesCZ/QEF9K5rNJYHRz+
7mE+8M6L/lTjHYIALCqB8yz3Yfpkkcgoy4yPMReVT+OSGKXZ+8BST0ZbsgLgfU0ukbNGnaKiwuzw
xCbgV4EPHI9hYDj9JsJo+bCrrUfN6lr4L6CnVq5WpKIvdM1wZtKRGsY4cA+6Q62h5M/9nHLmEH/D
9tg/BXPHoIZcNjE8TBD4HkcEj4H2UydFnVUclwWo7wrgtttxRgQvLic6/tu+eeuCJy7ujONcNPmF
5BiUaD4RSCZUmdBY/LjSalPP0027zmEutL1jK+QbVvMR9Z/p/BdLz3/vfD4ROkcsCJ8G9gPTgQHm
8XVytcmcQ8n4ecUp0NTAx/H6jYhGkcd93+wvC1fk2lT44cwgYPtWWxZMwhrq13x6ynZdD4uTns0B
aeYWSyXO8MkvlkzAkUjPCvZDQf156i3ozve41tYcdxn/zGqYj129U0QByMSBBSQt1Q0DLp8J7zxD
r/I85qyKmWfp9Y5u4PRMdo2hJzqfvhw4w51K1Rb1UEblefXi3EDQgW36/hhdouPxzw3D6APB4L00
UwberAUdldM1dX7doFrXBxY8loKMsYhBT9n1GtxSIBPXCdF5Z1e9K7VxWi9stvcQPaZKHVMpFxLq
e6bYaxcrtlyAfcQukoGxAJf+cPbNWatmhGT8L6kHFVWdWt8b9RKj9DLPfx7MVkO+jVG+YjC9XWPr
vXsqd49SxV0jhVUa2QH6ZuEukVEHZjz+eUPp63YVnplZHWWVWEWXEPkgnSJSX7gYOSzcmaK4x+s2
l1Jti/EcpJy2faZx945Ih6c49sr4OCIwNE2PpGUeONWl8mU2EAgZw8iGfgpHawJnyt9H6uw4lDBj
KTSZTt9IsICrIFVTfQsoboQib1OeV2xP7Jn76f7Y9anPGm0L0aO/YQJ1RN1t0fc9+R66WIR9uqdT
W5CXEr5U+Fiv7hOIWhzw7a63W6VO9hzv9m0wYvVPGXKKaNsZBRpDfkQ+hu655+ASTscLXr6YVEPa
jCASsoTYknIO28pgUWAqm9UXv4cJV5/LEefuGvDhFFvTs/3EG/H0vNQqWWONML0niW1eZD3clczO
G9FEVR/xYcBNeYoF3KSSeMZAGpHwz31WWw2W36oJXkeVw9wJhCCeY9WUEwx8JRAXpWanLJ9Ddb2o
GCzPVp1BlF5MRoQDC+pqD5B34vjne4GpmD9+5TuzSreOYsAD/OG51yX/3WqSKxeWW4BX4mUK5772
wRvCBPCwhhsonaFwm1dEcSxzEp1UYR1c70dGNXv0XYD3FqZRVnlicPa5227OSXMgiDShlHQjBO8t
E298p/g7OWIxwaAi+yWr+PGyHz+bzhMSiUSJVErxMJVacnTQ9S75AasQMRHTrB/d09MHBAC+KsuH
HMOoLacCS83umMBRHTfqiSNUvnbWBmzEIlr4/168AcK+uxBi2ZsVqFpBffQjIhTo9yj20+syFEFs
mdgUObx30fgl5/Fc9knGip3XT6BrYs6HiLFKNV4Z3J40QbjTcdgoLFTXi/2qjzZRuvSznxTu/1vX
9ppJy7K3fTIzSQDim+gqmI4TDCShvI3wVHsLhyPuqkR03c7stegOBExJhYoBHdSZ+yBMkUQ/9DKv
M+gdHPfl29/0W6+GFUAfnZsR1vVrFqeEd0NJKYQbq68/sp5uw4fWYnSrpVN9UWiwy0/w+LY1o0wL
5CpNFbieXNuvBCQVGE65enPxIx0USl+HxyGkYNmnNJD79QPsqVHq4+a872JMoyvZIXvgBoLXZnQr
F1ZPW01UAiKJmnyrqkkBkRrGX70vxA0cpxfaP1SnRUiue0MpyjXSbH04HTvAhcMEcTqor/r72By9
2lDA69zZBbQZeTk3O5dM5Lge3gh4rHcaHoJ9PaaZCyPfQNjUquhg91B9nreFbzLkmplhxnsqbUgr
KfLrX3tujMxK9gjmUomRxxd9E6pnhJ8mKMyJAcchb/vKRv86T6qM+62thFsWPmPhyS1Ivn7ysHPL
LOaI6wBSCmiCK8i/23719mRXJq+vtdWShoiWeFsiuNRwPfCNdWM2ZcCla/mvwY3n1tvLKQsMfc1O
cVo1NfgzO/eUMrHN+DJEiyDkPX6bmDsI7cdp3zfHJEo1WZJ50ITe9xFinaEJyv5NV4aY9DV3DJga
lmBVUhbVM/wkFoZHYcn6v2OQD3+GImXBIcNC3hIRgbsveUdfPr5fnilEeAGOAmvDd2muRKp3LtJj
M8BjPBVswhfJ6A01kKG2boaHMWwSb3QUFHMbcgQVZrq0PXhAbX6FG+v7858Wkg/z+/Sin1BVT2kS
HQco4M/Ua6lOUj6qLeGQBSH6xoKn4XsVFDiv5zY6zOJ0v4JG3PZXFoWWb/CXc7Q+ejV1namvEgaw
QY12ZidYAXcrLvuyoD7s4vH4TEPZMUjwscYXccKMv6xKQjA4OxIJlGY8W7+sJmorDcER/hsMDmfO
AqXazSQyNi8f3j1Fe3RiAdwmnrRKcOGzpYdNFh+ws99oo0rmd4qi2iy3zQdZCg15aw3e11MDopTK
JnNHjHUKypvqmJZGbC4xB41JBGcPn/tlBOBYYYNa7zBpsKyyHj16MibvnanFMQ9nz9R8y/HWePao
rmaciIMcU9p/4x/rdWlyTeP6RHlmsttnr/1MjWx1Givc3sNWmGez03WmLpNHgae9+nvAvyS42sWX
nQVldPXRWg3HPvI8fILLgbKujbPdcprNw52RYeAgq60UYKRazHAPxG3iTixfmmigVga0jBv4APJv
PZR4taTmrMdGGTYkJWB8uei45utWStOm70YoduD9Q5ojkFWTtMj4xhr8cTZ7+6oU9bgaejLdbeeN
3hWoe8eFsVQ1F7GdbtwRiSx0z7lbALeVkteWyq+AlkJAlFF6ik/1mDS1pgUx5Tlt4qs1nOcG7x9w
KLa1XUmmPD/RTfS5lkHCS1xpbs8DBuVwILA8aRq4oYs+DTCgtrTpvE5u4rmXa0wLceuleUBwieKN
8vCkK8N1Bx7CpBJDc2WpM+10WuyqN6nOrJTss5TmuLn7EyI/S3S1SPMba6bUJ1dekb9e0aBlCCU/
6xotQ3D6z5ER/CdPlgAK7ptOIaAhtZTTmZ/YHaoH0jg9Ca4KHoGyVOmLm4Ldq2z1TD89rVIdJeIE
cDBd5RBacturJj0vf9bLb3ZG0723ZotH/V1QLbjTdY/X2Skep6eZO6VaxHhlEbojGU/VoShT7zYH
zWEFE0quwLuXdz+gSWL/eB0SGl2jRVltFPwlC3Xl7pgLMkTm1XA+IgP3+Sj0yanKEh53mz9qY7PK
EKdGAVy9HwLGls2EtdN8Lxlnf+vAPmjZzAbEUj0KWOGzirPooL6PqhtnpLN1bBJIN0toLJNiNcVl
BcL6YL5KLtX0sjH4K4+4gOSBZss6reBOSwJ4Ju+7JjIa32HxAVPpfKpb43T9kWRFOm/BCHHtCC+C
7STSyz/I7pHCpshAwlpF4EFjlbjetWpUg8NTSXWP+zVwnstD+hmrUBd+FXswTeOjC/r5fkAyE/V/
H4Okua2qRzEHw37sUcrGWu4koCsRWDQR97ud1OhGbtbcX22EEcEWkkWbEm8LRdjAbxl8l9zakrD3
+VcTMjlLxyjH7OETU746ryPon2TGugJkpB0VlIBlX+ViDhf8zukX3Hh7hCMfgi39JNSh2V/XnaVw
j78luefyHc6iEJ+FSdP53JY6Fg3fP6bHKR/PpAeXLODvKQCP11rUpKK5k6vtBa9chKEECLhmgU0S
UeJkyWw6SwwB3RyX1vbtkL7K2S9rGl7Ay90cqQXXzfZcjG9Fy2SDYJChzUAJu5k+dO1+41yoRl/C
i0Aqn7Crd1xbxa4lVqphj82z4BvN9pYIVGOwKA/vuL02jP9KwnZesAXYxPPgPTamIDh+dDvhI8Jy
nFNG9HemzMzWSa6C8HwS4vuYjAnc3PN+IgQ/LNmWzDx/RLtGUgpqhaxd4qynHQI0ryxpsmZ6HA8a
DolYBgQ4cbOT1yXG/0/AHyvPcFTqXtsPpqIa8CGXrdARIzQ+UxB1+4/CWRDyjFqBbu0s8S1UsvB3
q/XB2I7LT7WtiZokdb6amvZjDtkpDwfKl3VBHYcYKzJcILTDgOwWBMh6SW/nz460EewAG19BvPrn
HWekCKUf9WMxz1zOvHkuwoGDfn1HmKe7jHdFAnBigpz1pvFzPTIW+3/xxjWmOR8B7PDvliuq7dpC
JNnkpXgc9LGDBfd100Lef0eSW036j5hAGjLJfF28Z7WI8tS0M45EPUX7fBWKXzHl5C5KFp5m8vfl
v5pUAY4Ety641M+QoQm9/3qw6+rcXZZfD4hl28WVP7WMTRf8QbNU4Fwv+UQP2fxYxo4D28zqxmJH
7QQn1kdRZy7Ig8QnigSb1l6vNskgMrY1BZ5Bqu1/1f9/oYmO1S8hfTpDPVEDoELqplPo83ZMcIln
1mc9KdwA5ujRSV38NzNWA7mqHq4sdY/v9GOtsk5r49bhUFxEK9CWPy0+0tXifh0ICSZmXRedLMtI
fOopY4Hbf/RtPfelUDeD+LPQG0W1Zl7kIWVu5/sWY2urp5ZjtAMYWTkX3mawWDh7DIU6bxWKrl7X
2n2U2zbJzoSLE5LUkgjlFF8sVMGzDt53TuiZTy4ZbkDPTGqwqV08TyVRzmxTkNGxs5Jl3Ii0D/vL
l5V7wYn5B96hHyLIJWBi3AIwOSIjmQzDYGZ/3J50yPjP2wCqY2nsOpSL5300Si1a608MP3izKhi5
4E4zAjyUzJXnxw2HV2Vuevk1khJZ2KCOhlzgkLRZL+bk5WDgTS5ffbDX8AupvPTGgB8ASMKZOItJ
UkNY4sxpN80Gv4/syqhg/562diJraU6J+6ow1DImga/AO+AeztG8k0M07WIeLQ6eBgwsWRuoav8L
z+l/UnciFyM1uVX0zC/9xuKW/rTFC4o+WkzeTdd5SAEi6DFnEftUXTsIRx3RK68FCeadHDuegrOG
wNRxQjx3LCTeoPxasS0fATxYZ/StBId5BGEg4KZ3FIhXTcozM77vC/pWoAdTRQrIzPS7/04xDVDD
+4Ca0FFlhGljtSYmn3U9YhhB/ZLm7xWiBd9aSJYlxEvy2wA0ZzoCDa0lAhIQTqsx98kxC0Zq/1Ul
VS/EzcImNPm1Om+6/DJ9/ASCYEr+1yMl4X7zJQrWs7JYo6AZ6nOtxSrGX0mnnHZqgviS+XG4IFeU
zFv0DxaVUvgJdvyhDRg2aDQdQpIF0kGk97ERWjAcBMeleK+iQP0cm2s/0ueLbNd6uSF7fpipbPIe
oEPABPAQAlXmEoToLwlyTV4JnvFIu9pvbU3uCD1MSewUmsThEzuvYa+/kMNsWsLe3btR3ydK94oQ
3ZN6XujU9uKG6epx5fWcO5fS0dFVAdgRQeEwRM6lY8LXMiqm3LECxNCNPXmx9GJ8dhun10ufpnKE
2dmjUGjyBQSjcID8YBlTdPp6yN2Lw0uLnmuYxpnXdiVk7MQ1C4egYbA9tEgpdjVRKHXN1fn1mEEb
pWVzeIgKLozb+vy9b8TfCd9husVZV6r8vYo8OSfOoxswBFBDDxzjNG0bSWuIfusrXnDKOFQ6qsSv
MM74dO7X59uFtfK2cjW+SmM2TQmMhvvt3umSVCBJsixHSLLh0cWezY35abOX/ViFsdP1zUWhv+6t
tMF+tgCkLhRC184tgLUAdf6ew+Ol2RnFfpNDZUaYKrEgNdY7aCgtcFRYSEXrPOJMHiHA8JUYVO4Z
m8UUeaNBpdh3UHvN2BxOAA0QMI7kwCStSs36Ql/1J1gsA9Nh1Kg46ghrxuhACUPaCJQHdT0h1ck3
yKCFywOrqd9Pjicogzi1arlu29/usaKF+O0fRXKO2O17yxAoQkyKIfQDW8hXuGbBw+o73G74K6Fq
Op9BYgWizaHWMkbjq3m48+TrzNV+skOVc0BR9ueD6zwU6CZmzHKy+9i4DGv+fdeNdbeKi72LM0AY
xcKLCwGjVdxYy3TkuSgFlV/dh8Edkj6cbqFffUqGSIfmEf9zlXmITZlm6wjfPqoaQf5Xs7HfQBeV
xVlIPM9bOL9xvOqiDpAntSgZpyQ2YrjRdgU+xErAgM+PEk2TMF3+6vJLTMs2CjjBoAWlFZ1c5Pvr
mP82EJUMJQiziuS+HmoQL9FUrvLhGgArPSpR1hjse3lqOXVvMe1QrJICFG+hDAThCL6G4RpevJmL
v74qC5yKSKysG9g3VuPu6Q1A1IMi2pPWlsY8EaFr3goMBbcBKVrkWgpyJs437IugkGH6QfhpuemZ
0Kj5j2jWjpMIIiE4QVAYSetC2Gi2bDKmWmuP/dNFxfaX4BF6K2piXJqP8ureYmpyHJfxsnPG0PE5
kBw6KQdGlT2QlTsd58lbpGgPV3XoGVb9vKgTBTmANnCqX1fZSJh9BVxE/Sn0K7qoku73qTtqQUy2
OPpalf53v1crJINwQNkoJOJxmrI0AakCj49bXbkkVmPRROEF4TA1TnROZy8zloF14Er3Oh3zOqW0
AO+mQXtvNyQ61KCIM19KYO07dXPDJE1PSsii+uouVZtojQ74Ttu8zss8woWcKYeSmw/NzezeTZYQ
J0DTZnD/goSM0Q7rDQ1LvGP5PwW7dEOkiYbNFw+PFEiDRJbBAiQmoXTJSynaXJAuoYeEBi5YEz2N
rtWVAkFJDfNqGu+IygVCgE+0FfJ/ppV1/p1KDKrG0hkBXoN/pdxKawoT9fNwSuMJsEjV71MbrvNU
UVh6WR4snAg4oj8kUaYVaOt5P0p/2XOMVXNsIYmljsQazDlTk3HwkMhgjq2jy5SdGAAFDTqyvKEj
ypRIt9R5aokrXiHaHvLYnwg2MHrQkEzIapbmWtor++bx0XYVjQ+MGfHXYgXR+KlyC2erAqK/cgqf
Oq8QKHWjVbTG06O3vgAIny6gp3w/jIocHcS8Io70Q8Jxh6bRuIdutRt1AbG+jBfkjwOlCYDE5bwD
pfCmlqHr8TlKCfiQ6tu22yzMk8AqirkHdM2oYRgmjFW9/23NP+4zDqrlKWu4t/DV2UBhPl4EfcVZ
ySXX/Iw2V+XeWYVrn/JHPFT8LnNGAsJGd4T+I9xKRoUxhICoime1V9hC75W0l80ScX3PeOLw9MxV
yzrIjRCjoozf4TB3dhik7XqgEbPFq/0Je8c3Pw+rhnxhyq/wB1PmbR/dEf2GEnGYbPtZn7B8enQx
BIt4DYwk7E5jkbCTcGNq35u5VejsP7EEZN1yGc0PeZTL0501SzOx8e76CW1EkEYgZdoAiAPVt/7s
jEeBCVq/msV/MMeP4aiFt8Vj5vUJ3a7PEwFdptO5L9Lae0aN+crIMnPqMmKyeAVZB9aTHO6m/axL
9zLFrEzi28uZyKOZgVfZm0hhb7ZczGWSrNltfhQ2bqNBqql65J/ZAe8SzV+ETlaf75/HrEAY3Xk8
cEcFUTSpuF6IezevA5cCuEm6FXLT+GVbA9Qc4ISKNE1qEZHodWsT/dE/8jniWB+U5LLqtDoHrzhP
oZPOK4obf3EmNG3d8wBgxIJi9u8tVw4L2T4M2WTIvxMKIk/uh2NREgQvapnn69vSrSAuQtxPxzTq
BVZQ+om/jOZNT79R6WMihAAqS0uTrqd0TpHJ3IaspNh/BXyTow8rnPvAROuAilXljLIylai7oh0b
OHUH0RiJF2yCHUlwVmhQi6HEEAx2/qEbR86FqTsSGDGn5fFGaI/+wFcPXZY0IuVVJZODk5dzbelV
rRXHL70t6VQ4nPSNUGbJZZItnPeZ/fb389KWhkw7bNN5qFXHKZdI0/D27pHvDFL1ZdK8BsyNCbcq
DBE1Ut/HiX0Tkx8DR4zKfi5fxkEyWWZRBclN3ePehjf6BnXiZQFBySCHbzN5YFtpvr1f1XCSXj/8
iw5l3QJrxwfonNLiSe0oEfhkKfRwlzMWm+UwfVni+IH0ZGhi2R6WS5VwFTISWYspuxUi6xvzy9fW
D29UqbHuGaQSvsNoGB36xUJ/yKDZtTdM03gP2MP0vHJfEzFRVZABbvtkwVsw0nSEsZ7Cwoz3PwgO
uODDJhbvHqtD7y0SeN6VjkuIZBZ3W7QkmLfEu749prTx0m1ysnlYk5bQvPv5sS5oyWwuMXVuGOSj
w6C8xcylzvPU+1bCOcku7MDly632HfM4Mr02fzrQXCEKAYllkTvvFCP5+GtG5MuzFcVhl2gPVu66
JVpL+wiKNhWlR/fxioCPFt42Aov8+NdJiYknB8X5sAYHnVGP49mBTzBoZJcqbSka5CEE9PIgswEv
g6IoOzLBXEy7KA/rXzzUeapSp2nK+e2LkiQDslHUd4n56rSO/c7169j/HVQTv/OB/sJIHVwobSo6
5NRZQZTWu8n0jZ0w+q9VIReFhIn3QjDUSN7MD5CfpUpvGpho9Kq09FTTV9hlQUEXUXpUc4iiFU4L
TowFl0SlVOVtbCfIU6AZiEE4iK0zCgIFDnL8UyPF99oT7Kk0lvjnA5OGU43MZXQYBvNE/hS3OC/G
3aSSmZ7Ph8Tq6Kon3d3YF3Tf1AfGUetA4Tn+qQFGAXxE876HXt57o3swaeQLU/Ng4RDi+QbX0AiH
kzWeKNH3ucM5IEfI5ipgtW5RJFUeulIRJXwkB5oBln37z8GxB/LU53uhctE9WInqTnAkaVRW8qiq
WBuMHJe+6A1kUdWBgiN1a9XqFor6H/FMiWtHfp1P4lmneOQwBLZgkmzFpKTgRCcsR9mVC6PqDaR/
OEg/RRy6FsW090cZLmYMWFj6Q7zda8nd8oZty4OhbnRLFD0Yb49J9PiWWEuAdZgB7XX2UaOwCM7p
uPgFQs/9Pn3qrCtGgeTrQ1Kq8j0d/OgkFtrKs1fv7M1ni6VH05+NY3hIOhs4EpccUrHAasrv2Bge
zonPoYNSJ2PoMeOTmg27f0qcR4QmqXE4k13eyNSKm7v3a4MqIhkjmDJZcQBjLNiqjQ+x/IpPi8qH
52yDhtRGp+KDuTbMPwK9oTujCeq1XPBGmlSdzLvmUucDq63MwY8RUh1siosZ5tz+uIPBOFWTcDZ1
HgzvfgzcTJwT4gOusZaRASOhqIq3Ya0sqwz6BD4ik4HIPbQ+kSyvYYY5T1mIszIjBbFeTY5yD2wG
kMSIiGVgTNt80xsWSv0GGwBjnQVEVrzyMLyGgU91Id/e4ze+0hUs04Cq6PXb/FHwfWrNRPHrugz7
HSMPJQnk63ltx/lUoMvsI3072++YsqG34w6ZACFUqwhGUiCIKJEGiTgNkVWUV2lyUxNBri3SAf/y
HTWPkhCVpcDmUO91NEhz2CzJWw3bKOz9xvvRWZvzaTYV/NantO2NKLV803EQVaDmOC/zMusRROKn
/Ce3L2RS1BXSQMETQ/mC8kMHyZIFu0A+/XxZJBjQkYBBMRhjMGZYfEbLnBXWuvtVZwYUDJHFT1M7
CtV+45yv56YMcOq85+9TmmAs2czHf1/9Vb/Jaytzl++O+J7tkhcKXQ0sRss/pC07u3GHYFZgfzav
U4URsq0HRldfKIEJ0pQWYpDHNe+jWYhl3g88XuV8SSczGfHv7nWSq28lblHEUJ1bnapTRzec0ECl
cFdqTsBtbvEk4MUAm9WGgShukihNaHtYHIN3RdoVdwwrPcofJbCf/VOLbPLhDG1jUxQ2aefyA7Pi
TowUhchETDpt84S4VhX9r/r0Q0qLGLCMQn/XsnxQUKRChEO/38GD8jTABowxCI+FfdhmC7i9Gqon
Y1V3A1lanPfpXT6e+LKzDBQ7balI0arE9MH49vMWa42wBv9MLNciN3aG+dH4ipZ4XgoqLR5/WoWL
reuva9dpj+lyccjWJJ0jXvQ56wRAn677CuX0aYP8xee1D1QrjnAN13LnEUJTsF8nt85JG4rivC8T
LwK704rzTWlX825Mh3siKUu+MZ5MYgRHvNAF3DPnhv/cTrSHVc/FVhycmsgVVQxJpdkxvcFdoeNO
XE5luGHfYRTzENgjjUH0tsHPffWa/yGMTEGu/17gfuhTk/BjCUQ/YCaLRzBfSNkMW3pG4ZGw/B+p
O+2zhHPiWL1d0QpcBs5jQqcp6kgEM0uhOROC6+Lvn+ClAoSqLVVNSDp5qIuHIze94gQeFfew1i9T
q2WdOVUuyDReUHyAt2Z7/8lg9wVpAWWbQVtUylXQbRJNIWKqbOS7SFqOD+oF5wL28Rb0L+f92lEc
T97sGl8wOAw+EC9ymco4Tz1EHEpVLVQYPjxQbHUpk9FekEXXDK+c9pxJDdTXi7kXlL0Gku5HtzyE
XKnW/C4pI8fbe7Y0zrM+kx9XOitrNJZkbPV2xg4DqIDwKqG7xsYBBHkYZi3UGNOlmPrWkhpPsm7u
ft+w+mVSUz+yIajbqkhgPapspSiiVTnXAxF3P1NWKT0ZgpLeWeSaKe9eavsm0uJ/0LfdCHpZvHkE
YQIp0nO3y5np5BjtYtgST9FQ8ByfIMWnQYdFZg86b7wHlm1Pwjmti3z50OKkk+abPTCH7KJIVzKs
7RPBYNE3zj4+2CMK07jEHaifQ9cGtatgrcfwSeteWKyDyQ6m34KvVDazzSrGPx4AUgp5k4nrVNEG
5OoKIIL1BHbykhcDH9IfK8atFkrZnXOXrtdEW9GbDleCR88cMhONh2sciqyBiPC8hlTa3sN1BO3O
X9QNxXA4TtWA5i049XpEfwA0BXVCt2j4omMtu2myAB1kM5r/l2o2dz8uZnspgcDoDASAOBG8P6Ya
xYzHSteBqNI+iWdU7UriDhzaHQxC74jHtelsXr6jL/H0soj0HJq1vjRMtUbluh2/3wo1oouDop8n
EYXMaifs19eQ5wJigGT/rrkHD4csLcaXveHY/8eHCBburjU2uDYONm8a+sdiJQpruAwJtyLKSUVX
YIjkW/EOMmEkIq/6JbRe/pFX3u/cwJS2xuo+rtHeW7nqy32G5Kv75/dlq0MiYsHmvxC3ElsxTgid
LIdOzxbJaLI604KjI1AoyV/jFK6AYmDfMZP9goaeouw+i6/V/4BHUEoO8tEwwik5DNVYq/P23Xoy
CuS7BIHDs5tqA2O87Ua3blYaSURgFHC4aLzVVhFR8X4Hh73eCwMRyZ2Mpqmwa1tWbKfjLCkzuy+l
7SsxFyPcvz4Cht8UEqF8LeX8uLTeGrxGqkUJ37E0YTUtDTrwgpw+syD43LLFQ5EYFXlmU/JHlK3O
mqNaMrc539yFg9I1VCHfq/75qXIcE/85N3Ygz26b173thHpBZY4RtQMizB7sn/H9TnU/F9pyHOiv
rzla4SpkA06QotZxRiPW1s3jUOhGp9pQ0ZK3QWva0QN496ESJPC0PBNKHjtl/YEuKNZNIuUpVYoj
jZPMhU9idpSfV3gOPEYiJR+jemCdGO2H5eLIjvGjGKYAIJz5fbIZF5IMXdgT3C2+wi787/F5MSoA
hczLcDJFFgftwhuDfj17oZHjTxVE/Zf8aoIj9oWQvb3vh862q7l7tixvQjh7OXkUcEzrbNkYOInT
s1J0ZxDAGwX4DQNKZzVVw3xyGj7XWqrgF0IMmn7cA6n3ioKjxSLYK7+JSamt4efsJplxIeAx3iNI
o9kqg65n3ux47SSAyTkBuon1OfzWa8tRYtOg4P4X5bm8qWPzpiqk2eePCp0IX69pvZgoENqp97gk
EqayA0hn48YASsg4ikUkvIAnpQj2twnPe/9jWQTYfmWwfHw/Wp2yDo6QK2k4vlnjKmrrdjODMQO2
YQW/5RGU4aFznvvGcLrRXiN+7urDpOrl98IlB8Nt8jj0U6T5AuPbFXma6uMHP9w2Qk/whwva1AiQ
GXpDxWr4vji5cuReJ5IlM35dQRGylC8rNI075nMzWUWsD6ZqYWPhndfv6B5lSVbaKe7+GbhWZwTQ
udZ6z+c/RRGw/mkDWC+t4hKVx1jHqvnji9EL5BIpyhKARX5uVD1Gesx0Gelo9V7VaOdzm5x0JQZo
4rjrY0iFLz1TS53j7sn6hJZlF6F+UR4VOUX3LCRj7xkMXR1+kPjC0XpzCC54RulNoo/sdEFKnXd1
KrRkGw3CRex5yG8Ubol2X1UiTPCkQX6xBVZcWFFFirKU25WHDsJQTBfNmXbUg+y7CwePBuCNcf2p
6gmTWhh5ikHUuRRxin6cHeEfDQOgeoEmamIDqJ9kGHdNwCOD74+wZXh5fNcDgWPRUedCwKV6siYK
CvOEjHEP9gQmmV6ER8aKyQnqnK3DkLyppS6Ld2zO9ieehTY7kZ4RbZZKZqOTwyJ5AxZ6q8lSjJqz
tD8ejpeMa82wm224l/43LqUfGW5AGoXP9hZMMZvF33Yl1UTsO045PZlr7HwOCdgm0umc3zj4Ryua
FOr61UQtNlVC4KahfymBK6CIn4sznSg1njq8glXE8ALZ2ZJpVR9PWuDIytoDGWzX8WHycQaQMFP5
xf32KGHCjbosZKDF4sD8UOy9DJ6Rs0yFKjTLG9GqMfN24AIIWD663Aq1HA/49l/35HmpCED8F/OA
k/irBVYG81rT5r3b/aeLnFcbtm6OvfZCAO8ZB+4noKaOCoLyrpKsEALvrcW/sBBBGehErV/3Gnmw
4t/dycyTOXAl0rpD3+bjHMP0PGfJNns1tsi9ZtESueixygt35spvSuHa04HxegCbuKlN7svKEx6w
LlQp/KNXVkrcD/toYLTppWr+RegNkqmcXNDcxO1gaAXIQ2MbIm/gx430TvQ36z0RyDtRSL3DabID
EplyF3tudVGybi+Fcpx3FQhXgbd6UI+xfsJ/UzP589uojmmYnmhnvTUZ1oE3PebsCmjRBugEu5Af
JFk5ISfVGeTAx9S47gUJ3bHY4n86aPjEzOhf0317sXenUAtYNp97pOzagdGdKtPONo/YGgydB6LI
o8BVfrhZ0j+WnNR9i8guCHKyNoQNNmEk3wiN4sxzom//BQUTmLnSrs6Qrxl6484ILVZ2wlu02M0X
Fnu7aR8j+0avko4nKYyeWY98AnchQXwfYIPhO7bDYA2eMYEm//q4UYVuIZJH4yuxI1h9/bEoEVIA
sn/4rjDriyAdiXXDwydwSdRwHMKXQ/yM0HhsM+Xqc3QvuKRNdbLwPloJJxYuSqZiljHO3+etYp/9
lkLpTmV87MjdMCt2ZjTCWQny/oAS/UzW31RsyTU4IyRA5uTP3GPTh3bWXYZv3RqtazRertN7THiD
C3QgXxTdRxGW2FYJH/R9WB4qeUIiEp7cBFp8SpRy3m1KriUjSY+FoaiD5YoEc+hzYmcUWpdNDY/M
pajcdZPh6G9VPIvlLocjIZyntbeXjk3MIE/tWr+2fq1S5LzKSYzeMl1SaL71QK8OhjLReDIjyaCb
Bc9txuMPYYF1A6TTLxxG1krMNzEtisdynQXv9h3NVVDXbWss1+cnGQ+9u1B2kV4zvo2RDMHXuFGu
AHIGsrCEFYUhMwQAlh35OPqMKQUyrnRz2l1zoK3pCVsYHP20+w/XUTB7TjvSn0YqG6RZa3jJMLbJ
uNVO1ASIHyYLL1QAsrWEAI3CyoQdTjuplJ8nE7jrUaePGsS7jQp+knUEeRb3kH88ipCsPOyzbDT3
bI+rkCqJHZwHtpRrTaSuY1xxu6X+dGUtyxNwfhFMzMuv+RFSnAS6t2lbTk7uAAJ9NgQ+yeroQDfN
9UHkg+7sc/Gr9o3y3L5sKDYlVMWkSsRGel3Tpm2HeYCJjCQCCyl85WR9RlrIDHR2atuoiV8Rwu3f
8JwGV50bNjyMEtSiNtMyhRSwZXYvDOYePIMMxLUryb/cYtSnvq55Dp9O9bMrt/HsGAFS2Q4O/WZd
5PuHSQxOuL5lZQRXfzMRo+A8rQhZugChwOJwhC0BZgPcOgatJFYMYaJYEmJN95/WJDd6DoxdSfyC
aCQ+Z2qIjoY08pPemV5KgPTgW5LIeJzxuiSURgJBFMcrh/REXC2xSasvFLUWE360OB86fNTnpHHf
r3m7Q6AnC1wmoNemHXTGZZE8qGP9ssvHBjK10UL1mqI8UmRwSORz/tvPJOcHy5lPdQsEwPuIoZtC
LB2z/xflZB9v1ZVUTbYJqlwSbt3RlLOo+QbHdEzVbgxTO7Bx3AO+pm/Ihx0DnPtvTGJNIJvlAyJn
ABD4YXmCHdl2rfbBQVnrQxF/7m+nIputlNnTPy1Py7A4Td5x7qoHc9bpqJCNanR7W1CZfQGekSTi
oQr3RtdGVmHkhm7ncbofHt0BUWp1t1ea5PpQp45Bs7FVqVXuWyxebNGovXyvvBRuozZAihLc6Ybv
jMy96wnswoPB1IOvt6v1sfgwNGVPPCtZJgGA3l95xBq6euNJylo9tFtmfPNCw7hQmOS6uFP7i/Rv
U4rre4z9Lv323VD8iOvgJ4eWGJA0+6aY8r96ZbNr9bEEkgXzCKZVg9fiByUEseufoedKsTJfkJZr
OLZm6fm74LLQ916nIElCplHKTeiJP9YBuDwi4XUtHyUrNBQis+AKmmISSXOjF7g+M0D4LkNOXP3w
sKtt6zUKjVUR55eDVEzo7KK2fUmOX8PtTFbJD/16kiEpjWnG6BeWG7cUf1T0Tgn8ufgwD/FZJK50
EtllSsqksjkHWv4ZIUvdKNfdjPGBzObADOvE+Xr5b22nb8zRk0YNIV/3rmWJQnpS4yjdJUnQYkpA
KcZvOLFk9vu2/aEQ+p2izyYQPxTyd+MvvZCE6bItCb31GulBrXGowR7fy2nvxARC2YLNn1TrNqLs
ekE5y9I6J7KWve4ksJ6U/WvayrOpCzwPkoKRgCSDC0pxEOPDQhVb4C0AwX+he3uoAG8zutxuHzES
aMx1jiLCJm7Htem1BxEZB7dSrWysVNwkDSkAt3Ricadzdh8EDE9YiQ+IiQiyVBFpwClNiutwNyA1
p1y+pjoQnex5afH2a04j48xcamjSTdfWauEDtUYGnhz2e/gNyntzg+VjnRrtC36g8AnWiPTu4lUT
ipLHG84c146leNGT5JQMos2al9j3vlHMZsiS0ht8C3Bz1J16uyXQDGOWK7xwADGA9Gfa5N+IXLEB
/N0zLzauqN/cqLZphuc/64GWQcMzPQA05lJnxfH8XPH/zityHojS/ZTurj79risLkw1VCUPeah7i
ExggnG+97b/xMHWcLMCkJ1OF5FFcWlh+6M3+th7bES8doxiAeBDhMHzh7YY38XYEutuVACsqNqnH
x4ok03RLSfU9prC5V62FmgXa+L9grAyudtmbf7XQsCPauZ8JpCkWpJi2m+U/WaGamiNEvBaIyIxz
Kd/KZy2968zojYvmX5zyfKbRUhz2nuLoVsq7NQubiOf5rwxJXr4X9w7S2N018YzFF3ygcW6pCq8b
uEHov4FedujDagYusJGCU17seLjciExUHLkEaRvKrMx0WGF1NU+4c829mVx9Un7MZ0sXW0eEtM7O
+DdiguSRwLYFCPFiCpODN908M4lWDgdOGNWBxVLBIYEpyU8U4MO5IiH6B/3Ob5M/yvn7tzILtXs5
7fA5Vv6hGPgwRy3ZEc/khJOAkA/knXHBPn7WPPHBDWZP+cIbT3C/Qlh3++h3uvhLa0fp1ofbGSr+
U/zodnGgWV5dQ8VTZ2Ap52ngkBNl0gLgnFPpLFJhUnu3bQDP4l0Y6PRYUT6OVDAhbc3Fg2B7uY0J
B3FT/v6kLDiSUv5x4xZPxYQirQeWhuK6SWoebH4kPK8dAoblfVVLK9BoEAiOwsyrQE0GKHyJZRDR
jU6I4NyFP2MF3AdfIWNfWgfjZamsyYOMTUUaF5kuD8QkrmpEq+nQBSSNe0dYA1ULGh+8oPCzhAGp
rOPpJ9onlXl/c77Ij2KgFDaFFOvaJBJP0keXovwhobQl/9bu6zbgLdRp07mZOUem9uifS/KTZuf5
Up7Q7H1+GeAW42yawIEWO1WcQHckfLcUtLmRsbiag70wy1Xrl9HLkPd1qhwlhXRusjGto/USqi9j
jMiwpVarYs9mEP3ktuPHXjsS3oYIfZpEThYSMkCTfUjjb4ufKqB3H7U7o1vICMxB7qw+VMOMCnIR
mqeDPMUloCwq4Yd0wcd5Fuq5JD9LF61rPYgSluDr+HiuSpIahgw7S87EJpd5pprRf5u6tRQO4SMh
dyV/vh63M8VNWURgpfDobQ2fgS0ay8uVkKTL0U5BjCPiuOyEmEht6R8Mbd7eS8iG6tVUUtnTEG0k
dJPjmpZ4QtQGFQXJK3GVzfbuT5ycT8rckZ6/ikaiWX17HuIotWWq0uVv+UFeBCVfblSGNXIVfiQ5
0luKH4UI66+4N+K4JqcRCMcLRnmcac5XTPS/jVfSpjkHonFEW0B0GLm5UvAtbSgb+svaMQBJHR27
MfFdIVOs6qnzuEadhBznRsIQ7JOp3KuSjc6u3E/G8P7oq0BU2jzVyxVVSrYa4ckmPqd1tiOf58Gj
qTrSAWjZSEsBAWNCGK7CaW7NF3AB+m5OW3/YEXcwovB8PmG4Q9y75H26C4bvQL3QfgiKi5/xtUGi
yzCLaoRShgFuEL53vzKIGmKGj7w4AWQ8Pa1AEj75Ot1QRZrSbjcu7Qp9/W5nDclMOOVelZRUnbMq
alj8fJO0cIRiY2LxN7sc9JUI0uaZRBF1SKn93F6iSUxRtRYEauKo/xbL2kfa6OjvFQDDKPqaARw1
PMdVHdjN8olZXyBhIvNIYHPIR9uZXdWcxjDzzZmVzObgXKoNkzylhoHA6OQzh4x12d33WPBSykPa
OXJXHh5oKjQzUgMU0VcB17imy7cH0uoYXbtsjyKsodm7riNPallOCOO0qd4XlPNIqXFTOpJCFnwv
TJMlIHE9fTXgcmAMVraSkcoQf0SFo7fYMg7dOnWBgTz8AL910/hJzGI9yG784Icwbf/vHRZGInr4
XzB9oEGNpJZE/ZhwMwoOp59I+AMpi3SAi2V11A46wHaWIkQqiWk6jIgrInLz3dKsebEZZEy7jsRV
1YGie/9axRTUQ/n7S77s4rKMWQLCkPBupK7hWOUq5cIGlgc50v9lvUr/0M1mfg+KwRZcOcFg2Yle
4gDxlEkfaTIArLHsbl7HFJ7Ff4fhBO2vMuwypbwL9H6J9fFocCz0OB8ET0yVIBYALx9rOKKUjczD
IbNIylG8IopiZuSgeL+EVFQA2Lki6UvEPYAdv6GH7+pMdGOWT738Wc7Y+Tj999QDubL5JhEqtiNx
xVgA6f8dzKvIKsc/ArBQm7G8SroyB1mjlGBMUBLbAjHBXhqNiP2oJ6Z/ldyq1Mrkcev2x65MwwBt
nNx7NxTCfqd+XtDUnmJH7CU1WIFdrnzl4WlVd4MuFg1OCQ7hRxXaBm1u29VxUPKDAhnlXu2TPWax
+g7XgKMvbp2zFJ0dwqUPYc7pkIcLuA56zDIUm1iBAPNWYA+ZWdn+bGFpeFJcQh1ulPdWKmaVsCFu
+USpQyNbB3gmoEkMzQIVLMXr2CV3O2AxFM2llP9cTfiPBwEAW2NQWo5FhZrkKR1NDNkvVAC4/EHQ
1mu+oB8MqZJge0QtczqgILnMLHAJMBA3N7lIQ0gzxFsw9UlHF/pkG+eD/wGjmvP4WMZUnsH7b5ez
tU/P/PZjURkaHscrQRj7SyY8Rrp1CcIHLDXofQCigdx2UqpYgpt9yPXMTzYenSUQMDLNYQcTARfw
bhB7MMo2Nxlc64DeDsogDyvMMRdFhnR8a+n4JoGp+DvvjOQiX5BES/83i1plchENWIt6Kg2VYCzM
x148/CMgoZtlf03N+inYBp0LMdpSBkTBMvn1tfZeV9IKlmYEMUyvsj0mGDmlh6nM70my8UT7M83S
BQq2ibTJv6/jjrseike3GjQTUWSXW/7x651sn53UjqirOfLzMLCR4vmT7MT/h3YPdRLDuWA+G2Tq
wwLn/XmGurTXbn2ioIRD+dYgq88AEb2NDZGK+bzPhjIk4Bnep5YLUe4fBU684tOQrvfuVCpuohQP
s8/kzZ1nZ8ZlV5AJ8H4Pq6Ej1jXDWi9FzDojabYdbjl7dr1VP/e/hdfUsVIWi7wsf9g809tGvIWs
cM0zS7yOk6c8QO9sTgmR+X5TjrM/mu6b6GzoS+AJgjOLt5cwARxaYnSW5JFipW0so9XVIk/J5B09
GsJFug9H2IqNhLvOoJBnLG5u8zRWnFQPkWgWU6VqT3609TwQNI+CFLiY8FJWSwt9qkvQNFpJCvn6
3nVMwjuJD2ujomklh7suNzsO+m5WYIiaXx/50R3DcnyfweCRfKz5pcGlPEzRMo1KUGHTrIb2wiL2
mb24OS0/87Rv9pFaau/0GM+1loiZZe5sQq4JYHEdgruNcbTnOVUZBT9RNh3bKOcq54XQN6evvFuB
d0Mi0aVbdB8G0xsUJU/vrcPaeXtZ0tkFw5APRuYQKdKBp4HhAOrBe2Kpgz5B7B2HQlAwr+OSPxQe
K9XYEMgE/bvOGISwwupSIbsNDqtPvMTN8iofmYlH1WJ+8VUBYb5Gfs2lTWRqrAf+NVQSHhhtjJCE
U0+Re6r6FFxHb+wv/EaLUBl+peLshSnyAJZLBvfLB/KZLowm4QPiz+ZbqWntsD1+KxDoS5XaMCSQ
DvYLW68KXMKf8X882PBOhosIjDXsQhTBogacSEJQha6f2rtxBXtAqpiZy6glIt+NG4kpQSolaTcQ
qZq7DmSFOb4HDudPssjEDggbDe/P3I//vpV459elR27yZN0jmpBBBx0/84rUZDGe6xtf7hd7lndA
FcyBlr16Jn87X9ocKr4ea08GmbJb/kaxBHfN3Z78O3RqWYcUFn0Yil5BnlFitAlZ827ld96mddHe
NPs2ynf1iDY1ZP91TkzLR0KcFQ76s732ZNM8b7tQ3CuxNzFYzJIwEhkvSKcKEcbIsXqNQMOi0k2V
YlWa+3lBQ3NBQwRC3sta/I2FfXesCigihSyJQ7ERcHdaGxk7I/K98HG3QxtR5bk3bZ+wi8ivRdKX
KblvTyf1BmrBK90BlHQtGVMv+DJsD1GlySk4PnUELsMmJhI3zURpK8JD94LYybGX3Jwg7UsSDh0S
L5JoWHgsY+cq4fVqRGXaqLIzdR6HO9JPu8kr7mh3aZ0N6LsLD4Jnf8zCBFNNHqnOiapD/vS3JqFd
8SZ523wyOan5JZmn6hAkeCpKObxS6rSQW3YRGJWEOhAPlLhPkMtsve/YpgHXe09lgakll/5fsdSY
lSIReWWgwE3Dz8RyOPrNM+3crIsMPJSMEOhrPpfh3MMOSEyKuhhcl967jJwcs1v751LaNuSFhnjf
8NjzZxIVxsTB/BC9gEJMF0RM3ckwUXxIwU3An/92+hAuupUny8qeU+pIgwwm5yH208iYhGjk4GXT
x8YcXSpD12NWVNGfTfbb67V4p4AY+p/4/ZJrW/9zxPKBoaEOt/lRyyhmyry9i80fu6EWx2YJWctN
96ZqnYtMRMw3zhOdZOmgTgmQw3pxGMEVM2NAxgjLGcCNUMNL6lpXQ/SQXJmv9lrHl9qmhaFh1oPk
MsX0ffQiSWF0Rzs6mOnExQerNpeG+sIdAp6MneBRIwMu1s9rsJDJIGWES9nv03j5x7WXH+TO3GVk
srYaIfI6FagbADp48WFJLzKUuwn38wEpb8vMrnJb4gz3orCWURfLGwuzur1Kfds6zsNhfB7YeZKL
/KofZ8x3+sLO0lEOkWbblDiQeKPOEC2RvlLnjDaj11pme01/gaXzlEiv5xrDddTpcg4M/TiWpwGF
GKfCa1UNYxN9T06adJaj78yAYP7tQHOrpD8Hm/uHfIfaTCq1GJyb/yLMRvMAb+Ulj8pbJpOoaKDH
rfbyVdxnLYPuS4x5XU3SMO6rLNLikvShP7TubiiAjzJjx5a2iPZ1vo2DsLCcCIDsNszV83/OSTPO
9r1c3tVAUsyURsbmFC8yBQLe9gWCJ0PbwIqAdKLRwFNIa85L3yb78LYlpRi+T7unjyVZmObiPsRz
NibD/8XfNVnpxwTykyA5z5d9Es/HraW71fcLhpcSLKdW+2YgpzB1RbZ76uF0ZGcbQgtHPwHQmwnW
04geTuqTMf9vxQq1OsfJxgWxx0bWW3/gKxLcRNoyQb0yQxX86TNxXnF5TvhC3JzAblTe00ieRg02
xv9xhITC80ox/cg9iP6qs+pWCLP6ZYII88tQ5jzuSsckUaQk4X3VLgxinJTeGwKjB1u5gM4sh00Q
NcVWR7p9NpnIaDOy8VyjitBSwfir6yWiAufzBqmgl+k4KDfsuyLHiEaY2OVXW+5tVtMqwgPXFuAG
0WAR9DhOyB8ti3LpW/Y6gGC/0PaUsEri+QhVm8XZH06LX1pORto71pBZqjv+70/E9gIHm0UvsnQk
9is/d8eAxlXUjqbFP5NhrQid/7b20jMKL1qZ2FxeU4lVZ4hHVyjPnX/up4JRWXs7C5JY8KfZQYwt
h9P01RxfghjxVF7nHBadquxASJ/TrkRI7JCpD6kiHDQWPpTSFcsg3i2WdspNsBjGc3+uS9whKdQJ
3lX6RCKbKDa1bUdkGpenqcZvEcWu341D86F4TBsM1nqv788jdxHqlz9Eht1SpX1YBv8VF44whBdv
S4SFlPcnRSnk5isvarIe6Sjs19Ed06eiGeWsj5RpD+gCWo+tMNhlYAQfO+JMtZkC1A2OpvujjLqs
3DUwS528a69iPzWxSRyncWluyMoZvZ0TY8xlf6+hMgazAGhH1Rj4BJRVnOc9jGo7DfR6SWZgPQim
vtV7yIcOKMwHE8GKffk1CFWsEG941AvGTUTdBturvNFr89/V02DiKW+qYdBmWM8NVwzdAk8m7WN4
BalcyTG2k1trBYfEPyeM+FpxR/YdZYtyvFsFDez0xby7XH/0sRReL6tjlisJnlvdU40Bez0PCGE6
zMn9c1EDjyyRyDwVetaCun078a/OFG2pfyZ5E98VVC0egGyIRvoS1SUJOoL49EhxJgRuqgzgufRp
B7rq040IwAsnbia02TQrQYP/XV732TQWGJaOVeVwS6C74KnTj7PdZ22nNyr4WiRb765hOypSZNYQ
9v22zmMcj+Nf/pmIjOs5HF6a4cvoP3KWPykX+gg7LlGvH+tXE+RYva3tuJEZer52lHBK+rvXXJ/I
tKgQ4P/btxNTIO7wNaMORfk17qsx80EJ05Tm8SWJcYc+7o5GTyg3blcD9NpwH2iYBD7pElDo6ZuE
ujEIqhdrcK33/NoIUkg9mQed5/56mEvnYB2a6EQlUIdAnc5e5kejKUrqA5FZkh2b8DbRY5LdT6E7
3KsN7+/g7KNhDTPn+rFPDx9bulcYxtfOi7ZFml0SisDDbOFGeS385rU0MeE94gSjrs4TaKOeIWUE
1mO4qcTHzfStXzTR/DMfi83hvNxHqxIewjvjTFlwDh8tuLkY71u82UFXul0/YunV9TWJHjoAPRsK
gSfIE0RbkZEHD1b7cz7+u0BAYRhwfkbYvxebfMS5kxy6/fyBh8czVlpTWlmUEJwXM+BFyiOM8jIl
bS7Mr17CWR7VA2iof3WyDB3Udl+m7clKNd+JjdthxYltxFSkrxvQBhTGZ3zJNkk/RNKYo8VYQu+7
bEQmsG1Rbib57i7N6nVex+rkPsirtZbG091nUrN/GAIhFu5UUY6g44BLxM/u+P1nAkuMIZINEVfa
vTEfw4qR/tQLFONiAxdOQZF+Apm3hrPReajg74wVOBHAruyriaqC6j/WWNCu7GFscFGXx8bso3+w
kZCY67nQ/g64kr+io1wj8US+dzntfQrSdrEzmMv3l+pqr8628o6YbwcmoV2+psTkuoKug2PQTfsm
1kJ+JafeLzzFhEuYPVYFIdZffRtgHO31hfqt/zyhiocFmbn33+5GcKnAyfj/GeGM0KI/WRjKuulh
zZKGAO3JCd7si2uxjwcKqHxl8/8rIpPLTZtTuThQ0WeksZOjLjs4Ns2lMF6b+RQNYEoVlayadxu1
xy1bBKwBTkoujIhZSpVRgVeJ2eF9AuzzPOhGqHnFStp9vCzRz+JyZ1agVvF9QW5ERwrzVc1ErEBE
flgv3uJtZj2nW7w382+NS3z6np5p+M/09+PL7BAfBtsb6ZkIj41MmA7ipgFu+AX8EVH5g6+N5If0
ybyI0aE7tzn+mHhYbENrJBXhgcOvEOZXMBi7HewEuSOHFec/nU2rDuPgW20urvHbjPip3p0z/AH3
dj6u/2rZdMAEixn8Gx0xHGN4yiZWPLPXxQfI8sQVYbzDsosqmM3x604F+cq5QRu6EekBukp4sblu
zp7C7lis+fl5kGJwzJ9T0xnHsLscaxvavOwBknCReJi6BoW9R0ek9PNeKKfA2iUnh7huxfTphyRQ
+TFAJca3otnHNA+q49iUS+OTOyDs8AEuKpTqTJHcLZxnXdiL9r0RZ8KazaXi14jW3iJlpsxJJPLK
LXAkubWxlXU3o6xftrQSi3rgUTsn2eoO24cD9dx8vSgNZ8U/cUtDD9L/X7FEd1cOWNnDzd5OBFrw
R+n6NWJXuJsWmQI8ZzwRMBMfvd+oCKYY1cRa+qh7lmStVNkR3vCE8HGm5oezwgk9FSoluMHxE3PA
dLH4wJQrRqQEVU4yZALPl/NN3viXdTyyytGiBCLySfX+rFCTPbEmLlZ9hqu/nL8jpb/2zUSN0iY+
Ozz0srdi6frHqDxeh0YKX881pSzSep6UkdnJJbXkAcde71QB1WcImWJyeSO+8ojXu59lLuGVn/4f
oIC4o0p6+6Qp36X2AArTVZNHEYFudNVbKSODNIKzzQL5QC7TJnAoTW3rqD7o38mLgScnMhsEB0b5
sSGpET0oTwhzLNxjssP3RfdPd+9s2fyYiguLOfuYhmoL66iAls9BxuRFMJrEY8fiOItXyOrzQiMp
mCOf78jMGeV58kClcmH34me1UrmDJYrD586Bf2AvdhaXGyqc6u8mZ+TKmTpQlzJL5uY5KKSh/iv4
+tnoq2mv9MoApFYAWQjpKf6KsYrFTMCf/damyoJpazOte+cigUouEz6GPknBiNqDchZmLgti6tUS
FsX8LVtylxQI40g+YRL9+3F0blb4GVZyfHK9reZ0VoqB3gKsXTJGg12x/tBV2c+Qfea0trtslg0H
cHmKpeB4jJ21Z7xIqx/D3Wn2lC03Ol8ffOas7YpZo6poL/mGW2HZPXIXFqrvMttKcyelhrDWH8UP
db+mOTwPEADZsBc0QQKkR/ecZ/F1lojrefdiR4I25NEpI5/QHOtxif9Fi/9u+20rUc9HWTvm1J8C
up28pgXX2TsU4p5gf1KxNktv4sLVphXCUOQCVBJ8eV7FzgQ1XMx8Cr3EVQC2llPSmi1XNEFuBmSY
Dc56qodtYZl2EHtY8LRK22aAfBg9B1dYGintPf4L8ZCP4+n3qRK++TneqTZK7dQr7w3aPX7ORd1y
rRlG819aahgbotdRpqVCdHvv7NbnnsntqLtzA1McKvghQi1lgSvi6Oz0+9Pprml0tH1cSzcHwWBS
03awQva+b/4UUmwc8Xf/L9gNXtcroXYgQLdaheCTd8frE1HxtsQVCyCULv9VZOUe9XTZuWzdlJQg
Amlx09QB7kLV1MYvaUK/rfiN2ru02Fami1KvkWW4Q8PnMtD1jaRt0WGQc7Xe8qvLQYSbewnR+LN4
swz/VFFFYBuZ5tbS7HGO8QKKn0X+rLtBcQ+WHpXzm4aENSHfvdH8uI2CiFqZi2QL8BEDfGks7d6b
Dr+JUU+CJoJ8/sOXGiQhHus2wQL2JNu/M8szfzdN22WgZlmq5TZrEomgai5PYCg/lrFEDW5l+UEZ
t/W5+HUS5hXgSmxl3QDwPAyBcqWBmfbQUPn7d0p3zlT1D9mnZuB6i75GQZwyZVAqRbHGquYdEGAd
T7OSvWU9b6k12grhIEloehjaxKoMhOErVlYAZCc4ktn1ieprQPpoX+I+DLhMqGhYn9mLHo1bSWmv
Gu3i0mhn2YuqrwAF5GhDcKJfo4W5y8kdlGaqUdnl0ZEg1Ks4OzvG08+Q5Q6MVDAc3ovg0tz4fHhv
fgii2RtRt69CvMRmX7/dHBdMd6B9MDOq/McyguGnuKBaKHmtgzFFuZcPemEkuAjeiJF8+QSx0rmH
hEsuLKt384EzQQohTrYyMqNUMaueARiQgYQnHeR+PWe9y+rg5QEK83wjzb1XTKCE3ty8ieTsp/5g
w+U+qgaBswhcLWtJL0EBa4xrhXO1Gan2o76W3Ns1i5EKF/8Z5YwYS4wwOcwmeJtRVVQYd6JoWpaO
CZBxASznrFW+AiMwYbwX6W1dlh5I4u3uyF5lHRNX5k6uFcPl52PH5BXMErvr2xveJmIgz4WRtrsp
jZLCm3NPmnOusblVwepim0P/bspJf6DuzdgfikSLt568/dlyXnMkA16rN0dLXyzpOp+Z8T07f/qt
Tygr219j4w/p2YqCSnx50sb7hQ2iXoQ0sji3Peq3GSXFual5pGslFTkUTTHdZXIouzOurM+KblmX
t8kZ24NshwUceim7zr6M9UldNWPTgAuW9AkGD9tVll5cZyZU/eHT2s7LJQ0v5nA4df49WP4OMixR
YtZaaYJ9fMmZatIMxan3ywgokIOw9koH4jzDcKwY7tedF0cGjndq/PFbdXL1DxC9ZV7a75US4l/o
BpxRLnNnVac+RCqiAwz6yoIjVs8U9tooP+KZnaAjWtsTr1XZZW8cwCMxs3Qv//frPDoyjkvVmJxc
aWk2JPKSt8+GnGc62sKCOq1zWZk3LLWt9CTqQipsQQGwyUjGS3lvWp7lo9E097y5kUswhjsa9ZRu
X5CQ+FfUDuMSCzfSe+ZXqPXG/2yj0UrnNtvXp8VZFu4ISNpzYSnfjEkVlSdqSX9JRldwSSKSlqTc
wbevpcMasFdxNt6GkdXhLLi3T5XWGLSuHx7bZYjA2M/0z7vsrCwAPB5G40ifn5PiEoGp8Dmgv/kL
6LGCaoLyDXhLzrABrZW6OPzl9/od2eMIrV4CGseC+iBg1bdqGkSUkj/oF3Ym3lE4DnLY3R8DUc0K
rhORJqhjZ95Qjkk7ZYpYG/ICiR3VMTCqGbuDNnPMcpg4wqbSDAE9ArmdRphP0blBcosf1rE+DH6a
/Rn0bwExYbJtTeZf6Hosr7S36LHAwUBBSOKHDWPygCDWo5GYfXINaG81ZLt+0vdIO0JNCKjntIbl
tn0Z1o1B46pVQ3NMBJMjTg73le8S1PcZgtfbLcwe+5W4ZJujuIVS3Cnii9C7zlDlh/x1QZUzwqD9
7eRoOTBr62q3XpvQuz4oKtoTnlofJCbEgegihHxp0hLYMIhuIIn8j+cMlzPYEVsyYuNgIj8udfus
bG4HtHm3avg1Ltye/zuciEnzFIV4rEnHQOJa1bnxD3E3fXhLrkvxHXgqvYo9pD8CD44O6ghjdhC6
UpZ516WxFeerePEXga+0Pbp1KVYDLP9lsY369rgnLYf0yLOqmw6Elaiu0f3vQk9yNgPN9ZMsuF8S
qC2AB0O4LV2tFs0yfq9984f5IX7Q2kHsdFI0z05HrOr8hMwgIdtOyHBAfkr1d9S85zTmNqSh3ZNM
AK65GD0Y8blks6F63O5txTsvULJ7RVehEMa02lXqzgrwZK7uEtACb6Z0BzkmjTMLD4wh33Yob99A
t/yjURIF+31W9oVuPsODHfKMOSOMMb1STpK5EAKedV/3NSwOG0sKldKWMpNfCehdElZf3a+7QPdw
4MXsDR9ZjIHx9I8dtvUC7DPmK/p0/ZOXyNfXqbmJ7SpuVmTBkBsy6yle8Rpq+oO99JqxRkmz9Ye1
tuxP1tQARr2E8AxDnMVCh7QI4z6z3GyFxpiFNdSvP+Uf9b/3Vm3OOOvKclO8JNwaTUrO8NxTyqW4
c5EVzYpKsNck8+ZRKTJCW7AucATaUru9SFbPKUa7NxfkAugPnGD0t1sY5S09eoUvd7+cGIxnDXlw
M896+B3qL7uXDqOjqIErvEVdHQxYnMS2ALIzWkQ/8gKf691qeGtwP0b8NcidzST7y1tAoGu8Bp40
Jl9/6zgoDNuGsuEY/7fQzY/nXkj+u6oWRjgNgMztsQ1r2YmD6cAHFAS0lUfDrubyr6T5iYRfNxkM
mXgIsbbV32WciJrWpaDUzd/SyNvrmNXAwW80xGKNRMBHKWQ0ZniXgGjAsdffrp6gDUrUvQlnu3uy
kKHHMXTCarDdKzOYJR4VOrZfhPu+koGKXY6lqazT2oEhZWLlQc99oULx7NRvR//CMml/OQ0FEJW2
7Xoh/YAi+5ZiP01iedMMTwBdHoz95e0BnkISACyh93TQ2zDdHEpVUzeCM9B735Hz21XPP7CQubkM
vxVBuVQBgvuCcDvLRGTbDpWkZylBuR2cWq2RAOfdpDGpqNx8ohBvaKFUWbSDZK9k4KM23OqEcjlK
6qiQLDc5uiI0E0pBh3LKLNbhlFXtGcdXNm+LTHO/FlPX3g3l1x+dojAYzBsd2oprijVyRbMmGFKB
ksNlsEoe2xoYAsJXALcUX5lWocTc1O3KGC27IeWi2+I+s9GwdXm6W/k6EEceelCIIVVnGB99D+cm
smq82pZbechDQrS/55olZkqvROqEvTKJiXPrOgv5G9ao8VA8GoxlKELfT/e/q1mFa+41LrX3hpcK
AFz4+HWljVNWYAi4AJdhE+RjKSQEAsnWpJBxM5h3caliyNNcqfuOTvaUpO/k5aQDJvXo7vaPAX1F
SB5+dZhSOFINbkHGbwqovz303krrU+AHA68Je5EaivPV9i5F1EE6qcidLOXcoRGQ9Oln0fbz3NXl
iMS3uKnI6UwyGegbd5vdUNdgoIJ6XfBJoTXv/x325zwoPgxGeFQA2L+chxjxWepg47yWUzD6qfX0
KadmFr3DEn8Vkzl+QCEw6DbLvUsMm2yAAtQSBtoYiLGzE44z3TcQJrRBoounwDDDCpdtJpNcs1jL
KbqbFXCJZQ/Nx4gMJsZwG6fzvnta65nuTnYSmnDqvtyLAQOipvAGPOlPYMfs+1PhkGInsR+sqNky
ptIbVdLcdPl8Dtss8WmHnqDH+FxZHjkErtDvhRHhYE/Fx4JWgoDUS5cRxh+3z4byWooVaqhBHbpz
zW1lfxUBuJCRL0zdFTskqSoqD6W+BAWKLfw9XP1xtfg8yOd82mvFNUeMh8/6hJTReyBvo0mXeNwv
10/UrqEdlJhJdu8cME/SHT+LJZwCi7M9K3PPTPgMiqrE0vgC9Bheh0/UvMUCHatohnn6aIDvanjr
0cJzzIj0xXLqEcR31v8rF4tsgdxwvhidTTb2d+gMIVwY0REc+AgtbSt9UYNgmjK+LZ6/LE31Yyz1
1oOxlIfdwFB1FN3uLHwDzkK5p3LyaB+I/Dt+RHs0qAjTRUyFLNou6nWNGLMY7h2gwXbL3cbBqp3D
ipi2AaTjdTCFeequjEFi50eEkdjMJd2rP93g57hX13yW2vazHKhmksSzdfBIknz6Tkoy/YDUm8xq
2FWA8TktoDvT/6sOZap5WXHRLskOc3Qh4oKHlnGOJVVHeBRTR0gn0y7urJ77s6hcNdfLmoiNOudu
Z/e5qeJxRkoZNODGsEW0HdCD1nAr3XJXZyUHoyc0mPrDsOqKD97ozjk50r8sbfdWPXUf38YT51Yf
tRIW9ggeR4HWURmCGTvPkYeXVVjzdTQQNsztbzL/xNQtrqvrC6cgL4ekg/ZVVKT2HLjMBeK0rJp0
uUY5Q/CYQP6ImPbeauxO3ml2BbeF5y0wJYtSTLM6cIU1HPbrbj9+/FwAjeGhXICaoKGuTHvLJUiN
+w2JYfWqqVYyzaq5y6tJvyNCDQg391eSEmjm16Ozlv97KG6bJl68JkHQPJ4jLId0ef3/JetdjxxU
8us33Q9BuA7dcHQA2Gbfupls/ekcJpY0Xr9rZsPZ86yZs8wfeslDZw8JzjbcuDawXasuh9HsjiV4
8ReGfJqwTJ8ey5HGPXY3BvXUyaZByNgBQif73Y+pLTpFLibggT+rlKvESSKzTcQg5Vk6baNdOPgy
dG+Zs62S53SEJgqnTG0pznizpvA8/+pkMz2uvn/dAFRBpVmcK6z3g5x+MHJM8CcG+qIuaS2wdVV+
MhiUdNUkZjpKci1wwhAh6dnakBienMroAVibh8Rk+rUpjoQsR+wo7FN9psMCFRiBXmOOUcjHcUsD
YsAQR08xROlj5goM7VEWGa99J7IBZZxiy5nf5juJLiAsyu9wFfC4P/VHMgJj5aF4KbuKLuzruNLF
Ph08EJEFJApgNwNeOMPVQqikIO+tfOboZ4ZiyF73+ulOwB03V71rPLbUOqLFPHmcRJKGT9y2R7oE
g0J8+3pXVhDwB+KVuvTeq3c1h8Ft8MWu36ryMYXZCbaw2FhhburRzRwk6+FsS0Z8QPeGhaPLrUNV
lKKeYILmISKpaDS1tR8W7VQtvhb5yjzARBwKg6zVD2CNeAWVxNRmiDAFgV+JwfJCtaiFIRcxt94O
Xt4NlWMPB0+/hjS16nNSYb8c500ZehnSWtJkFRtnhf0rqPbYlehO85987WKGaEnosgMzxDJwMEIF
JhHVrl/za11jfgWs+wsE8v8owgn03jVHXfBBqEP+NHCYVNUkipinBMJLzcI51vaEjl6OpMt+a3zN
pNCQ2s2WMW1GgCr+sGWaa5GiJq/Z9mBi38fWBXriNPDjy5A2nsozDmgwCZbArmgWmMms01aluH4d
3VCiymE7A4y4nBnoZZ5rTngqXgJcFZuqz3PqKwKTrGPvBvO5WDi4rQvxLryZZX7Hj3zCuOvMCiYO
MlML4aW1gRzXtMc8T1YB2C3xtFFtH315SgoJaG2Bm7xOSb+bauJDxeGB+xnfbtpKD2SQRl0KAfFC
cUay1wZQWpQLJdlWHRCHxmOzE8Bn7GHF0kKcPg939ZJooL9OBlwR9M8a1yqAZjl6n8lL8k1mycqh
GgJ/+okMGUzj6dOYj9kaG7rU6MfsU5EjvSBK9cnhkMyLZsGwk1pIYVjuBdVdpjtRl3QV7AgQcuug
4ZfOai0hknk6dbX7GIPWuqMB7e1Z8nSTe4wuFQMt7cA5TD9uY4RTnZ4yM0mgq8nOve+161QOzuvV
YHK8VCmgjrisE3Ftel10g41wFZcwqBIDEhV7zrFRUJ/QhinzVllf1Tu2igaaQRxBnaF0Mgc0MNmC
wBYeCeIBWeHltSOAb71UL9ukDMF2dPYhM7cH3mOcrNFyzC6GRRHFyXaqhmgAbNMEV3FO1YSjnVTR
d0CnMz0zfc0xztGcBbxocVWmMzqC+vZhQX6N6gEq2uYE0c/e3uxUJpAF+nFezW4+y2+fR6wUVAfV
j5Yt/05j++ZpaIj6cSG4Awf4zEqQvDAft1LwXtqJTKJ/PPZNwLYKuJvIRZxOd90i2lwt4dWOtH1w
6n89n5tWfA3qPmKbR46v6Qv1yEVS8oyYwumuLQ/wgzWM42sJKa7fGFgK64a6wmk9rJeeRdn4MoiJ
lSwpHz497QZ+8WjLXK4f08uVHrbaC7jBFabzFjdqaC+c2G/Hsl2TAZ/OwNN26yHTbo0pkvXQkaSV
iIAlzKHo1UNiIbgko1reyAkgMdEywRGyP4+DlC5/E6oXfmOVGmEgdlMsdxcT1/uE31gkEA3cXy0K
2DpfN+2YuasXKgAv5GxVJHQx0c89AHifu71qwUjGEu3wzXUVqRweVY4J0bSqUf85brUZtDjzmN6I
woLsr2D+GVXSQC6jAkhmVbaw+c/nP57kAMY1dQXhr8P6U9xLEAWMeDohd0pM1XoFBvhnlrKBq7FH
V6tiKJ1pFJUJi0eHRUxNBPmculVm3jazBoG8f5GCwqJvFpozmhMpOawr85qV3Ala6Jwox7DKxxz/
vbDvLvbwO3JS0b5jxpdj1/gSb9unS6kUg0ntgV52Xe1u4gjkrBhuGAwlt1uIFzirzlTZStZbMM29
+7fGbcpRtdbnWPjr9e/DIwOTFmJRvqC+FpuZ/n/PEayyLmIHWmPEef6Kuw8YrMqLroKYpt9ieyhW
9nmaMGmMEEueEbBmvfDfpK5PKRbuZRmv+F0uCPDn+VUPwnlF5f7AWNGwgWiIvLFMLprk1pYCgGG8
Ro5l85w4Igmau4HadXtqHyXarxor5YUoYy7DL+IaOwXgSTk5k7XLymQGiBuKwG1Vvkupg7F3EsYz
BdjxqeIZDknIzfLcQnNGmHlPGWd4lnbRJAbWpi2IsrcajEEVEju3wGuzuW6nymkWejCuiZMzZWJJ
J6L2bTx/sLs+JuuC14NHEf8oaNzVZKM1fdv0bG+uApChFDyZPOYqfkbCM0ozs3OFO95zqB+yK5TR
Rutm+wlcM2nzMn1LVTW0CXQRVPIMHQ2rTtetPZ2WAvJL+NOUn9OJ1kCr+WDFB0VsDEL3GA77oUG+
wjlWHmFXpegWp2DUJQCxa/k+Gqva2XUtG0aaieq8ZvuQCnDYb7o2xRVs+gWv+P+NULdhQIxqeWMH
vhZzr9q0+zNUOYELkRaXFIi6W2QNwH3kGi0jlc4iYKphx9ptQ/UlWuXv1dTxIpXpqMr4M5Pv6dRr
szUYyixKCfucg1GEp1ctEP/iF1pTcbNIJ33Ov5rvJyUgCM53HM/0hVhHukne6zxgQh92hA3lnq+Z
siDJAykhQOx1vU9LvWM54yP251JqZAdANp3APMAyzswdy+Z9enLnoyqu9cEMMa6I4BgQ3qahUOMN
CgDqB8C/fG0Ex+y27sfOkTmD0vysbEPYF2FvFM0YOqw6hFWhaivv3J3+6BqLtUIlaqi6ymQyHfoK
2Sc2H6wAgvD9ovyCjLvRSQISoi0Wko+haBKQqXDNt6zQfwoi281ZSWRh1lPDpLAaVgF0bamTzl7E
n5cWV6dUQjLKUEwvxRJGYjmFZ6q0BMZqPstuozfrMKRzd/29PI1KmnHS/o/JALJKmEICw1oJ9w1T
BdB29UlWQ/xtHdmW4IkByIHXfSsX8Y37IyXUhcK+a7IGZ3hJbdxq9vGZ8I1yf3l+6NIGG8s3xeRA
eblcxvEmbxdCj8Ckhqp7p3HjUJ5jzmzjk0DJRZSCV2+sNcecxjmNx6NAwf9Kt1byVF90zWS+41fw
vuQ/oI3Q/wp6yYkthpBwYKpF55mSlFYhbNX3Tpu+nxhNfHL39t0oSlJd9+f846O/RFoVrEXawmmO
NMlkBtlEXfu/m00Gwwff+r8OFyaDaXY/BUBjm3L8ZQEZmcMmYGkMplMZnN4pWYZqmNfFkc+UyEnC
i41E2+s1acKfqD2DXNMP5fjmPhITSoQeOGRow5ocLXli8QzoZN/6jFOG34hrzNqbcBTUHFH9acL7
sl4bTCWlsbHkMMdT6DyhF7kyNdjFSpOcWWPhdXbY15CDWuiCPAiIMnsipHvHQ6Z/VyQ+x5yaBAkS
WpxWlwq8/iSL72PCH/38KWBQPuEf3+qa9X8qonPrL+uyI4zdVOLh+rEXEyI9BaE6T23ait3+M7eh
CEJ4ZxIB5Qj2emZrzM+v1Hv01OUZXrDUOWvqKk7OsDATNS+KRUBU7aH5vznwDVOrE8i/XNWIwCZK
eYqVOurWfB/4PCVH7QW2vtBC3vBPEGtOfNooJ7bnoBB0DDt0fm8oQp2GqoxpwLytLZBsWujH82mE
Wi47QxdtT54gd2QE5nzOgikXE+y6o17yDginG19phLTwh1CuqP2iZDb2RLiBkl+M1hM/b27Xx1me
RF2Se6a9nAqCOxqfOi+Vd4P4RmylXIgti77t23LlfrrJFaPbAM+YkGOXIneio05WkVKNucTsuJV0
Cc/JMYUz5qwMGYqDSHoThvzqMLIstWx1nsLMJcF9t8vb3sk4ADliKEi3Jz6Xgum8fUKZe+GcpyMm
EkGpIMf7l9BjTq+TueORc+EbK37UMbXhPpkVyOOHl5iQE+74TPAq8TPUjTzCZL6IKyEw2nV/w2Nw
wlYftm6PLiCnUkXpxS0oHFm9wT7d3ZJiKjelw8ER+hCXZjlQbzsyJzgyWhOxtqZtQxB9oqIMJUoJ
j0JVDltz/a43LATxXf2JcvenMT7iSvaEPbGINyGxND78DdruezygTIeDFrxkBx0b5FK/qqzZtyER
EWoQr4h0KUG0KMfkNl4WHMu2EFP8k5CM3ILDjQNAs7aSq1I0Hqks6oVzK+x+BvVoEKTfN3Y+j2DO
7aO+LdfnUrui/QicVGoD2ubrATlXSW+8ikgyB9eekL3cqJdp9K5xCUpOiR6zsfvYM+rp/ffuT2+o
cw2zBBzmmuY5C1hmt36FGeLMAJOieaTjPT5NV01Pe/5iWBfTBrUumG+kGTeiNfxLqdMNqiqKVdMs
eDFmCy1eJkrh199/89IcK0p/bJVKlGyz7PDOnOxUgQtybEwdHSn25ojWBmVRPGhXMDSF4Bb/XQsC
sPpqlkC1oZqqwrljuQALJsZy6ixD0mE4UVT4OImwo7dz/yFJmQc2oTVorZF6JqB3BQMcr11dQwSA
uPWVXBS0vaVU3bbd67Jeg26T9FexaopFm6SMRZ3Ee5V/WB9gwc0rxHVKMdkolkiJKl4avS4ydkvx
B0rSmwusWHWMQ1BY5KBWoAQ700AjGaniczCrMeLWN8tuo0LIeQ2HkXioJn+oyn4GTbZbQvjwpUgT
N+NYD3/1hLOkfSZDmdC+w9GYThcB7XPXEAyL86UcpEN70ft5fw9W6WWIu9rHRWTkye38eQbfu5bS
Lfddnyn6/LopR2B6oKPst06RI5a/MUf2RzvWKAz68xf92GF2kaFa1KLNlkgTmARVgORa7sCkj4tG
7b+5H8aF6bhK1ByFLe5MWTXI9W0tzKmDKsA4ASabc5BmZpuxY81/L5PYDPCn3CdkEvExXQjn20U8
5E6Nnwp+lKbWkCVpv6oXDPYoWNa7U5e2NRYTwEme27B90i2rILrDPxIuFS0fpsqi5UbnC3FQdug6
dLkPK5yI8oXNwpI3taQwCp17boYyxr6ELRfSNOjNWcz0oO8RFfK+u+qTYDno2BngkE8AWg9YL6WA
gLqjl+D8lMlMwwSxHG9Hp3I8fjVIcrYuIaGKR4EjPni2VCbv5moLSQKgGZFIkfDEgB/wHWr4pYJ+
ZRGttlpKFxxCWriKFSuY7rhGPrURUbQI2gY4A12GXsuvkzeai4Jx8Bdmjdz/5zTL3uHdw+b7xmI5
agUN0stjTJqY8AslzVzZmhIXL6rxjhl3q/yFJE6Y6nK7mfxEOmeL1+wV6xNFKmlKF9AbXvMj4HD0
3ScP5c+Gcm2oUNEs/u+nElx3zLL+2s0QnZ6xazEiZue10OES/mzarUs/GfoZEjzqrp5WUXc9BfwJ
2JmC3W9OZKCteP9b2CzoASbiNcX0WxCh2jZaEIfdmp62v1oV/YuKddwNlIq0ZJahj5/40WzorgIm
cucJQeh1UeiDxHlNsPQF39HusL5pXBH4cTPIZtTX6z7+h0eOJrEijU0Y9UNJVLad3+B6IbV3TU7R
CrzE+rggoNYbV9w3i1H3Do0oeUSjIR82XIYOSJAS/WkTWE4htjkQuQ5v5PiDuKs+rKcrsx9gF9fW
6Q6q3HAIROQLE3DON82KiFMj0BYbvkYDkln3XfmYSkbTekfhgkUlIsBg7+G2i8YSsywziNuBqpIO
h9KM+LFgoAw952ZO+6ERxcMa0c4Hjlgo02pfnt/LZjEdr2wHkgxn8N/Po9vHsMaMAuYbaIylVtBd
Kmsk4bOLZ81T4uqPVo+VQ8kZyR+wQOWDXjxBAUUbgW9fnTSKnCFnAkQhrwTh1mjAiHRAvKBljkZW
2U25O2Bw1DXt0ISgWM5P2gLLnCoGA0m3QY/13zke39aXtCVi3UP3qLC7VIAme1iyYxSMsm6HQlS1
56hEfVdizun1EttKnrFtDnJCHXwVJ0xSxiNjlxYLaYOrZEgTIy6Ly53Gkcd6YIOqkpkfYKMN4uoM
52o/pj7Ncy46Vp2KNbqn67exqDNYuqOA51GIfM4CUtOXmG15oxrJ2hUgqwnRlvi/8jNOT/2rqC/L
5/1pyBq3+P5Jy9f1UjIXEmlzszKN1SCVK+RrGr6iNX8RqdU446ovTCyK4/RrKA5gJYXC6gC55x8L
nwAIX7OENdp26E/WT8nq3jm0RPQ03FyptABNSeuBB9BZa48e/SiqWJccv2mIhwXHMK8j5a7P07fl
4v2z0B/5vIhOipdlcymt5sjCLAPL0AMLc0w+aOoPGLbhXegOByDk4/DkfelynZgslavo/awsDjph
WYGGk1rjN4V1ZWTtcV08SUuKRDdfWqzG0Ur5PAwnR3YCSwrRsOt/5c1x3Qf2FlGcKLZuW2bW1omy
v5lhjss/lpKKVoHA97faZja8dWF7Tv7IapoFyyLI2A7RuoQwShsAO8n6W5NhaH7uSGE4XsnrdtpC
RxBItyxHniaLn9W02ajJ/Tzhr7quGVSwYPmEDlz0frfxIJx35kgtnV5F+kCtUmsVF2pBTMCtUzzU
hIjLaDq0QVnXxq7IVB4SPj2O9O1OfwP9ZKbQwBQFL+p3n7opXpv5Wi6rklxdcCCkeQlOeGnlJ/lh
R6WRpSdeka6mtjIIJIUD941ZiMAYg0fEeftU/LdgmupsfOtAXDrrJFwW1+wSIHnS3eLI2JZoA60h
onPidAcjxQd3DX0WS6qRo4+VdsAZ50FueMbwJsOO5aZ77PDdBRJ78Xudc6QXkYIVBNc27QniCHAp
+rkdKmd3Zz0M2u8GExQugptV+9MJZGxuTGnM3G4/Y0+DNtIatSneRpbEfXsOACCVkqSMlAqYGQXb
oJTWOb85Ep+z6cvaQoTwTNcLur2sXiFrXzsE3qsPZazTLmUtN+/YPLDApRlfIkAqexCKScEXWwT1
CUt1azfdYJ/MlrC8rOfj9P5hEjJ4o0/CNtAar0huoXQayDwUeW4UtrkYVKrDxlDbVa0dpYZ+SZrq
gT/GA5ZaZ69BE2oGpWKtqe44AyZrDlROJEUfNXlccl84s/AOHRm4L4YJ7GcvmHvFBYZHJ73p8WrK
MGT2aXq8PjZGWRf0YvbTrOpv9GypbSB+V5lAwbWUX4mOCSDa0k56gAaR3PXikE8pifgrbP/Qud3f
5KccD4zfhSTjbMfkCegZJ298E0kR5XxN+5YwzgoRFs+l3wg372xPu6eUiDYTID3abh38XXJ0XC25
aeb5skW9s/AtFbz3vKhD3ZIy0iVKbIVSqo2wWe0/AczTFbo3rA/cLFUMeLFfubJmRtouMVXqUpPf
/x+pBOth1ezKJmgzoSOGyNa4oO2ex8WAkP0I7dLQYDDCjTgLKHnp4IZlDNt0KM4R15pczmX438yG
1iZepJdE3N/L0rT/IRM6zNUYmdyD44Qva7xfIQtCTaQjIrthTOpK4vm9CHmiBFSBorC65xYPasRb
anbIJfwSx/310MqAAy1zlKe2YaluRCYvRZHPTEznLs5P1MoxlOK/nMbnc+ernptVc8WMrYslhdqJ
h5VYqckmvE3S0TEnSaPZc83sFCTYT6Na6p+Q0ywKBb7ozUS+Eqs5XQ+QsDDwoS83SKVRQapN3Ro+
JTsTAxn+65jqSK7i24pdk9Jd5/9JOsmCDAR4HvLY5HX6vRTvHgjfvRzPeZvFfzVDL5Jru6HGu7P/
zqcvzwT0LeKJo38/mPJfZmYsScsy9UUZEE9nx5aaCS64gUN9RxwvqiE2T0qmKzOdZtC/V35DrhNd
BH+ZBjraEProj2nMeu1QIssvm0OZ8sewlhKF/t7GRZJOF3YsHIzfz5Zz2ZbDQQwD/cb0ue4AAOHa
ghfTstsSUZgJKlFKsAauMKSFjr+1EuYfRx1NhPbgkbs2JDEcUqBNgg5qmZFmBaHDuSys4c1f8U1H
XGmXHzt1gTok2d2UiPobQDzTA7Ne3sn64zT5XnMilWmqjV90ZdbXmuRZr49dXLitMXdnuBXMFT3v
zt8Ua2mqdy479gOzCF2utzbDhDBzNpFgsDWwyHGbvTBJHay3oyPXvI/xnIKHI6lszZJCr0FfFyUh
gJcCAW9z1TnRDQ2RJJe0MGYhHhnxIaLVyqRLSIlDEj+61l74z401MScLWzcaqP7/lElVnhGy+ijg
jx5X+xFJk3uAZT5pmDNw+ANri48QsmF80cK9fStCCCycBCcavHNkm7JhZkcbXWscanwo6TjQ5e9A
q0NSeYgDNbAB5vgftGfXqHu/iladEI9Nyl4q+RvuqgwEJdh/87Y9Xq3WRTxwmOSbLG+zq6oVWvzx
lkorE5bTcREuxhgYlabrtJi921AROG3WJKdPaxZyB/Pcey2r1INEYWontnlRn+bjZ8Mv1Y7GWSFC
n7Gl5ZjiADS5W+GGxbchR7ZFOYPhcuc6i9nnJ9jb5LkWKacrgXqj1rsOZ/LHx7LRQJYkKQx4+tu0
Smd0bIaqmqDeYoH50dnLm1w1cQYLdFjpBel3ixNi/1G/vM3dpa6g+hraifNc9oX7yfz0BhJ50eIi
IX2XYxfLVNi1OCQAujeSLBtvIaKpIjcLm2ecu2yI6RdTc97eqLlS3SJk6t2DvlzR+W5FdSdvE8/B
5Tq8rs4onDjcW1yLR9MJ7i1WiEXhh6+6oD1XQ2x3z8p4s7VQuJSKNHZEgA4swJkiBtSdXyMiZp3w
d8aRxHyUEaKYrmjkF1rWFOA6r6VHC8oPY+2NSPId1RaqHBq9Arhq0ldIjSmO0FsLUoJzLIS3N+jc
F/9ovEqhDPLBxTaM/1/b/6LND+M18M01237gWXoYCgUVmxd5rFPojgRHpSEO+phBsep3pd1Xy+NO
jLeFXYdX4SB9rP37VCzv+OMcO2OHqWF6iFuljOQc0SogOUokXFsT2+Hg4TbN6Lsf3wE4kjbv42bE
aNzk7NFQemU2SsJA1YCyJXzWPMOYeqf7FLQb1HQQttk4RAego9U1yk66PJH0vk/C0u5v7LWQBnN3
Crk7+aSK6HBN209cUdw17Trhgb5C8XxkWaqA51AgzdY3qMOT8wAG5Z1+yNW40EHbMsJ9y/e6Pnzu
q35KCu7ZvzgSaZn93hw9x8vY8omaOzlLJSPNRallnAff9JfzWpBVu1cDNNFq1Ywugzf52dNlAhql
aFmxKzBzeWwtHGa7zzxKETn56AQAve+E7uKk5McRrfrGZ7wGA2gvdiotoDTUdwYksT9KV8P5akce
a7H9S0TgQSoEpirjkrQGz94LthSNDXZ6PwLaKSIssezPpVLmj0HwImhAF3irwZcfHMRv/z0cwEi+
GaXi6OaFl+/YdIW0vei0iuxGgC0S7cF1SPDgBRGs2ALJyo45O717pauJ/IRpWDTZANQT6HhdMgXT
ZJgiuLnDl1epTRb2ISXWsSqdfrA3LJ9B/diEtPCcBn6uFmiPTbt8KKfn+SxtqJwd4GM8XjirOtFA
xlLw3VJLXvveNNVL6yuYfLkJa3OkmRGYnXr90zFH8/POZWFo85tZRNOQWzDae+/v3H/ixGObeeQW
LMQAfPtYZ5ZonjNzJCcZEP7wKMN4Qfy3vhVq/QZh4SRch7g/cmGxhV22LThayb+wV2xfN73q7ISl
zXF2bS8Ry/ugkOwaiVBwYLxFBeKsxBYIhz4eQLCFltdtZ+mCzdLZPqQ/2ywm0NOIdiKdQIUkXAQ4
iomtXIJM80fH+lHzpMdJVmhMXCgF0sSG4WYL9DIV/aMn92YtbYQCBpwx20S2zBE4bJWP6Y2284lG
3PPHAQlZK9Q2FC66Df5GLWBEEJf/+Rf/D3YtuM7fsW7bHYIXb2AUQovcJi0tBvBGjbnBCqmzKfuF
qpLNvs/kZPSkOdnN4z8CDEvx3rH6QKio+vvkG4U/fkN63F/rFYFRBKNqB4sqA/oA7lc3Wcx7tlqV
JBmlvt021LLxV2ktzj7/vseNNqyKsnyCpU6RjugooeU3o9LRZ77ut15B2BZJcSuJhrEz4ey5b+Cj
U9LtY1ngZhl5edgZZW0ZgIpr49UCN/dfGOyp7WVX2vxZipZVhJGFTYyGrxpASzgc8ZNZQsoEdebk
e4Cugd3unkrCG30IfDwDHKq+aZDWX8+vYdlKf5aWuh2HLwEuliT3WiKjR34LK70gUYl2Rj0udSda
A2IkO6IKz3nGtU8NJt2Yd6mg5yovCsoQEWw7WQX3JrBja0WX+922w3aLcu7A0wjEkvmIhHtV4pWO
u1HNNqlabbEE4QHGitTfnd9ky7Z9ujSFcVELy9fG45NiPqpT3w320qQ9on3jK8GgYw2bDTmARMhO
J7gzqpO/Z+XVbwFDrhgu79JNe6qY0c/S/t1XQJgmAtfTMPGHyx2CqhmrwywCEcDO1vX9pNI3pXwz
cEV0KHHZjvr657FHYYbJpls1IjyB8g+sAB75bo/kZCEhiQizEj/HghEMhkZypFMaV+wPMRl7Yej/
Z0HBiMUWBzdHU1/dgjgA+RTNU4Vnp7p7delPi6oPpdH8v/TvWtxicazo9syM1/NyhGn+wvP5wzhM
T9Euvbyg0hnhMoHExkSL2OIuj4IBOzQ969SS+ge2scC26LbAlxzZgTfUCwHJvRq2UKjT5Hs+hHqg
352/MxrrvBAkRPO9xIy8hGsitGoiBpDeMoLtL8XdrTtyIvGpVyaIxzh8A0ZESk+F6L33DHT8bbxU
JFckZCDHJ0sdHbverDMtryoB8vShVKXtH3IGmLyfcHeWoiPy3O0wXIEPvlVCUjrcjoI40m6yzshv
LGEPHeiex95sVckjIlDnXM+Us1B2wlMW+rvvBCz8dBO/JBRWP5zJAy3pxtaf1oyGMiy66ZoCML+z
Z3TIMUvaJusBjVxsDW80PExckmTi5ZcEQnghngBuwEN6XFVEw8BkAWjdvy5/Cmk3UonYFBCGB9Ry
Dlm7CW2NyGk7jai/ZGbJStFK4SyXrNBxG2W5omBoNbw2V20n9BPoNBjNcLCeocBD+NP5b8nJgLrT
00FYwCsedul2I3DTCDW6K2Ge+R59vpndsR/I5V+bEI5/oT51MHjNtpCv8ssOcRwXwIjlUh2foUGw
yY1TuZ7y/S2DXTjBo9sc0ogepf8noL+CmGHuAdcaGxfIlJNpYalSvR3wOoAeI7FmnCGhVm5SLKmB
wEe/m3lV1VVdrtIpetamvdJ0ETw+Q/mbAD3KZdbQassEzUE4hcCrAiiFLOvt9kK2Qm670b/pQeKu
KxicxVKJGAdKPKWBgclEhH3EfLwMEPZrVMvTmoc9cF7ZhmMY4RcYwXQ5WC8tEPc6QL8Jj3qwAdaF
mTW4dG4e97N3DM03ExS+2wpjLGkalYby/xtIa5/wUgP0LAr9LMdURdCWDWtVi7ZSwg0KRR3ac5FR
JBcVpGBd5U6sYql381ZIiv4QEXMXHa5tZvrUrCr6oGvdWDL1JaQkQ52WWb6ZrogoWWHwNuMETG5w
ky1h6acF8IL2IK+WsUHNEsvYBduS50ctMZrA8X48Tw5PN6s7KdQfM10RAE519YaU+x17erc6fVzt
s4lgX0Zp0aKorfmOyge2Z+oAozvE/nPiIkzN3h8SZXWR0ptr1+W8PFOjAmH6Hp6XD5iDiQPpo3U3
nCYyyF5KfXYP2c2yH4r+eXUmAsJH1r06fk0cX3uWSpfR4LQ2pP5VC8lGg4qTzHT3Eci+QvN3siDq
POXOm/x6nozlSkaIehQyh100vdxITEHlMvbF1hXotTPD+WX9NGeYd8zzi+S5tgRrun4hIkzH+zwx
+cp75R4ogfUn8EEvQ4YynUFVUE/yrziYEcbKGbze436ceGVIv30SI2JivCk8GFOzCMMnr27M6EP0
OltbB35l+cbG1qhknvjRnBJe45zzzLSHVZqUgv72cRaurA/TRmOwf6TAZsOI3V/4bTtYA5KILZVg
6UPNlKTN3L/E34yfw4rxXg6aHBJnmsXUdKWiHu5F4b3IfltW4uENAOtW9ZwRKtvtkb9BKbKr9ogf
tRcU+qbVk9yQ2DpMppS0zqC4a8M2vxpWtO31PMKVclnfO0HCAjrddlOx9E17HB9173k3dj28eT/i
GuWbjHkncBUk5uQKCI4Tgobwp79+1tP2sLQq9zaMs6D4TZC9w+lw090OrirhtiW9LAlwoB094SCj
IFk+exOUf2nf52fTmqP62OyUVGeO6ZNqU+DwaXNBB18vxz3yKXV5f4bZEUQkPVpP76XgVMwXNO57
f455Jk/cgAcbw5z3YBcfK5YbPgk24Y5puT3yhwrRENdqqJcNh+szpzimiHpOP6khZz5alR28jyqU
aoD3cQ1wg3DuEQmvOnbNkp0O2X3pbQ50tSNdz17JKYh7z816wJcgmheoBhr+ly7kXinK5M52zFa/
3E/Btf0gA6KFSbZ1He1lJOOVsr9DrrKf/giPXKrIVpI+AdeiSgSedYrp6T091ftA8v8pyAOGe12k
eNVW8fKfZUE9sLmU5AM7SjAN4jRq1yI/D/MRhq2hoQEOTbu18WSRit9bmOa+3pe1LPVIGmy8qC0U
iDNUBwoetri5FTXFszNsDXXD4PvPdaZUXncJwR/O2eJwW90oa/7Ih/unIXtAgAPeg5WnuLqDwpIq
q883SK7aCkQBZpFGNVoDESpPgwhf4vjnlRm/tuFgISxnjK847BjUVma7NEgy+PnojDADsVA8FPsC
CaAobyL0pMK7E5eg47fh87xAWbt49WONBCIfdONUW0oLbQx1HRgkUGjJinYjg1+h9wuV3DCb3lgb
FCi71HRzPXgTmSNAZacJ0KYGqS1CK+vHmYef0Kq2qnc3s4u8JGyMaSszdBgMsRM7udQTVimDlFka
JUIA0jYIISsJnunF65j/+2RBZd4GvtUj83P65RKipSEBEh+P/reKtBn7YtRRMkYBx93ur+HlWxS4
JQgm/btl0r8+fgZheb0TGVOR+rdJEjyg/kgPpdm/Cc1fB+QTecyAHDHYJ/p1sj2y6qLfM5QP7+bW
sZKDdXuI4sybVFIy+7/VPOgXLWT9X89f2+26g0Ja1b/a8ZuVn35WPsRMgl0Pq40pgn5dSlf5RoFT
r5xgsY6lZmOqisC/Ai8OuwKHbVTyc4jIJ0yFFyreEcLIuP7O8hkV+wfs4b8Z6HQym1hCRGnyEpr9
TzTDaWk0a9b2l/lfJgTx+I/nfN8FRFECzN1NFTkM9BJbiY/TncvBJb/3ZYC4TWKbEzFVb3bBg/Z/
aXqqH44bMRQJisvJPWHi4d05wXlFF+r6LXND/cH+ujjwOm6P9eaH/7Lru9m/GsDvG0v8acQ2F9gV
hRsrHTm6J49bRwZY5JjnqymFXPQfyCwF/YZeToGe2bIym7mdIclHejygzDZC/6BuW4qgiw314xOi
DXi66Q0AOaSo736kok8U19osYKv7V1RqXXehha1xkwPVm0v2i0aEgcxYboPCsBjsIRXM45B+YqLx
ekhLPKIDQd3gWIEsE4ZgpveC/c+Ex64QjkHl8+77QNhIuynxxrV80G8/af3C07wfi+C1uc+0ASlj
paGBK8mtbZVg+OiM6EEvgdaTuwglvlkJudXDs4xc0n/1MXjhYcUnlJb//jU8hYBjU4tHOJwjxg5j
FegnMaM9TssWJ4OwbCERljo+pH3mRfT7EZYyQmZUZWdbKjxzrERb7HIf6zdXr2bcBvgM3eQeZig3
H4Um/I60G0Uv9+soRqEKA/G5iP2N5N94rbg822TF6dg3inm6Ia3VZfh+ABAfrSpOqbA3IcsivEXB
Nzkf9aFObq3QlYfvdSKOp//aGEXVZT1cwBgNj5KEJLxy8dAugzOmxvelCLxa8T1I7pnRHa+1QPa5
C0dLTxhgm8XqAQPE9rDvfAiwEzYSetvCGMwEOqoXg9lwA6vRkeRK0QH1YjUB3JtmmuxzGXTWS55c
q8UxT9gGmkancKgYa2g+5sH2MHeeLwA/rrISIMalfM1fkBM5geWW373yVL6oNs6xlaHZsdL+UDAa
Tdv+VkMMdAk1CcH5mqDL4Vvk1/xspFyJpf+mhN+EFsw9tzibkW8VohyteYiYtCLEpPgE8pQfqZwY
AdEaD2/xTWO8ANwPdKXPwPEPdi39y6cdz4UrEt8EvAWdDMjLJD2CIBQJSLtukbR8Vx038LMBPa/i
FJj2VieIKRbjCygt23Ov0eZdXYtU6Iz1P7qQgDlqjwnseWUmHLCbMZ9D8P1l0IpFSPncJ4mo+JQO
C0l5ARS9FI+bU+zvn2Zo0d2TkkcKGbn5M5OT7lcPrLbjxQmeIO77ywbvs2ugPDFrp8lE0R/wqST+
QMhJAq5VcewfD9QH0dVoOmGd7y/nfSLZP/H7CTpTL1RmsQiv4wWSDLKX5e1GOzespXLmsvmXbb4d
E/btZ22N2xf+5dBlavfHy9pBcYdv4WxLVPLNXhqrp33TEVxm/jzqBWT8NUPiBYVDQjPGbHWKmuu9
6Svw3I33lZcziFnNVSjGu3ACI3ksj7fl4Cy091qU+EJTUoTRLqYqLgJ9Zb6i8In7WZopQuk8X2q+
HYagFF/J3qOEkj/roYgoSllWnrc4+oJvzPlgE0IRBgHg0RdOdSq6E8cbsm1T6lwOvsiIEbh0km7G
qYTg7BFT8mT7Hw7FqstffeS/hWPXILIK1UuZ7is2K5sQoRpZYBpvOrRJYn/hzEvyxwNRn86ihoHx
XEQYurjzExFzYEW06M1dLC3gpfwk4xLtdmsprjDCjRksanFX4TxUQZalza5oId0c3ZxhIuEPwRpz
lppJgen791dqDwUa9B1pGGDWb3bJiApp7CK0dlO3nTCaSlkSa4RgQvaJ6rzrIqFG/398cPgjwvjE
ho9Z/HMJtWs5s3eVY/5DryeQdR/MFFZsW13ZsOM3YQ/vxbkuqcOi9TCdt2Dk2BBmBuMEFp3p2/5X
+xwLQezJxUUQMw4DD2U46o7NRiSvqhkiU0H0hbh9kHuViiIJPkfXQ2iitVjegPwNzO0FPH33yfK4
5mFpFk5eZEAZSqHLDUKkMxUvRpSU92cKAPuN0be14xxWJQPCsDDmgWlv6kNSe7pplE/6MM8NfKYo
1myoq6o8eIZkqSBQpbbdAXA3+BTDwKpNTC12lQo9gqXE73p2HmsJtvo2eM7OldHH4p2dySb/zugh
QYeX1yCz5lb5dO6zyhqTXC3BpaxhSNClPLO82qEk+8FEzqY8pYH+DOlha1QsIfgjk97GRn2QXhte
6KhlhzqgwOqf5DOXZwGDS+LzEU2jsZPJpMYnoxQbfBBpUYuUbqC+1fFj3OwFpFWNJbp7mVYgBZ5k
0KFH0Uo4MNeUbLuRmbyXIp72YKccbonHv7jIPvCrt5cPchfKsz38C+jsOqWyRI78YX1+nio6vgB+
RV8leE8I6SC9hxuO4hbBCD9YxzaZ41TxO9r94PlIbYt+6e2zEIwQpbhDsK9A4JcvLRNIP1L7bOhk
pmCJjYvylyUrdQWuXHcCFtHwONYLZ8z6X+IUF/rzNOxAYJ7KnEGXDoyVx0QKZi2lWPP3rEOwbd3h
wjlMguYctcf6EWXlzCgCL+iMlTzVg8ck1Yr3TmzI/pTw0oqqnbNEhe9qaj9jjwNCMUJydaGtaL+g
2S1z1nMNX0UrUryLzLUPlm2b7C1C0/rxnmxOjR0p8/Y/+GyXNxM6AXZwVi5r/WjBCYDcmOvhW6tE
uCM0Ed6tPlrXbhFElIn9/sW/glfr38FhBihZlPmm0ayIoJJmiUf6TRlpcM6Kq3Cx2N6mG5ii3CP+
KV1kjbxvSz1B9FKXBH8Y3SXQB2FkJXFef+GTP6s2TLQ5fVAMUl5p9R3RIOjXI0dawXRaSaNinU9E
fQIDypsO0VRIhU6+i+eYJW9Yn3XBBkGX7bRSl/Ebt2kUqupgzeD/uoI1s5CK5AZUp4iFgg0m1bhr
oJJxKxNd7JEN4zRq0Tnl37Cji63Qk2Q9gTJp5esQaovSrCPc+3Y4ANw3TfEyM6kDrksjltTEuJRV
4yC283BuZub8/svElotBe3KJOwesyvTlCr4h+zxGMgfP7ppDDVfuYrygLYXaHDKf9v4P5t3IRgSQ
8eBPAaRg71Y6NcjBr6Ii1g3k4hjBk9qUfxsTH6cxeMuLrSJeBFIfpnl2TOZNGCJPeIVVX2oZBrnT
FsO7SZsIbjINffJ2FyeDB2j/ADlkrEqQ8lK5msrp9O5D4VTo5sXZ3AtkdEzgaQDHwBvFWOuUhQi2
Uox7hKAC9OVeKqgIE6qx04PrJ3aEDljNVMbCrmsqaBWnrdsgK6QKZtw7rElfuD2EM/P0vEsPX15A
OVfcOnlwXvlxtnMNn05D9BOcoS7JdiKjA3yLw82KVhhYpeoh9fx12vK+VofZ3Y+NNwIc4VaJNFJO
i+n2t1xBCuTrKJrYs5NV2wlB2GAFvFruKCc8rP8cUwosuep+MIoH15P/qLMzYfhR+T1QwlIFwzSP
CqKJ1cVji8jt4CiDB+itJRjriJdb0WttQdjzKLbjI/th0+fdo4gE8sbFqEfPn9oBiy3g7s8oMzzg
41HR9/VHyAXHtlhJRh4Q4kugBlR3GaCWL5KL3zgbS/bpnU/+JyVFAKzfwcCB2rSMmEnkK0t6ZZhp
DuxdFGbKS0ZWMiQPGLbUuq1RPC1t1iko5utyovIEU9rcqAUkxXLzxMFHq+WC13m8km1lcJrcbNYF
m+ejS3W4xNkmNIMoWjgt16d8opAm5zAvaEeMju3r6r4N5pIDNIvYrZ5gz+9zsj4JFOCc8B0CCGPC
jgwrH9EOeHXoGnpD4jMU4tL6eXTzE4cWEd/u4lQneeKS/1cIJdvFMK3dNHd3s1TWKLtCwBEXMQWM
JXWufJI2GHW7EFOzAo2/6q1NYpN15sSVt+RK4I7cPUwsHRb6seZKa7JO6DVRfI5+VoRhgzwIaXec
RssLEDkwDmAkgIxc9m6Jz+UYHThlKnjlIf74Boxq7Z3u+SS1ZqQtPzDx7IadvTfhrT2NAyzfQSL/
rXRCXqd0QYgXieK1LDSOq3ReBW5P/cChdfYECRWqnv0vt6WVhoYxrk+6MBke7ukGfxirBhaz8Vws
Sx0N+52w7TyarjM8D6UhlSexomirKcAvDjvmBVCJzoGAEbtPKAEDfZOe+zO/cZ/2l+AaSekAK7yS
XL/Kgn3kD8FEh/KU7FoCux5zLDE/07n/VRqpqfO1QOKaQaYwnWehD3TPanZ4u/eibtpK6Dwxua6/
CFwtXOJvDGf7Kv45L0eIhpt3r8emMgD+nDu5HqvVhhnxBAf7OvXx022h3Zy6AAtsk0uxfcHl/Wrb
MpvAQ4gEJaDg7/aMF7z6y89FNnhukjbpn6LFcQpzssw4sAf2FMyJmShX2CZUVaPKiEZGjP+gHNlQ
wW5O9pDM2jg8vOmA9YbiWIRLu2HX2Q+NCXOETuuhTolqnUBfTt20QRcLRs0yt4iN1P2k+B07qeED
LKgWPWKiR3sH4/JPBZgxdRE8cmwzTRZe+FWtOE7hqGejBRBGibR4r+xTW7s7gMaVjhhZLbNH31mM
fC55qZUafac6JtiY7MY/Y+6DeRhUHdecBLFgpbyQVHH4fVGjLhq5wDpCn2hZFcCy4bKbTbhL1Dwp
74M/av1846i72yGMTnyQ12wLLO9DPi5aes/UjCjlrLkiW7iDULD9wEj3xAXt922RBm9NjA2Xwdeg
Y1GwpqBE25Y42kCPLTwjDu/xsfJ43KBGgsXYEDT1yGUEDlnwK+EKmeMYXu6Dee8ax5frSg1lhd8S
MTkNFCTPz7Ou/226TStyN30DrZQ+TVMtMfDFVPQ3oEEgLmOpOzdOzKHKDaH6Rn3VLL2a6k7wboaK
OBDkLml6p+hJGM7wfsZzGhWmNyBFap+nXPKuHF82zouef19jH53p/1B2qbs08By6dDpzaoMRs9vc
tRjX/bPo7me4fOMEXmoozFYV+GzofpodQObt8DaZwT/2RfNt6yTYrHLe5Vb0DXI8GplCFQlxU8XS
mXm6qap+M+7LUQusAbn/SPPeVhBu5VvK+6F5oo9QaJRoMrUVC9A9Rh4phXc1zJ5Of0lGqlrZjGyA
OTGw2LV0YULhkMpiNCLdx2fNnIe83KKIxHiLNx9xydM07jx8iMKlWufKuz0K/K9u3jezCxE3/FWM
R2SE69dIpjuwYBg05ExyuuiwkWg6d2QDwpE0UO9tZW7o+/f693mtXIHIJFD5wcHelYFWERp+EZ9P
tgpE08LAaH68YVy92oPCcArFB5v+kUpZwkhfeb7b6mRV2FKKESIiUgsg/xqW8UmIIH/YYN2gi5dh
vP1lm0fs+5bIYf8bMevO8elC4BOaWLfWTZMGN4VZhMunp9AUbyd6rW96rbAFlmHCdh/eXchxMNca
yCRVYAnZrGScR2IOEVn2QAdeX37EqLdjZ3tcoZ3ybVfAz8xDhmHyh0rCTyuN2VKo50b5NBH2kKcm
4gfEcGvrxNR4GZTpWBIxGjKfJrxfqNwZZK7Sk802Ljvb4H5D3PKA62JZ846x4BY3sGbTUBorOE3V
S2aj3fFULkwvZnU8ZFSfmM5jTbyAtAHtsfqlhYwURUMayW3XrAj6jcrEVPuQUPdJksTwEYxPd021
OI+7p3NTgne0w7zRj8oBhxxsBBUt1vGwI4OLgmevmkXHOKIBGr01Ggwrxw+lzTqY5FL81xn3cUqs
nvtmAtOWvEHowNcZQa9bI2HKeYyNWFa01xTh5jneaIG6dDsJJi7OKfcy9nKX1qrtp83ij2bBQhyN
Rnrp8u82lDtC+HCwQLMMgeRNnnJQaz1f8xzs56hY0hsloPaxa/WIScVtf+rQopZjaD7gVlMp3cgX
GbkKdrDSKU5upGDWfKYhiyPCqQU1roPXRb+Wrv99zlsP1+L3vSivDxsW/FDapcv+9eL3ZEFklWnh
mGWlx99dJHo+ET1qUmWwU4oIyf6njtIh7Fy5aAX6QrhWorMAvyiv7G4SDgZuHMm4HllB9dRtJ3om
30Er59ed6fjfblNQF7OqVSdyZDVnxpWlhYcctSiZYcUQ6Gk+9NXyHlhRgnoV5+6AslVboRvVV7ti
9+15BEnfLiAz1eZn/Goy//QfM7ttkNvcDxBhF8nUoIAepVI8m2nVSNRYgcFVmRGUCsLNmekE1VKG
IP2wfLCSKiQru8qzWaukzv2B5dLZtuvRwNs/FtkE1HPuK5GoZfNNdz2qqUHIuH7inko8NI4obzIv
gzIk7IyxdhIaAYdSVyLN2UqwY/TvtvWJJN8mwQSDHyKILnrpBBrGDlvfOzDJVzutwsSi8w65LbSg
oCf3oMAwiLxpILPoiBCcb58OPNeLccoSFNsZmeGyPfP5NqR+bPUk0ct3UK1fpa+L5L1antQXdDef
L/2LV8ABYl9d9hxK8eVdK4UXZuxaqG8zxY5K+tJ+fYxzZgWqECChNbEuHAt5anXCG22TYsJmshE4
qPJiIVExDhdx6uzd9xDUuYNeoA35XX4A4FlceACGulw++UgUU9PE/FZW+3/hnwJTa4kqbI0t7RFC
vTae28XNRWB3g9W5p+6Oxq8BrQkKYO3eHYfZ05l/UsUT0gPv5nw0SYcW5UdVAq/4QFqYxBfxS+aj
f0ies99hiPXNeRFSPt4FsK/fT6g6yYhshth8jNb9iqA1fqILXynAmZ+OSusCDKv0+er6g3yXCuc5
TycWhRc0wZJRXn0LlVlVekkpfe5z/l7p90oi6QQh4obzIXxQJupkoxVajBBgz7DIQwJ8MC2XjSJL
IijgzfLJCGCOd8pjkg64t19ZbZWJTHRBQxpV/wbIFAEFNIlFPBkyCnDPbniiHEOtWGjHzv2+gCiW
rLsdVqbjASWvld3s35OlUKaOIHRboCRptrrnqB7lysOLo8Me/yDD9dRquMObyiA67pVCYoo+N1Hg
qrTlvZy1/jRtnDk5EFzj6L2pAaS/0yhgtShBiA7AYr/Q7h9KkPSxPV+z73UTkKmaxRS6/XngUtpN
sVqjLIZMGNjoMf4DgHxFMCB0pHqY4U2RrokEHKGjDkWVq0taJHWVzzh5BofZAw+0uibBYIFqKEzO
8EQ6nigpsSKKQzAVADDwNvzYAQ66tAbPmHyB5bNa/7dam68iFXoGj6xiMQcVvFZ5dGzqV6HuLrho
JdLX8U+EBkn0jojLCwDtuCqTSpUsnKxrCeLrufpSgO/b2xpvMTwLu2QBynEGCm588kqN4Os1oQNr
0Xvp/5mpcnIQh1EQMI2XOs4X0aZUImJrdkFE7PGdGpZUR8Dpw7lTVnUmXBUq05Bp94HsOpjCw4cD
oCLN6F4pjmRxgS7gLiU7C3SlQkD0GaS6nN+r9WIv9D08u79XCAn2tvjX60lzdg+9yWJxWGe/TGxy
YP13WJKRs5W+8uUpffZC2U/H0u82LsTsg/YGlCqt9P3hM4zllWvGyL5qK5ZZcfyfXWI2xO7dWZqL
fF7FEMNetadYukbikoLBMTZm70M4ftGzO1Fh9NFpXp6niu966QFb1pZAmdTHUeRwlhVl5nX8v1AF
lqzyDFwc4m9hKvtNo5r2NhFvSDPErvIrCYCMdD9vyeLwZ99KgeNXV/rXJAxEAIytdabIoJvSEfzp
GmrpXSaFG53985NPNBh9/1+Rh/RCzZCUNraI3sd364RWfEAWm2904YmfJ1hNi7pfI1mZI8ugxp1i
FvXPvah+tsAhySTnOyLaDMO9dJcyjydryTwAAL5LbEuO8f9VxrnBirAuNEWxS0KS5HdlKJBmEwNG
WdYBP+WzXTbrGYuLNkeCEnE5YnUT/79cjGLhCjVNvTGm4gFLWw7yPg3IHrM/Aar9HeN/mPg0j7jp
Ro/tbtrtFfW+nqFrUVZeGrN3EFIO2OVUHnk1+Y8K00bYLvq2+TX3lDHeRs6e1+FC+p35yzZ7PWmv
yqxu1V3xmS7FeHgrULxtoY9NDmDbC7OLoxWKpi1dvNOlZeRDeXToG+4mIyG2o/+/pMfXocV4gsse
LOoOTMxP2GmGK5dV+jsPLP3Gd5oUoOZIWAwnp1a6dDfbfw4wFUmIj8KHcZw5ihU8RTEUowq2TyL0
kyMP090HpGNXuHccKXt/4brQY+MIUGuajXQdMQQByZg2CPoDCLi5kaU0h3gMEqhAErWjDDW3usg9
BYbejNNjEu8xudtWlC6I/qG4+/N/XiWnB9JOzpDekMe7YMKN7LvpL5uB6AebQtArJJovod5xmyu7
etau/giW6ImgaOjZrtN3VW1w6e5sBYhrRAbSj8POFHd63YrCYOakD5YUt7wa7Gq0nvzOkJ09gGGf
mU5MEhNnWGjuyDMgMRoUcYwKhTo6jaRKkNFY88yhTHHAkPtlEyXatJ/T6fnigmOAkovLS3rVrZbn
2Te3nC7ghJIwJear7Hyg7z7mKStmc9TnsX/8Q1YZlSaCFUSeRB+kgvaag5zPS8fR/hssPFsT7RLA
jFld3/rEplP1oG0mV4SgrzSHjxfP1YQ7CcTUvVkpWtaO6952CUbXmMASk2kcF8CIcOQuxbUO5b6S
yc873zdA4Hb1Gtx5LCx92ukbi+/uUFmXaSU4zc1UwVqZ036I+zb6FwR9n2BLUnOyHdB4W9AqNqML
1qTcHXkwQl5agFxS33todrX5xx9nJlphbDSUfLheVMve8eKDiHmafXk9cXu+BZVOeuyi/Tk1/hm6
/z0S/VTr6zE0ZHy9OxUfRe5NGf3sf2pddCtVHKskKKPxc7B1me3+VKOR0ecc5hJxfRco9K3ZvCwE
thziSLuyVtqfIZwbiAs5wJ4BBtuwOXeu8PUcvA5dpM7Tl5d1oc0ewfirrCMqFu2Q+c8OILT65fJ7
xEB7nHcKweSGDVzFmlDqSKJkQvcQKcQjeaXNJ+XlV995QZxRMBnUfdef7+ZdYAU/a6zI4oUDpEOs
F825TCBmw9DHO8aeLkJKIwG8LAPC1RHngnMI62rYx2ZeZ7qZGMKQonoRl6ATPPWXUFa13McBUb3C
pn61Q2LVouy4WIAIEgC4o29YatskdVCRsc2SsG907QUA14PVGM04wx26xtCeWi2UEYulhZNVl/TW
8vFwg7FIMnaYmZynJ8+P3V1nAB9Ce7Ws+AQq/b5L6jzpbXeu5akJIVmkBLyLV+ZtRWe1cskJEwNf
LJL4KdjbamHSU6hsCdGxR6rw7OHFajTjbAncdANnuqnxEdKtMDNBvjAlaP+Up+KpVKQGjkjVRgTp
XZjFGWYI/9zmd6MAmanGO1T5d2zFdWAfChFQxg5Q+Otn4vVOAquyml7MWAnilqBcMw5pXXaONTP5
ZcIvgZ+vg1YhFhBhRbc6/6ZpOlf5IUIMRmKoMtoDPdMGwrlcpuXNFZr+chditjsrepmbgo4OHfT3
pmfsl42pnvEP+gmCsZsUfV1IETyeJr/GpAPjxOivUwKOGnN4tZZlElw2wVa7cq4BmqxJeZ89wZau
sv0SBIWkrrgGJlO8ErWGEErodMZpBHrS8rKg67wX/6uDsj4rKWMEiv3FYy2EhHc7LPEnMAcqlZqo
Mz8uK7NTo5Aig8X+0ydMH+Fv8QHM9bdK6MyZg8JVFpA6Pi09m2V4tiBf60o69tOqpNp/y9DldZaF
kpv2BFptzK6ZBEIGLH+ZEBaugQhpT324El9sb/kk90R524NhFhJWBF+2aTQUtGbIzAo6R/+jaFBN
Ff5qzrRHopMUkvc8vb62LFTHPBY1ntdvUHp/Vfqne6FdXJU653ui98iDTN+J8ZqYvzNsQizSXVj9
5FnD8LN16IsViVcIh+0OwPLJRidd15OLsxwRyNltssPvakw5nqiAmRYF+VJ4AbYBb9R7bOzFmqOM
9x6ARWZuJ/1NSmNIZ4uHLgvgJHi02kJa7TtWdI2RxE3uVznegMiaF9fSwhcGYOc8+l3mf+j7Ll/D
yxi0v0ELzwezXomb06Nb6ahttX7LcdZFidqhPAlcQjFX2lRckyVCCin5aH6gTr2lp0ARlzdkHBSd
L7Pc+5FzqoVvS7k7CwjtPJnWdRJj0TQiMzsmH5Y5sQldnqi6JUSP7P49Uk4IiRAsjhsDXj9AaUpp
Y+GG8X8lR95zDj/PXkLpzLB/ICRSlX67NzIDhTlcl1qUqyJy5iN1oJ01HxRrx/pBQrC/Vgj+Cydo
4UQMbqybiz1XTJ2vWXe7vHuwGOvVuTXMOf1gmUm9JLGSkDpcJWVwOGP6grj/cBJZqYJSr8WQq6+R
iTBYmVxP9NvY1lsc0Wl4d/5C3jWSbu03NwtbxVmlOT4+MokegY8vRhTug0g+lS7c0CD/DnDrZ/Fj
4R6PiBEQiVako94d8GZWoWdlW5Tg3ngtnqz4uy114ckWcZEL4GzYy5bZ3cRyAP1dhoSaz4i3g7Js
IwzVuHq5hTHChS8AnJap09eRmX3Z0L1N7WZiZ6iouUpAnmtKWbP1HW9Ra58OwBaHSMIFcPhuUELs
3ZVx2kKOx2I4w+RtTlQghtiIzkvD4on/U64ulAqF6+L+ypB5FwuFYjfLHWCvCtWGC9nDWIY159PN
TQIVBoNy8NeHmiR1Q7IizTrcaIOnpjQzmZV1iUzyNYg1WNicWI6jvd7gJ7mYzisZpFrxFzJE7PZS
w1ktTlVvF3Q+i8HlpaBuQ3KKqEJhqQRBlOkz08OmbTxItxB+NvLpFSBILzozPFoYGGsqzVzpcMTr
eXqUMsX33f4I0SIKGeh9xeio3SwOKjIbMmjWN78/kvnkri4jBLl/yZXxrInH8TxRq78gu8HsQWJk
tStIxelth3Vm3gpPts8b8sa/W/uy6QlDDkGsgi0olMOfv18MKAWzs0X6U4a6K194+QtvUC/Ax9yi
jWLNuMACpIsR3bkydMP73QQwXKY37/gMsmTSvjWsWcEJOceyMJMJevZ5oNMd7wVEpCqysBNn+tZo
ARVuwwo7h22wymmXDklJ5z5YmNv7sTSCinXU/gvA8lJ2mj83HY3RAZsfk8ZEdz3a7yGXUUR6Jot9
xUwaaTH3BaxSjqXUM8dNAjAUOkeByXhWk6BDvmShqRGsIiGT8NDhMTTQ9UBZk167gN1Yuo16M/tA
4Gp8Qg4bCCq+o7RwISdKpuBmC8ywuuy9Ghz1EjRtSVNRQ5c80S3yNQH5Uq+1LKSdqRXhNY0XrXvl
HthkaSk6UBXfii32USbFKx0QYCufJwh93YYupLAQgLviVg3U7UoZzT1TZl12Cd0RNozy5SaTZBCF
DA5qnNOa0US0plMQDQPeREJmZcpHqk2aVlN3wdy+02QiHFJ97Xm7rHmwWI/3B7SNk2I92Ek9V7Ni
UJlwFxnY+FXO0kbCHTFn1gz1enwPNQgckfDCZUNIWhKLxlpjUi+H/ATPgVALPzZzKIsuPx/cRYSs
MpknpzRKbW1+8HG33PbQ1Z14PrMxcW+yUGd25dxeb5Q0DKOiAbH154FsPfXB0tDYEycQbE72gqG7
4OaKGsFIxmVe2iIYXn3Qvx6soVJAzORJKcMU4x+DyQCgzHFynSVh6Y5HnioDAq3uqMrug2jIhctn
RYFFPPvvyXH94H//OI1sulmlfRhy79roXZnc1iTZuq85N+bVHSCEnG7RA58yfqYf6os/jTzExtyZ
bMQRXaSFz+eN9GzhZ+lq36wD3e6eEJvc4GtoPsqStYQ91mA+MNmZY+YQhV8G5SoLDaiKSd8ieCrx
pCKyzsy/Hxga8Z0xwx0WwXFW6eI95HN4QFAA9EI7HtRlBdHTDQNlKPteBnswj84UAV7WpOfAojKY
Op5qo1Qagx9w+Ry+nK1fe9b/5pD8f0KTTLDmNnYl6i2Bj8V1CgOzTGMDiNxpsnMTIBbWHmLMoEDb
x8qVFduYcmZs9EVtEKbmON0F9P7GdXiyaQxoAYF9Knp1tiNzK4qBSEcu2wbZnZ2zOdlwIE9I/3Y8
fHcIDK+BCzkb5vla0H7MVzvp70DL05i11cD68e5HtMjCiVrXPj+l/4F6+J6KR8+guldzH4wyNrcE
hFVGAm7Gnnj8Cc+N9ADMtptS6a6pjd3hMyGXBO+DVV4E0PaywaJKvdOu1tSBwlowThTBEjEhyZX5
ON1BtjBc/U/N2i5KbExhrCKtEM2V6p9wHulDeZwn7gQfvfS7l8zTG1MqE3seLIDbU2QDX3M2g225
6y3sTmJ9XAczNYMVb0joS4qPVT4PITdp4nUVQCQAYttHV18pmR35C4CNj4S27uUHMuS4LzcU6vjf
hW9yUspXsT9FrUdzMeXY0eDj/pPqpt0UUdquxVgyFZEzQZpaYc/MweWpb3btiblPJa5/Gf1QUVHf
ZaKuGSV7JRTJqdn5UNES0Q6Lb0dKBBVuyGNrlEtFHm8pU9HYhZZOKULC3FsoMCL0XyzYWbN5Ayib
wtcE2I17uM33oXE98BLO4cp5qBT6t9+2tL0mI806YhjJ3rV/t/npjd89//ji95qfEtSJ4C7oHw+X
0eUBN9+Nemma7gmLYUcEA2nMDHoOtoMryZRdDysRpeVCnv1RX9rem80By5soVirkzpKXMTJedxBA
a+xDlxU3i9ZW9s7O8a/jddXnMoOQLD2SG3Bar7omlHxVYMhzcJA93gJxW8yt5vkH1v6JY13Xc3w4
gBNyGSwEC/RklEhcdHzjPwci3ZaUkjCzvejIMtzZZK0vR3jZEnotgazoZrFeuNeurbJxfbkpJOMH
clV9NSSGyiGhUTIpjr2c9etgMtITBxiDs6xbvB1g94NjOlKrvpagrVVQLAq8ZAjsn88cuswbrrL9
y0xmwrnkS9yYwkxWXohsxbDzXRasdBlH3bZgSD9fR0GdcA7MvRuYE8I0EWIoKVK1h/Wwp5m/OtrU
smzXYt8AEgtzvSurBxspve6qFHka229hqhguvqkTz0bC7foazYdBDRQCjJWn44zm9Oz1wXFrfbJf
v2Vqhtjk6HZHJX29ie8yErKQoA9P4AGcKg5cvjcbbMZQOAoSASnUoPkd6xN5epEcKrhzo4DkK7sJ
iqaUQuod70Mx0hOIirBrKszDRBv1t31cW1yTMmjLx2gyP0DxyHY2d1wJtVA2ra26XxsKGppiP2qp
VKiQX6bqyzqFuJJLAo7wg/PdG3HqQjmYTkw7fPcCDBVmdH6XeJGTrpvm+0A0V2vD36hZqErrERLt
2JtVHH0X3YhIEy9mAwoVlKgZ7HbdX7X96i1c0B4sEI2XqnFFjOQd52UVNQJsp9rSr8yGEcSe6q6C
opV4OcOOpH1ebLX1KYObHK5PiGLaBfd4VZUIv3YtXZ1IGWpvstjuTJeL2t5sDOjGLGLKt38YFskV
eWR9xx4kVdX7u3Npj9MgWY2XZI/wFUPu/cNAg6ESRAXu5hPou/mCngApBJiqXDsaLN21vBZRAwM0
x6HJEpEpS3zv9QY9xaHjmALKvlr5QsewA8YdLES1oOcsoRLx6EYGftJaTz56EPGI31TiP8o2QA6d
wHFeUcpQRWYyv3bd22iOQj6pwjxUTeYW3vqO1UXMiX9m8EDgTXeYuw+kUiqTZQkwCT43ZzQlomDq
zu5dvqlsTNODwja4a2m8VJUqn+Hq/nRPmQXXsa7MMWzduMe5mJ5t566QnSv0ooMH3Y/atTsj7Rsd
YvOMwZs3bZQeOtrBibm0ZgXi2VUc7vABDx/Jdh2adEVHPL8Xe4Nd+qaAWL5ghEFd+5NEDo0xv7kM
itQ1KhZ1N06SuuYWm9O+b1dMrXpF4XjiaEiVYWLiseelgLpqLmh8VdfxX6ISbnpV3x7ZmvGQHpND
J6tw2e0BiglODlTLDzu82mfhF1G5TyqcWBMt78HHMU4LlQpx8FqHC0GFDGS3Ov2viFwEpCVhIWPA
lXRLAIWxiWcSxTP6khf57G05SQ0Setyix4HWFGbinvd7fw4/twtPRIciBzeIVvSBb0pMIHRbbaWD
n/aw2YdZrpAEgIYSClh9wBOdpWgT9CiDgd5s15U6oBYwJx03GHSQeOzNyWVmK8t09a/ZyDo5moWT
N8F/TKiIraYvmWmyjrsBrVVM90kCpNyy5kvny5Ml334iqBOp9lfheChi86xrpBijtxqVc6+XCZCD
J6xpoEvPEPDm8eT8X3a81DdW5KkwmHLZspjnERZhbiEESyGM1vlFHuy+YH2R28R8cYuiGnWE9VR9
kOtF5hbqKceIhTYhJW6rFeWp2L1yV4h3vIiDmynOI5hLbrbOF++G0oT9e2SxBJCKl6/tYpUDRebt
O5GQeaygFON1VZ9wUM2FVx2WCuUXuhAYepAROXGqDccn5MnGa25I+b1cSQsFnggZ0dK36MowaYNg
0WOvLkpRGFC5FBEZR+hkb3/ITbWUGm/OWPas0BSkq4mvFIsz3PIwc71A+EvW4qd/ZKQ7STGA28E6
/gX9OwxJnpkUACxcxftreGcFoxXEXNTSESP5Td6OSrSzBVM4wVQf2JOt5nIWeJAkjDDjmF3ZQPC6
kjwV5/54fAQG8okci+fZTvWEeuC7QGKOjd57dRuGxxJAiPz5+DCx7VdIWVhGS69Muxl6zKti9kjg
dEGzAMDok/kfzmgtiAVgaWWr0iRwiulmL7E+0UBF3TSUg6Db5qwe67uZ9YScB40YrmqDSgDT7RCU
ss3thhrFmOfs0D55ZuVPYBTZ8LzgTmWSbX9Z3lJX8iQbSdIoSIfSg7dhHX8SV3pox8hOWbArMuLH
SRksKTF4okvGXbU2Tw4a0bVEfuP2WnYSDVACXLqW6HMsOfIFEWS//Gcp0smA3LiTlrYaRPGj+Tk5
4Bcg4/4+RbzoyV+JDsDVZDHhcZJQ9ILqj08jwQEV1qCsz8PF/Pw2Gf6BwTzG75r1dS94JAly6AUH
TlX/AWD6N9kzrod5uwGKPQWnsFM/IhP72iwwSFBwOa+Pb7abc3S/3fUxmqhfEnxHlpH92SpAKUQp
CJkJ9S8CYPLIcBxNH3+qzrRIZNtOOt0tpPLBv7LKJ5gpJAN0RfZPKy4g4bhs3Ss1gzZPjAZtYAEU
AqkA0IHRr4kc+jyqDV5PtjQ/ZF7U8y5vNSA/hLnFOQ+WkCBpyb40CfGDncu1jJiudB9CtGTOFR+A
QmOj2xfJudNzbk0NNJkX/q75s8xiHBjPEvwN5vLMRpAetvo3zCgZElUfIzhmSf9v94wK+xew2DUj
TUFxNKF1lWNFUh1oR4EzUanUjquUDtu6mZI2KM0ikC5KTIcKa5B7qsze/4QDu6pbQZje6nFIp/Ai
vHtpWXvQHY5mS9syQykeMFhCMaL4DnbhyOdE01CnjWzT28zrUO3yO0nHXF6DORyqakSqCRbpZXxs
MfvIfv7KzypDnWJrS5jNHajJO7Tq+L6/GE5iAE+EGMFBb/JVtNiWdKUDjZzhiOhpayMqZ3CAuO6R
h4lOvUvCpB7ZTaJHrwiRFcmwi9kJRYpHopOxR5+1hNeehfq3FKlOsp/UwLRrZlalP6isrHMkWhLg
8ruHPLedkBzWD+9nDgmWMp8jj9GrHun3MwGYYe05yO623hYqehsWpO5/eIRsAKD/rEfIGnjhN3jw
h81JL/9J8s9Hygvjwy4vjHrRt24gzPJHdWYQywfwGxyMd36k+zDG6DKmf07uzEWSVvBUbJsk3nij
pPrYeQvdyq2C5jftOKZK8P8GJ7WSn6JaBGg9A580kqf6pUk7QfORZwiA41YT2Xy1ptih1n+ds7yz
LRuyDG9szHmen1LJvp5Z9YHfXsEseqBVw1uixCLXwAnjaB/yoGnZnXgb833n5A9pcmhlEaIEt+Jk
VgfDFwvoOemaFTGSwYX7qumzaYxHdlhgSJEhaNk47EhDo2CjBQHVauMPO9w08aWF0ojwg0pzCJMO
4lcg8c3rO3ApxzaOxJX9FQq6LpRNAPzuz5BK5rpzrXfDqDrcomKApZZqZp8NxhyvEeOs5B2C4KI9
rrWf+lst1w6eADqUzYlOJktnfVJs+Tp8DDJYhDVhpsQ8EWQyvGtJKy7NsoyKGX/ZDCp9z6BikoUG
b8OOAH65m96E1k4/Fs4Enwp3BBxJduTyGSp13f3eMRxgEiI59CgaPZWZU7ol5wYJHI6jCN7VIuxR
xyNmyMArmjI+xspRx5zCPXS6EZdWuDiKbtLKVvajSidCCnNLSyacJ9Edayi4JwXspeDAE+BojeMc
C84an4wg9j7uMvr7aJ9WQzF1xEkE7GCp8savrKfq1Ry1wH/WoStTCxGHiWqd8p2XHTTyW2ltKnAC
6qH/Nccx/Ib9mggbQjyMl7kC7xK/K7xSnD5Ih5XfAAMjEkx6YenFvvadQwDr+MEQPg9yohiRYFNy
ySDp8Gu54p+WrULJIRd2a5VOUNveJ7fvVelPTaaJlG+Ggam4tlao+scRVGBO1N7rC+paabKz2nh9
zQp5d66pULSJXNFEI097uYP5jbVwdrrVCKiZ4YSY+soU1mUtRHRqKDAxmYWe4To4dOnxbQoPA4dl
7fECE0Lc0/A9lMYDEy6Kn//UCWai/Ortx7D8lySSFg2db7OCj/VcKXVndOY1mcBFgprhL0wL0/Fm
1ReMYI+nbifjT/gGARcsbT0aPl70bFoOHwV5Q74XUOK5OngPjbUXGsfqQdh/DpJNe2FgP4zPhk+a
CMB0l6nT3XRDKuYlJfFWu5BFKMAtDa4R6RD5Ri5x+h6WN44f3XKh3HAVhX/YcxvfqwX0PPy2L5/k
QjTnbFP8SpMo2fAP53nLrNlJR18u+Af3A++PXx9I1eHAOgjh0hJ/dFhTAMNnnb+LgGeU0oWuco6K
HQe0QAqTFBlwK4iqvUKv5c59kSnoNlzKOu36HxalECf5CHJqTQ13bJU52NOfzhGZDcWx4S0EH0J/
+zOgYJO/NUy3Yku/8QtqPlu4HCDixakNSq5bp+yDtLCjdRvNMLYz93mRuBT+643arbxFB61Zp3Qo
GpBEHwcluyRqXBsauXbmy4BIJSXeWMtRsZbvXZYUK+5NemQba+v3iBUgmhWSfoN7arq73DSRk9IW
4BxAjInsiNRScJYKgCPX49MeBKRZHhsnwmmfxqEzlVMae2OM5wqXtZAL7p6XX2BjD33cXfO0k5OC
cfpcLh+UV+sdWJu2VEnns9pDslIEaV7iUOSSV2r3tQblWcxo8ScIbOJATCuZht2kSXjau0qXkF8n
tveXJEoN1VDfnmTTa37lknEytj9cwrwClSibQeUZJuJCbTKxK0lS/xO354/14tYTSZXl6+YrWGZk
tAMxoOQ9H8Ir3/52G5wVnDWS0PGhI1DK6gjvbQ9rHCsNDKCmdpuG+vZLMJaLpJX7Ll/74kJcIPIB
HiUuej62IyveZ8ZAjohMbYAWWrjZjxJr+Up6KCRqeNgdS9tMVr83FucPqHmpC0zE2S8hdHBX7IxQ
d4OtnVvwCQHZAIT+ED6b4UomCtMRgLUtkxd2JgXRbtBV1qIX9RL/s0l6hwlSA7YU0UFSvdwE2M3X
lrANEyu1xW43nY2hoEr9hUmKN2XJuRG1XlN3tLayK73cjBKcxWfkn7u+aSWaAROX7iJkQ0m8RscK
5mgCwDMy9jAtCtcXTPen8rb3cpKtsFaYPG0Tp+OVfbMpOCDlCxzfk8pf1LmXW8ahIEEm8nF+qIWF
A6GdYgYLrBnkFMts+j5gTlaFUsHcqtVb/M9x42QyZ7g6hK45MtEp1nlfs/jvnZW3K4Ry3MEr3dG0
0tFwrC1817vwhFcmklC61BjjiJveq5wPM9nhZUl4hh5b0CoMwBxuJWacx2LjSblPGzs532ZtBaTo
ORSD3Ko2cUxI8iJSDcKCHBM3UmrSZ59s+z4nFZWbPwsI940dTnOED0cDzChGJ2NXvldKAGrZsY8z
TU36iFActy8PnwBQlULz/CQ2Pcw+ts06fd9Cm5HVROvs7qDA7GX7IXvhdhpwjt83ZwfX3v97KcsT
py5xumG1JtpldYeqzhzVvofFdD7Qx5qQyDfkjXRJJyZpfdvRdAzpSIoU1CsCL5dR+hcHlZGSyOCg
ZTi530VV6ic969TevJC/OLCALftB1HHduU4B8GjCT0KV9OVJF9QZ5BgkBCvi1Mf/Yf5HbHER9W14
kYpDDjFatMhkJfsELxQSMPfocD3FA+2rhsm7FoL2h5KrmcbhJtoSBxfW5lCjP/QWDCnbK6TERhn3
vXj0XnPT3IlBrqzS/H990VUG/jR4sW4mMl1kZ1OFGpwPlRQmUonb2tPn/5GNS4f+gxsJ6zEZEUED
126tGKFlkph4KScuimnnZtvqM1Rw5t32r5hYq0VzIayfNpxOoXhXPDCD/rqR/14Ga4i/otaFhYW7
oLGa5Oq6c2Ebx/YPvQamou7lCxNzm0gUwiXpcCqgBlDcRYTImGH7CXQUFca2dYyEdWJ+mjOIGCHq
n1CjalTT+pd5jyyrgA+oFQbUyANSTv70ddhUfu3kNeRlr+krvs4S8s9KRR2pp83gYWyTYxWh/L89
9ZiicCDSQ53Uo82wZFnvpSr4PLbr4GWeuACycqEl0NMQBQXIjhiwyJr5uwBmiVzYMInTDmDfPnlH
xCDWhAkGDYUGT4c1dBu4vU6y+fhkkBqXMMSVIlu+/gXfa5pMQeFKq7xBo/z80hbhO2EAIuY9ABnA
85YaBeruAuq+do++sAzqJf7FAOWyngOC+IXmh2fJ/WNYWTkTSvDWoTv7MZvTp6+2bFYF3+9+jf+q
STgMe9ZtPNRqZDWoqF9kbZFB6f3NF3kWe9w4esBKCrdHRr4yTLIeM/bONJwoD7w/nfhVm0han1Zk
H3oLMIDnE1NeRQRUWO4mAusvin8WxoOqQleW0H/C4FZZQgXdFfPMpMEZBJ7XJzUAzOouOIxaLTf+
27wwLu3qTip6kGyglbWKdOBajm5x3KL+GwN+CXBK4fpdE3K2OnXUyPmqt9NmRz7G5zsXqpzHN4Ui
lyI85K76YWDe1CfwNzoQRbMOEFPxkbDmbmjlP3CCJBjkLC33ES3s54aRL9vgfJzfBzQWI+eYqYv/
EB5jGZCwNEJkOd3k69QDLXRJUTpFR4rXPnWhb7r7xKjJjs/Xtn4ha9rcDar6XpFVg/wEObr8W0Tc
ueFnCtXt6P/a1jyCNS76posi/oTLJkwoErSwTLVgzGg97Np09zyvnPx0GzxK1B+uXjZbU0WufF4B
41XfTCtDePfZ8d7kC1v6r8GuaAVg5IbVa+pOq1JetTyiqJ1EUXGbYcUoNLzw8brD9E5CkZ4h3aB+
GZQYqFH3zAgjhtVIw7bXb//97Be92aXxjOK0w2H8TYL/jYLpslUL8prdQ/uCmjEGX4C3r4PzYL6/
BruImKKZ/PgnKBD+Hql9mBK5p/zi+B1UqxPZwvw4z8w+WLfpoMWOxVY95vt/6Ire7mBCHstEvmF8
cP+VsFEeOLPcsujTolRGPcYbEnOKEGNwWFNX1aI+547nypf+EtREOukgIVJgucn4z8y7Hwu7YQ6X
kP3lO4MXyxAO2wiCadwI5MSm1qI5Ovse6NhwCc5LsO24dWJ8AjyAAaBh/HtNbLepERpx7TtVDoeP
BO84J6Q8aV+4mxtiFxtpEUMTnSf1jYbNqDiu5h89q5Si4u04WAFu7wXKVskiWQwb1A6TmSR00gIA
8T0IonlDtKQxTA5HKyVWiFAmUzhlFpz6E3zw3j+6WAo+Z95KHatKMdMXAVNTNdNdcZIRyUL2n1PQ
hKzfPmFnAGaJtLEGk9iIaFqu9GiUpnMHd6wfEVthNMapLMTDU7uRAFSS8XxByPs9PRMOqb2YsrA+
hOBDcUyeHlq5Ea6Qgrs5ZUclbybNgQu8yxb3R7v86SgyU8byWi4D1XrhLMJ+zl3n2goaulbTJXoq
bTszDlen+E8R1LbJ7kTzcSBc3tCsW5xhVHJZvf6mJFNqHQaYNygWnjdAP7mqXnXhksrpafUlMb3Q
uIcmT5ePRiZB5T4aM/eQwFE5fXnCOdCC3oURKZOjTqEyH75L/9xlVCw3QwwcKwkPtsb0DfIBX7R5
PbgMhAnnC9EQiKK8rgagIgyEN5+cjyN0+4pivv4P0ymZn7H7NP7/HwBxRsrmoKYQo8r9QUAZquJ9
EJC1c1XgVlPkceFGlOBWoaRmc1JSJBZUZPvfjzZoIrqpJDQ8S+m/nQgXs6s3jw2QStiVgzd7wTe+
rTOsD8o5ewnFh6yvOS7w86x4valYOc5KgfxhuF8pVFssJhnwuFpxn4sugwEtOiaDXUjVtjaB7B/d
ezplzS0g3BWXtxKv/QqQd37803hW7+Wn/Q1L67gRllnXfmohtuySA7Ca3KMXu7vx3KyynAxkpMMw
z+HOibLXw0ffmDk+bKXqRVVtYsQWHbd4HY9YOGVh79SG9qVhzSsQ2SgMIis73sQvv79cfUZhD7Dy
QhEqC66cbG2l5RJ9qRWKCKac0mdsUby/hZgo96FOkD1o35xPPOCLU9mgpW9Bpqau+hA/RNXtOhHG
WT34jwwFWwqqDuQlH/HG3DWzlDL2HMO5jzR604n5e7Nk6jTUPz31t1NkHNmXhA2P0z7h2UxheBi7
RF+qieYgv0OlBYdYBU+nRPIJJNEbpNODld8L42fD1EfdhJN0EdcHHAlfa85y3vEALB5SbJmLeem2
k0xZWphMIYLHTaoxykyFVRtpYpb2A9vDn67MvtMREN/3Mw26jB9u2I6/REEWYjGf1XRsdIUJ39Gg
jSV78ASafDp1ArIe19ufLHYg7OUd48IzJhPv6clCY0WmWTOD3KhVSKm7uHTQg+O8B7+hDAi2EP4t
+sZrBTwn0GsfQrrcW36eCpmYT2EMdrx9/nepsEU6nHDwzZ/Ebq2XrGc7pwpQmKsAbSWRaVTYmL/g
HbvxDN2a+4VqdvCB+ucmGGOnf9QPY8CsDGJNXJRYkB3t/bCtp0ipEjr4V/QZ4eBsqLB+ml1uUOtJ
N0new4rHKhQIf6hUd/m42WWNYTrQ6f+ERMZkfNM2/M/KhobxPzyhFg+OZPQ0Edfp0idgObc6M/Xf
GV95bYF+Chqcz1C3jVZcAmQO2rzBi33RBZhEc71YJS4nGsUBldy0by997fnsm4BNDgUdIZ2bNa71
MwVuU2pCfWUhL60sYMue+8iTbatIhDj6mqvDz5Go528d412sWC+v8+dRjOawLKBPjDvKEjJTVXo0
1iBCInV3wa1bMMbOTu9WDkVatR/URWj1z2+LJBIfUtnjN7QyFBWstjpOAgL7P3md8xzAsroSfKvd
Rf8KfVHMaLAcdHINr1cBXaJpsYtYQKC72nHGx/hLeU4JbiLsN8gIwruhI+yguf8jwX9kbWJ9VsKM
A9byZuHD1+VkxwJnRl3KQzQQ2Kv71UId0rh1wHBj0/GNhvR0JpVUA5iDoyFWVwBxnwUFzWo85ICn
pPlmYBTfES8tUrFOPSV9lS9v/TLBgQdCIHvhn3YZpbi8QPZrZSpZ2pD4YfBgCiq5J/Fh1z2kesE8
55IjL0n3N0zAoFdswaiQJl/e5D7Lg/DfzIkTh46DoqpwywfC5cSPvEn5G6RHbUpvfLja/1Ck4xZH
3zFr5Iw2DMCSbdPpH42Z6MpxtezjsOfua6gz7ctnrtHTG24i3D7HoErs+WAF8k0qEv4yikxxPl3B
27mCjYPbH0GZhCArRbj1VbqHaox8draBO6AjrLuZPnChqrtVibHrnK6vwWO9KmBCYcT40JpuAlxF
OvrmpyNGUHIrcXLM5neHV2P6wZTqF2W5iskowgVZXSA9bP+UuFYP1AUnW/PL7FSs3c7Xr5TuU6bu
VdrFS4L6Z2WAHii/T6NlZOAYS2d62jOtKo1XMNpDcENCQO0IoTWc9VVo+xpVrbPsTwv5+mG5CmJb
9tV9B10p26MoP1fevSd8MBh46k6ZQJ+pxTZ3ZVmoCoQbKNg+WRJx34SjjZflfRN2vFGw8hYZ3VP3
9i6By+BZgQK0GTbHUXS+/xqhgPcaMK9ohHgv23lVEXqT5SLinW4UkTpgc1kGb3nvotQdMuvbMnwf
l6d7k/2mROO9mret64zmolVOHv7zx/OnAhug/Q40jFjQoGH7ZwKsoUW56hhvrwLw5AAszoPt1ZEE
IB3f9lS6QQEkjouW5jT9hr0OvxVuxJnOhYiZfevY6q5MtxEXnLw/YdTrnCC3qJU/W5AlaEcJ1Xiu
D3msZkqHk/fnuKmZblAwq1IYP38UIUCsJAKdlankHSRp99Z0c3hoeWTJdIicr0kP4vuSKIejrcoW
o+gznMoe0e9xl1p44U3f40FwYj0W+oZPQYqNLhZrHDY7NpljMIOru2kC60LWym0b4PnPUrNSQ9t9
P/HtasZ6QoOOREMC/dcfUjRTibmk1ZoDYS2hVWCXE7Z1TZxHM5YBXUDDJIqDRBi9saj+YdAjb04l
hsmpckeDLTSpiQ0zDrQ1KdzDIrzIOWk3FHE8RUP3bjMcTyFW2coEsnonfPX5CKJzoF18S53nd1pL
PIcrYiUY0eZb2Q9hjwb55BP/2/quIAdfsuh8TQGatOZydZjN4M4nMj6H2d4Fm87rFZUo4yjlkVv+
/sZ8aYm0H8YReKZm1Wd3bUfYoH0MDn3JgVXYA4zaojHVE0dQvmUDJaK3JbbERvvxk53f2vdQVRFK
EkQ3zji16VrImBhD7HzGVRpqP90blIlSq33NP9R3jHvk/gOsMlgcvMxJtH7FMDalCQCYQAdOjU47
fEfE1si8FoVrYLjU2J3gy/3r+2XNmO2GNZKkeK0ghBYHwgcYdLnGbbvGkwykkDuDyB+wxv5d7zV1
g3YSI4Hk+63jnN6gPL52NP6MktSIoFJqumw+kD1xMNfhnu4SWPYV8r/C3zw7CWkZC0Ly6vT7owic
WyAv1AlCHAVSOIqxdH1fNBT+DCgJZkxIL/RFWhelElOucpoGBY2bVrWnvF2V0uwsksvUT5xa3xbu
AK02ChokI4/gn2xGtko82fvD0OxOcVjb5h5W3vyIe2oXycPsAKuSp7dshBe8ZvkPsrQArkBoEFcs
6xoqvN5DVUWzP5/RYR6NaiKk+YMRLuJZ8CnCrVObH6hOV4mkYZz8+WmirN/EaPEZ8fTW0z2KbzPX
kVrdlsplNpGVk2S6tMR9T+SN0LPguJnTyOBa6TNoqD/SnNEXiiz2MGCdY8cyMCA9YuA+kqwAZBiE
/02Q+MW7V6AcuiHROZbhd6tNz60Ueku5HqwXhVBa9doYlkRbT818LLF4zQf7WfDQyJEC3L3Brrfz
MFI/1oQzoD5uL77hR0W/z5EMC/HzsPSoOxvQdSFZBvUrx8DtJ/c6C5KHk6vMaAWttQ7zZsM231Gh
Vyg13W3eSQL9UxivSfO9DehyXx/YtvNM+BKCai1B0lrZ46Idb23UHXhvxrPIMyZmoxuvXghnB6JU
JVndvjig8u4la+qCXyd1PX88su65xW06VzEq8lxVvVqR/lF0i6ya5NeTSqWuqP9s/kqdqF1E4WUI
VASVKkr0si4MF13DjK5G3OWrnu8gDBWa5a5ZqmW+/7sENGRd74ugoy/eMpKIQGiJKcNcN6/J0mht
bCfJCcsmKuMVKBihJ/CYYtAybtn+fDs35A/nBnSRFRhrgvjOq5WVVQyfwtmDda0SlfDQDyICdhQb
DHAd6Bq57ApEiR9CZSv0uZ0O+V+nArILwMMdT4Y+aX3apaam4NS2vmpFVHhVMOoerAPwJt+oQ3Pv
NfibIhprmF6gt5sj0T1kXVXSXOiMiTWYeFSkXd0lXNI6bhHT0IncY6hSGcbUmfsvB9iQa3myq/Zc
fZMj0fRzUuhlDw1sZJNS8JEjO+t/BIIhFjiYqI32kCJNwUDi+rHKOC67eTkV47C7mK6YbsnLrvTw
QZqniGy4Ve8RO1sdmIYPDoqvxhZ3icZVsdTCC5PdYqnhc/TZmFpkXyb4+ZoQI69zhvmu9G60u62X
Evf6Bt/5BNWtd+DDm35SOETQms0ru841VRR2YSUuFHdK/sRVMpNYV8LCX4Rjwd+LxyUAjSDJdmil
ouQtsTfTMfuZvAEqynVLOj0JZfYC95SU8APwzH27XbFNCpZVvu23nqY/PluubpRr9jVx2TCtntZN
5B+JyvVW9UfweXwPHAgJr1KSqrxGUeYuNcySj81bcjVIX9IVUJ+5yrmOWYbUscX3L4qcraX34Kgw
i0n30SWx3md159rA10eYlZam8iF+KnF+OqaneX4r2RUMHaKVHaX1a7eccQSoKWKBddD3v+4ggHLp
s1A128wCrCtocMTO1uui//tDaaOm4WX6EvL4makzfIOv2fWzqD2x1ICQLaTthggGasVomy6urrSJ
ZMe3LVi7sBS7E0BIly1+D+2IHQJZsm/7obJWJiAtqk216n7jKQ4flif2Op8Xm//XIHgmDiieobkV
Z8iSMx2ABwl+x9QNPU+Uz6Mq2YMmIZXj0Cmq7K6Uy9XLLa0YHovN8Sa3pceuJdn4a/pGIGtotfPu
ByarmO4E5dQjvskoGo2bulCqgPlVCtx2kZey3oqGNJ1rxPK5Ho9DKvYWYTV/cnzMU+zM8/KnHIcl
+k6meBvSlF/TR7Zv3zGcWbX5cekDmv+D0hSslM1vPkM6HnwviyBjmGKqPCEJnWa6Vmqy3pXjpbMW
IiuEx309tSZxITTUk9hBT+baDPf6rpbKhOxoKqxvVLjHOPGBhI1WnFXI4DJNV38wEhqsvQLa65FJ
kGyIJbp35+M+lCPgNDOoDBjVSwTWz2CCKHPD4OvCD+ox2tZz6m1bG57FmCl4M5r/RKcj9EP2wiqt
RTUE/gFVc9LBiMz6JNCVyU8zOHLYT3Gk+JBjHizbFWnzqzV3nQSTcvylaArfhWpUfG7Z+Gk02uNF
dW+Qmuckt/jYO/dZi9YhEfgwaxLGQ9u5qdy17d+az5CGnwhGrACZlcB+vEuJ8Mtr4rpycVxhO7hM
yVth/FFrL9Am26Yjol/PubFlJ7hUDm+mKh94lloxGahBP8K5ZT3jO8NGf8ywEKOidkN+HKGXTi2c
VkZmU0xESTpzmxf731AJ43U9V8AbX0M32JDq7OPRyFBzw7rqLMtAZR795tUH+tyz1HUhRuFEBM5e
CQyR8cj3HhCzx316CVGIFx+ruP1+EpdDk5kyWAIEpC7JXX8yMcIR1hH5MLwIK2D4WolcuYeQ9rnx
BnHS1U5ujSink8aMJI5j1W8kH0mUjgmT5Xkvzt4UWryt4WOjaX64AohDf4lQ+U/6y5+wUHa3NXFd
SfnGDS2KUBLO+la/HtL/NkMUyydm+7KzmVJAQJv7DDwSzESKkl/wtGjGtp2dW/It0F3XWoViNR86
rxyMq4JCiXuJD8IXptJX5swb/bnd9jh2ovhrlmZ5CTZdoYj6MTLBGPEjCayVxoAh30EgvPIXeASt
EUCm0j4zLYfAF+huvqH4C8/Edak3p1hZCQqXfaEdC8AlJqwFxjJ9vIF0YMZL/ZzNT2Fgd/uILew0
F6U2kf7RiE3kh+zD+qagc8PQ5P675/XMstpT9iyLAiFEaqAnViW9p3utJO5aNuK3wtfj6jXLrpls
C6MBNBkpndaX+8QymYGD1aKdwXaSq+qvTkAsKpHl5FTUydH7nD2k5Q7314pKW877JfyO3yYF/6U6
21Nb9M75k8yc+sHJM4Kp2vAPMUzFkALTuiJOS5AkCfiDUuQAcnSBY2TsIY9pesGDUlu6JINLT9sG
fGtkxJKHFiD8lc+ua4fOqEdD7dHg5lNzgmw07HqVLu+h7lP7aC/wAAfVE9oYE3P6JtsrJ09szmfC
LhLHxlIicKuhWwR3IT/0Tnf308bK0U6whlVh4zLHlsFgMGptPzo/uoUTj7JJ0LXZ3ThkBRFCjLE+
xD0wnTCGsDGFjSvPot0TnFQekJncqvQKGW1lbF0YDoW/HD8mWqACenFxKNlts+R91ZqV3dHr5KSg
L9K+Ya5GNs2b4wZetJl/g/bjEkNcx4cR5GqiZdRLZM+LPnwIqsFAA4zMLR8YTsR1JasX/g4JsFXB
IT3YTJmD+bfv1pcW/2yXjny1LYfkRe3eOMDD7KR7SYBBc6K32r2LKGLRqO3GchjdhM5AlZJGs16R
6QSyYOy8YUb8U4gBhFiv0p930GYFqH77V37E0av3oJLcVvJ8uXlPkUtXBmzZ6wXWSZoDnbGP34DB
Xf4J9UfHBaXue06JpqTYbDCwS+nFucmdqfaIw1p9h9gjDErlqWFHXF6FGZKnHaSr6eu1R7VUN+M+
lZC/3LWgIGtddwnhKcADpF4ms2Bt0pAUeSJ+jXJUEqYHbOSUPLYBLTxtH+7Z3PttamTTwymc8UmO
R+V6r1NSLv+pLeyAu7rbYnt/JKqmiUf0j+kbszOe7BfTEkR0Ac0z6FI7b9iNRdHCgWtSBOdfwAOk
Gj36o8rr4YIpHn3WeegPP09H0VsNODiPfWD7gp8W5p3j43xuXC53TaKPkGmB38A0KqNongR1mWbz
zOKGAkcqp47g4vwPAw7V+jcI7+Bfgw64aoD/IkyICZ/6IDc/31BkPP5uHeWpLpXgO+zoQJBBZxjo
2LvZFtQNo7AcNZAuJ3+xDghPnJidFfuKPM8FatyQ7n8Tv8PVdmzIioPdWi2K++LXcUdJH3VV5jG6
icn5t61d+81fph+fMHdaJ7tDfF9T70OzFCAXXEbOa+pPr50nNuD35FZ1pSyIvXrCER6AFtBuBYgq
e1NkdvSOa4Lxt31RRKinSN0S+HotKfNP45/yZFxXMGVU5lKURj911uF7Lz2xH5qjh06nBKfMl5r3
HOpAL6bDcvMnfE/BrYRm/aGyZf8l+/QeU1Xi+gwrdgltv1M8LmvmYpI+HqU1UWxPUpU/MJoWrJX3
iDaNsBrdrQuMY2uFphEW4sF1C6WmLMOdcUDPuVOdu82P08Qlzlp4B9piv1JVTxEX/OaV393ahWLT
Cjx50l6Cib9x0Wpw+fq4BGmH+LMAJpoTIVaZN27smK2RhgHAKPonqBgB94m2vzKxFGFufg2/0P+K
tKeEtEwQ7yBCQBvhXiK3cmOAERjEJwGVNd1wwDKk7VGowi0l2YpD9M1811QM/R3RyOlepnWIMnpY
zgHAxkn/yK2TLtGTv0WgH5FFZEqdoWCZGIo1aZyPeLs8tFIt4dzjuAc2/FX1r4JcQRMpVEx9qKpN
+o9/js+vEAl6TQZe5rQqGT0yISX/md/Yaq2jQiavh/hqHjGhOWtb4Rr7l4I74517XRbG/KFXEGh5
TVV75EYlkoQOs3/6SYakVgYiDLF8XQwFHRJWJHbjPffT6EH8ZAyF5uvX9wUUq1Uj0JDiUoybsfjY
W0kuw+Mhb6E3jHvq1LmPk+5Dw5OG+2ZmXWKe8fSftc2yB49yRvZaetWhIUUT3WGiQF7C0QvjdUyn
AVQ33mXkHiwxV2QNQYjhyWSwAGZ52ryv+q8AlG1nIw7s6fLP5+o85h5UdlQ1FgyMP4VIF9FjksSV
3UK82x/qO/NbCiqpF+gzwCcAahunTZ8AVnYg93yej+9YVhN8crnp8SLzglvG0ebc408hZlhnQ1UR
G6zLIJUphFaWg32YldQQ+UmefYNcdAOwz/Yz93X997PYEvSjNxYIfpUIKagBZ+VzxphZ4CfL4pvU
8SW/Y6eInZyIG3xsKX3lP+cBNHOHBDKYLxxFvXjWXXNcJ2rjA6pPE9iEt5CAGtmR8ID/sxdcZr4E
bBFXwjxLlv0VbUncXZNDCiafzwyyIrD+gASK01Fuh03NdokZps8Xq2AcwbeLEWTybm/W8cDHJadd
Vxw+GG85uYqHu3u4gTagX0h1DaHcqax4buFa/UQQ954x+oKxldMl0m7YJk+MLvHiinvtLhiUW7lC
cLhDTzAaH/8+uHWJNbrGdj0OQ/6VT1VrVhz8bCWBuJ6iw0xf+w355hQfvShzw8HCTopS6TMqNY+a
8Vo75C5YD2YrUyFYcKTQpB1zah3KuJ2YI/MTC5p5CTZUUcAIa8jFAXmv/yvYtE9yqszFkUYHCPx+
qz6QlzJLxHgZ9S7PzsssmO2smgvU9FPc5EOsman7r2q2g7xIcd233fuLKQRPd+6fl8Fmu/newVD9
ck23EECcMN7m/VG4kXqSRsu9yk48ReaNJR0hIkBVz/yExoWGP3Ij82sxTD1Y3IAUaFrZvaRdQbRe
FHx+o/IG3ZezznrF72J4ALbCyh9ZopiGUjtxCVIW29+282+1q/UdNxuqKBKmkCAoujKSq/OVm0mA
lMbIoO4s5ExM4PZmZgG79mzTJVjtnBWOWQBlLMV9bR0PA6C7uNE888z4N+Y6Nt3EqKTorRSyXFVw
XxBO6PxIDWqo1MQ3djRI/xX/RBGZwpF/EmiLu88kOOLwI0kt7W5Qs6CMVEiI/GfE2x31Jl5slUwi
pO0HtcvCkI0z2gjszg6uxrgGVM5VZOvp5N59pGFybZkjaLmL44BYbje+DfXyFI+obvXhSTMqVR0E
kjVQm4lSbgymdYXfP/wBbvhu/LBVxNwClRD3tEpBZjgOeFbIe9qKwAqi26jpsjbAWYWs1dcCSxWR
/nVpCsJ/em51f/yWuZaF/EtTmkJknHXZmg7QBzE2PU7zJ7vLAQp9cOn1bcgA8LewcL4OwLb0LVJs
HYOEOThn7XYKSOcvbcOV47a6LjqmB3yX9EYK4mleI+E1S8Qty3TiOfSpQiZOhlA5Q8fzGaP0nqpa
H8p8OY/yDeuIg0JBYIdobmNV6B8RHT5Dnh+Nu1LkjTbsriVaWQkA7Hz5kcOdqsyTdkiAM4OpgobZ
uX1+YcSXgBtC4W999guoYO3Y6xTBslUxe/b6EDM6U8ESVbTHCHgyMaMBqkXafy7z+w6sa5uao8Wa
9MdcCH2MFTQTZFuJFWAZsruHF+/fpA1w3f+X2IJVnfyfa6TlpdRoZsoelrITB+B4CLuKQbaubXmV
lN8GS5MDrCKwM/e6ZCDpm/iOvf/I/Jso0xEw0ujvdbhcf2Bpg47lAnp7TeFE6vdlQF1Lm1wVumWK
HkHz4wpwahRgch7d9Y7UiMVxah7VNtdqXP18jkBGPO4ArCz9cqYdt/U4CgWrwcdAw19ttRRW0/rK
5i8CJd5h4ZCYUMwmH2i41Idtq8nfS7hV/TC7ymQ9iTDGAKtjZZzaa7/2Q5n2UPoSpRXnxrbqj692
s0GMzFcAWUVbYskLAXC3AfNSxpP9fmRYwZtN97UbjOxqdHSPnlaBLPpmhH1i71nUjqTZaU2wL2Xf
lznZLFglBD123vhsQQyU7kXFKwj0/b7uY3BzxebFfH2oqc+0WVNPtK9pm/Dh9vh/iFobGXlA7fsm
dAQ2cAj3vyX1BOdzE8oVATG4AGKJlJVQqo1ldmRpErHQLssjx6gojQc0YhuyoOAlYSPdXBpXQd8U
jMmsP67b3tP5cgFvnqu5S5qzgooeNWGr7OP1wgw7TIIexO72jpk+LXDq8bWyJwZSGnV6Husvirvg
ORSwsO2WuiZGLHHNFnMHu0qPrNnQv8+IAVxGdUntM2yecyBWDwBJWuJmpnfR+2B/xIX7/8wGYKcU
rDaoB2wPEwMWDTa4HoAytafqePtjBzgO8QqvE1Beqb2rxbDTjY7czR6wmfqQhwGVVswkR/MbgeR7
x7hBJVOp0ehjCQwC+FyBwDhqpHv620Sr7n6+Zzlucsa9utQumkreGBasQjCwJWPkSbSzE9UXzAr3
Fnsw6RLqnVxj7EGzB5cbxdprdcfHk/savsDNqHzSVG6Fjh3ov9+zF2gI20QVv2i+cEdeTVmapD8q
mYmqeOD0dSQ50K9gdESbJKrGY/ATryzFHLqNcTiLuqPy31tRWd38jw22Tuxcww2l3ENfGi+vH+E8
majsHA0G3doYhU47SDDGuBvMR1gGPiX13XzP6r6vfiCKmukR0lZVFWmrX3lPjcnDcQkijQptt+jO
yKtaLLJyweXV11H8NUHVNLKWB/SGCvQQCSXUDSnUw+mWzIbSkqAJ3OLXzOdEDMF92M9rTvFMO7wH
M8T4RCKOLluHSmnYbLSH4lboP7k6IjBKSBQPWIUfWMmNZv9oHPAodAlihTOanxCy9UYCA/LTYA8H
67sao5a8Tjeh6qKTXMo0cu2W9b1mpOHNH/w5b7udo4dhITl5/QVUgHF6IckmEjS8yo0xHBxcbXvn
qf4xJupakt14+jUQt3QI1wJVVuynCbKNyxXLuhoEcwpmYRwF1eEOsoPvJTvHg0mhpusoNq2NEOph
gujgprEhqQA3X54sn0O2V1C09CHF/Hd+TF45a0VxiTgiwCnRHUyNrJ6QWBrM6G28Tz+P2VnWMQRn
8NACNbFFC4s3w5+8Ics+QIs6ujuurYh+MbXUxdIPR5P1zceDQdmRG0kL3DELT37SeO8jzqj9Vdy0
ChXR8aA66lpT16xwi8uX9p8KeFwKLc6VpURR3rR4t+fxWRnypAxp8odVSuWG6LJgS8XlJph4YhzA
pKJIiHB2KmxkN+BseJO6UxjzBqPfAfkfGrfp8gYJBI4TAR4mE58Rw7GBmQQ+CTN8FxtfvIouOLpF
/XTuivtHDZnQyCfrU7ajyJrXcGKn15n8MclPK6jOUnS90CVvH3/u4cdMZKDAu4Yr6i2lpw2YwCsv
nXxie7oGJQUSHPKo5Yzfy78FUcAIbxec+dW3nt7UbbBe/Bj51LnyVWyf83cwXXcBY5XPEZTQpsx+
ihegUklmMJiKefX2q1fz4vhRXX/E1mLspPi1Zbb5QbXYHwkaWchNCLiTRMWF5v0zYMVYh5/HlpGY
57LUyTVKc0gUN+asApgxkXx0nKuZZpK1jfD6kYeOp+eTwcM9y4T0X7CzNReFzISDsF4B10psoT9Q
s7lrut+vWr4gFNrwyxMpom1XahpUJgvqDbsy//hl+1vMBQZiQR8Zyv+WsoUhr8R1lLWsHxp3l7ra
pfC8gz26nA68+uVlE/lv15+5rzM2uHDQG0oY89CqYJVl17RFrEAW1Xed5SU19uWycqyhShupA4nW
6Jm2TUOgydr6X4rWEd72DukbBys8rlvOYmxP48ifSwiongrhh+vNmhm+HdrXbrYsl4iE2VZ9e+3o
VWVNQMY6nm1RrgAk1ko4zUZ7mexM9mCuPT3cobVvs/CJAswVIO3m8qVLFEYvbL2kxpYAGhxZfyRO
pbpQd0aWZSqR43vFR6xuAAE9Z4DFlI1/fLQWcdiFmY9CmrGJEgqOM4PwO8mbONR9MW6eiT8wg/M2
hyOngk34KGden96CuCphRaavNemwc/mH33T71LZX1cDC96TpyQvFeydaNYUgFYQz7y/nK/4wKmrQ
AzNzjqKJ9cIY0iS4xG0zhfocmtedz3ixxMk+/DlAFNIAztnX7kguOtSrOXPCPveLVAeIWXPosrue
8fpJQzocWnCYLKWtQxJ36QmeSk0JbM43cDM8Bcnv4R7XvbEy5XoFm/YppXJZmKTJCGTD45m+8Pkp
H1YPWnMihawWI+tIj1Q9+qm78YZqMTSACSV7Y1xNK+JDrFId9P+YI4j3VENRSPRFOcClFzbhegCe
BAZU79C0IiC4aDrmrOSR9uIKINYDcSRJl9EefPkmf8aBrBL+Oo9GGpGYoDEPqvwaKRou1tXxd7w3
pEGMa71qPR8GPZ5EYKCEKlkZqlx7DImSmClCw1LXGobP/kVe06xvpYGhqy4QBlqsTBWoJPDEft9o
Sykr/f6O1oENEFD95mr1OP2r0H/xYKtlcQIGH6LSiRLHRFJ79NVnG1JbAk3BzDJPgM0XbL6hA9Ty
vng6AdQk/FnCKzZcKR/cK1AnSbm06q15YiFYeQLvff/9nn2F2MDqyguT2xxyl+sUZ6RZHpfFTFWK
gtyE02gcqm/hp3tNmIbCLjA/8xzTgHCOQkDPYMth4HcIa3EwDhH3zUlatnZmoHgWdCHHqYaPkg4S
3H1p0VtkSRUvtLcQdSYsNdcCpsUvqdIFRhCh13r78wEU+jTJpghLzD3FpiZ1zulRQjmwdtkLHzur
dFDL6bQnJeTEJ0X9awIANa1HBwa5NnDKGqNCxN2fB4IrYQVaNifuROIY2ZS/EZoAxi+cXDRdnphp
+ULk1q6AV+zK1n6WR7mSQccQbJTDchJ18Bpd5MfB16S6bK9lzmH02gb8B8a2hput5zfH10eASmqF
Zdbkn8no36H3CEC/kYZY8k7pM9vl0o4tvzwh0U/15Oe3RkKCjW3dEZS8n1HKT28zE2KI1VamIor8
tzSy8sgHH38lXvQ/PKIihnn3UbWdnzNmGXBlsL11F2Omh8o5KEug2wo41/UMjntGi67FELjbWHgX
Dh4FEhLljjwfgzpVtqhIzFwung9SZNFA3xr4l5yk4387be2F444PSIXzW3kO4+Ws+WKIxMUwZ80k
gbCV2IeCTHTPJDSKx//2VGzAS2WWU9zYJDShARdgSs5dfVQ44zFfsnOpEOULSm/lz4tOIpTErLRz
xv+RCa8zfeXh3+6IDzPNGDScIG5V1ULoejToMizmRDcGZW8hj0sQgTa2kOsyPgw49rKi3IlI+Yt+
y2dnHjP59zahrulAZyDrlXC3ACXqn7pbIcRRlpvnb4hyZK+rE7yXO4W7rtf9I2/vwxPj+gIke9mJ
l8qza/M828rfmDeus6ikMVV46Ch9h9S8398qG5tN92b8BpddPhujXXX/9OUe8QNVyiU2DYZZd1cg
d1zFlm5oG8zFVykXE2AeYjeoQ3bs/45wvo8iPA/QoQcLlXBxUrxvk1LpoTDpedZYT5dwB7KZdoqr
WIExNaZrgrc8y2ynPE4G1EvdrorBxfeYZ6sMhMA1deM/nAmWF23aLZqO6JTQte/LUJ3G26ZkiBI4
RSN4nlqwEQA9GBtYYkjdzG/1mDmnx6QR9dmX4c6xpj/e6XYUWR/hvSxOqJUQWLe/iWOaeXALhecL
2wd5jsZdsqic/toCF43p1FAzLxW8emwpwnxUgkLx9HXhwUlIH/fH2wcUeaEMvCJq+xVMEq6nVny4
EHYKvBS/Irz2m7YKHwyp0kIqJJiotHsEGh/yuUsMBl79o2dSdKAEXgdxsFq9OCqgAt+AFcJ/TMLe
em0w8U6+8CszWbM31ZB8pabgcXBkFrdy37YGvZWBPoMYSmGPTB/IfLBWiH5E6ddmVgYGNyHhrXqZ
aludDbFFe5p79Xm5gH+ANpGd4PDhNT1mnO0kBjugCQxfXVIWcq5qEHsY8gzpbIxN0JUdGqWHRQWF
sVyLpsDi7yVbFIX1pEXxQheDMBja12FXnl8jFP+K1f3DLU3BwV65rLzaC1cc0+/X7souml1bDKU0
+dyjuzca7Ben306PzONDA0exGEzkt2KGSOX7abPZVOS/zqzzGS+ZWSEBF8bgoZLNQ1LdcXRRjWRM
yxdR1asxT5bYzGY0E6bNqPHzSYcl7KUMo/lG4DLao+LP3DB9yVr4FKfmLvWw1AmiN+U8Hw1nVWZq
2D7DGN2NA8qWtf0hArbbMCJRZ+7TejAFUtGCdAiV7giTLnwEU4IW97OHeXtPMGImnHg9WZSqvRy0
LPv1st7mNIlcjqdrgusJVKzQPU5MuzUf2yoROL9I8eH+/ICM1N6T+ebVKVA4z+hSHag0SuUqwmrC
P3NhB9KIpAIk78oF0J4cweDrqzc2iOy8GmIALiTB1sdHUG8nMkG8mwAhv7ItkWcF3/7+9qIltqNs
0Q5UwJfLng86/cSZn7Sf6li4aPkprdfpjmbfO8iZ9zNI2We1iwLzmsVZMRFsS0ToAxXQnHl5ftNO
ooJFdpauzXZJONyFWWj0g04MWZrhCGLRfsjuTSF5NqsUhWTchKYHERinUXmkx8fg8MAmYSHVbSCl
pD6Mjiq/NHA+mIKGBfwsJjc7wZ4X02L5/KEjuBlclNyNUwQF/x9KGWgNnTjm0+8JYO9IGoLsExBq
n2ZjZB17S9sFj6PMoKzgr2xeFxT94vBZLF2gUghdfDbhERr4ofqbFbBCH6NxKDFysoKNmWjdaqHo
ehH856pi9uqr7mE2sYP1VhPfDfb9/PKwY5B1cFySruCNEKdp1H5UGHOG+S/CZjF5l4smQoUZIFgs
LcFARXWFkxV5dGe5tED6i4PLOg0FcBSHLRtHSVurOXC5u8zNeFg0ThXRVTZSGtKtrUIzwGNE+PVg
F3moLzHgl8kpe8PFXDqFWGJppcffGwW95tLR8bK0GKMxHW44qWkjabU55BYe2NIU+ZDwLwKVdCne
iZmyVNJQ+u18JIgaVx6ZgRTZSeD3vtsTS/k/bel8elUWm4TgqNy4i4yr7jCtMqXcwSYKke9oE+R3
DZdcz99tniyfn179CTT5jw2ORZ7M5Kvnqez0MVy/LN7XgaUwmsVSisNI5L+OUYsxCcNTqP14F2lN
Uir/I2O51pPiGym/M8BkhKakBHAxZV3e9dhFhmMaUPXKBZfZpnequPGn6XvPef5Ro1DbIKAAB+Sq
ZYvkDEwkugiotFpJcordWiKRb01oggvbO3p2L91vES+73wdIlaDih4t0x+qyHxMzk6SJc7A1qi84
6s2YWo18VE3lTx4mCtQASg+lj2DvczNpJ3W3t3umfxgi1JCLyKROmfQxzOcXaXcRon+aWo+qO3oU
VzHXw+r8z6cahr6525mZDxqYT5lwp8NOj+Ame+xmZ899HR6aEzhwfhSi5twN0u54oOd1onW4DFmg
R9nfEewX3MspuhlcPeBFEJOeRNWjtBpeqXdXNCD1iRHN4gjp+QU6QGrOIVbRox0Rk9qji3Y7hdV1
XiGEcsqnyadaBylEhUxA++anU8rlvMrhlfhKdgtGdhGKZOUlPCZvEYOeJbJIHpPKeBXCz7PJrlPP
C7/p/7Tg13+mZswW/gu7O7HKi5qrZKB0Br+GBXZaVO5VlITDY1UKQVmO60gnV9hq7D25+4WQfv+O
HCX2RkZfvZDoVIdXXEnwevFkvrrWEdVE9xgtfRsnEe+rmNmwZ3I0VyhviPIJDMD2QIPzvI/hxS5z
bciAFjIrTdXmAmOhpDsPBPRISgNdj/nPks1eisacp91eLW3x2ORaa6x4ZCTrpdDhNBvOXb7rV9oi
M5NcCNVz6TGXDybjZxyPhsXLfdWVvDOmh9M7YGZCunYerqoFMhZFTMqtrTqg3XeeNGqMX4V45TDi
RcADHocNy75pj9lOdN6QsJUS9okEkgDLCtWKXkaaR0eE5QmPHgHyKILU951kDu7qaaitUARBrju8
10XZ9hlbSUWeXyT2iiuEN7bcu0vSD5+4mkqy4nNyql2XOlpFbUTIrEivZ+tlbGKQniNZDfFn32VM
ps2DIEt6R0Hj8K0rPU4wRX07k+lX6x+ms+K1+f8dIUGoU8J+Ry0SM937u4z2185ouF92w/I0jd87
ilcXyYIL0lNqYXoFr4A1HnKHOblNjK5H9VM84sTuoRux/XfBk3XDbteK9pP3LURyDWG21q+0Rv+Y
W+1WTYaoKoB5JpuuECHTlZgNO9SrtJ4LATZPcFn7kL5fWeF4L8WvVIJOmeydRD4/IGq4pXssBOjx
YWZCWee/dAsxCmGuajd/chS/Dd8IpM33t0fuFbzD0W1US6CgxVRGh7VQF49wk4MzB2V1wR9DdLxB
D4/T4PvVGnsoB1WMlam9ilpf/HUwZQlOTmxL0GcQNplw8x9YhdP+1j/oeqhrt4vrNbE8sbzplYVw
3PC9Qtl71GEb9oDoz4zjsA7RP1lyzL7acRqrqW7PCi5pmCoOD5Eg8QkoWddfnUZbOYO0tg7czOuv
T/HmvEHuUK8z/BriVFW+suqwJJHpv7MwvZf8/4F79LrIkpyqYGqB6o6J07f5m7kJoe2vadSty2W+
KmMlm95vklEZSD7/Kwt2pHGxOR2+OZwz/ztymqoDUwdsNXJAARy+9lZgwc7fYO0UbO8gk5QtTFFS
YKOy/U3hbV4aHgCv4XMQ3tI/cVN3h7dw8WgxPQFN0rkOoakRS0rw1XqxsgF0EbCjJd7i7xzuh9Oq
9aM+/dlvC7E69ImaDM22TGAWA/tECxQY075h9dH1AgkXwrFUhbvvAR8dDxAFSTSVpidnmhfBhdw9
yF8+sNsYfqHXyl/UYW0jUzyFg3sPgKL1OYTF75LUUw7GXIJ6ytB0rzeXLw1nkYWOAL+aiT7CMsPy
uyeRHZ5evbRkjRhTnmKBLOt9/oKHrke0wByj2POAeeNUEWpCIdiYx+7nQYL8GJnu1tnATKi1cVDr
v0B3W7KTQro6Uq9QI+8cF+PajzPl5R/oDGfoPrmTs68+2OUtpcm/Kl67/ZRS9Ahj+cPzqdrtos/5
CEYp3Wr6lYnw8C4NoldVBLifR4OB+1fxn63fY6kz/A5EmTYYCUez1zqPzBZfphagyFL5Ch4plAzW
e1MaCeranqtcChdumY16T7mQ2WyjFTA8SmdoTX09yscreUdIw9/pHwI2pgr1fzUAbm8NcZW5tJOt
MZgTW7a5DUGtkE/NDz2V/yOr57yGw4YtM4zn9ZGWktVqe9AwWAJK3attGY96uhG9jNKwGW0y3fZr
auDSfhfvdW7Mujrq4lC2pGD/DOaA9xA/ljS+q2GCDKL9yvW2g7FohM92VmyQArWUGRd44RZRhBys
a8K851VSPY3wHrB5qZIGDmzbgr89bnJEBypkkOWrq4juz/EpVmw3aVVx8qxZPj3VNWKKTlyaVlpd
/VTPSR5nZjNp4EMZ5Xdhyio7ANjQ0F1FTfkgcxhkhHReagmgbr8oyw9zDaqLQqxIInBHQ+Ugio28
jzlZLWqIbDDn796RPW1yoT7iA4epGSBNK6I2de1bRfsbpiE0WZQlgS4ApN2vBLeUFKuuxFj/Rmkt
5CpXCEyxaswlk4NK1R7FWjfdRgm9QSddxk1x3Tz6ey0fvBeTmhJerQ7YMMjWii8UiUBV+REwpcx+
VnmJpbu6q25Dq25eOCjNiLi1f64PLhVgvJH+9Y9yr46qKvFiuG8EbpRfnX2OGftXEhJ4FYS7OF9P
nPsw6fvvupkv3d+sBSvCsUf6Ynw/HSHkrrzPoEqeQaRk0gySXH+W9qYZMFwSQWrbTLJ8CeMP3jl2
cX6VdBvw8fFweoukXTqGeGWv3XrX0U+rr661hwrql8vZqfY/Rwmc7OCa03VtnJCi1qZYg7OndUiS
YI8RaEgXvVMU0fpG6haff5hlslUNnWpsthnxBsz95xxFIO04gtkqEMQgbq3oVEkBOgpB1oTilAdo
t3vdg2U6/MZDkPVYE9LOUW8fOLYZJs/TRPKm08CGxj43SYNb/wmCMJ4PC3+TCAj1LoHHcU4lZEWR
YKXfXikWpbLNsIazpVKeKWjKzXMItZlio/V8FIfeC03hFxlmmSEZMySYFjgBAmnfgwETNVE47QGc
rK0Q30SvZZ0iKHQvy88qqkF9DnmBTM5m8yZb9Tgtqsx8f+xdcdm7GGxgoSYD4b5R+qUrR56lXDKz
kON6ZLXFhZVWyWqjPz7TiIvS/QqnkBKfC1p63o8Y1oEjafhZbOhZYsYNoIsxNHqN5f9byIY2FDwF
9B730FRqkWICfoXgbTQ1rzl5XYI2XjG+8FDgyLuAUz32tZE8zkWPZspq7Ko/uS6dmHkofi/m3136
V3u9vOx5YabSIPIhV5N7JKWsUZEMrm/G7qWZN1ZI0UryLEB3++G8h5sb8DwaOnnr99d/i9J04Lri
qvhxxYVmqdqE0wngHJrB3WiAKaK1AqiJ2j/aGhN6XVnaipPzB5u8NL1mTqE28ocAkGlO+wuJlmm4
WdbFDxcSxHnPpzJTlvKA1Y8lmNlFM7t9CLMiE5Sjf7xHNVeHUQgSfkXY16ZbVDubmoxg3T/IM7gr
bg6/p3S/lj0xMcG8bKQmNPZgo/xEE9pw/5VnsMH68nuevzDw0mznAqDX1Z2HX+FeT5tdiyATn3rH
f1HM31JaY2OX1Uob4m8Dn04SIVzInVjRiz6zfZc+8z/wXux6g7pL0qI5HzZTXOUEi2yRS3B/lEit
4LQo/E+lxr6h6YdFT4MArWt9blOYnFttQLK5kBWzwRU8599MUWtAOAgPpr4skjbKrg3djJUYltZC
L0Wt9yWag2ZphHfnA0oCB+6axdmMKEgbbLQeJ/ucQURDmVSFdbjk7XuA2FheVajO3W7qLCP9Xcqd
qXDECwSsRT/mWYdjdE8O65ZYNXMSV/A5MySs6s0Yr9t3uw4eEcRCVLhJe7cTF/aTk4JhxvHQnR+w
SMqNtZ7Sz+l/6XNTjoV7A+ShrWcpSE6O3IK97EBE7A1+5SczAwb7bepMKmGgWIXVWz6QgCgWMBdJ
l4JDYeXbcHFicEiQMjjxgO3Q0qI+MIQfMF7wsNzwZaRawIjNpXM5O9DUIJMDZAvO5sK0nUtFtUX2
6hIZMwvb6Y5/ir8u973NrQ2oPid1amJAvNZpSWovDpG8NrLqH3R3ZBav/HYZwxhqUs0Y91KAze9d
W0DZ57TS+8jrUna31VFxmJ/b/ui3o6ay+jKFxZW7APJr99ZMoknDMcNQNKng/aKk2/qWNGkL7NBw
lDvD/H55taquYJvDNoRftxP6M3531mEb+4+2CWBT6YfOsqhL0rZxSl7K3gALVJEP8G61PGIjS7Y3
dpAb4e++FR72pC4sMk3+IOG8qXqGDEfSe8eVhErGUEWRNaJR7B+1dcTu7N1c8M5K/iLF8lRcumj2
jLETbMlaAbgAuTmBaaBm04urw/5X5cGIywxI2hn9TeHExT/lZCuZqyAqLdz7kv7PDtP+Svtx8Tpf
D5s4yxZGAhE7ipkcI2RNEMUUdJSonSP4f2AuzL71FJ34E9j3xOCfk7SlrsvjFXIFYbn4F0s++QQD
iEk800MoMa+9VIgMYZn9+7+b2Ewu+rMJyeuAQiDdaGVI4PiZnst4QMktouS+pxrVe/zZGButzEsx
5/zesAV4NWV1LqtBt9juKKpIr3MuqTNb429dJDzfJdD41gfNfHooidTUgaViK5kPw+/2iQXnvrVJ
OO2wkjo58ZEzyE91Vo6bWzFCrw22Al15S5doSFtNI0zaB7ieECm0Lt2B9iYUolFS0PdOx60zkJgP
CJAtBF6X1KpSqSX+UU4Cv6LIiHg3QAi3v5hbO9BQ70CVCluwmssoaaJeNsoA5EbSuzq8EXrAXFqy
/74dAA3hZBvVPubeNKTw5kHHhswC3imEf3J6k/itMkXrrzqTh8CdVnEcDHigx+cE+vsssLhg+ihK
rS/kuiNUGifLWEHv9zxebYHQqDzqn7H4QQzeGwiCWwrUeftdeuvnsOugoNbf/JFTK8WBlfsP2cT3
U4iq18NgeMjDtOEN0HQgkxWxpSbR96rRfSiUQehr7gUW2QVSuTxVONLvNJRQiHPpmFj9C4kr2t3l
9I3SWD5SeOj26CWGlaQH9aQXBh6LIsL1Oo/DaDK6+3Z820FwnT8POIHUvmXy8hgrmRoVwT3nRXFL
9yzzviNYGrbMr+8KB/nrippk2fhBcHpfjKySJuPE8LVlbdOEjOWASr4R6smFozrxYRXec+g8INre
2DOWuCOj94Y/vQ+CMLuni3LpermQ14B5spm95do1bbQ6fxT+UPuxzGr3A3kzC5B0IQcVAbfYTXEX
4j+dwWoU5u7wvx+U7/dzxkII/9ZL2dIKkookndNNzk2gDpQ9jPp9RidG5DP5D5IhgCy6FfZSMIOQ
V+1bPQhdTLMLLkOimVGQtryw2c4IBqnQTb8Dc6HiuHakJLzZEFtCwZ1oWzayHrgfhAAvADM0QP1q
0kaBopH/oMWZQkuS00+t2Gdchvp7cn4x7GivrRHkK3lqlXEN8xtbYJvol0a7Hv/r8dwLpWfxoU3A
L66+OofGzwVuxUNgw9zPdhv/vacG3XYwf5henOxo4qLQxIfhH1YjoG2Ws+1rTcaMePNHme+5SNk8
f1JgK/wLLV+2qj32OxDTEsqlDyFzT102TGBYSM7I/54Xu6A0vghpZ2v5tFlhgqX5b730WkseK7+N
1mhQVcA11A9dWZBTBGGL0HxfdTLq+CacbPYqoP2QSXkgJYMKZH0CRlSMpinfTf2lPzoi0lHzZ6TU
TIwTkoof34+Wl89eNsLWHuj1Vzg+CjNsa1uocy36FZyHFF+7Ia+KV/PTdjDz4AtiXKBZmueJJbZA
S+Q/C+l4NrcV4gNeJLSFF0QX7+k/f6fXCtZopDcr9zVm5r5ACC0oXMA+97YZQ9N/LTL0h/q/QhZZ
zjO9hjRqhJ5ohBoynWtwKNyzpF6iJcxuwbJoFu4sGP3Uwq3vaCRTEC2NlqLDzoHjl+LjAn8OyCsx
X+4EIM6Htlbwc6LAAeNvi89ZSK4taHkWXFSSMi96j2ch67arosMws9P1qvw02310BZSlPRRr7bDB
ioZH1EpWIzzVwpve+qtJkIk65jrIwInxb7Qz/Gema15+4aNtYY744/uBu8NPxRbZ7jBE4GqW0/kl
g224m8W7+gcOqcd3/n6k7L991IRQ/Ro0wkYC+GvEiBOxjES9gNxbdWD+SKb4ZHOgfFtVMnW1vbMN
vDTmCVrKS0wwMk6V65EXf9HqJMGohWHbDVGP3S93BU+08DkKo0iTjdnvdQb5zbhz77j4Jv4/1Yme
ZqZuDUa1cghdoTfiN15xGQczHf5IaPRcFeeOCUWUuyniB8u34XTDRhP+Wpjv1XqXe6Iw3K+dIQ8+
+feoTKeQLGUVsEJey5n1LMQSB7gCqpusLu9WkjECtglYKRwh0OhiX/nY0EHZhtoBHq9qBOapZiTe
bal9IMKSEbCqV1QER7g160xd2nSL5eM3/QVIDvDo+d6tAdWhBnPwX8ZJ/JN1AnOz2LTFTX0MX3Ht
BxkS5FB9W138zB3tlX1l/P9zKIUfYM6HV743YtmDcqJxbUV11LsVgHeCmSzE+xgJQJ6pqlmn4cTM
J0TLIsMDjrFr7qUk+nvf2h/1iKdcnVUyCKSkGjk90tu4cYgOOBi7Ui/9vW5SGESXAlx4yxn3V2Nx
r8wJ8tKpwsNb2ChxeCAYDBAayadwIn8gAL5kj1ATqspuo62IcJcpy7X+kwxTkj8VgsiwJptARbGN
0FgqtmMez7bzMDX+LCkEQolMOiA6+uAsBmwZx17HIIgKCtH7S7zkp/PpiaMTJ2RXeumJtcQgwsfM
XRarqBzgncmY+J/HGGetPPNCvxS1MJnb3LpDeHsbwF5N8nJT4s86EOo+sHAn81//OsKJlTQjzj6c
vpsEBXklzdwKhzIP45T0b7LdNmqegxi+TlvO/Hx1L0XL/XOCFDHXRyp2X7Moga0E+Yjvfy46usl/
Mz3qkjw1t3wJosEfIMyYbTAiUafM8KpnEuYgl69cm0LRo6taUhr6Y9OLVEJnwV/VfOjmYabwgTw1
Mbugr/+yXjv75CnWYu3kHoevpDw5CVI8uPuojosMsDzyhSuzDehXK3fiIbjzHlW7hKohzUuk6gJy
PlIFylqHnPGhre82zCiO+h0DyiYre+Gp+F/HJn/FtGkoCF3o7JtYbm+7MDCIUFiHjwwGoTptzSg3
sfNRg/YVdj8Q318/35oNm6CA3CUaSc8oTjNyoPtl4COKuB5mgr1m/xYbTrZKgRBilnHGQ2ZBwWip
20AQKlDoSOu6oxjakHRKMxCssAVBFwAMl2jWMIzFVrf3Uo7ix6fIVvkPqRA4ab6H/sX8Jb3z6IYY
ekgz4381Fnu5nvdJ8MdG5vEIy+kFQ78zGJiuwrn8gvkf2sbrpgM/zls7f4zCv+109rR5vgCnQD5z
4CmS+Me7qebuo73Nk6CSdjIsmrfsSqDP6rSWbTSBgLwMo+fPZHEOin+Dg7IosFNBqhjihSAW9Sm/
/XIirmu5EODua4qJn2DoKjf2m4jSjdR4+wHk23PVKlXph99q+cG7YZ8siN41WzP3E8qE8+CERoaT
npu51TALgjM8U6vzeh7MGC+/4ErsMX+jd+onFrDeBfG8a9H+rkY8Srakpn6H+s7T7u0u7NU1IuIw
CF2OYAVyqvCVc2upWJHhwwDZhColFw0qKKGWlYxONnFn9jTkkl7oJrgP1lRcUw/+LrC/dXydLcsF
t60l2sYlQ3s9UvkuiIOAGupxlJ5oTFQQO6k9+QkAFvZdCJlaCercNrwUpmZsuxz+Q8Al70QLBTo2
JYyF2HJ+UspQTC4mK0e6VGQzR6PAQxagIX9DqagJYcWWeTUujo8ZaVi3+J97O07/oPcL1tVayK/E
sTC6vhA+iFz2XYk/nfX3Bkfrv0aesLCgnQb6PfvmYwJJG6QbcZe0MMUCLurETL0XXfGBZ6Rlo0yZ
gAdSPUQ6ThKfGw4caesRzPkyl2Xqc0pFpRV+99H1lpiiwDQvw96mqiA9u5YI20xXObSBdbavvEGl
1sd/DrCTyVtvknRA1WIAmu91csDOQcIVVMo6WJoTEehqP8WfdOXhsSosgHvxdvsqCDNCvMu5Wqm6
0ELbvA3ewby8xILIPV269XREw9dHrJmCGD48X7JAkF21L1YYBkqi1DhiOUnU8hTFPQFimCYazqwn
9AtJAIa2G6rqLtXMUhzmAvvMT62sLgRko0uuDjlXSWnZYwuqq/o/MsLirv0WWfBfeceSbhy/9DYP
1Q93LRqCfbBh+8CEnGIBRJHfDAqIQQVq72IY6C7m+dwnDMs7x0ydir9mL0R/e/ks9Jxdj1DEKQx6
FyU2ByiWezii2+It+t7xwGeX7wxNWWEYMGN3EBzbj2ayD0QstBp4B4OCPWzpEjlJAdeU5sPcf6Ql
N+JmARiVetR5a8qp3tf+MURYLbBFIanFVSZc97DFNoOhphtNesc9UvbuFH/vLdGdPwdTzQhPFK17
yic0GWZZR1712OplSEWTYvwraDvFpKIh7/YqvptwKIsf/ybQ5hBoQBCZi0JipdF/yvzZM4qN/UW8
il/W6Gx2o47L8uXSA8Pl9Bv1Vtd/e84iHiKGB868bJFyuTgF5s4ggmIxdC4moi0UyHfHB2tNuPnV
x6ZgkLJahqgfogXJf3VsP5qFRVfxQDe/wgTMBeZuSD4hQJXc8mh+ZxmqMHlG60F/wIVTQpqhWh1L
6hOEtvlc1r2/Yu0gi2cyEM/ipzky11O8ct5kkrP20AivNaWR8BiuOL+3t8p2h89hbvRiEBoWbM1K
GpsaOcLNCLadVXYXwZg+ueNaipZOyjI2Ff+JdYBG13q/66ytWHrdcURba9sav0rMqpJb58dwc8gn
2vK4lYARIuHUoxLruq19v5T+AXBHWNYI//PsE+UqajnDtMGIdHXPoVC3cep3MWIRUzzwhinUdvf0
TocPhqdKZn3xvl84mUByxf31z4lVCguCxatsuZf/3mxJ0Ljsa4gv+CI02g8AdUM+YrLiwpKf6Wnv
GZ/Ng4yIYRKm9Vc3Wyk/Z1/WLCaQqXG9LzaU44Oxf2Up7YiZ/vdPoa0/erY4UY09XaZun9cI0ELJ
14HyZlx7GWpaxVNahbtAKebjvahBaP/2tIg0XGie4jvX4noLQqGjXoYfcl3j7yibu6wWvJIZiuN3
G/lP6Ne8f+FVxfgo8Q+2rPzTa87Rrk8EhX3NXNhkfQj9hVfB1cHoN5D5QaPscKtcNQcLDaufhz6Y
1MLtmb+Mj29vjfG5tAucDBuSbogKcyIrccglser+6bLx5DADmLZkXXly3aikw11h2cdmfTDi+4PK
6fWeQNODVdDc/m7nhPTOY5VmqXfRch0XRVMbigThPym41odYLu98iTqDnUgjyQLuSXoe4QFBDdyx
ZBLVFKCxqSTxOgag/a4j2rMaTndr2u163Eiox/jpLpM9WoG8xoD3SrlggO8KrRv4ROWVt6mbpYNI
wQC7Y6DVi+1U+8Lv0LA4SpmgAGHhXLu9sGwLBGOVSyoGBVVVtq2fCEFj2ytT14jdMRhqYf9EpvKk
ObeQXz1cw3RK7OL0xAEdmvQhYwAVMzu7/1LME3a4AZ1cw0pWdjW5OmfG3mqEz50Yp5wMfEC5OIyD
30FXQoDHLX/a6mEm49EprruCEZW2AObEaqQ87PRYJ8oLtFmHFaUj1l7D1M2uk5RVX6sZBK5hssYw
Q2uruD1brefoti94OswUoGIGZCmNUXFSi64p81p2FUxeokF4VS0eqXWIWLYtZplg+RuCtFEL2RDH
9Tjx1zwoQsj4t9ZYfkvYzZlbqJ8kUjeYAUqMwv3poQkwD2/1Fo2cjZqf1ZB3K/nXLfFciawHwuBn
mzzB/+UipENYBiKWgHaRdSq2enbDgwxmQiIQ99S3w61bSdbHoeWG/ImqxVYslkMQTKeeYb+GygN3
L+Mc/+XgM6Cw6R+WE2cUlDHoMuTNiOBgh3rzULK6fnxguxxIDuOBCYC/QZhgOht+CDgcMwPlkPBS
2yGDd4fBf9AZHbYlrLdAh5CwvU/xf510XCOk6r5DZzGWZzitmssqzzkTSaKjgT4q2JK33HAXabmG
lA7LXwL8l+KlaFEQ8DlMeBaa/lh1PmcUdjVi0cfNRDqqerwvrlE6Yrf47+gRCidsOem+uScTrGsQ
j7ZzMUlf5pyb+vSSUOhMiQgz+raY81Y04j3cvW3JYTvkXWNC86N7ihVzrosWFWQlxSLY4SZX/vhf
AMEMPwwtCJn3d3IkS99R+U4V1niiq5d90WXqaQdlebBJfb3WEonSDiZxGAuMgLFaRl4H4ruBPDiF
fWZOX8NOpxpccLStJSlZ0WuQpeoIekA3NjjZ58HpvddQsClQhpGId70Sy1ePcwKUgJ3ROznAK50Y
++ByUj27jdct2KgvRFwifI9gbBepKl3xYIeybZdN9N0ULU1zzUqMk9ahWHLNtskLGqtyqsqSaR7T
FFLqDRkdaBxynU0vSKPQ1aouug2gAyB9yPJcKTQhc0GKhO07i47ylF2OT9Tmtoh8ExkvaMqShjbj
uS53nh8yT+WCnfwHc6wymn6cB5Xa4lb8GxN34mTQmnyr6aXJ0+PGMO8OkbpHLCEJmJdeCifrgnnl
9xHBm2U7fMJ1KayfrEwnek/bq1HWUz4ERjxFfRzYe5GAmRjIjvH8zS7cgCWP/EfzzhGVGgrUx4eU
QyAKodPQ2smbu1Xx4PJDpal7xHzM3MiFeQ95ujQfB4GKm9AzAAfAxOmB5lZsjGUkEpyqUgf8/Jvh
KjyiLkT49doCbvNjWF+e3MWX7GSqOn10Lp1agxqfEXRVZZ3QrgIXaGjJJt6Z7p0tOhSweqBZIWGl
xigjZC6wweos7NCCdlKB9rSU4h9URpbMEOy54jl1MnxK5BNtE0vJKU4I/Eau+Qja4+KDddB7Z3ao
Vg/DJJ2o1Y2a5g4hSnLkJqG9nDb7y7B5pdYAgoG447rV2puPrY2q0ygjwykQAkISQoJMbLcwh00W
sMeNSzP4DrBNSc32Uek8W5C1sOCdd+n6x47KLGXYPyf0MfRZX11u6BbPgwF/qrwOChEKtQsZjokt
d0BL2ilnYCPBdkyFJTRYTbNCwxikPjkCAPrB1h3uXLD8uqofwS1GDnnib9G+NKcSeo/6j0YIqQZw
YDzou2LxsMPpFJN0WWDNW1ea1zlKXd+VNwrXwQ840thHC7oBYPKRDHnGTcXCJrsb5vroQDJZtUqd
ULAfAxXqvurOj8Y0hIJRZFGniRoSp6/mHRYj1YfTb5QcZWCusqAn01kTNyXxnEN4HrFovT9Ro5Gq
+I88Mg4bPeWni2V6/lZfyGGNT6Tzsy7MUA0WxPxBXoknjQhppkWlMJbXx5IKFHbLRKVfJwj0bL2h
DzXJW/TTJZy+0Zx1V06NK/YSgCCd+cac+sxyWDQ62qJn0sJBvIWvU67cZ0E7F5j1dGZTrrzpzqpJ
MWYco6cgmCjIQ9JRSZBxpF5Zm/d2G3g2WiTHy2pozpKSYWtyH1U6zEcifL8+8XosSVYb52HwzChH
+1U0sELGZ0W80obujg5obH6tZLOYljCKoLS+bDB3QQunS9xsZv4PxJrYYNGQGfDbCMN1LQAbiQIF
TTt49qdh1JlMwsxM8clEo/+Ug4+sPYEUBez2HMC/Sv7HaNx7Gvmq6kq6YE0iYHijZ7sGlcXPHNx2
s0BpgVI3xJdJv8YP7O1H7XwzHLb2PiAKwatPzalU6tu79vrLQSqFVJXvEPX0JkL3mgt78IYCsaAw
6akIFvMmJ2/0m49ePmN2Y0QIVmy/078gLE3x4PDqa4t0ijxI+tQh9lBpjRvx3kQuhjog8/jnnfSX
RRBxvl2T58v2Iobntgdp03A3v1KdBjhciT+BQ8wKzUCcz57Jk6QJwxYxSlvrIUCRCVtyenn1roSn
JUNKGjIMdYnea7TP8+IUpNDPUyp4aMqknPbq2OyYhWatW043DH++Zh667woBgx44SfwG2wUVvvUN
bo2YsyZshp+z0OppVX1AyI2uIQnrGKzk48rBpf4VYnAxV0rcRjhp7zzNAmtai/c7f4ijjptpl2Hz
X/RspC8kmrX5HbVDOfi0TGD0nVK+ZOrhRWVapux/s2AyHCQzWla2TFLDwD9ToqruH6RKsAEwTiZt
xnzVVdezvaPi56BRQXgO6eiwaahbq66E6xQvEz5jEca/Wqv3iWNd5fe5b3YqABBmpWba7LRpA7A0
9YcV5++4wKAfVXgoT+yJQKW4HbWdoIINC9nqhF+GikVwFzbzeihTuAwEYWVNMzSnF8rzDNYk1tOG
SYNS6KQB3BNIj0GVt+8lRWsiK5IWa/qEA5VRjkY0yI3OVmT2u/oYOJyWgMO4y5118iLqlspDr1Kn
RPvpx8+DTMqzK/Y5Dabr2TrJUq9+/ukqr96oquldwKeZR8wb3c+ByP6S5YgkvPCMd62LNQZGBcL1
6bJNj/BLHmpuQ2xQUFtGUysD6bKYqcpJ19evPnL6W8NoIWTd7CuRPGhioIHwaQl47RkO+SLAwCKc
h8YvkWakACQ8po/nf8bxscI+6gIlSunhAiwLZyOAt44E7jraT34wJ2t8BjPiTM2eG8M3YxhDgBDf
T13Oinfoc/KtuG+brgKHJjBzhuPDgCdoYl596sX31WOaCIDAPckQKmmcPaemR4AwcD+y+gSSUa/F
dRsifxdkNg5ecjDDR4CWUBwdCxUH4yH6ALknvMnDzBaSBiZt+2CT8LkxWxQ1Pl5mgIQk6fVRm2//
7ZlBS0ytqEoUtzNvxXYZuKL8MgXDu1Gaw+iEwZ6AvBZm5eJXofI3cx+jpWxBYF1ThtmxXwmv2LPy
e1fStsXJB/Yzsh88G+b3Us1IEvHz7arVBdg09+nUMitIP1WBRC410ZQIKjYZcmTGITMLOhNcXVwy
IKWWypZrl25oJvto9OfRF0BrAW0Vm4/vZN0DBpyA6114PCWRjUMXvdw2ePk2FpCyvlDC44d2maYs
bDqfmwF/lwSVCcXdeVqXtOxmAUcMtp/bcPWY9eziNIFc+ZEka7afcR/yeGm4p0SyRMgO6ITPN7QP
J3c9Pm51ySP9a81nwTewm6buRUEx7/m9lyatwO5W9bgDn/PP1hTXwccSD1zK5eo1kp6OGHrTjE5W
X/BE1dvEQDFS8r6GBQd9Buj+hrxtFdeL/5RzjLuyme20BnPBKPYnBSzcXlJv87Ui/A2sUzKxWyov
V6bOhYLGn8EqBFR/ILwl3uD+JvUvRTJF2qOC5nmZfpJFTADbOpsit3/z6Opgporx9mvkifiF62rZ
IvP4/ucEc1aFswdTU8OeXBGQQGMw1k9yHEAioKscKR665M6aFjcavA/As+Y3I5esa2q4a/lA5sl2
g8Stqar/CPdsf5TR0vM7nZAt3cO+D5boJaca3KGoIZHatqFYgQeIgmqyc/fEePJR300DNe6IEzpO
XAuxSMn3xeQkVohsBqRcbhvAmrr7cdtxhkaYGdVhZkDtM++R9HpFx4wvNTyv9ky5OMj5ohSnZxOq
FE/nfGpoZAOFYm9y5mo5Q9G18nTJcDPc3Ho91Pb9k35JFmE/Oysu+d/EAeN4MOWYLmubImGbWqbz
avqYgBlUD32EBff6EiAbLiCQtuPasKw1fvUXaB7njGkODALJiyx2Dt+k669UFJQB6KqaqqXJnnkn
vHrLzKbGhJSGI0y0trCn2DOuuiwD6CTJQAtIOTh+qaPzR7CQrQrCwea44VRJQMSh3kWROUU0O7zw
vneejMk8bSY8m9xFx5cp9GWPlIV7Hj9uwpPHbyX1w21iX/qQKSWALjIbVoXe0Jlubb0RZVCGe/38
5MWH2YRWXrm9aqlwJrlBnMzgtSWw/uGpIB+Rpufm00JDinmvsIfPn5X6w3rXFi0+XBzFG/0z2NUI
oVYIx4yvmjmRnNVmEj9dXdpR7UQ94oHT+wOuBfD/1lKU4ktHxKmEb+6NiyksjEdAprUVnf8J5Hht
1y9QBQBkvQ5JZBogXkVJFmvvYPRyzw47VE3K/ijVIMdSTZNwINfXtEn83Wod6kIi3S/cNomY2WXc
FDwxI4XChEnkkiwcg0/3ZDKxNONnWu7KvO+a9bcXXtDX0/MTNwS8r6J24Uxwz2QUhFafv+JDugo+
8nA+uwzRyxDBIGdSAcL1AXJfeMdGUfx4JIF2iWHLT+DcGsHNkMK7GCOQzwK7YHYvdxbkx78bOVZQ
HgV/C+vI9vg7w8KKOJGSgB+AjJFseFNIRFVI+PGjI8H2xg8XEvWLXrpPJZfUUFxUZoL8iJrhP214
IQ2TnDqE5zwi19vbOT0kQYxtxxVyd3/x4ujg86JVZo9iPtma//EnNWonbEC3h2dZKKDitH7Isakd
AkONrwPRlGAHtEKcgEqGOo3PY/F8o83fIoScgSSQH8I6kTbabT/k4UJL80ZZuEtg0fYAkkVPJyhM
JJIfTN+ekyVBc00BTWz81+1bRhICGdwiZtmk4HupPYnP0sUPxjvVU0hHq2Kr1kUgMfBb5Ymzwq+A
Dmwhas3IHhU4PZMEi2/3PPY89ewm0I5zRP2+ZM35sJqVRlz5irqMaB3zJ36bU8gh+N8bvKzvPfMj
7w13dzpTcdnhZADYgIn/vLAEUIoGgBmaH50gbXFuBFeCuNVDdFVIQTE9DBmSozjh8ncY0QFiQF6v
Bk7XOQq+h/b2PxUbsCeIiAephvxcepPos/eeohrhhB++Od3SgoXMCnB5cUpvNlJr9JF1XPfojR9S
pmJ7R39RgwMk4CjeWZvZt/BdnDDREtX3bC5WYSvEVgw1eWyApfc966OM6LLMtgxRFIAY8/b+9aZ2
76rkUzGhKjkNl7H6v6YDGRLtldyeklw0n9OHe8cwlntDYO8Xmk+3Uue8NAttB+BQobDMXwNPoL0K
gcAZvign5c9wjBNg/oE9L1r7Zmoa7bFeZ8ZkPQ4MCNIcHrkly3X6oZArUoAGjd/Pk0tDApwT2I0z
478bkiAKzGrpwVArGBzgv9NrFHc32rwddGONh5hc+bgTMmYOYlPPmxFKHfjXjhC5lQSt+A3t5NMx
ujcNdVcDuWkHtsrsQxEj+4dHV+oC0Zq4DNhSB+5SXHc5EF1LnARgn9Hu8OI8VkyGSbZ2UU2k4cpq
pQn4eIR85mL2t/O+zS/znyg0FCZ9xs/0h0ZhIiVRhaQnF7it1ydKxugx8PPVu8Xr8akq1BFCe7rX
Wqzd0gah75qHvhLTIhAh23y5BdVBhN6bNa3Kq7PZNaZSQ0eTGwuuCWomFr00F5LGc3IxIsXpWyrv
XTRCyhCT9MpCN5buVRUn0F9wh6VRunIkhvoB+QuiFT3TDxEWaBNrc1jzX6R/qFr1ztCEeoIMi7xV
HJSSkyrNMkvnI3n3YWNPMbhHc8wZlCDGXPhV8pwLsfmFESg4eQnULypNacRHW6/30uUTwaZusYJo
s3vOMwd2ZnMyK4T+5DK3LFNIeJStz0RzDmc+6rhtvdfuKiTbSeZgFO9tWrfp0XWDsdtD6GUwiJcw
5KtVwdg9Nb38BB8ka9ILGnRRs8XJb1oIs+KO6XYYWYD2WPDLVnwC8ikWh424FdgfI52JlHPCuw55
n36H8qThIgD4jpPZdccVkWRb3r26JMDkAhO00kM54pJIssSFrYKNgB0Xh8+aP13CHkPedMRKh0kL
RY+qX1HZlMroZ65zJvbbSl6GiJ7nAWtZmEnstDXwsrq8/OiG62OktHMKibENqjY4Ec2cxLhhGUfI
Y9treBh3RxLrTVkA1oL9EhDbmvnmskJZVnYM6NJRpMJJW3dK7eHcuGarfmsIvEhbXToe53vkfdR3
4yeoGXa9zZozzOjVPFWKeiNwX/okjYZMRKFDWXyEhhnz3fedipZVv7wvMsNCaa5X25B/ZaTyRPPO
sd6HfEX/i8z5gr/8lhfG+ei5X+WTWzc64EaTm0PUHXILL6cnCKj6dCf7gHIozlpFgpynWSRjybMx
kXgQqCgcIimEK0pzjq7Cy5pgOXabz/zPmL6to0xFIDCte0D933e2hat45G8ivQGk+wUYF7VgH79q
Pz+xA2Pq9NHxg1oQwQMNcsM6YaJz7061SujnAO1+oLK4bspV6hxz6xxYiermDvI0virtAs80kc/a
CUw8u7xAuwo4nrzYyu1vQHdpOC8RR0/VtV26MYjoGPWDVO35XZxEG/sngfHz6NgLGjKwybho7l0i
nh1r7eeQhSWbUipqbP+wa9he5uSDxGs8ySauzdrp5mJ8VouTmDG3W2RtPkHrYqDEwqJF2NbBA0uz
AD0zzCfopGgsJf1F3kwLFwrUdiIuKvtYPyu9rcXN/xL2XCLHE6KRHNjJjIiylANgBi6DMAjHTmqG
kCxR+ofWjzi8ScXTE2ucpGrV5tl9yrCJlpudplrzp3zDv16kLteos+p5R2eoi8CDGDHko87MKffI
Bx2/bUfpjxju9r261SIC6iDC9jxvIsUWcAHPHXpTTnQTPzZYO6FO+DVzAK6cdbO0kFTuplTXPnjg
R/dUs4hM1a5eGzHVclx0AM5zNv74plYZWcx0YPwkaNUayPJS3CfFbMWafgDFHyYS6QyiXAiMmUaL
HoNAM2wAtcB9cEnV1lAy40ZS42/JIKnIbmgJSkbXDYOA8azCHlEHERT4qaBjrrh59uxvczHThWdu
s2dssvUwucsMgZbhmurglAgP+Pd4Zg367SoGZnKSFLOIxk7uwo/2ASlrq9jqOzR85EhjDFxvWfXJ
Y96owDGQ8evZWs5UwNPVL+8UjlonfJUoV+BiL4f7Z6HRXEGshtgQC9y29xMebhTi+wRrVIixTDIk
NxxduChbp5tofb8/cEInPjJdm5PcofUnKtEb4y2AZTKHXsp37MPQjaHtaVWx9ZAA/DO+L6Xcl747
S+M4E33Ev2AgEAlg77r0meFkL1t4hji+i9phNWL/6w7QsoR8n8DWYuMG/Zxqwk4fc0CaSXAvISnX
44veliSoHhU6CdBwDuWtHfUSCuX/na30ypVi8ZDxnAxAtAQ3k0sYEktjMfFeqjk+jo/K7CW8/2G4
muaH+2UzMKLSEtBtdHZSBjPy+pQORrs7DW3pso7GJo29Bi15Vyel/Kdw8Eg8JANWQgD0SVgyXTN/
HuNqYO7ivdA07v0ij2htw/vcqxTJXAmcadBm+vPPrOvIKtQ62FDkYOCqPDKjPeKGNUyfN/wjikYo
7xxwo9prTUOB5F7HCOdzdiPD2p0zljmWTA7TGiduzKDxRsmhAPFDf2coPFdSe/vmf6pqaEnfMduv
pphzvroOskkcSSyW5p84V+4/hW5/02azKxD6U0MOESeZJSbfT8VkdhEuEbcxYRyIGNbpypIu/Kw3
tCN0v6aUGUmy0DrTWSTreWf/yG0rIGHTt+KwMoSdeCvOxK6fe/i0ut2idtyYjc9DMpoMRAwLR6nv
rOQIh3lcRAjMtfFOLNu6gDKTrs7a59h3GqChAXt5UE9or7ejx1ABHf2lzRu045Ih8FhIB6OSiYU0
CFu/JGb6iRDi2wZ3FjZug531Zp5TXbbTqVn97Yxko4fqTKa1zCfTqrmobVKkt5waBK901Dpu17XQ
IDwhDMlUQ/mBPtDKyI85DZNoYMdK09quYH9aC3APvmgSV8uJV4XdoB4EDsVSGOSxXF2KJxv5s4pz
V1Jmi6K6paXPhRDik1EMCduH41IRBY6vGMOnebVfAfacFSsnbGbwKJRa0bMud1didegYh5LQqRve
WJd3XLYiJ/6QECTk7T0YXCmnWDsZBpQqftTTgy+PtueOqvw7b2y55eoLzBy0eic1ayEPhkesGV9c
flaJS7v18uDPSOOzkndXw70ERiEsAoa2teKKucM6DFPBSwX7KHwzpBIwa4/iU+Wvzw3YDcDnCsdI
tF+UWQOvDSJTjd6VRxrXTzCWuPm+ywRPEiYAGmkvN1D6DC6ci7RE1NSgarsP90lT+D/p1kN9gaGv
4hYDs7tp96OQNez53x95PbLZeViObLqg8mQZt5QUxa5SbWmNG1f88VAL2cif5Z0SDqDfCWqZnC3w
MQ4w/I+WT1/GoMqUKfOglXv5i/eUmKMRAgCvKUwSEbQTGfewLfEYmqZhXSuhwifE8rnNaBw4nc1U
S8NSJDc4gWbMdgMUtnTC0Q6lKKaeq/q4T+VTsNJZBwqUD75/M0AIZw7KTSVMCyxLXckyf106XBMe
M0FJe7A1SXph7ZUQLJLllc7ejQzgqxg44VrMaxxYklrTAvL1fLQ62PagFsWXXmQ1/NJNtoanb2Zs
s34G/aMU1z5znhyGfIh1eFiMCixLGruw4hdgc0CcqUx5ZyGPqkmGw+jJTweegwSsxBbx2zFifekX
/Ty7ZP7UJnmFdF0OF3ueqqVvzvq1o2zJPndjbaj9TjU8A7GxtcSHZNL1NTuN5AUzOyPTu2+Iu6Pl
xmZr1r6uvE/InI3B6Gy7y3Jo5dFdsT58/X6TW0H6JhqV7eiGYKsFsSH3F7omy706Bkju3lBRgAfW
izWFcjoHmBw8MM+i0Ly3SGo9p5xVBnlkd6jo4egB+MLkvx7WOB+G+IcLZ78wy9EctUwUL2sBOQp/
h6d99Iwf6KuOReJlFgx7DR49v6gehJV0wCagMpng0hItHiJlM7LYikjsoiZ+8d7oAhLwGLYwFA/j
dCk+Y1VmocJN+Nkk1MGKbDwhPhIXoOi96VkyzpLPiZSTLb/XiBQZxrOVnoQDtpF3bFhKY3OJYq0J
623NdCf3itPECd2rDutiBFnu3buuTYJo2VfcZWYSABQB082yCFokGxr3bYKCV3LdPAr+o8sBvJ3E
RF2DRl1RyLr5S7xOTCOOdLzOK0Qkv9tG1HhLE9goqV24TVxt4jAowMZXzfzg23HnSp7E26ZS1vC9
HmnRjp9DO18Pp7kg864DKtJln9FDt5UxvFo1x6ULkOluyV+71zI7Ee+3gbkdEs8SrC+vDrwOWEmh
x5l2iIT0JP1s+0TqP2LPU9SR5P2n9q+9hAPfD9HO8wRVjqPns6piCCmyTHLLlSu9Oa4hN64Z9hGV
JqjZph6lYNntFEkcfL1i0O5RjNymODd9C0PsY2MZVTzUtiF1ISYxyCJPaG0SKFeGlimQ3JJXWwNi
t6/nfbsCmerKblHJVWhznr3cPfQhYp2L0LC1xLyIwdxtlWidpeJEBWFQvXFSeP3q/NLFQrNSI8Ub
MQ8bRLAjDcuobJKYK+7CNxG1eVePDtygxvGzsAjYepj0k0McptEBA8DrjRtaPbsqmlAhq5iDuiRk
7QDsBZyMWczQUQ+C169wQ5JlKWfNtw3vMQVk4oY2l+Cnfg5U7mC9UBCt9MwxgGOQhidkrmeyVcls
Yb+Hlk1xCH7BlFmlUCn2y838yI0MuAcR1FxOn8wjjMx+sQQ4fsZgEze8bSHe9/HbQC0L5JEkqgme
abUMTvreiiZy2dSzzurQjvjZq3GlpZ8kkl7BL0QUilWJXfp4v6Q8nMUsgEHEu0ad5LqX9kF02FyP
fhnBto7IaRKRfG0a8X3Qb3gHTghGicIAsqMoRQMT8m1bP2HspbMfveGBjdHHI3ZaLaEPyrxfozWK
0kunuDiyu+zw+hEtix063LkEVMW7yuezSHXTNPxCwBJ2rfwzgk8mLpPEsbN6/C77qwLUGnlLxJvp
SHfmu8Wvyi5jJVNoDbY1+g3HgY0UaKLg4OqdVjoa21d8TKmVrpOXHSUhvnXe21tWO3Flan9d4H9c
gZx1dlLvivCiZa5uxIoXqqOFy7qaGbkU1udN2bRxXGiT0mP2UXiZossFNq8H28+f22yRjWaV05Ta
QnXo4qvVGc44Dm9ki4CrN+PJveelSkv9HoZtcDIT6Yp0YL0McVDdW8wsgcftCUTrfBF/IlnUKdas
W2Xv1szkAx0MuTUmwDHFX0T7oAwYVguq3iyJWME/faKrp8qF2Oi5eOmfJqoC+ciJcaYJsTphGw8j
AH1Sn5WoSE8gIdleS0oKx6i5LU54OUbTbp1VCXfPl1UJ2sMHPRjTW/WRW5UVdLvnHrebdO2uLCBL
Zo/feE3bQ2xohjWEusmVCUZMMzS1Qft1sMyEPxIiZATt80QH2C7OjXf+yGlFIDIcGWkXgol891lD
ZTisj5agZN1V2nj2gAtk3cLd0sGlOOALfY0B8dnf4l23Fo79lW3Uzm2QWDa4dXRhIwOiWs9578Sy
LXwKQKRRTdHVt/6IM+uov+fxNK/W1/IRUi2A/98YkqDvmz3uxYcfkK0R1ttkfl3C5QZwP3QcSJkd
ur89g79lslPYu7wdTG3cO9ZvI/NOsBJZKzbrBIOfnPJBZpZADOoZ3P5cYNADVe4LE1ByWTspt2S/
Eem6kpo4zLqcu+BZL42U9rc4RglxjEs/0UUH48Sc99QK0pY1SZijLh3Xde02lIFcsAjz3Ncg7A5I
hwV0XHXu8qUj4gfZgsMY2T06Zv8Kn2j6xFWkN7bkUaZ1XvyaWOEvM6M75AaXrT5fhpqzgBbkAKWT
ihMWIsfDSNvlcD1VmK4p6lJ5nRwMnsVZxbOWXpZUHrjJffwkGwMMSDpX2iTElvFRhiVP+SSLN/ae
uyEGdXP7VudoCV9p67hgA4yV5HMN3qRMP/qQiZFtE4oDIP+taP4bawOPPyPh+8d5mQmT/aRAVN/3
hG/JeZhxhof4sehZSjd+kmHh4m8AGxXW22GNcfZZ8/DQPuJhutl3Yi+ise0kvJIAmDAi4IMRpnSV
q2UJ29ZIXTE6aBEwC9qKKIGlEdZaYyyLBmoiDiJ5q14QT8E5wUw1IGfC3qH3MgPvUhblCyuYX+IH
ixmbuUGbV1lejhZ0txvZXf+13lUTOWEiRPtXtAc9O5Xx3EShwCUCX+fyC8BvZ+PH8cwnjmeTh1qD
ubpN0ThMiWWK9GAtmSsVVJ4eZt3R3rQwQ5EKtMpUjSKbn41L6rzUUIr/wL57BYzTClJiGyxgTU0o
XuyXIChvokm7HESwRN+z1NsIBqMULU84oeYnNF19fWPqBg2mW9/o2dltoDEglZ2hZ0PE8FgeLUPp
ApZYYAQUwlEW81pTbaaUpTVAHYWe5r3nzaRE2bguuNKfDGwTiNptbgUkShLrf++vX+Y5FqyteBfV
a4PII19jzJSR2NPtRsksqbRTstz+3NDgOE9gtGUci9eHOJfu7fY0etY1xzRrLggJyaeG4vI9vFrC
DWOG1iAk6+rGIKGze5MtGzcHb47Tz076QgX6umrp6GVny4Jauua6aSJY9+P0aZYjjcTTBRCFy9zr
jb/pzC8lYk6fzmpvTeoqB3Q3spFgn0AYI39FAdRTvCjfWPzi1m7LH29PDhIvjk9/OgpKGUjNgzy3
69F5R5u+qkh34dqjlrncyK0MNzGxne1IMa9Gy5zWhZ48sJoyfW8Sbuyhzz3iaJrJ/O6PJb0B9Q7b
Pz5RLo5UNFCrkdwfqOBLnUgJn/hk7Q4qwEx6IJn+3PfO7U1yZT3FPel6JCuBkN0lW3yObEpNd/5r
3B5BDWDdoOQ0cshWeVS3V70fyNU9GlW0Is/vphJdpDocBmoIMH5HOynNYYJN72Ri3q9uzB39OY/Q
UoI3AM2cGZwKbRW9tJa/CXxD2rrHXisXhaekeXRq3xaJ2wL5+skA+QOrxFQJBRozSZmSTsoZ6ED6
Ie9pPplg21SjRTsU9uRtynqIAziqnZyrbwQpYrPg5DdnCg0GQfCweI2r9T1q8BfmJDWRq83jyKTh
ApFTeg82QzgI+vU1lydDEBSCY2ZdjXE3VceLYwCAsKOxB8OZiEF0mKXPqTC56al8qQuG1/+CGZCh
VvEs8FERqWvEaW912J1P84mByDcHW0OaqDuPW4J8WYb+7mb7PBDFCEJwXsaH3F7CEnMjxKQwZBVC
Q4vo963bs40aBLyS1IuiN/ZJ10dD1njdTmIketkGaEra1y5Aty6IH1enjRZ9ieEdXhc8hFHWBDjj
r2P8Fny8v6N7kvgjDtwdf/6+sXBQ5ICkzxX7Bq+bysmw1QavaDDhRFm+56ZFdJbGTWdoCkbYZ/zw
4VV7nF+GdaEJ7rf1GRKe6FNs3ddZ/U7gRxo1vycc7hpJ5EpzyUZ4QXr7UcV/8A8GbL+G3PItq6S2
DRcNe+VUMQR81xUXeDdPeHG2hOIQ80e+zmhVFrmJanoy/kZZ3yt5wjS2niKhtWb1mINhmS9RnZHq
BlUeaQm3m33sd5CCpPaN6lMfl00oonj/jOp7LwIaYxcDlcI5c9l8241Uu/p63tCKA2kIqlqvOWHc
ibKanbUsjCNjgaen2H15CbX3F1Vs15JU8YnC1+RjunBiox79sW1PzsYhzqNVcZJY3rrG4VCE13sI
GhigpQjugT15oo7PcmBsniaCNYcLw53d3Esnc1ZaEOJ7bTjqXVZ1v773Ejzbbl0vJA3nMzKeIWSS
7xaK9jRZCb/yHseXEgQEyyWDFpu4zUOSvQPulLsffmNEy1bYSRPEha7RmILgcYxTGp7zCypMPjFl
ke98413q42L9UsVuGGFQUJO75pZOeMJhJyyzL9LpLTXlNgHbdU5QECLNdLQlvNdGPTf1i/BnOkTg
YhY0FhZf0gGgI5TBMG8XFFXvdazqzGXGJOtkI+6Vgf3SS9F9H8CXeky1WeNajeGaQxzdEsuuzykZ
91Sfu1/B0YgnCODt89Qvq6BAZmU1JhTYpnKDpQ1aFUwGID3S2pIItst3fB0RDqKsKL1ZWNFimi+5
guYyMMKZa9/BH1OueduwjYrGKlPac2ZbmlzRUE9mLhmGX3hQ4BfDNCviZE4/gBD7seCHJUN5GvWf
jS5hofK2PsOiMAU/sWs7TBjrRWMx+y/ocrEz7CUJvpO9Ym4grgJKqbADZ4hPo7uEZmapBLMMG2sa
ByCKOkoqDfGWWFAjGyZXybhtzornD+LrgrpDi83YHc8IjsnGhjFxH2+BHpQGZ0vh9hW1ddq/9PeQ
Y7rN89Atr7wgKWxql1wyI9yD+FWQMTucFXeSU5towaIP8RvSqlRT47Jh6A5hhsQd5fGrhR1f0G8A
5zlQO9KZFjGIyz4qFaDPR7N9Wod33/8t7UMD/x5l3FbEmicy3eqqi4Gb64kQxYP6hWvTuqMtQmIE
kco3oSyx5dNdn583kUNRuI85FRIviFbwUd33/ILuasVpjPnc/uEa4W1PLQbzM45kCEYCl0OX6elL
4OliL9TSMCX5EzwugCl0TG6cNyefVyVp0YxogxmgWmFnPAasvO7Yjvlqo1Nb9tKtU0BlhAT/OCnm
xYvuQCe0pD8czyT9s+ZYaONzmZ20QMvQ9N5rluHmCLzCIBwO7HVM3L0MadLPHTt9Z3Psy5vQnG5K
oz9TjlTaUIUKZd/vN+RCPsATlxhD9ZJh5JjOZ5istnBgRxgZcMSFkRx/avxVgiF+Wrx0PfZBFxb9
zPMA5J8CcKl3e+QVZ30VKbwYHeX+C0zFNhoM5fGrCvt1171SKt4/TcLpwHrRja6Y4fZ37xYBy3q5
vHvW/0T2CTiwxfdfLVrPg60uqKlD0zqyrPCI+SAIccg9vYmCKbNRc4eFdmgsBBmTRXvEkZiSGst+
7mitQu+Uc38u8RePvbl2BAmQCCEui0Spgw9/yf0539Sfj8yU6AZ/K6PqtoGHET7yTX9cWt9nb3lb
uCQeOrCQ3ABerhbJHhiehLx3qJvFlih00FeF0HEnw/bgLZr7cLolFL7BNL6YfxmeQtXIaT6zCJps
JoANxSJSoe7gOji/iP2hMrOSkClsGTuOWyYI16rxV0uyP79tjS79cWEaUQ9sm/7vMg+mctO5iOD9
RFVQaTMIJgXXZoJ6WZI0fBNSbyGRhTg7b59mKi1Kn7Ev2Z2VBxZtL0q+ib+ma7lkl7KlBf7wJAg6
uldNmGL36cWpiXvmrIkOUeMJnrdZNYTpZgUW5FdOL8AFbqeFBP6bzf64eanmrOVviWVyyxEheJdi
RBNU6KCT+Eedo4H6ZKb1Qt3jwnvd9Lk0Quc0W3CwkPVRsYjNeZRxZXLNEKuoRm9quW529UezzTu/
U64/4L4Rp9/70ssQNinEvwilEPokK6467PLusXdPi9Up+vfu57iIaiDA0ZMLI/uBVLtmvghnLxqL
uA9E9idWJLXvnmTrXLiLmuCsby6Jn7BoFeSttBvb3qQHpW7w2+zUwCbCliQosT56ECl66k/kP2ZB
zjqp0S+ViGtq+TJO7zXMeUCau3n79/pCo/6VGBvciOLZBVfSvnMOCD5GxbsfZPgXv29PPuufTnyt
06WwvW+rjzzMDGRLfaiMy5RiudMh11jamo4D/zmOcBP5sPj0C2nv+o7I/MBvnNcKcoxTd86JEw2d
AfkOkfnQD/ul8DauZnh4YRtYK+2RiRTBaUuPR+Y8saz1fLjLP1qaRzxZebYEFjaOPmt4sGKYCsBE
mT0RVyARurGNxDOY0JtH5FpiZTxuch3U9EWMKotz+QllbOeutcVCLCbz67V8uqIPZnoN9iZrd6wv
zpQuyLimvRBpTPAdLjZSee1OHakX4YQDkQLzpIp7sAzW/TFaaUlwn3WTUp+xkf1aiEhNbqODUmzM
SUB3tZIjZa85I5RVIe91nMas/3leH/H2VoUZ6AR36Up6IGR1BtftWQzdqeIivhaLCgPJ98OlUbad
ih1VgzuQ17IyawMzku1jWc7W2e1SuklR530soFCY/rAZ9bWF1eie53IANWdiPXTYj7iyalVkNd8c
rN8gx7efSvOskK6U05++tHAKJk+ENyNcBTbneoK+ftKTQONAEcSnWmSws2dtAnH9bGHAqFkJwYEw
SmRXWN3gTFGL930+EWWSfWqrdoh70G3Hfw7HaZD6NJaFeyHgeDNks0Dx012DcCVcPmHxzTFcJtua
b2HUgbJ1gpdqhZu6X3pm6BjY5Qf8jCpWXZqr1DEa5eeOqOev8c6TVL7ueKEngDZLsJG4DZjOoPGB
QV2bExgOEy953ah41+DXIXhVmMezMpfeUVa3GsuD4UZxAGM7/sUcBt4Q+ApRj0w7kFKW6PxJhqf1
kWXWtfa8njAY0qUCK5+uXHvjtHONJpjkYagnQsLX5QQkB3tC2UcAKg09tQ4nRg0+6VrauZ+qB8kY
arGLiFohV3IhyG3Aq283EpPNwhJCaAfcQ8w1PGY1MkwDIFpESVMyGwZqKCD/H3D6Lux1JJdUQcEW
dC+bZCN/6klG43yJqZvqjVbf3UZSrt8GvxWNCvNLJHonQYoyuR8e83kRpf00rwvYY0paI4U3w0uZ
AT26od4uc2gG6ANsqhCZleMU1WIu6A02BL4GvWJyYrUwSX8XoN2qvec96yDmqEVZGIwrMlACAPO6
oTDLPtodgAXy+PcEvq2+dxyOKKX+2q7WKmiFpube32YEpnbd3LwiMfTT0SsC9KfZXQOh/jZcuQ5B
Sk8uoVt8t6o4qEuMF0dPcgEygT9SR4KnA8Jr2yO8V/on10Fn++VTdmrHwMBUSdflQwYlWrcKJbQF
f3E9nZqXAcifOpVIsG6nL9lBHGAudkosZpWSfQbp1GNWZb7x6HA5efwnExe0O+RYc0sJV8QybjQn
xRQW7XNdV1Ejs2dg8r3tfzPzfT8z3ayVzBT8JybIvX+7xpCcEO5mnP7Ldzy7Mfe/tJ+rafOEsijH
FQwQC/Hln6B6qndIBbBC2QQeEitGzTGZAfZDJACbBBT4xin2YWH36TBcNN8S9ijz54gZNtE4zYTK
p/2PkVqovExKs7bewltwryzm80p0Po7ZjXh4xqjBepc5Y4Nb2j8LCOk0kies/wltclyPU0wXrori
yNkhZsjLUXVVlv4hTguMjfC4+1vUZ337LdhlW1AWIKbAcPQT0qBA7yJzObYhP9yw2g1chfd5v8ix
ZuLKaLLL4kTEyfhiHVXY+FGQIN24IRKPkkqMKEtPj/Xw7VhXl/WFPWwkOEtaAv4SbSbLOFOx/gpI
mHMpZmq9AmKeN/hKsjyuuuKp1LcGicHOebpoDvMGZMJjpHvr7QA4UHvR1b17cSEia5cAD3kftUpo
pDC0R4zaQWOAbOwJmKNrWfdXMJbmbkjQGJbH0Agnzaq3DeFs77T2on8s8mO/7dzp2NWGFY/0KdH7
98rAC218vmycvuXsODKl/EAB/A65Z32bccJbWkW2MEXJCtVtD2M960MruUZkkVLyb8MBdF5Zk2f2
dm3gpHaDzKuO8R9OrVh9RUkk+POspduWAquYZCaxI2FWWQSsGNmPj/vAzX9wP+rpa5wh2SmWWUJ7
6WJPawrHcvrpgksuS96Y1tusi5UnaFmMw8yxxkW8r9/uFh1lufIkQHFwpCxMUGndy+e+aumTJHCz
t8cf0aTQbTKTTy99bDFgWpZr8+ZHPgYn6+R3hKfhUTYKgZGi4MD0C3hHrSONawjURuiS6Vh5koj2
r0CinuZ/dpfeFsZRNqLXAgWZVoV/iI6CnPeAd7ArMmRM/niVOXdV9qk+3ZuWbEcF+lHErHh5doNb
bkDlEL3v8I3MeOzZwPahD0DqrrJ+E9ZkIMh/zjjqTMgpBKZhjUiiI6o/p3/rk1cZE5APKQ2CK4dr
ub/feDWeiWCjBZnUQjdg4hT+xoTko5h75NCUFOx24UgvqrY5cwXgpSXnGMxTMx+S3P15AOA8R5Nc
0JxszlsRaVEbCzfcSVt9Yxv+NbqNUrtAJUiHxfWVjSCPtgjery9bbCNXJK6LTctN7LJQIunnQt3g
v6FLn/qSDDd8r1Ti0AoQ61dGGnpAx7ETlUVq9pWK9evnCS27Xy4yHVdtPmflYU/Oww/Uvz5P5Eez
mrindXVkZ/YIkBmshidybynn6VETrzeH2t9BwSA4oR+O/KC7pHg+ETCYZU5gUqZ9sH2NtF19vSbs
pM24PIu2J5K8FzfQzh3yFlI2quRgvBxu9RSzomFBZT70QwkXhcbws+JsEbkn8j7kGr6VaagrrKmh
dwYjXyEwDcGVJS9T/HSyIyEmg+itm6fz+thuEIxRSiIsvg27RX370g1vHxTFaulepwa02/++cwzy
gdfwyytr/aB37ViE6TCNYuWZE/fCRgdVsaJ+touBo3CdsezwQNe4YbDkhfyYO2zXMT4B57gL6hsG
zY02El50xSK8/Dj8yqA8uEnZpdZTEE+1i2lN6jlkajJoP3K84zYuZVwWRpSAZghTDeXud3sLmDHV
9M0xNEAyHk0S78dowV4Jy2RYDxJZTvT3BL5D9auMKIW1w4SFKBuSIB9SsA9dUDFg+YEuhxA97oph
BI6j0WFrbZE5TVqE63GbmCIqcG+VUKSNq67lEmFWctL3yP81VSzV8gjAjYkiRjXtk4MqxFRA45/x
pOhj6cVTXqfmFA2x6dY4fpoq58HQlDjw6qWLnslBnMWcjC1lkJyFswDsDbnnL4PS2FpkpC2+imjx
aGORVDmPAwEUG/pCmzzA1/wx++77DRRAGzgWLOg8Ucj6RqyJyLj/vVMXM3bWOMGcr6eu+2Z30v5/
YwdNydz7vjBZtGXic5sqIWb3DUMKw9HA0uIEozFRaHRjoDXf8PYTwL5I60WdYJ0KVgOxJXkwrHFh
myrZKBmaz6htZO78bGT4T9GekFyzrZr7Iv4ei//7VftatgGjYdztMQQGC2Kpt3rCZ23mllfD0iaK
9dn55+a0bI+mJLL0H4WNoC7Q1GVpTTlQaNIJ8iQddGDhuXFfml3InXCq5Hrlh0R2gaja9v+/N5ya
r45MChX9Ttq14yiF+ahGf7/FqtT4r9qYl0wNDMuQeJ2VMbiZDgwMlOuNhI9/pm4CaxRAW+LPs4dW
0fvKjatOu6+Q+PE3bWxY6RCDf/Q5gDiL2vS9ltBJ/B/nWa+4jL/n2btvgtKqNEW+8F3jYi/IuqeD
wOP23IITG7SIAzhwkMxCIB1J1yB9TZ91Q1P2VW4l9JIwuOSdWvTLzSjXvtopUAs/E/fwD11s2T8S
wCJqdYUJo7mBa0mr9Fs74fDSz+6WjZ6ITw+woRx73ui4exGWj5mw8vmIplimVeug10wNTJKqonq2
4YPGjTtH8rJc8NP9vwWpNNPkQ9XoIJQbL4rMyNqPQUib1voy/eOTmrsn6y4707ETYZznhDDZvVmH
eE3xCNtFQCUafcJiqcTTejNEP54jPSk+I18/WCsrNfI6+nIDo55VEdKR12nFfPztHbHQNGo4UQQe
DcBKTOWkG8YcUpICxeITupO9w9pLg53EmUaz0URJhDrIl8BSzh52ReqLjR2RfgynWduz3dZyqUTQ
QX/sURo+xtpQw95DmDwAIEQetFbFo7sAdMCqVE9VnI3O5trahlBlb1gE16io8a4ULafrDcub3RmA
P6mC6zZ1ZyalwSKQ5VU1ATDTLCoij8lzQsKhR9ZrChkYQJ3WjG63I///rjzADR0im3ve9SvFK8ZA
i57p+RmCfQl0+EFGozyc/XlmNqKsWj1ktYvmHRT0g3fMMrmSSAfwvQ9OGZdae2QP2iijlO9Qz9KS
C15sP15xa7zHWvJd99oo/aUMnOLeXGHjHZKvMVwsOd76eCnaupEhRZvPPqP5mSx46bB09+8QWyUw
G3yoBgPeQ4Lr4UH3l7K8qGNOF15J3zUsGp/8P8IHT3vjqMYpbFear1h4kKbZNCmSfMEKAyL1Cq3s
cHLX5hPzSJ76g5vD1ASopJlivpPdw+ZA3qTQOxve2Koph8VTztz107UCD0qn9E1eaRPfKd+c/jtI
Vm0ps1egranLE1ZuZcD3uUBBsTiS2bTsLrX/QDkYtTEldSBk2FlCfoPUfZnWzSOPfDklSkcqmHIY
uLXyJY4+tSQH30787D1hTTmNROn+wcUhueFcTBVbwH0X0InmddXTewU27B+zcmoCStLLlMaA+LNa
vxB4Eq5h0BeP24lOlIjuGc7lVQfqOpLGUTDH1CDQLS9iSD/nif6ZRXek2QoBzzL/GdJxD62alWqy
Tfcrpn+j9iLm4YpkUAr8Gbq+ba2C8FGb+WNpZNH1qnr/bQTm1wwVZDVOPYDMVq6cyX1C/rgG0969
RlEmz/dZXC8wLZdthkMEt4tQJGOulMsioBOqdoH9GxodBlVD1yvM9o3NcRLKP21Ja15beK6Ejogl
1+r4QcJghrG4vziNe+/kYbl4Y3IUn76oRYCAywqiMQ/HWb4vaWsWcsUfQ8OZmiZdR5d6BfeHk5lr
9x+p1tcH/LA7bboCFeFYrS9kjgLPqNa6VrCWzyKllGuUc2BZVfBKMEQlK+uWzay18j0EoDB+h059
E/a9Fr6efJDt4A3m1hxhDSK+CqTKLMq8UOr9BjLjr3utun997m26wB0HFn1er5SkSdThtZtd9VCx
H9ah5vX+hxs9nCU+8gxkrzzotsikiGKbDeIZ5EoKuoD9JPlOfgDDiI4hEA4U76eTXb9CgKPIJLBS
Ebq2XzsEi36Dqxt0diF4dQHB53JQpEiAFIVwDr7HeoyW3utH+4exy/SYM7SunyMM8ZJXLcrhb7wM
iOPJ9gPvzITVvGahHCq52e48Z04YJmM82fi6eNs6PYcm+47NhvYoqf1FM9lQtWOLzzp1KfrB8w2f
kCvJZ7LQdD8JB6oI4Qv9T7s9blWpQKIyoGhuUslop2T6XTN9C9u4v9xa9QXAf54rvNu9Jm9jAros
uDA9Kgk1oo7+J9ZiXvURMhDEn4E2mwvOuBMVcwSDMSf57wty7aNVvPtfGHqbz2jWe6o2SkqFdm6A
RkGxoszs4qXVVY1jc2dIrgr8+zhraHSJYCpqLliK7wUx+umT384010eANcuLFwjx91OmXovEGSSr
0FLzwQbqHMrJuCVEtaN7Yt2bg3rRhn7xQ6msJqDYVdZDdYZ2Epdl82SxpVginp0dn+XizrS8C65v
VgXyL1mtPrEp8UeLTPdtIibjQWlQGFm+xfJLh7+34aazbauWEhyp1d6y5IzIkdg+fRUetP04E8Wk
7ers5BwiJj1IvNOpejoeuRvO9Fmb82/5xxnMynX/wz3YLUc1Z4zhwyIZr/5jV8nGUZRxN9xqaJvJ
CbD6YlIJi94IIQVVKnfAqzJeQzXhlunsekFjKs7lxeTIV8qI3hrsjjXc82+RQ+Trr59qgnCuPw83
Jgudv0a+RCt3cbGKZW1uI1d7amMnExBQhrfxJP38NIpB4nk+YVt/IOKGhKziyfqu44bI6vdllqAQ
o9Vaqg2KES4AhP996uUaWrLnXIz7ek5VdpWfeq0LT9tD8bZP2mKmOFUt8faehdI4LwyDm6k4TOOk
g3hM27bVJgqc1ax3dnlzZjDkO6aIht4ClbYVDw+bIaI0KuZPLo8669Hyv+IzlPNdgutXphAf+3mf
KVCFCTuIdEbX0xfZyKfn9s4ZfU3ZtIhcMxK6LGZq6RsxTf9zAnxJdFsFoweBIl9fMoASGYtenGQM
zyhZStoonEGqZIiEcmNM+dp/Ff/CklfiJ9/4m94mwenxRziFwde6NPFzjdGVTdvUV3xgdJgUwrfu
g/tQjCVXiUifINca3MlDZmzVf3PWLIpOePgiIhns5/oo5jIxs4U2IDDKjFffqZXz1bniejbLMCfn
w3hvTOMmHW05AX9Abz36iEATrCvi9Ovs+nXgBaxgx+Hc2uEChYD9Y20ViQYRStQgReHyNFUqaTgS
g4vg4CqKm7bL2TTNGjw+4pfN6yMMEy9qEIq9DJL6G+Qf042ToWF3JKCR/oUfn4TxO1z6eQXRINkv
KmvpLzwuVPENagKaULnu4VkjAyTgxZeRkDHgSj/+L5SPKLazwmKxWQ5qBMFMGieKh4RlynHhA/Nh
teaseuP18OmvMCsqkXqCgOpCcI55FzTcSZGHvej99w9GdizMPdAMN2aVMHMlI5L/0EbgO8iA1Y9M
S33B9UrQw9UBHXNgmXs/53cWnWtcmGWtsXIvNk5WOm/Twkq32t8X2/8HGvA+O2omhPJt8eufPjSO
eIT0eXgKg/juUob1tGFCyLhriO7gjXTr7hpZ6k4SQ+leN5WQk+wL4BRH2s7PimgRkQViUNLQx+yV
PfnTf3gMKc4nvow4rGrQg0v0l2PVrhzAvBTZmVB3cerkkqYTKHPlD7VL36MmssB2I2j7kz+53gu9
4wM6PYpu2MqCu0NJ96EpY7jDO82jeRG2QlgdoneJ8jTR+RwXUWqgC6uInpneJhFVps0M3uxuTDu6
7W3Q5IPLjib+8D+NxuYpgUdC2gBBrSk/tlkaKyi7eLd3bNpJuagaHAsE6Pk/rJLLJwhhGLsrsWSk
a2y6PJrNZrQ2MGapNXdRnlz17nBPhPjSDW5drIkqfrvtOGw9PKjetXf0iHXElHWR5o7cAsATJT7u
6SS/XfYjHDww5X5TVsXkPt/3EnfWIpeGWkww5T9VH1DeVNLfEmETb63yqiUDOTRnKrUGAPoNpD0U
Q5GWPEbrdMZfqeHXWLfN4KvI9kurfeQABSgQCek2J/n3KQGSxw/Qq9FYT8lEZdqbjwLV5RQVGbV0
LyTLbORo/DgPLXd/hEeB9YXIazz+QBY9xsvK3QDhWk+2fmHjjy5qzkatKbIE3+8f2C4KgfEcWN41
b3W++s4HN4aCoVay7JpfQ09JawX5kf20vbWGkJ2OyLDG/CapAuFYpF0lCm3Mr4UhXxh8N/RLNbgc
99XiMlWiHkx1H9mNZJUuLzyTUDL5t7nYsMkkLTGFh93RBGhYG4LXtT0hjBTU5m4daS+x+F2BoV5z
RM18xzxpNcMTA/g77dB8mY1tD8RRpCyBB2YMNfGXVMBfycoCb1gIK1IRmRMxpasQfzf1uVqqSi5a
H3khWjqCE9IunZZul8hykXkak6RpR8x4st0oHWbpo/sfGqntLmEgQoxgO9PkWzGaRcPZZVm29eit
KQKSYVyFPcuP6APcT9YRvubTgGmH+g0Ex4xE9KfChr4yUgyJGQDpQ7h+377NXT5Qtxf9IheQ6D5s
9qx0aP2hOS8OGGr/MBAVp9BJDHFPgse3VSkQh9HtY/065tGrxSrKr/QdtmO68T/EJ0+aw6LEZ3ea
LiUeZXfcw/JAswxq9KOs+cpjl7cf3gKeCPxkpoOvEyAom5sX8HpzOD72LbVhhcD5oluWMCE7pHaQ
4dcMEB1YgWyG9+5rCbhrffkBpTDiiUm1EpYQH1RDEuHF17EdTKmaz9kSHv0dfVZOA1v9w+xJPOqA
vBxwFV6KulLuDcVexDM4Tb+uPDtFfyXc+nYEfbmn9JHSTKIi93weoAYON2WQCE1RM3L3foED2EV9
kH/3VcYgb2Zner7Vn7oiEhKU/IP9fK40cycIxnV/OurpZyDRNunfd24wt5NrNuQ0MSEysIrIpdD7
V+6MQOgdwZD3ojeuSDtHuXGt0Mga4L4HXqOv6bgOVcfS+9Dbym4iMbfyLUWwgKhBcNaHSopbtuLk
Fmfrlw395sP8HnRocSdoonHLgck8UwuddageN/B6WQcB5Ie8lNQZ6AWs+iMvCokOL10sRedsCeTM
C4PkBZKqcfZhkSDpgSKoacfavOuumQxjp90VyeQLJEKzDjMoLZxqqcaUOTarPPAVqym1fwdqTzuK
xhMcYD5VWiarhek0Q80qz9CA+gvOokXJddppG9i+yrY601jd1yAnZyJIwl2TTWQAjY/3Avsqr8SG
f4YUa60GBAu2RmcFTKQmeZ28AdJgaIsw984CRIB3zsqmjlr7Qp8h0moyMaGhG3Y7fy6ShFSDLSMX
jmf8S1dRPFk2Hn33rBXet+EB95y9WJXTSpkKrI6WQ/qWUcgLvZqpQN+2LLmwcBzxISQ408Csn2wC
xjXVF4qMUrkw35CTAuwBeAtHW5ctihMalCJhDwWW8JgWBBqwrfGeQZHiCdLsKOgrRkR4pWUfckJT
On+tEz4v1FN+sNH2vBJNNt+3Rad6JdQRITyoW51p5Y/Tlkq/0PIkBnBsf76YnE0A3/cKrPNRxI3Q
B6XYxm8aJt6AoNKUXRcYRH2WKRq3AAax/9MILvv0CUe5HD2ed7Tz+rLSX4zLqHcrD7MUBakyUIAv
xwgefHzscBu6wWOgTn2VnzIHDNwIVommZjtvVpGKNqmajjgr1q6SeCf0cy0yEFYAzkbHB9PTFLLF
+nXiRuu9c59gfKfL8sztVS/+2lgC5CvZ3HkZ6BI1s0MqVC1IgQ1Rm1me2vqMVyuVwbnzP+pdtTw2
lXEWyCf3rIAA1FcAYWc92/ZEBxbOPxbMA+6DjZiOPkSiw6GlX5iZaar++H3+G3y9dJ2nubIB5jsz
o45Z/lOd247WP/G53oPIA5oCpfMLmoicM1Jm7TM93peLK+Hdm5/bqPc8HG3tDpOiiouV1o4JjwQo
AlsoCzYPKkAZEEoKz3qhXt3Gog1sWGJAt89bvBoedIMomzf87VdZwov/uT6OnW8j4O+r6tUQOXVj
CVYt78XEdyA4JkLpnt4cZ5Tve2RzkG1NkqHtw9Ojrx3gs1wR+vqcbV3G+FQxFr5lxEucFL2yjatN
zASIQBSPXfCtw/tbBUTV9PAwU8Bjtca+venFcRSqcPdT7MAqOOtjGRA/k+zN03qoo3N7WKbivawd
61j2JNF8YpJ2SeGpOsI7tWc/fEeUOWIr+/1riIpz0px00Kc95WpIyZRtGISX4MSNnv965YYYovBS
6gkI/MUjOaMiTlc1wFqsE41vvj8MNRLk5l4jh600YC3GV6juJD5eOYZNuwNWGV61kKphsr1D30ak
gxiHeW09gpY78rmqP1yeXwP4rlcMbErHJtCIpyrvH8J13Hzedzz34HdVNuhTnbuElTzxzP6DerjJ
aGoqOU/xiZdCx75o97z3NjhL0LTEgI7Yj9OjWyb7i2t4Q/XTclmTVVk2mhV4mY3/VIPbbPa7NTsK
jkkORnAh1oxkUti75fhLesEI+QmZhLM+J6eLm8Q1bKMHaWhq3ghcVLqC7UrZF9TFdUYs+jF+6JBU
mDdI4HWYsA+YaE6OWPcKpLx1jrD3oZsIkRTrH0ekuBmRXqpV8HPDtKoZ7ySUV5U4+ddVyaD2McXs
QomNmqRFdURauZ3aE8WstdPTF3rhLP4Y9mw2W7trYVrL248NnwU+7rDeX5fG5EC8NwLenqVIH+zp
7XpfljboOewis7JQK7LIVQGCm9+emHEPiF5C11ugiOFb+ZJn9aLy6YrQQqtOukT9SqIWxeniW5hb
chAOmdoWRdEHzVxpiSqO5iO03HUA9/qf3BGq4dKx6mvnTTuU2aA70OJ3+En5xMoU4Fx6T2XF3MGs
hA1Tf8c3YOPA7EjpglO0hY4dBPH3PcUolOhr4Qyr0hBkF54YATM15Rzusf5b4DAy5/FMCx3uVYVm
XkAUtul2FQq5Qjsz2FOhLtWqzm6PDGnh1NT5vdrQpqUuK2VmGFhi+rq/pu+Jb2vX7G9ZXq0SLwDe
WK3eM9SBmrEdERsHutDq2L1APKiQG8LqKlIrcb3CmU4tyhIqspouDYKkEzqx9aOSnLxHuI1gEhXh
hgtBzRgTgauGKX+IOsBSQSdnhQnEpEzc/dnM6yiBvRyWG9eUAGp6wq1+N+v0cOP78z4freqGXP+4
+kDWsbWmz+o/gilB4qTW4L1u8XYN3r+zKZ+tnDOEHifQ1w/AQNsLOfirPkuoNOWk/vaQUBofM+K6
tC1v004RUmfQ2Lx87Mu9jsyQrRXnoMJir/St54XBRJuZWJI8RqRg/9Ma+BU2G9FxCMecQDVxcLS7
boFulGkUC1ltcamJjc7xouBmd6UtvrGV+otU5m/WskVl0wiHRMZmLrY5T9v/0qAUhRZdUIudQlbN
gLGOVGwlb/GQ/YmwBkT0OUkDubTPqkjYiEgxzNLr7dJpffRWCUizkyQ1uPG5RkTiu8CedL3fsXMp
nKxc1EKWgg9HL0sy4eb5Sq3KM+8cJSE/z9lM63gu2ia/qf0gNSyo8qTcIxVB7UJ9fPcFXVa4DEtO
D7Et5Pw8PiftAaBEMmR3Tsml0gL9aQXwLFzoMuWZNbokWrcZ2JfRx7UkOFxgW/rntev7XVkG/aSv
oXMkK//+KqcZk2mSorVDTSZlT6Wn4xsNhXoCyOIxIkV6+jpfZyd/QqIhBLlH7eZGMrU8yL/5RsxC
bJVT5zsO918/CM++yFgNn9SbcpENCpRhj9FB4l2jAw995Ln+l/33GPLe39xaG8j1aZz/JEcAQWpt
yc7nWL4usQtAuhqPc/7U9ZjHfvCMaWJQMgp0TeHbjbCJhLBqoC1pzQ6dvJGu0kP9LTSnLv/VZG4Y
uQ3Dd9zk1hEg8M6HBIbErtp4lt05fwXa2AQAIprU8ik9FyUhJF/XBx3a8KkQXwoadeWromObNsL7
ylap1NDnOgrin8+JTULMkWNlS5o5iKuuBdM0kGK6ky8xnwfW79N959loUuOO71Y/KSptsOPtqqMJ
hRdaPitbz9C1KDHowvX2eExgWPOgu6bxYUM6+0CxAzG+vtama4I3VskQeC/I48Q7xv1sjirxsHSK
ro8cbk9mLEKsdwRD/GikqgLxgR/BitJ4MwatKgxX7s6w3zMZ231TKkN3rKEP/kCEhjgyUvBFUQEY
U8xXn/C1qJhPlntGEjuvveVg8xprtCk61GDTO9IuQ9Ju/9qbGtCWsg8x3+jaFobrbxN9voSPjq7m
wweQSFGXKZbkCBvMzBz2p5pBVYe+00YaVMHwpmQSjuPU0VdjJ29jAo+a3ropWX3/oExpvq0/Iij5
Balkods4VNapoPjOOskWukHU1ytSar9Kyxf5MmtwHLsImbR2v2kd0LUzfDtUnV1ibbvbJUbbOB9v
xGGwRxOa+lmyQbNdbbOml46ZJt4BdrsV20csib6bKrICAn5pq3JlggwFlZwnRcfRm7PIrVNiIpLY
RnAu5j15zOKhpxDPgGC6eSDMajaZcmidgSmsDOhCjrVlISIGDi9bUOFjnk1I6kAZEf3/5E1i0OVT
k4+SeaGcqY37Vrfquah2hMxx0JcBY2Xs11yWRXkWAeNGzMbyFIvScv32txFEdFiImSIhP3kTbpa2
JH23ps4E1TwTCqBGtDg+O5lkXxZwjEWv9J603lVxFehCbIje010oa0T/1NaSclQmw/A9yh95/C0e
1EctLg9sX+BPcDJDJWWYIxryNun5+3QdUnzpaUTDkvQXYSVl4Yl3URq8dA1XKHBBRFD5LaN2yVz2
7sKtlD2AWXTfWfLRwBtEJlfN4EuqfKdXIiMBcbfgH0cwcQ3uyRtQhKUBr6v5WqozwI5rfno4hgil
zMVSiyYN7c87CkvatUvLVmoDyC2MWYQS/0ZjJySmnvc8oStCt8h0FisqOA+ArGNIitsvdjMocaX5
EDa1AFx5Hv8rXtRH48DNgM0oprGzgNElLKBIKaAD33x+3KA1rxkPTIyOtblgHtGlcQRrgrJJJs3A
LfMaS5tTfOQp2J2sJSbuW514ZB1vfiZxwmKh3MLfNfJOLpmLSyakojnL5eFFYDDPgVSocew4/zGL
mofBb99YH12qXGGwSO9nTxBVm8CM067v2dkXGucyVaFG20ypMyw/6gUplmHR6CftuOoFkh4E8s/+
JmTo/G5H6U60PRK7AodBsmKcctzKCuoUhoKlOnYdst4UrXkWVQIDJKBWEddOSvREwhl5kGqqEbFV
oNnKmtK9BF0lC1IB074Nni+7AZgVBdtE8SdEEDMyOo0Tm3MsAQ/N3nQUVUCkWPF/59Af+WpTE7QM
S9GCqxaSi01aolHP1WxFh2T3Ov1v2XCLv7VITIm7SZplStuRfpIA+oRr1dDaQjVRjS8mwAv1RMI0
a2gMCjOsdQRTijswlEjWYDULmjEd74+bznI+c/+3+wwfK/RXKN/7mfKJ/aQ8qKd44DyWw/N7bM73
mJACB7umTRtT3xMxJ6JhlS8KzWGw7P+IMrtBgY8ZlY/FoaD0ypINXMBl3MA8Yi7uLWpD49c/XtwX
7BZ89cSDIWYa9Cg+g0vj12hvqXjI/bP1CpOmdKVI+/JWBiSSOjM8jbp9xBs/bQjpCr8KOMzUh7Wj
N63aMEd7BQlopSoT08HXrRW4dZ7RVapJ+dr8oN8bt8n3D/y2+rbFDkCTZNR5g4S0xjpfPS8OuGTP
I0LP/15CAVJQKBgfK7yp7Qt3pjL5P3+FRds2CL5Tm/mr4IEnSNoXRFGFepPJH/TGe5fKcDSmrubY
hf4rrmJvckz77f1+zNPOGSTLFeD/RvdWCAiVfsc11r8Rtr85C3u0Zt0YX7MKBaiDaeR31JQdBK8x
QPsaKd+1ups1TzSFItU46ASd9O/PdA5b+WmMwbdmc+vNyc0w8bnXry3N+U+nSuEBqIu5pyl33nuF
slyUYBi5Vs2a2kwx7fMT2PSzdDl0584dRDHfbKE2bqfLQmlFjMWEStMs4HXRmFCamnmuNaMDyS+m
SWPHSUvKzWG+bfq9WwDHQaHOm8X2qUUkPr2cLjt7aAhGQEn6wsicVZqoyDgN/zm6zcD2Z+u22wdF
33baUX+GsIiU7B+Lu+QB1Gl0aXocKZ+/U3+QjYr03pUT2ca+D/bM3KO1/su4hg6/PYN0v5pvkq25
TXCp0nVWbYSRXaH9u33RAzJJXJrCU4bvLtA5QyoRbCJqnY9dTyKiIcKllcbrjRnheD3szkTGZcRK
uqDd2fwge/mUs21onUSKJB/CaViUgxwrgPEVJ59rjKy+YLpbXtDje6o59HzZbey6lq2cGj4qvXTx
Z3tAZTWQpmQ+8RJKrJyrn4/2u1hLhoS5k6p2nySvSEvCzPROBW/Ko1fDRocXCsY5USPNX6vkYzD0
y2DJT2tYrDgQPjCe3GtuinaF7ZlN5pzgKeN+SJPD5Y+g64pVSQXNrwiH2iCpSlqIT/AHCN2IulZ+
OOh/d8dGsQ1sh8dYRWbVhlB0h8zXRNfZ6ughlgXvCGiE0+tFd6vMwMfuociZVZaCNogYAXQmIQf5
gOMcGmFk5zJrKIF3te5fESgQAlB4Gh7zk+ALGp/jmy4HrweRMizSJu0ye2WUAKQ/o/aOc+Brk9XU
pCvnwQG7gCBx1ph0mDYihsuw5ryq/It26JBQPzRu6fBJVXXNyFusyK0Nk7GaKX/iRFMk/pwwHdsS
0UKhEX+vQtTnMi8q3VdaKYpy6kmaQoZrgCIzBwO/uP7DRVPSAMrtu7iJ0/9rlMkItLjNFubuIAbU
vqKPS1zHzb5r0qeGDyHsTCEiD3rgxQV0/PPnCoOaYJCPh5nI6zlj59gwWK2xSSdtLef/278cfnVf
0IcaQGRSH+0k7IVOQiEEgI9bomFLv/kdiaDNI++/Q05fLc0dXkhKS1Xt2mRqlLfVHo6ZJ+yx8yqz
wnQuBnKh95Nfw75hgjPvPHqZRc7WaipWkCb/ka+q4tnjbtfwIbqdp7qkrWUndE4vguBQFbKCo2rF
S2L2cwei8PLkvqmY30CYvPYNnfjzojPocgdXpzgKoCNwivR7aLZKGOeegsmXY/Cv1b1hcggQ9RiD
AG3oSxPLy+K9Gpbab9KngFUxfFgFkdsBuNaCsvwL81+kaesiXAiMWRBniMhEzzQBGosyBTwd7LNt
eDMejxCxpfBmgMnqAxUxUn0Da9V3KUfzLGVqac8McFypAlb83L4iaTjeqsUCIoVO8hZ+/EulA1uY
cr81up7qibRgMxdlZXQNkkh0dFD2jXEXsmqghQ0zSkfTLqeH/ZIKskp1INtpeMydFIs6L5q7ZUMA
ZXvwgpmxRxGu4vnHC9oiE1CywptlJNvCRqiJx2KV13+HOTDSpndQSG+oEsthEJqcr62Kg5dVUYIF
wUPMahuwa2ZVxT9Mdhm4eqFS6jsPneuY98t6BbSz48rpK7ansQA1/N6EWW5yL9wGEWpS9n9aPuz6
zscai5QwdZtHKUxgHm3ZBoYR+24XQfCeyqxGys0iuBLq/vLjgQ1JXC9Csm3PLB9Olo2NDI7EAXjd
x8H+lD5VGBTD+sPxOEMQ+IKpyaIvryKn/fXWlnxD6NrMvjqDvhcc2uuS1TkhOFNbvBUtZpYdcuOa
ZFaFpjldwObdq3TdLtWvF99JdCREoA7qBFborFmBIS0ebfc/W1pWYToJPb64u6zmle17fOy8ytYz
D3haOC5WqIbrNvmfdM1R9Y1kyXGBWxIroK/2Hv9Gkmad5Bfv+LGxFlonGY2hBH1cEn7fy8BcoxwL
SyDY2GD+XkcbG+L3uA1YbaSLPhX1imIgzg3C6ayUBamWzHb5NRtjaZCdtY5TxxEZ1UjjwoI3/8az
uEsAQyP3GqHAiQqeoR5N3s0ZW3tVzNP99a66V5paeDZIz5m/WShfa+pUZub4B0/oJ1B5aORq6kO3
SBlBxkjtQS8vwfsMr48oJcHLltPmpE+F0YqWNBapjC5S9/zP9canNF33h+3BmIbOSf2Yz84dOvUA
HMHL8WwcE/yZqq2Gav9N8bKBHVqTpXVeI4dUpnIfaRhBDOF814OXMJDedy5ttKN5b5Lut3WstyTd
4fGA3dFL1xQ4JqhYpgLpS5A7TmDaMkS4NKkQQsYlDwMGnBPPNjiDCR5vAtJQMzRk0U/SNnJH+TFX
XQvpbbUqGr0qcx4vtyYCxBYQvEMt+cDd2V2ErX517XVcXKhFMAGkfrRLuYGySLV7+UZ4i9Di/+mW
O2GVkjN76eRo5WewKb7qNjp2aChvEGx6umlJAzeAWZj7WQqoN1gpYRnTBgt7qleB25LWiB2HqIEM
3gdqwaCCPbJlypPbUsrswKoSTJMH6VrUSgLnImn9tQJOsJyQ3vL/jdlUKh+jT9KkaGkwDDKHVtAk
++0ofoltu2uZ2hfR9jfTYoOSUCitrwFIdtx7pUV4LMVLnpFhBc4yrKkHl54K83Njqa1e0jo+1mD5
7AqId/IZfRQm0zIdJXAsb8YUNYN2Ugcg8DDGhmOFay7XjfHbK6z7YcnlT5n2fxvPo0GtiHtSb9ZS
C24ajeX6hQUaBQwpyMFJidGnG98fjOzMYzaXTLqvRIfd1YmGYYzTOIAYnFGyyZVxZxRzeTGXy4o5
vv4eNYNWpM6IBl1BUng3gxSZPy47RDevKyEOSVRukYgelt45gRejZwQq05/RyOB0fwzY16XCA+bY
tSTU5b5oxsFltbIrrSqz8BJczMjeeXtFc6La3Q3B1hBVGckTBE2y5GWQhduMOUEd3Mps5YecemtB
+unVRhzcqW/hqn1FSJ9WG7EhjTwRB78HDDbcWJp/f1KAEpo4zT1I0R6fv8NuDBDwKVAC8yYAKvIT
yw3ySoklsnXZbhR2rBpqLFfCsz1FqUgT8WvDygBo97KkyZMQwEJ8tbnPjlxgleELEEiui1NrZSPQ
zHHGviM4kgEIHgT8cuepSxrnFxPuhcwoTdAxpMhUvwjlUwqKFDdB6vg8meq60ai0lklMh9CVXcM+
mJDcOsm4G80DrcX/syCY9PWK2Jljf08xL2E11XtV5UYbT++uRnjV76yTSxPASg/L+lUEpd/Y4ccv
AZL2jv/xVdLsCLb6qa4FkAy/m6J3C5J42PSU0Pjmksp6HlU8SOuM+k1Tcx9vji2MR6hR0dGMgGNn
hZyu7+h7rXT07wGUyH9rWMkAkqpY9ihd9H1TjpgU5YGiRGI+4TyfXJHHnZfB/vSzYgEvTeDi2TMF
pXwtGaOOVTx9hZ5GpMWh13dPUrJ3c2Hm1GQu7yAaLYL+jhBPoRGJUw9GbfVv4AdcKB8BpvNTPSIb
LdYJbdTMgTm1bNipoNfBC4QfD6I26WvAFdvUTC54VnAKmDhG1nMzQGnXs9gApiXWxmMyIzGMtLA2
g1/ALO4bQSXB4DVNschTqckSdNVRXOiA05CWsoa8OnsO87bDu/skV/rfgI0nXHFOCh3OrFsKtHiX
2UUQvzWSVNfrayBe5Xkl1xvyHYIbI3WcUdI8XU2+EEOoEBUy0hGyKXPWkSpmv8glPCIH5ZJYf5t4
FPIIeXYIZ8m8DqoC5U2uJLItRJ8JV2GTZkA2RZgrQFFo/FfuCSRzQw5GfOMmgjryPBMVzt63D4Pb
fkf2Ayw0y+/mVBiVrwguei7lgVkVro9AVPDk/EYdzKrEvgtvqNRA0nGt/GnXr7sT/PKRMNk46NHS
0+rXbInD1dE9vhHVZRPe2anmtghFgx0VFQi3UsDAjV7YwkjWZ2J6IAHnRZ/C7jpwz34uB98QVzWq
eYmdY0k0vZvHz8WLcgLL9HUJxZclNeloGN9YHe0Uf00+C2uryVfbSAlQIZCKl4H+F+6/eVhe2Lwz
+PgmTv44F4UEx4S3eN496D47jeLQe56FaXoYvmW82mBx/HRxw/LBEVkU/qOEj1CrWQgfP5UIQPaA
4rEndog2UGiLu86CwskCGJFD6i2sHl4jE9YgAhitLB4Cz/u3GWshub44S90jLPSNRTx/Q8nM/yPl
eP14gKFbseLSKCUYYFTO61NMgiDCOaa1gH9oXho+79mXJ9rswS08MhyqJoleYx0iNoLz0UtDjHOl
psN+xP0/z1/u/t1X2m5z/S5dhMzHZI4l+wJfDg+TTSRizaRIGp/hHiA6ard16kK1xexvG03FaLAo
E0LXrIYVFoRO6RWlo+xq5VztJlypcSeRG6+sgC4SbIyKdwlFHDgTY4vidDTiKIWRjdvEVeJgZCd8
Cev0uTRcJZ14mpY0GPLtwxZz5Pb6/y1XGWCcSv3vwC7ab0h3PLwNd4jmtGrmxo2tfa4pSAPrfgQB
QTSJXT/t3gRb77Ab4SvcNlvV5K387ZPh3HQR0LRkHLy26q2BsU2R4CZTx5s8dK4UcetM7R0Ph/OS
Cxqu896VH1UdmqqwakeaOwdfLNNvAFMACsqIc8taDsZ4qQcSGfC8XuT55cC9mebf4WdIgcYRuXWM
E7IScMcj5otLPrRPg7VtmCp3FOQ0NoLYNnDRSF8iioGwCn4X5TIp7QdhuIUX+U/FTsvVOWjMOLqR
SIk8YFBfgBp7ZS12cre6lFzg8zbmMWgjxrV8Sfqbeedc7ptUZoGkO9N4exKVHAUl7KpAJevcNd79
7bSRYuEtV5Xmprlb9V2Lq/BVWGg1yhBlte2VSJi/QSDs8g3gTu+i1LOo0HMLU7PgJjgML9eVEqNn
zZS3mYBr2ZGeCZexLR1ryOaEpjtnzWyeCzsR1evX9Ee6hSNmZWxtoi/LEpCr2TKvWx+ok7qdzGmW
8D0VHCyI/a83MXzD//cZVdvIx2+zBsSOGXvxWyKVMokrKMIFBhYige4GD1H0WhfCyuyX0xe4mXpq
ZL26EfvjNJtYmao51fu/Xjv5Ga+liroFpaVj6xNwd3b5Icbi+G+e9Myg6gZzAHrimwE0LwSRqPQh
jhrmBfmghxZwKKloJFTmEKAPygff5dIzxPDhB9gwnFuGb+SxBFFb1kSNxYyUlCYM1e2RzjOkE2Hp
zcynPh6YRbFRpE2dHaA0YoOnFP84E5c9wal3hX0/ZK4bpEI6S1RakZiU4U+H4U/NjFwC3upNqtr9
n+KRSqKXWJMCkRJEcfO2gUT60SJJKsEA9px9ut0px+FKL5pD1sSwv7f/250ss5dX1D/nqBOy4ucG
yNt+qoLevsB58grTrj2FoAtIgLm9wE9JydGXGcRDg8L1ezht8VIBgkJJ5JKmEBtEA244syLUQWQN
yjvssP0WFKYBCdsyYtdCMTr7CfjjH4/QBU1DJBrfaiOsXFBbYX8IbRDNnNAhbuanjJwbQKV2lRh8
NtivazAabJsLOqBKRW8xeWdwjEKwueHbjwA2HIegOmVZJsKvSHDv5+1lrwRggs899mL1UcEXjki7
hceVq6HW7d3V0Vyc0ubTw1q30zRLnv9qYNYoQUyiHaBuDKyqoaJleeEAQzPV1zpiwwUvOwsGm/v0
tnV3BeiUXRPh1XrDQ7RjXA+gcmfBKMdZUI6e7zGyBknRLgTEpySDUkMg6mjwCILXnbwvA0C44AYh
AraW9KgWYJr0K8EGFl1Fklki29wyisixV7XMmSO/ABjpYG2xFm2GrZSTAc3ayeSwUW0wLOZRI1dA
MXQISSRsw7za09LkEMJwPX7LqbFlfOM49KnW+AyU7AwFYng0rwADAQprVeeXUkDa9zBZynUTqaNd
eQm4LSRCCxnW8eGtJ65nsjrCVRpL1aIiUbjlw2jStOE+w/WHKIMESEHY/E5gL9xgx60FCDkqeeJJ
2+iFfRyrgGsTJSWayjRxZy/pH5yj+yV4nBf8bEuKyhVLm0+h7w/wT7MZ+gpCV7nQz0Nysxy2DORq
vE6w7Ig/feb1JjkmxE6AYEHpr+OS+xUnK3MOCEISUPs79V3F2JYMh0DAyo+E8WXz4xgMTYgHXpGu
IgLr44fY71OjrD17E+xozPKjZcrpZGf9J8J6nU0SyD6dcYShWpj/Z0u1SjsFTY2ARgCyfNnnnMqC
YrRm7zR6Tm2AYtTvvRNr8DJT+C1WPMkNMAaIT+qs+VcORPXnLE1YKgjlPgKJOvz0Kmc/8U2WtjLA
kJnL6GH5GtsM5pHJmdrQEkIar3fscHnMGrA3N1CcHWbmB1OMZWqlZ660O/Pww/KfvePSoLO7/0o/
ySZe8ZyEQr5GIB9HTXIBoE4pl1mjMmVSyIprnFwhO1xCnVUsPTcUO2FWVkgSKoqa1vpl37CU2O2n
AyAtWg1IduN23DQOqmu6ptZ4z6VNyti9ZQ/bzkMgmy1xM0KUDWxCbpBramSeXYjc70zGh7zhR3lL
2690QYa9wlItRHfZrr8xCER+i+NHAMuwAA859WRRFPj4J+RcWOeqC8M1HQ3TrLmAzcRGe54Wvnk0
b6bUAaxdsGvPUvOLba/uqZwnjCud6pqz+t6l5makz0jzj01gi8vHQ/u1JVYBWSNy4Grev/j9ullx
TQfyfvOg8qRO1liSiE46OL510g5I1Lxfg5BifMRG/aLGEfRZYjxACmQvbMKX1YQyHiYU7pjSeJNu
frKlXzejX0J9fwzLXWB04KXIUVR1vjZ007fl3N2asfuOqx1fe2rhD7d3jFP0BTEr1jb6d4Q9vpZH
qYZ+y7pLtXgwd7M2aPKDjvyoQvkro1CWt95jVjqkB1B/3Clo3AgvCYG3mJgR0NZGCtuZZFnL09h6
Htsp25jfxuGmO9+ytPXd4ebjMjUX1sVPXpcec4ezNWNkNFtxDLvspcfB3dLf5GLPNALZbT+BiXY7
DimvBTP41M7Z6MACzFeOwlFrFrMuhoP7QO8Q2RSAR/EWbWxsrFAc1WK78FI9zF2P84/7/dLsV0cU
p39dkLcZ39zKB+x3PtgiCKa4cqWHPqqlurgo51BKiVIsNB7tpLHbqQT4c13uhgiOmkunPdNkv8k0
E/YHFPBllD5LdA5FbI62j1WcTEnRbRLHpWUO1SdPi9reV3PAJ3yrtXBDvz1M8LGS9IHZ1hYXL5Do
CxEJ5aGJBHVy74ZhK5vHyFInG+JzchHdAe77whDYvr51bWS3DPu78EpZVqldhjzF2JT8c8XaBgJb
WbJ6cn87XXNfakt90Rf1czX6NW2aPYG9RcDRxLW7MEYRMBWFk110zDd3LKQ5oERSV5Ro2XuqbIW6
fLLXOz10qTMV1LoxY6SbmFvu8WNx7EQnC0v+GhONXXVMZkeTTtEW8FfL2fAD2uLtZL/vLioV0ezW
vY8oJ93hm5gjmFbODPhOkfz5ZlkZhL3ewpcMw1cBXc9qSVK4KKQHPwL3DS//+TwC8zyEkcbSP40s
0Edx4Ggmcn8yM+UAOROODUq/m5YgmUBKdJYahfPN19EOS72QErz+N76zfbf5sHKts81Op0JZzxpe
eNQJKo366PdsdD5mK2i1MMqHPggFajc85EWoBU9aWg6jABL0wZ6pgTbjCmO6NBcXJpVVr6cxnR60
TfGOObALlPAuk4i8N9qLvdo4cJy2Byy5HxsZ5PX5QVKs1tRDPwyu1GH2d+KmHJlOsjwjbQYEpHNe
YgRXviETyVLswdfA3PNPdzXjU4LARTFkxPtLYufZZnpySE/IBa7lZ2g0mPmv0TNlPDi3LfFzv4Sk
vVJkZspVg4CrCS8BlFx7GK3IS7jqUdgv8f+wVlArlW4HpXZtLkL1CFwlX42GxQ7VUvPjzfle/fEL
TCKygISHkOT7Y8edKnjRteL8NFBn1yk6Q6ufiSR9qbFKDOmSKK1sKrhNWoXfP6cyC6q2Vs4qGuYe
PFMURI8hCBJ0iSdYN1gj8xVbAaOALZjQ/5T49iEomIqBXIJOKyOPkrGkpmZRJ+N6VnEWRKuIwMOK
HWsDZ69KMvYcIcBSI/1uDXyty4erOyRXprhtb88xoGPNSEQXVe4DQuyxVCvNbpoyfO2Hpe9P5LU6
DF1CKVEecueDdITCgVNoyv7ZVPjmdo5wwgtgW105i4sIPqy0FDTCZAv5v8iugIYTxjVe8GZ0RlIW
qNtSatOol3luJyemeMeepvWxIjoC4WusfNnva7MhWZ4rBI585EqxtakAeCscxjWYXwVflSeWtw1T
w86Aj7SlEiE9/lFJSlGrLpItoSCTFlG/VhFb04s/la7c3IE//3KpWUOWSSPSKKXCUc0R1NQStQkx
l6g1Jh3eDL5Ohm97r/VjrV6TiShBSU/aw7dCOLnN5N2GGGdrs+Mn+sxN8TaeJTIUZS9WvewCiBqh
CpnhPihm4PWaArT5NWVYs9t0vJy0QrTYUGC2lk2C4V+7CsDImYzkaPlGZFkYgAdpyc9HhRsOREeh
H0Z8+ZRUjwzpFaQF8Kc+7n8odSOx2wgr3oIqhSbkyEY86QjyhxOCJMNLcRESqqXontgmugwoIRaT
PXBjhkt5qTU/8Jb53y1288sDiCQLbF8caJDFmRohSMMV6DPeFsS1v74O9vyH+7AwTge6DfdGwgAI
gG3ZMafi2BMQkL7/8E8gedAXMxi8UPw+vo0PpZ5CRQ/aUridl1MDZU7EkliD7vloK4xVCgwApWFo
J2J7GQ5QFztbalnqgXDe1CQihtpKfsTre428pjYKYUZK7tFrlOV+q5MFCmS5NNdQlUwb4lOmBZb4
LYhsEFpdTYCPBAukM4yHcSMJapIQK7DvoeHGSwSx1G575SN7ER+3Icz+V85acVWtqlZU/uBr6Q/U
ipDuIwgNyN8yDuH3WOITILG1lhspRokx6RS4RtlY6cttYq8Avouvxn+yW6echJnneILKcMdNQy7u
M6mLUUDDDn68YIYFg2BllZC1h+Qy9XpUDGO2+E5ndaAyXviui3tyN42rUX0Yy+7/qb0kDEItFV75
DOwErl+CHD8D/JIdEF/K59YwS0XbUj/RYWYwgGwi07pcm+SLlmed9dqpkZU+F/6r7Fp6g9oz5o6L
+/1WKPBBPPepSpSmw1rsNQCGaf5T1hrhzD1HxAPzBhtH6xs5pCM+x+K9g11JiQNWbof/eNj+CYOb
s2CQbY0olkHLPQ/3wL3bA93Q9+wnyRTws5ei9LrRwEDcjYslphL9zKk84qacbBFDgtAg9m7OeGs6
8xj3M63qX3EcYHO+i2apCNrucG2f7IhjXz6lfvkumktjE5q8ufb3j+opOdzs53oSIaVv1EdsJaxr
/lbr3orkJmcAmaXvt4hV1Cc4GSydBKpMm2K7VGZSVHFVbPE0FQVq2uURxEtY1zEqkW4MgI+24PPK
hoixEdeM1cTtMxrsXrN4s9ku68I1EX5kl+i+6mxioDEdbt7rB9DAhEniJtXhesA1KowEoG0Nx+we
UNfhgV2glkfaBc5rqZl6zynKFdXMmsWNjXEWAvb3Ot3MDd7ZqFwRU9N56jmz8Z3cyn+JEZt+31oG
j72s4eMZamp3xLTr1IodvhL5a8fNlYnfDDWanJ4FmU8SuGdjLR8b2UpxGDd5BDVfazuAGPUNh1rz
apMgvcl6gj43uanughXWhuJOn7pSP+ZOYQ5XfGgRmLwymL4bT1AUPTzlvtLYKq/JN+tC91Ir8rbO
iIyrUM01d2vU4//wC8BJPX93wyzd+digLjPMS58u7o8DxxFduhGGfSbhA2qJbacAeUSe243V+1k7
GK4SLgHBxCKKbLLGjY/3HZa6l4IZa00jMXZYHVpHbyZmi3jlyWQ0m38inXVKBndFVggMXEZ4SYh6
hk96dOilvf30Nm0OwHDllOvmnZJpnRBKozQMhuBYZFakhc1XuuhPrEzGMFvKoA446IGB4pvP6JHI
WpzW7WT7USA62jUqFBJ7GD+BDKRwwnoR1Z/iZalVSQbC3c9k/uhPniORXGRXJdT725dqLn0Bf/3w
hghpl4aiZVuXwg+s0UGpwf8ulZltJyu28Cswv9fuoWKqHjbp9i22J7kHHgpyR5cR1NP66tXxC2pU
ldWNeRZDKTGDDLitucC9afxWNi6J2d0DlH5ShYUtbJ4Y+yy99PKQy0+TnjEaBw0KEgyQtVwAU7Ah
blMifi+7+k8ZyVyyh8PM1kD6rBMa407mjliC8TtEUgIfpBw8uWXEOkNPos7Y6kbaCP5w5Jj3MWjz
Noc7Q1slo2i1vzb/rnGyMFaxwavJ9e08o1DT42wgkg+QweJIDM6HgTfqzl/xglv0VWP6upErE17O
7mHsx6kjkNrB9TyL2B7JmdhRD5IL1ggRBciHnkwBiEANOI1B0enc9opHE4BAznriIfxjscgXvW+w
2wotsxRZ/YpEk9kWKsonf243a/6xg9hvgY6vCdoAhF9gKqirwtGXEb2qS1NYQav4ZTh3PEq+oyfa
jcdDAtwMxi/I7c8NRsiS2VBIFZeoURdUlCbR59tPTp8aB85aGN71QcALP3pur8nt9zYnGfjlO1kR
fVhaX2qwdi2qto+I9w9+htM6VbgvbwtV0ejEbiA1CTWvK3QAJaPRAckH6uWA3em3CK7lmYd2yPYB
jK8I6fZAjlPYCYXq/UYYyVPLrW/vmHi8ezSwtnS83tNZ7gUDMkEs2PmStZDm/be/5R8jzudJ3+nB
CBzlCQu9UFovE2u4SevS6s64vO83ZAQO7hZSeovYnH7kN1WrBpCE9jCYux5j1J0YrISNCaQxDt31
uTdN55IMnIx5p8XQj9J4hx0ykwmB8dqCMYOhsVOMUVmt/Btd6p1KGvLBOTnnBqox7Co4eFBuFWd8
NQRqr4UrLm4ZSX3FLb+SHCl3ciV1eDPCLondyIBuC4/dH4bc8OkGXGY6Z+7ek428jsQBYD49H7jy
Q+FJq7RgXa4GEXt5Ph0j3iLOvw9/cotW1UIajmw739b5iaw7ZrHbtc3nzZqMxa66zQgf84pLMFwt
SLlomhIGtATutn05v1xMxyA88F5WHp3aLBB7OZTwMdXIEv7+0mC1ZPS15Ji0ucjWzM93/9fP1td4
3muiPTXRDj0v3cYMsgyj5oAD840HsXh1mNI9PbCzGlN4dT0YnCgvRP4NQy0VlXJ91ZJ3IFruGeCd
3TZDp4f0ocD+uaNugQb6yCoQ758fXyRfiT4QH8l+PTq0N1m3G/waxjYqvHrpPMEWOw7DtvJgjwW+
pZACdiu5cLoM/qsZRePBOELRhsvpkb5kMfUMtDyxtQr4I0KQK2x+GfggDaT9fm37FHrYNUUpKEYl
8RwX+RwVnHAjkjdSmnLpMGaRgmapr7OD6DJV/Xhd3p8WFltdPCCS5nO10MZuccgqNH42nc5JUxWj
S3t+xsLFOuvVmHAxNNz3bs8vp2ICORu0YxnQNy4iRwltGV/l4u1k63GPkyHUHDYyEKg7r7XLtTwa
94KwKAetBJtx/rrSoYC/ZzyVaUr2clWvoB8lHJijNHoqRx4GpbVdFuNDV8HM+oCklYtbhTjSyMWg
e1htlMLRBf+EVkvxByXKw2PTNj8xVcAUrjV/EtJ1+gcWE3sAxOxPqVlx5ZPlkRUExNV2hx85fvzS
Ytewm/EvdLt8WQhQ38oJ/osBM6jB6LIBuPtFuH7nF4ENhPeommppHFLS53iqSqKVW6btnRg9hXqe
Nx/NhjnXe0O8Gy4fdHAKm/uywm2bRQy3BD1KsPAg7j+yETpbHTCKmcxRdKziMJO1TN2f+VrX5DQL
62ZSqKGRGT+abB+fOYZWD8bZLMqDm70/oicRPbXFkIcIa0OhBAdYwqzzXehYAoTKJ6R8hHt+hHi5
Z7cxUhRbh8Mt+dTkQ/UK7SBE/b0+cFwYrPh/0CK5RatVI4ywKN6fFN7d9VS1bvSH8fIJF6t1fmFR
WsvcNnTtSNnj2btcU7xEB2fbbS7FVx4mlfINIxxed3eptEWKuVBqbE6pzKmafIdUJVZakKPHHzj9
Zq1mbSJWfWwm/hiIpu5WZw/CYun0HcAVy5z/aGoWcf4CxpNsuSsCNS7cvPsklokkFOdSMuA8t/8A
r0NFxeTZAcSSDkhVGjiQJHjmK2EzvhXZAec1k6wZA/+w3ZRqm9AOQ+LFOec9xzkkMMpz/RJutJ05
yWYzNlmUMYMZzZwzKqln/YimK341slAohKh0oDOrdVMYtLo7j1q3IFnMBqWYIuqtG3iUs+J7cFkE
VYEQyLMYKkvdOUqVfoQA+Cydocm98Yg+y4UM7z5MuPMp3+0ku1f2WGuMkybc48UnWSHjLHk/cJ3e
HkrmIOHkhxy4t/CHaS0wlHsqS/hvC9KeunnGLJEEs+0sdJdiTesJ/MQHvqTPUPWcg2fWd4kg9g7U
NA7nHg6mNKwmKRL+KbdsYPdcQDaotnhwkruQWv6NIEFt27YnJKYpBxRQdB/PY0HRxMSekcBsnvLM
Gl6IYWoYbuKE+FrOtuadYnkl99kdAFTQzDPijZI2lCPccR7hazXmgLiFVHNVupPJOUwLOeH3Wp0m
ckSZAVSG6N8+xCaK4JBba/kePyHcLYGw+Hr+YAi8JNmG3WoI0z9jTI+xupPiBdPbSNSsSzsgRK3A
u7p3NiXonIGHJr2cMnDIHko+vkEikvR1ct1g8/4Ek89NcyiL6orZgBpK8JRzfhF7zCb+3F+JVO82
itKykgsdcLQypLjWK9A5X2xeTdcK8y57eXoBEsS+rNFKVLK/76NqQzP9bsFIHVuNx0lMYLz88SmW
VE0vRMKRb0ZwdRSqbndBLm34GYnv76MB0Vm5YEYw+zPFqeoWM6CWIjkjOaf7VLnNEJe10de9wF7s
0lcDrjIYMaQe8/HuDoousDHDEGZTgSrAQOwZAdaZiQK4RDDnOw3zwuHcryPaON3HTiQWx0kmRA4/
iRrWddo9V9IFgOQQsRxwm8TBJfsfTJ+/oFPCxA81Gqw/OxUuYhxaWZJvtzCt2GDoz7ahzhZNFan3
A6spaVyo8io0ncz8klMJNINvKhmRuuOkglT6XNZ81EWO0GOzF0QQDbZQ6LcbMZ2dZa7try+7wgR0
nTkb5Dawgw1c+c/5j48JjhhD31fH8Sm26K0KAslf1awD5nuysSpjF19stlmwy5Y1f0/4tXKpY8ZK
LFCJy43nI0PAwex88NgSQ9E1KFvSg3DW7A7fMqKGX/ZdE44QqfrRn/Mj6BaLRdei5H3RZquyS+f1
mGVs1C4/VG6RfbUbrKl+0P3Sbfg47PZQ7FCNn80BPj11RlgpY+6LEH//mqK4XYnTz7pcm4DmPGz8
yZjkRM95+iudbYR7EYp3AsK3XpUKmYWXdrDrF7F2K4Cuo1VxLDWzrUeEzhePRB+WISvL5orJCqGk
C4wxjMg8ZuRnDXROMVbDn+RcmaymAPN5kZcZhvLqNBYFj5Q6/OxUX9MP5mHakzu3Y2LwAXwOL365
pEn33SyiFet6k7dRyxylMuuO6YYVq3avxoa2WKMQpGiREdltRXsGRH0xtEG8NaRE2dqmKxIa8980
3R1eKzFyEIsnMnCowIgvu16qL7JEpw3VYkJZgl2/UG/99exkdPhbzRkE6ntTwPF84EANSl/Zqb22
7JX2E66u+UKpmV2r6EUPxrqQDMFZKzCtj5wgsEUNOIZSGY4Sf+HXBvqWDTjARsNVNU8crZSuPjBz
ImtbnnM3T1Q1xKlYOUJhEcI4SMT0UFSQCDUMdr4CvHgGXx7hEEcs2yqowvJBk351FwDaSH85UGxm
IPA5Vxnsk19Cw/GPawXJBfb5T2/MtLuprADKEq/VRI2SUcmY/HM0Wg+oT8fQfJd51/NaKEzVbH4H
erxkdVmfaW3meMWGRFg8BC6Ku+cbHA2PKyyQmiCXUa0e1zJ+My9ZfB02pG3K2S5FVT/YzkWO0zVR
K9Y5mO6Ae3hkO82lMottHvBHRbTiaGC38ezaKHXOb8yfEtRVDGs99hGgnnGKJ54MZZt1dQ07Bw6v
554pSqozf7hnkbrqRAFDaZDWo0RDRgAX/EQv5w1JDH79RmzqyFY5bSYAYDTaHfRRa15c4JpRoieV
hEXE3C0ybOu6NBE8ANe2MrA4qsjUVp9+ng2IYSATDY3TnfPX09kPTH8GNpqEDVnjHom5rHSOo8df
ZAvPqJlhiBucCmyUcm2N/Wzm5XIo++RDbigLb6H0hKaSpZBDOzqvsFGit+Pl3JjSyZUwtBKtyxdk
yGGzsqp3+qvl11Pwm6tDlxdo5QXAPjoIynoIlUgcgE4F83mc2UpFs4c5H55dMuIxs6GuN/RWFezj
s/n1xMIDTeBlNMbLx1N6kV71p1+gPYYTvF8Co3YtH4ofd4Y7e+tLMVjbq6+n7butf6tuFuHSU3sg
OUnM0DUchsByHjmNLTp8Pizg2xDG3NZ/BS+CK4gOf3kBE2m6Zm1vIMZTb9dwAy7+7SFPCELmm5Xe
kwwple0dq+4G16tonsCS3xuGZx1ANk/Iwrh/P2k8h59KkLsj/DDrkGrTgyRarpOWXOmaQYh3FGvl
8ROxV2P1mRJm4USqXndIYeclhu84nZxmsTw01K10yZcGrP7pV7UeRrDZS03BhnhICf27i0c9g/tf
NckTb9NInew6XnK2nPA2C9Vpjo4BJKPgJdmbOLKE28jc+iis5+o5xwjlUqpuxuexS7JTiUNbQexN
kPUwSBcZyxwhZUTs509I34s1I/15Wpb5e1Ku54J5BxDXIVbDTE+i05Ba3PZO3Hh3I1RcYWNZFD/k
fyrUuhFZ9P4/f/XeeF9c8P/prvWAvBhD9h3AxCt7+x6GKehgzjaNgLNmzsvyB2ZYE2JxtThysE70
wIBydp8LhXUwqC7mEcdhOU4gpaDl51XmPZhsKgIqib2nDv4R5AANpHrVNRrgpnX1hSVqPsLbS/Aw
D5lkk+HqcbcVjVkeER1SJoSll0uWYhV16tHf5uqgyQTFEKlsODlYKkgdyzuBpRgrNM7Wy99Fq1sK
fLpPMIvk2KGeZAzFqkLP9FBcx98X5Px4QSL27qAHa2c0NHuh0qEauNselq1Xj3M3kStGckYilQLh
oXzlIJpRe6vxpf0Q9KomfKP32gVstOXbpmqIMi/+58dvPDyZ1/o7pgP3hGUihwFzjWJrlJ7HlpXO
4gH0cM9rFzjZ6VYvpBiD0nIlA6tteCeE5ejS6EohJ+yPPtOVUkt2+lG9Uho/7TzpR5aazYlUbvDA
mV7k0hc12MiegNgobc/m0in5EA4TlCAwEC96r9iv7SHfljauRvpmJLBxkCw1redoR2+5z/f7D8yy
ZqDcRJMSVMItl3V/IR6gMvG410lm4ZKN96YJRTdmJcBYWtvLe4m88dQRDsEK2N/VXZ2g+DODyt6t
XQQXrDuCxUGmMGM7iuS/pOpD4PeZfCxPlrNsAFTqDlbFQhCEJP0gB0/Dlp695tucq+xQwdB6l1+d
dO47NU5pRVuWEvRzJtCe9bKoVdnlIHQdsrBK/QFDPoeVpvwUAFFvy++uHqgLIHfW8wLJ7VNdgS21
iMh1HrrfvWCVLc6UVKkhz9ya/dEGkkTqy+c7otUi/Eb4fYwCY64bpAB7E8pDolUURUghBA/okorI
SmieL6phuoleUwAkBro0frajgSorJvlLOCrEIzDyseG19G0U2RvibUT9sWvF6ISuNYIWF9qN/KyU
gpoYZIUDixOmworClWTrqT0DEE3EKNdNPROUT4uaguA1g9mcGmsEa8b/Vq1cT6rBKbx4k5RLj8lT
G0fN/hDWp77kbENW3aad+IspqqeespFWyKvED54TN//jbty53TYL9objexkvawMJxC81EUytS344
oZI7n/ajdeHMsGFKCnkTTPmwEnrURNEbI2U/mvx8CnJt0m0oecKJ3CfctQTXJOAT4ahq51WoqbiJ
7qhIeg95iNfDMpTfNGI+BlE3M0dhJ7WgANISvN1RiFAjgwFRoKcqT1xRy2ecYrm9scP6d6r8vZ1Q
mcO8odhdH1gELHXkj9oDZHHf6pdNCwoRFu4PWi8q/M6F5sdY4BmDq4PZkcjluYkLsD2ybnNkEvbe
pNOsCswrwMCDU7PLDPuKgwvFeudB1I+1GnhkXzx43003MipCoHrppJ1GCAkhkPAc2eXANeYHX/Xm
NxAbtO0BXFhdk2Kbl8HnIvFTA+v1bsBv6NZRCBEqpvxXHeWbu3FfTOU5j5lextDm5pncrs6Y7UkB
PZIhskAoE0CCD7Xcgk17pmhE8UDT118oczuweLBkZoE3Z8qP+vpMgENwNINCXigibQ5cmXlcIBEw
z03o2ZfK2z2ZClKoRRMdrqzJZGqQJ/bV3TNqQodROVE2izM9u5WiO/raINU3lgOg+oOFnVgVM3Ip
s4//tPK6bou2KBBFfK6gJtwPNtq/DwmeS4FyIio4GDzYIwHXCuYnRYeT836BzG0qd2JWZhpsitJf
Mop0/Wkmnb2UDdpGgzR8yZRTgIodwcHz6YhY3r9PwrW1x6HtyvEPchprZgmLnCXAhnkmwfAFkVQC
E+BQXYW1XoShjZYzyumvrhtcT85x/eJxHpLoBrmhNDB6ZwasECXiSIS5iWOj9DdKugKZRMdvzXNs
9R73hskc/DTO6TwlJix7RZkpFkW2CW9CxE48eCevifXTn99gZOOJmcS2+L4cVx46RP3u0aJP3x1C
kywG6MDhipZRo3Z3jtyKLQEPdwqWi1IXhAyhye+/Hd43Oh51TDzOK3d0eGMbqat16FuzjHHZmmwD
s0jrzOFUfnypHSGluz7lvXhHyr1m2PywLiiMI6GcOpgJnJ2xAWJpxdvU+uLwCEOhoKJ7p2aS6trC
E3j397VibhV7Ye2rOEMvioX5lrwmnW8DalIBE6NWAsds/JvV3+Aew5WF40nTi07prSWRzVxDJEMj
2MC4vpAvzBU+dDj/jPtNWsjD2EZWcJQPPc+UzIxEjFpvHQodtVswiitX1VSsRcyobjaQ3NAaITml
XWfF/RauUSPuxEjdfBlWN12CNvKHcJwPOle6lVlb29t7OHvRDlNR/b9c3fSK/ExLIMO8SU/KLiAr
+A1RYj1X5zT3Bn7Fktf7Iq6LF75jL8Zlgcm1Rlp3uPH9+W9Fau6SgLQdfeY0oAMAdZXAlZR/hx0o
VcorJZhJuGnonjJsSRPZRXrqppCI/2FjUEBSuug35NLBH3x4/SL3afQqzxnQSLaUMrDkDqzqC8vw
pYz5dTxWtAdhQPkwZuo8vN7XSYJhFHDrVnc+iRG6+8m5MqhH26sjXbOJaZuBmsp6MS0N9Of4bbB4
K8u4XD1iRX8kuaLPfwTl2ywksn+hcl7DM9gwT0S2HqbNQRqN8fz3wjl49efaPJqYPmVnbjWNbQF7
Y6kd+nHduis7K0+19X7tbL0Ige4EG+2LfTo/U+1okHS53cY7hiaLUQpVgixzzfs4Da230K+yForo
iDMGw+VMpKzq1hFJVfC6q8WTExLuYxxcbMrhOZQaq0GIV3TGnGW7/FnVOIwkG1wF4nY8wRxniDAA
xml3hMRXlqCBS8oeIKpgEEBGuNyw+u7urdEmLVKBBq991tix9rGP10g6xlfxSe3EGoLC8cgE+gWR
ra5l5/Yve1v85rfkyw+rYavii5B8fhV3kNVCYFTNRqUjdtDG/bKb84pumz3RYUhBbiQwvZpUInYj
thNWOzmXwvB1iGTJR5u40FzS/CkTxAjwQwmE8plPB3dw9xf52jqzOaq0HVhc9UaGVV/UgmW8EJeP
pdhsb+y2siHYo6Ug/PrPJsXhDx96cwaWutHY5bT3/gKaZ54+92RnnYYeTRsZ7OvxXbjN/I3gg0bw
jzTL5ugUDR9OTi/FE6taiCLi36J/Y916tByz5oBwN44M3EKNjyV5e8T5JMK2eeS8SQu2QqjYDWNf
YNDjE1G3oEiNSBKh3vAqK+Eg7sMG/dhmuRo1asCbDvN4EwUT/Qt+DKJGPajc4cWVtw81RbBEvu6W
avTPHmPTQ/W/6udUC9Yq4RypYnnQ6GsdUf5wE1CLj4fUrv4iAc4F2WBjs4ARWB27kL/Cs+eSSB0K
f95fxTFu3gGc2URmopD9lbeCMa/dYiCI3qOogYBonAoxTGYjf9ZPqM0rb1+62jrz+xkBVopk7dQA
7n04iPpS0k83yuWD8OWJbvs3dP+7hk3W5PK02XydZh/nJ1UL8vbF8UNM9RnozXZ/cNUR/ekSWgzw
JAeuPWXdArSFqqX3rComL1HtkYgK4Xs6eSMliebokmxGBag1SUwjTBlI1/Lbh46broqUbvRoz0E0
1NjroIFqV44Yh3dFqpZit40EdG5CcgwBuwMEwl01VUTJnBxBsaAjHi91IOm2yD8xprUWm4tbuy/0
qGN+0QSiFyLwQzubHoPFy2Qlvf/dJDbgBHBxmKSD/4RhteI0q/JJKqyUd905Ccq3hsYrflLOJ0T3
zwz0CBwmAvx5DDsaYw9H+SSTv92UxTAQKqKh1b4gk89pgT3pGBwvC2uuX2SUM1305Ko9IO2BgXv0
c1+ob6D7GoWjbjwWkei9HQpIgp4O5xCDMYU3zruAlOWEQA6iy431KZ7ERW+oRRRjoEdEShrNmtDv
ZzpTZhsgRuHN1jV0/nj4F1wKM7jhEBlds9hlai8BUpO9ysgA5sUShOk4jmXbLpFkHptLUw+5J/FJ
i59JW4sa4sHSC4Q0uVUCeFKl9qyAL4i1zjVE9B/CLpoO2oM6Tw0PtFfXr7wym1gcTbCe7zGoRtzW
ZvAtX1i26m7vCeYpGGvJmAiGagDDD/Icj1Jcqz7i8LY8jqqKpDboYKfxini2y0RkuW5ozRkNUXuU
MwMW2ZLh3JHgROxsS8Az52NxGzEZjpqOn4StfPH7UGN3UXRNeuN1QKjCm1CKRtCzY2DhLJJ92T3J
gmP3RQOLRcFhiGKOCbzyXavADiK/77e/xN0E3E1eiyNwb59m9eN0JZba26RfteBJ502K/xpPZtOV
vY7jul6qkIgQFqxGoj2cJWMd40b23/j+Z76shZ64OGI5wLVI/XTU2xIFJXCr3tVxBhp9indOWeF+
D5+Xp8mBvDIDArPHsql4J71HcCVCBgRF+o3DMUEDoM4VvxlXzGsld7/5FjpACICiscincx86ov4Q
AbvRI52zn1eU+t2CvUe+gt6Z4VTeK1NuMfKjQQwYpm5K2pV63B2nfcmzcx/aYrbnCYVsXuO1T2Kz
DEJEbGzyi5Tyb1zuzrABT5yozYO3fDRKJOJBDK9xfwnLk7z37kpbbe8y6zanZ5lLmz1maIqE2CD+
6DoNNieFL0brWHQopcNd5DKhJiWcOysCPh9uU7zW7DFTMQApyA/Jo8sCNlOd/aFhkY+DUg9aX2sw
taVDiHAKhwmqCvXYI9AQ9/7HPe2TJdjwePiIGyXUE5ELtu0UfQKzmu48xMLC/R1jHRZTxipzNB0X
qcpAJ+ozLIfoJ8qjY0Gdob0766e1z2XPC5fwTBoo7WB6skf7XS0HVyiH6ZY9PpUHJ5D6wAffROD6
YSOs0YlYNK1Sj7h0JTB72dAlk/O3u3yF1/J1H4axmPWGGPmS963ttmidAqLM/dkBIYW+X3nmUJRa
KrXo7YDyi1s6LeBuSrFs6eHiNs3CR/IF4Ekg9Gd2qAlT/4I5wOdHim7SmaJgzF1ZUU5TrSksX1QY
crlnfH46NNQtbKOr4RHqwZ9AG49iGRag2tmcrAcPd8Y4aEGvhbkZ+CtvKE8z/eOks06/mw8eCHp0
/IT7WCsDxYBHbatn1Q2T0OfChXLNgfeK14FcK+Dch8pHLA823RJZsE/Mf/S6YbLOfchkPiS9s89H
N10NWcG7hecaNBgUpqtN5xnYY4ipSzA0AUzI46xl5Sy/B8yUdPaZMJilt1wjTmkQTVB1QFdYUnT2
H4fn0Rop6LIeFmEwUOB6stupXd5Nul19bA0X7Tq56QReHucf6A0A+MLhInX9TX38eUwmw6H1jXVQ
vSP7BC5TDNXwl0EfHA95GQq9fLLk98pXOGn616z3YfJCv18HCXmDgo3Rcl6vLxCjZVOZsBgXRA6S
Is31LvLWvW21dbS1jHKaxwoZxlOJMd2vy3hVQKw1yrTJJz43oNWF7msNPzuv+EaN9KVUBnb2DLNS
fIavF0a7wLshMEaBdQqcsj0+2g1jaJCPU1slS+0ks41r+eGzAfpLlSKcNn6cfYvcsWrGLLCGEuaL
q9CMgOqDUYqDqan/dLmEGh/7yUgdLANzqWiKcGXqKDsomvX8T3kGv8h5W/2cc5WKbph1+KrvGf7D
uVhZ0rqNpwQgVofA7Zuy6xSr8Ejh7r7WBgoDukbg3IKcofp8Jb0+0zFjLSA3ldDLrvVDpaXU+pu6
DkGg1jYQDgHx7xPRO2thfXnw+VEtW2Rv2DMsn00mlptQg8PlYFtYD8y3FYiytXzQDRVyc7qkH7Qd
vsaGZfSb84qeJfqqVgLJ0QLlGhGLGYMuVHgvoYUEHUelQb6QW2ddrj3gwKX/6gbeiWlh4IhM/gk1
71pfKVEv7RxKTf0AYWOwpQSPkL8xVfJst2wjlzAUTCgCtighdqTHpwQcjxhS0iWEwbCzkkXReciT
Z9QA05OQcJBXnOn+ezqjtA4joI6XxoFLHWW/J1WcFHdrWYMWRdhDA2UIysVr06Oswau1pkLT8hy9
i4Jv/QOWl3pstDtiz8TS6wuLgDrQ4/1v8aFgstDV00Dg1l/oOPPGcawu5xEESeOpBba94agkCDWg
iFdSyCugDYlIHSwEaB2MPtO5cN3JRLraiFZOn6EJSLeM15fVMiaWH3iLK4o1NjI8InP3C/vcQ6P/
PF7W6vJy9vMx/52g4OPk6YGDC+pqbnIzUnqUcN34l0uMTNrHwD1gaHGWk8QJYisDDmKFwGVqKXbe
TQYQh9/D7jub9na6M3MLvNfdSovFJUwCKmCVWlwwIHNTYCu/I4ESaqtbYqfNJxUXsBrLumeFsjr9
2Kpyi3xZi70gXJGNn1l0usqV85LNOhbxGBDPoPIwBkewtEEGRSgv0ec2OIhNB4EEcTti0AA1Gymc
OQK/ZMOlcYcllpWVOp2Wc+wIAGHl4LXbr1LQc7ItyriT2dxe1/44gDc9V7xMEPsPo7wPUn+bDrWX
cSvq0yhMpPajjIhJwTCDQcv5LWL9mEtTcjZgTB+LIGiC5jvaJK1YY0RNj8jgWUZAZY2dSOQr8Rbk
XK9kOsGS3WSNXb5GTfXmGET4y+wV3hIG330UZzETxJCekvBbbk5U1/kRQwsuwqhMx5hfL5U0ywHh
EA0RpQIJqCr2/uJ6Ap6gJrgwCTi5hJDxqiLlFmKAnpM5ZJnKtMKaogUyI0cyWC/S0KfNkd+HQ/yx
c4CdTrCNHt83dKk/CfSPWkzyZfSFBUGTSC/z9CVqlFYe1RRAgVTh85hs5vptM3LnpKMtt1QSeurA
e34hOLyHSk8XzS6UxWyaDf6561MXcLDv4DcTyQq15D2sTIRbnUduY14EHTlw/ctWAFKLaJzmVNeW
9bCdqCHwLW/IeGRSUij1F+r7NJ28gNk6QAyc0R+Afh2cRDGD0obwjfUoRdmGp6QiF4xT+1knxVrk
Lh7vpj4BYvMfU7TAgjYY25zPCq4B3Z64cnt5Ww+VGXXrILBg2ijSkdYVDXF//3R1ofAoyMFTrDkJ
lMxCC+9whhICqNK+z8wE4UkUjtdTje48CcpKUGls1sIA8FwMMv29FQXgNgi1H2Z7MuaprT1f/Pz2
Xvqfhw7Bl+/rdpG3VlWvtrl/65UsYrciSd05N7cbXA2HUNDaLwd+rNEub92aMOEu3iuHQnWah8cv
P8cSlqvL5n5Ww46h3m+Diry01+7WDuN8T0pmFLwR8eH3EQKK5kUMGz4ZDj07N0nmrusYChhqybix
RvkUjB1Fj94mvoz4nOoVqg/JlFAK1Swx0bbTnt5OVs5/qAbCIyLjjZzBjVRTb/ilKMxmEmcmjCkS
sSsp0cUcgtcwcv7l6XMNiT5/DUdJnm2/HvjBuAO7D+bL7ANm/19+9m9A5Sc7WphlSE7Vusz3Nx8m
l3jrnjrlG+j0H4bJ3aY6y+0xQ9G9l+U0w2jvG7d+zIXDCY+gxfqMKbqwQKN9IQ6x3WSl6ac5cHRY
PCIH/bV6V+0u6n92Z8Fb3CqK1UPzat7O2dwFthJBzx5wCpy6cXAlVHKArnw0EuV00JXM0Q7IEdJD
NqVyCxEli8aqr22qNdujGTXBx1GHoyfLu3zzpc5zcSI4Krh7eOCwMnD51P3f4dfjw3XEr+G1p1TC
2V7ueNnBsEImsO+Q7WIWkzk86eSaK0bTi1kyVH/rWiebch15IiLC++3V0eF6dr/PUsTg1OWNwdcn
48cPzkbPmeQRRBMacKazUQAUmrWoJRlBCA595bbKBZS5XvXXaZOovZcYGjw6qEtjexmoW9fxMOxo
smPN1RAlyunMg4TqmKj5gwAcslhf17CFKpwykpT/TaIVBhFxH/fHXlGvK+OS4jNhlicPhRraCmE7
uZjFwQgyPPmp5ta1oBtkSHHMYDXivpuc8Rh+bECEardw408mtgWqmA17Pq0QcEkRjI+yb+yFaTDQ
Nw4+i0oEac2/pJhiHDYrd1wJ+nEVxynzxlZbB4Jwe6UgavZiFwP5WTDm3nA4PDgJotvrP/kNHZPC
DDUCLYkdcY2JuRbTGeUc05xZq0mBD4NBFqILPwm4F494RF9BrxbpV/NrMutePq2pVIhyZ9XFNpr3
TMu8TrUFQho+86zrA90MLLFPQ5DZOMYQQnM2mxgOhZ3Bt73knJ3qqijEWbP3yxnq69pQebeLVX/P
0vNGVzJT1XzRuxtX8BDDqgb19t1MAGLWr1gsOs9ZbRgE5Ep1XpnjjPFGiZiqX60VgpW9s5B4xIns
oYLrKV5peMuqUoPnlcaG5FTXF/jQQa9fuLWlLOtyF7DKZqQ50Izj3f9iK/1MMH2MfwJn6E11Vpcs
eu4koaD+Sw3ZBWTqVoDiw1h/tbkb0nJ3mTy3w3ntILPH6SfNJw3ngDyIb4b3kdNkhwchj7GlKXyV
ZzRbxTIhNHaZVTiX/1G5eNZ6O98UNg4wQSE5gmUS//6pWfCTlaS5TYhNWnNs9iSTD+qSv+Rcld6d
zUSq44dZpH7lnkU2/t43Oqkj08SSbsyukocJ4MvfmbE6IApuzsnZr2t/sOPRyeu+wROoe58BGbaJ
Wp0Xrlm1NNMsafLuEbdqHNQaznb4TFUrO2QycSWQV0l/7clx0cMKmEVOD/1X9XcsLvClPpLws8l2
od0bPthTBSeO3EjH46DLTTs8Z1fP1EvU2VFPwdHG9Uwxu6mqDvTekWCjOafWXHkEQILntEK5X0CU
hhAsNHS6h1Z5u4JVq2jgdRfCNzX0RKoH/1llInLgarTq7je6/fWE9i7C9o15dSSKrBD1YNZYyw2i
ZXSZft/ODsk8nHZXVWuthg45F2p17GL+UJQxs9+6MlC8H0viChY3icQYZYYxDcrsehpO2niVgJz0
Kxq95FUvKXpIpAvvtComKgFQ++KFZcYoOoz796UVKV2sQUH0G9+n2egimLDfLCiMwa7ixGXaGB2a
rkOeNx/A2xBAYKW4XTXO/KGqYMNuojTyuZkyrBBkCCqOVSa7HNDwgsYLTvnjqCQzjtAZmHrdb96G
Ub1rT2LTBDQ9zlZ1yjCGhA0H3mjzTKCre/ksK4hOvp22EX4weYO09ZwXsw9jrtajzR8WCea3eWdE
ISCO8Knppnkfg+xig5Bg/bygu98JsxnuH6dhwMiEYHXjBk92bf06E9bodhChgR/8G9oBLQV4YFxa
N1Rsdva1EmxrY39JJuzFHqw19b5zOhyRPf3S0kysCp2I+MYvXFh/3NLh4OjZtjCdP43aM9yIstrO
FDnoussaqw+wIU0Iviof30sBbKuy7rXMogvru220XbQWul3suAIgJF2EfdZxY2n/BYUhYYCf2mjF
rWS4H61s+SoMv7Ov9ZG+mKf++iGTxH/JPIYJM5WP+I5UwXZ6A0FElpWeNON5fzF62mCp8Xi42Uqy
cwJmF5kEjCEFIabW+sqn2pZZikke+SUOAUC15LFH8CJN6lAB8zobUt3eo4xRzxLcUWifJs7jenEP
5jQl2I2iTfT6BfTRv27npgksPLo325z+BoaL2JnAq1gb2r5rkUf+mYxtWDr4eWUNpZ7CWYbgAo8b
hdqwUufdUVEJoTV2LuLC06qXtlSl7DfiUwS1tPviqU9lpw9OVc/UQO4lh+gQW6UI26NDiJm6pAT9
QemPjyhG86cQ11HxD8w0HZa8LdZjPCYEQzearx8zX/7KuhrsSWYZSZzHURlc2RhR1BfjveuA3svk
7AXxt9Yel9+zO8o1/njC7ItoihyTL2HI3iAP/6AfjTFKbMVaptCdzuqXhbBWLf3DsiIYaOX7V8Sz
goVdrEFGrkJ8aAcLSOkSPz+KGYlw5i1qbH0w+fRHzGv9pTKW4O+qOhSMdsF8CTvthjTRuU+s07Ru
L6tFrNtoXAvqsaOmZ+eB4kcNgepGRUXlY8ZKxka1YLlqVl6r4d2n/A0aaXzZZl3RsbUSmJJgTAc0
Vu9Qfy9b88KqrBcfvu4M6Hw5pV4VB5D4U/0ujMpQKVzGnXMF9FiGaxdpfBJxxgyVFMsS6kzl6+3L
Tg74Cp6Zj+1MVAlFy8gNFdeleO/MdkM9hDc5739TT5EBYBVGFwmh9QyECI18Vka6745jtUjQLOhw
ERLbyznExT48ngwEm+KwzM5Wob3r2VGEFOGWqTEgxUOcaqzFm9xwSBiuA+KANt9fZHFUWNX48pkA
A+pXsRrHNrhqZwd2AkRYhNxCENKQ5ZVIdtk1Ob+Nhrlae9j+4X8ZBapp4h/SQ0QMD87bUE9wqKUQ
qEREJnL2DbeIlL6+ShE96q7RHjT0esUf7pqUftrJXXCwBM7mPe63dS+h4vHaE7gexAtZ3PgFdtaE
Pj0S8PZfHib+nJd/r2GVvJIJM2BwrVmtNxASKKgf2gnfH+7nFEJ9lryaXIlA94/vhHdSVML/CTwd
ISeWxAuwjiafrhDRda2ZW5swDtSHBB3QdFcP4hlkpmLZUBlVy3qDwzt8uyy4kG3EU5FyxpqR8xPX
aNzFIhIDhLZFq+0ue8sciyDX2u/AeYpvtfDADvHOgOXFcWArbCeqPKiekmj4Zesd/aJAyUM5gnHP
fOxerwnBUlV2hY4wuaxuwN4i0R5o7YjDEzx7FWhcov71QtkwVyyP59THsz5bBqLXnH1AiubWHtFF
Nv5LNRwkxO/dsqX1LjcX9v5vaTOFtNr1i4hvSXYF1GKJISNYHOuGuGv5yUhOgfDkSfgmXsXkbk0T
Lfexg7C/IzC1AEsOw8ARsOuusCjMbzaar8PTGlu53BmSZP9AjhXfg3/wruSVVkrxkQ3sPbupqTfV
1lN+spIyW/6F+MU3Get6Gyzm1HZePgLmOkXW0D70cOg8+0eIaLvKaXvaTip+vKIY+6sKvNEhGSN1
evY2TTPECpbhqYV9hbsfysEMXH4pg2eAY3xyx13W3fDV4JR745OGVVBWVu7P2uju69CkTIP/KqUG
/ZET24FuzNzPdRB9Qn3r9w2L0AwBsbjcPAnh+eUUVkqwW9L6mxhwQ0u6iC80JtMy1v5iTNs5RDlB
etC2yls37A5EuuWuyZI+he/FMSA4T+7ZuqLzZd6XpDcr04M453kdrHQkzQyrHEwZeqb3Z30lmmDa
jPkPNyVcpaoIVXufUAhBXkWCIPrwl1GHw3hPmuUjFZ9MMym5ztaHDXsV1jeVW8KnEjjX8mFe1SHc
nXlzF8FnVIHDBDii0tMN8PuyU3hnmekvL/etlPU8hw0DMsR8LpPqD91zV4oan44Wqyuu7IEndMVO
W6niC38hgFGeWaubPK0WAXaCpsii6TURB9ihYl+2i02hK8L7t3vxL/XFI6eSx63A0v3Jc6/k7a7p
ENBQN7SO+juLwXElzf3HicfSPeKPpFrqjQSZDnFf7ZqzGBou3dLKOGMSTxwoc4tWcW1dGVsd7SWL
LOdfma21te6LIah8GYaZU5MilmGiE+bs4jG/TyqmAMrNKdMDen/0GAJA8zK+BAx2SuMYcCm1HzyZ
Qd9TZPpnWtbC2TbxvulD0yEL1rdhDsX7ro3aYftdp2zE/qsG1VXt4N58Bgt2Omjlu3OkgzF6QmB+
3ovnYBvvONeJhLbbwCNRb0ulO4eKH23KMOWmgHofXUT/2Ngxg98e9xEYmVQ0LS23xX5qTAqlqdVH
2mbtUKhUchmRrsqKMX5kK351H9NW26VNtaY5I105rJ1zweS+wEV/ltmUiiigXHerPPKONFQ14x+R
PNJKcV28UBXyp5Ad3PG1v7f/6ZHGL/2YqI583I0kWurFpbGYqRBwHyHSwEfl/1zv72sCRSokwnJ+
ehNYtdQMEOZ4dd8ADL/jWUJqNKIXZueMJY/qmyeOUbn/ZQes2xXdBqz4ahuK0gQjzdSSaivZqJ2k
ZaEE600F1bmRCt5Ge3RpABk5tA+f8NQbhYqTcOR63KZP+bBNUkbuzrOVNCFcYK1nzOHBrUCtMddl
Y3lJckC5lcaMsgBb6IBFNra3Lzp0KJaz63whd/8I4KVknM7ZKErCchA4L+SrIuDAuLAx77YaV+KY
NodpbUMAzo1rnG3VPddKY3UAYHcnBbs1WppBEQ6vBrqN4ZxZZ6iZ37b6/lMZyK8oDK/h6bIpSkk8
axA4JznSHbxcNvNCbIv/k5E2pyqdUeStW3EEVIIxGVFu6VpC12Mwv/F72USyJ0zqqPVnlYfRhRcw
7cmjztDe6mAJGaCwWFpG3M5+wjkVzLy1PRaOXgXNCgV/nQDskn/bQwgV48obI4TMVrkJq9Cz8cMX
PJayPWd4/hdpfjBPDp4Y0axkNNnlL2rNvmMkmRoyotZEcSE91tAAmNdo9zZu/RoiyxcvZ+BJahDW
AiaBS4jSexCaThgwLh7CUv3F78leNJIVnxcilNBoeR67Oip6nq8evJZefVmrp/46i6LJxkJHgV74
tUmQmd+cXzNKgeSqIiXFzTOW5Xit4IdzIku00UJh1AYZX007NrShWF30bDY8nWIvcpJokf6rlAZq
wQamw2+eJx0qpM1DuKH3yYjFMDarI9EWvmlxwzEKUoEx5X3j4kCin0UYz0kwNoblQjO0My13MjCU
+ENsSjH45aPy9pq3RU1bYcPj/+G4wJ5jp2vmYWKn0Jc2v9lFxyp1ejPvAA6myKESKDRcFfV0z1Kr
mP4LSg22a6OHV4F45nvlnw1Iy6ecPUoUsNMMkpnGR3oYf4LP5FldEQW3tCs7KcdIkEtwvAdd+2DY
eInuU29YecBO4AdFs/wpAHRt+fgUdDIjWisuekP1GokJbTCQtcrdyFPZVRUjD8fj/DiykfnrCYjN
sSScAe9TlJl8r9hs/eAbWMJM8wMq4bU3OxagcPHOZukj9nSPTNM/uv8t0SjACn4UVfIwiE+JVAov
5npIvruUmdGbVdVEzDO8q/uPShLLX/sHN2JPkU0GjBhiAehYEHK61KPTiLNZpdW9WUmqQ4Vp4xF+
9c+WNsSRkeQLYKiw4IDPU2Q/jhy3yMi6yN/9Ogqj9mc6c77Ylw1aOPJzh+BEBgJ/LHQeKuEw1oVi
yvZd1s8XHwHKTUepA1j+zy2rQHLI7CVRLHB58oWUdG16WLKLSJH83CKr4snKLfQ66Kpo3IYFcVvz
spQgl2TCnV1z412OGbKFGTMeVYfNIWUtogPgOTH8vB44NpZk23zd6og23t91sdoVejEVPy+bGJsW
TfbjkFD8CIQslEyO9rapHMjVO7OHxkXmtoMVkxJ91dSiunTCuaUMYPUls+LaiAG80qVDqwURDfB1
GhmVAjOb22p1fPFPnzwpysNLVNG34rpgWMwBxRRQrI+x/xpGXXyP1MLJlT+pC2fkXlwiFuTSu0Vy
RHz3Ho58UJygcotEqtranHYO8vbdYrkFcZSzEppXfK3Ae8qd0jlKAp79oW3/svaXSK7ceV0zXzMF
QXLtcXrHrB4K17Kbr+mut4lbRYw1q30OlQaGMkisgUR+4tJmllKuVTD8czUzKTKQcdE92OOBexQg
nBWarI8u4+0L5m2I1VMXPhRwrFuwz6i/MhWQxHnzkTPIWBQ+G0Nnyk1UBkZ6vXPRmVr0ZfQ8xJy0
k6r71CcEF+bUkOk7xo6YHXr75JLtX4NpKZ+lOdLU0nkGndbFmTVfrvvCw1u6mXaOXSSaD+45xQXN
FA5N7Z0Qp+ifHTGwsNKWlN3xM+nVuwFBeaOUsZko2jl7WRc5dXYKPqVQi6MBDtk7ABnOUqKo+Oc0
oSkgZ58ZGfj+Owec3NEl5+X7wzMALytpX92Kg9QajoB1L1aJm9CSDxmdaRR6W3ruIENHFqjHT6dB
CZkyfmIrVCoRgGUEkKBo1dLO/L8wILOh7MzuVjv9WKLj9QHI3Z/BNiO979dsgP9ccnosp8kp6ocX
w1TY3R5JKyEm2VLwq1tFW+cFAzrwkon7H+P9zphFj4xnUlBCTsYSkregdjEWwcUKJGiM+B44FK82
R4zxRR3KqOVRrV++Jd7jf3xerwv8KjAQB/Uc+j00SGBVw4I14AFXFZO81v6z2eVk24AhyZdNcQ2V
U7JsLxlj4kjjQ/uW4kuo63hrIz05KReiLU88CyqQewksVXXrTteVS4D9O3mEebk5pB1uIVpd3lHF
NIt5P4i+YfmUc+/CcbUJnFxgbAq7PgWOiM8CUIdAQxkGQMmDhg430SMqh/xYWo+IELNtff/PGKbu
usx5+P0UBA2zeVWXTnVKS5W4DvLNSJ475HJcw1QM1j4WxXPUjQC8xe1s0jQSUfiybj9EivJxRrLz
Ewbbq1JLiV5ydrSJ8Lqw4KD0eBx+cCrKHf95bXHKRVWT86Dk7bddlftgIzEwtSsJ5UMsM1NVghDA
XyBKIiIYgBD1MWgfj1e64Q2DKl6JK7CDDw5nzLHkQTrOrThW/xkxCzWi/r3G271wEyJ0Isj1EZS6
Xcv6bYULyOKxNnK0YJAC/iudlazA6f9Bxr6suna1U9uCfjs6a2nLcyFwsnRRFRaNwzSf95Svz2IY
ush6zA/M1w7jMAoq3Y04DgX1wDBS+MA2+08D31OJUgEMVFWiJvFXJQbE2LFdZcK6jGO/ErayUQVx
ecQzhSVLIYGixqAtYaKqba4QvSXFw489nbpVgWGfnE2dGqmwZSQVTHjRU7gRa7PzJ+a29f7U1E+A
hnxTEDl3Vyv1lvVm/eNViah6SZ6d/PJw2Qjnr8crQ4JXRFSmKrciyD/7e8vXh++dRYMCWrHGKUt7
tqFAvbByYRxQiKbuYQpm2/s2/AzzJla4l5NOFc6ZKTQsP70KpMKsMUH/fxOEayJOT+e+rkX1XHQ6
3KJvjfn/aFznMURkB8jDDU+fIUiNrQGAr9LbhjSXDfvQTPTHL5BAdyd051f1dfpluKDLoqm43bCU
IQXDuDdQJExgOiDpwW2Uy7ibx2iJDF/GH8mmDUSOgtFm4OVWLUXoK6W1K3jATGGoDKfW+Ro7bk/U
/MlHV850SwnvsKqphNTPjA0mQO1z8OF55+w1NCjlTp6Q5GAm62pe7kKJKFA59YlFWF7ys8eTTfWx
GfAvlYgnmWYVE2H+ebGtNEFwMjt0eWZZUiy+ZHHcaYycyCnpqdfv3e0qf88PRlb1Qhg09gYXHOUp
smMhKF0bQcdKywJy1qSVzD7oq9AM/wDVReIxic0dpn20+X1d4H75N4fPRJbOEqjxRyMy8JX/4nWW
G//5qh7RVQVZbX8/aN1p3bhhkaz00Dw/SnZVk+c4yNGHImffF/ef7K7Nmhkkr/SltwO0Qo3YNDVS
b+unx0hbrG0167eUasgs2xACdJdbX2E1XcFEXRxh2ZHicp5+QTC2O8cU/UiAWogX922XJmhaa3L5
d46K+gyaF239tEbrCifXYcvGIINWfWwg3P0VY9LX57/IclN0Iz1jaznaJuXS2erBShcWDb7xQq7p
8TWbIJfl2YIhjrjH2vEp/PvdgxAFvzXfvOfpPwc/gW1LRfdsu3WIk9gFG/o2OoI0hUU0djafWazG
rE2JFYQ07/Tzep4Q1eHIChwm/11AUy6ydhcfaxfhk85PMIuEw6Eu2J0lQJsQsyonSYorbSDKnZ1t
e4G3aX+GDyM6B0veAXbEC68wsgyiNquq7tyBK4xfxrRbHwlb0xwlJTNnY8uce+wMWIpMzYqdYpQh
TuQQ7IA9Po0AxQm6qwMSNvu4MH9qTT5TYR6OVkLpguoTMZxH8TOyritBqG4dRRhEses/tW0cXmoX
pSBMNKby/Goqy7smkF2qBUlTfhzPJO4kDQrCeaDldBzQZanJ6m8n9Zxkresm6q7ZLfQWyyPsoAdE
I+rG22ICHRQXUIx/F+uJunKmlr+Yt0XRPNRzLVBhApPdy9h2bW/Uc2l6V+2wtAVS7n0Qgi0sJ9Fv
aebIr3/E8hPIxgamQbORoMjD8jKY7GvdT18o0nLsxTPIQ6wXgaXWAb+Yo5rufLbSUwt8RGtWH2Pr
jLUDLGLuy6kUrdhduwU05aPPniRlRCs1djPtWAA15UYlMgFfTmAGSmXawLEOKzhmpRAFq8eLWTZD
jjD7x4NVCqsObhTjFg2ZDtY/Val8O4yFQytjH4OKkHdwd8xVbif9iVppXY+nYEMLy04Lox028rtW
ZTZ8w4/wS3zSBO/vvx1TOxiZCO6f1A7TwE2QO8vmfB6k2aYYw8qBT6n53C8MTr8LnkEa/jh0sflU
EhtLgvfCTjBGuHUbAdlH3/pVAYVRvrExZxGaF70T6bOk1bf7TNUQPnpZiyL790gJSU5JiFB/MD+a
LyfIrUQH5vmxwsEdkFtp73QExwBuT2e8hsTO4dWLli3cEfS5djuFpbGC/LzWpbtE82TBFeCPpP5F
yeKjI/fO2B5AZoUDsKjABUdk6K1z6oR3xEcVZsQJCEO8zgRYUZkWu09X04il0KyGUdZR0rtGJRc7
rJTnInGk+3hiAQXO+spCQjNov4yc4fOtf9nQ4OBmNn+CBXxZwWLXILH6CBi5QleOBn1KuUJ/FLDm
G3i000Ej9ME0VLUBSI3cmboJLRJL+SF+CHPD5y02npgyW9FMjhcMEy99OwtsGW/fux4W6SeMNcpP
TiJBML2x35VAHdRu6I+0Ba+gd/MGYqXWXkHLoUf14nbmtOHgXMIwUQOTPeuD0Ipoc/D3w2iJdHBF
qZMIgzvQsjl9X98yIqag9Ja6nNVmYGGejiojANooqPKL2BHW4SjYjZK0N7ztQR8by4dOcVWzBRiH
aWYu47WmCSfD7oSGE6VJBdUfLbE1pr7uf40YzhGUbArwIDNQRa5CIhAf96tMdQZADMv0Nznmu5Q4
O3PlpKdC1jcHguwWE82nEhqsur6enMHWxWCzBji9Ts4an9rhpL6PtarZlI0pm7VCKmAWavHXOOHh
lGy3xUaynJ9L/3UozaAl+SSL42yU+Mi7YM0Q8X3l8njXkMcK6s1Us1+iq2l0s9jMlfHI1S46ofv9
jJUV28ltxdb4tQemhjfhhds5maallHatDDh1VML/FHmk/Qmt46dIu97bzNuBjxujraZfJ6LT/pTh
CGXtUyO6senSwMVUkUQum6AnEOJj6DWLuBTMbuZLP5H+k9HPIvRhRrwYsVD0Ckw/QfV3OJsMqHeU
iIkL5tT/xEwcWKRiarMqwOFsMIgdIpqWGGlcNIZtoxPqrqn5NcH+nlnGiDhS4xh198Q2WqskHeID
d1KWjnO0KA2gE4oaLRSlWG/5p65T5/QxHvloY2TOFLlaaJIwlFNFce8PkH+hHhpCtL6g3GWtsJro
5trTbSlHIZXee/SEIq4iUgxVi4OAGpAFMVxsBfWwHs10Me43hIgKbigO4tjeuaFflRyamzkKnawG
qrcHnJmMrS9/wR1r9RlHbZ56wjjlQ6vhD4PdtnUp3cd2JeZC55Kp2y3npMUUoSG8k40eACD0nBPo
JkB0pI3PntzuTn5Nh08FjlIdqNiJwR9t5ImuVgjKZw6DjJGFojw4SYQOgSWO22x7nbA6ShhsJPQl
LnCfGxJnNKd0u8RNPzFGSxs4t+Xp6KFR6SiKr19vq8UmISsj7v/a95fQRj5m/igN/wrdvtsXk9px
Rog2zG86TQJb29TpoiZoPHySOPd1N3BoklBwE9Cx0T1puT4BMZQiIsy9M0eXm2qgugdpv1MWsEfr
HlkM/XhoWBnCqWGIMiKBey2lupV/AFJ0kxuNiHz9pHOqqkbhuITfFHOKmiGH1Hri5qQp6PuVmHAy
BO9mYyWiVN3Vw183QBODXbw4VrBgIgNPV8/D6ZT+rtl5Dapxcgikd3KTJTgVk0OtufWP+DLQ+9zw
nbYQs+0IjEthvTPHRbzWEolnn+zsjONRbZc0ImYa2cSyprunr1gxW80kvByMh6uGj5YYHDQViTcE
FzlmIee55/z1t5Hbfw5xh3Nnq27TiLkTYvsE5Re7FAQKsaQIeO0TFsUZ/YXO7/htagmS24CsFAUT
3PSP3SZVZN5VMvCtpR9Ce203KC7ZMJwQm+qKD4DQN8Kx7HRBhZBdQ1+ORS7Z7jeAm7P//7fjjNF+
EKdSZ5dMZSC6Hq2Kmv0QigvQzUXaw9yHjRcIgCiTVfy3wACpWlbdohF0rQKIwBoK0BYjOMDsB0ic
hRt6NM5uYIvvdj23Euqe5kXUiEMczN3J7nVebcdmPaaO4URUDlmNCRpT39V4KdhvUJCKB9cyUe8k
IvgyjnXikYntXo8bf7VSLksMkMjBTzVkXS2cIDnuxC0MIWanFqAXBg0Nl9XPSwmDG++zGQO5EVJx
mezaNsc+i1wLwqgkz+vkbizBjDmeGgsVXoBhv/47pWJNvDwWSE94GuVE9OE4ryythj8kaQidGsmO
N5BTRfHCSsJvjkrdVci6//a/HL8l1JNtK41G3W95c/Y4G200Iv9vPte1AarxTPs8JetEu+CILcHw
qKK2wThi+k9rwEwkusJJa4gFi4O/3JdgIiZSYKKwiFRFIPqeaH9AbD+rGWqTD6wyLmg9DNIxOj5d
PuK2oc/w/+4z2N0wpicUMnHawMmjr3wFaMbYySRbjdp4+q0RBergDc8cUOMEF2pRUWjcnGYKcKlS
+J5xBSQlhwvcXZpDc5jOCxDMndD3HJxO4+M7bwl3QoRP1hf6ab6mMfAZZbgnP9ahGbMUtYRP0mJH
nkkfFA6UpCyzK4Uu1T9uPvZo5uWVT8hsXKBUiCK1QWig9iocAFFMEXvKpzeumxecVkI1kPnz4Gpc
QH6Tr+RHSkUuvNrRkKb0JglVZggOPaqXStEBcfq0a8kbjcDS5WsW5+MUz5W+7oOLajf7gUfDU27N
3xwop63A6pqy2RVgtBqnFN5dL+eE601EDOM0ogcchtqcG2ncrvh32RV97lnL+F2/us8G6yXEg3zU
qVoevz0T/ubVwR5p+wVsf/hvqFY0ytQx5fXW9PJSJi3/S/+7l+h2CRSMPQVM/SMQqmnFim15k1Cx
o/DJMLYC1vmM027NSd+N/2iUdB6cVB4uM+vVKgcI0ML6It06tCMBql/uCVXfSXyvZvNO1tFadshc
qNbQ0rX0ZaXrIRJgTFQ8GF/6I8LhHFTaveLJ2yzfsKJJOAs6TG+M8uw++vGrvt+SqirayPWFDEbp
kWHOZ4AmHGNi8lht8Dmcfzhq30vR2fqGG2F+1m6o0CZ02PlwFMikVhkWsGBRONj8Sk4ovYWQQ35N
SW+OTrxbbd2UdRE6Enkt3w0ixS3gb6Xb3u97CIM0/whGo/vLEqewPQBVgF59dcWSUHoZRGZTZWia
9qprToCOBqzQzCNlVDrs078DB1G8EXb9rGeu0REiEktkcQeYmUQqEr1H92uYVz2dSjXUxspvRwf7
8OaMSwUQW2SK1+WwaawvyRBWo/twcIxdoSTLwjc9wPo/m3yfVdY3Dl0N+4cTdeCYw3hqAresauHC
WSyWcWP3AlrAVn1qRFY8KR1XxPrzdkVYIlJgWtm7YpF9r3DXb1dEPBiJ98YuRk9S05AaeePJL2QW
Tvck1TRrZ3t+ULKDvsVBpyjtV2Q885symdRFV61Bm8niZbsjLuTRibyb4VmOH61E5k14Qix1FB+9
UqAUFOHj90rfkY+fe124OMLPlJyc2XVf/TnjdAtEuHbF5XAuGtic4c1b1vWK3GjnVAmkujKDX8ar
ok2Vt6XtmiphrqhIpF5j/7zgNer/alaOa06cLZjFUVsP+6hgivNJkFesCWTD2QYeH4NJey6TtUI2
lxIy+dZ3iK78F5Zw10OMOetjJLuH78rU7oFSRwz2DDjgJ6IButcUuA9RO6ZBORU5XDWx9J9eXStX
tQkn1jYFx/S4K+lB4+aXqaRDRwIvWUWBVFZ4te6/U7cI5S4CqFgr6Z4Eu7nb4iz2LHcyP8jyJAXe
a3XECrF2QP2OnBIu9p6SXQN/H3+LAP5VlhKzL3YtZaV46NJVZ+dskZDLS8RRrYgu4UemiWxbDflR
RnHK12dP4+MgZa6UbhKYOAEREjOHZqxNyD6ocAOYfLxr+bG4LMOmIssSFxoEARei+c0xVwcm0lpW
Iz4mY6cb+Iyf6tnW8HAcZUhMOtHA3lTcfvdEnPYCJeW/HLptpuC9IN/upSr7sBxhl1A94Hh5ZjV6
KbNKZl5JJXnMdYJmG4PyKzRKCWey55PZsPD2OkIgP1di4+Xwx3Fx2f4ec+cHNz9SvooVejXgo1hk
EzEAyKWABw/4urWpfFW7Z0S09yzAQlI2jdgAEZ8CqEyqkqx4eAKcw2mKsPAA2VP/od9veTMT5g1z
X5FrGDmZZSws2m3b0ykS1lHRyyMLdRjoMlxWjkBaCKe1T82JnzATWRAvTN4TwDs6AHuV1fZ+CsK5
PXpGoA1lcKzcuqC0SWSU4tfoy6rTMuF4or5WlD7prVK6xLDutLo6ZE4cdQNTBx0aDIIsvuMPO2g/
lOK/p+U6Fw+VpraPaBW9H5SV34yDU9pDkss+6tYUaS/UF48MqW8dbLD9spqMvkIEmNF+QncQajj+
vmBXb6LiIuO5iVLFrAULw+xDMKwZBB9vaSoStR8ukVHIdT/UNRSmY2EW8KDyr6jYZqCsohGNcs6W
NKdbhnYCZQ2f5enVSI7IkSIvahcflyaMhqPLTlKJWpOzl4ODpbJv7Wku/P+xkOBR0rimmDdr2WmN
pYGLPxpHZNvgF7RQBJg02SRF2uxF6vf6hPjObVraOirNSCfaHw/ShG35txIbLPXa/Fav7P+Xyktw
tRCZ8yTK63vkMJCztcFyuPUIxwNHOuTgybXX1vPpihDHdVDrWzl5ZYvZxJr5meZZE/7OiDxlJSKL
/yv74ogWIjt94HXh0uoQxPoe5W16LzCuS3eF2/ZWsbDlzJ4Vy1pyHdbn/SdbncwJGsictu4fZx5m
7pL5rhANCnzTwnbsFg5EMT0ChQPgIxNG1G/e8T41cQCgaQbK3HMXkYcOnl3HdYUKjsBlt2hvCrfX
LaxxFxgfwvpbyna0+Z9RxeEvHx6mUXjuPGOwDuFGHZZlsKBd0Cn/rCjFUqMVqYvDcBsPgvTzb0pr
XPLKNbBLov92pCjbg54kHnO6zAVbznsP+1qFG2OHphXMEO/CGPPGmn0y3xdjdVPmqM6z1RstH4KP
T7eEfz6RP7iDK1pLVV0RF1TUwdy7okcNGaU8vvEJICw0jHgTURu+Rzlp8ENFCS31/WobAiCkVDBQ
ksu8P7JJrzP9wxQD+UQFPs0lxeKGXuc+U4w3yazCrx/hP13u8egFgAW1cji8w0Q0t0iaBSzNyadz
NtCLVD3vedi5/eFLQjTz+YwDwwcZHnPJL0RV1DJd3i8b2xndLC9HZA6V5Pq2FrlXSAr5lCY624wd
qzaKIcx6+4S9i5biqLnMn4QSP9WzeiXQEt7BzVn6L7lEaM/Ah56LzXoLPj/XnSCQC/OlU8EPGPz1
nMsT76nBP9n03RBOdMoWosKRRcGz/rDoFP8TmQQN7tG/FbTndWWwiRVJTyLbBKHKD1qnPH2PgUPz
0pdMo9WkmyCxoQytNFUf+z91TgasdKfuROkXK8rV8SGSdmFWWNWMgMrESKrvTXitfTs+qcnMbjrE
jUUpnnx/FknK6EE7T+NItZLPXZhVFQWAyhqTVBsVGokGJj/LWImCbOShGVjOQY4MpmchMYfzNljl
Y0dYP39F/V3Xa4LcJ42uyrEF4MN80d/McUgu/JTIwH4Ta/9SKN119QCroldQ254B5UnaTmOM8GLZ
2/AD54MlBvZBsLvlZfxiAqTw9iQMvpArC2iu4F4gQj5vWgTxuHULjCY9GzPE24LRNrdI7D2mg3AG
tQW8+1UnMRe0ZHegVlvUgC+Mz2G7JkmGOR3zSDOAIvwyJwRBmNxlDZquG6sh4CtVVMl6IdeFWTbf
q9RIhUl5tYvT8zL9sK2IWoduaJnyAaIXciCeEmMd0drPBg+P0UT4gKRo7ZPjhZKWOCCIqkfdCSsu
PDo+qAYeWhBlySE3zA5+CT0lPC8dSUitDIyQ4MDHk4bKBR7PU6aOTeTh435Uozdp5cGiUDt0LyJa
Rsp/UZGKXhQwMksTEIL2qn+QwVkru31yqpqJl/3kVfXVlYVeLxOxG2qeujlWRpWyjSKp7cl2a5e9
zNwfiNEUzi5l2LQNEPCuhD5Hts2aCLtXJ74IWFQYjJ/vTBROzc6c/kFY5QdIRbH4rlp6b/FSmHL7
RukHG7Z2OaaIl9IIPQq9t8spNgyxUwCuA6lhzhwr/+vvynT3UrWzrAmNryPZ4WI+T24ps5+8H5UT
vX6FVT7D50+j1XyyF9FIAmBh+OAx1flm5uKdeED7emHuUoRedCm196S5GWs64IPFufU6wqRGYUAG
cgZf2q/OHzx3wLxcuz+RVSd8hj4Qu/eHd8eQwnLaRWXZDirRz3gl6yV44Y28fvJCfO7ABYjcRpnK
vTFbDGHRWl6A00LEnhsVJv35v2jlSdlqlPm/GT9+DZMINPa3qh2Q9NPtZ/nky9iRNlmR7nhlxYdM
8NG4qsS8swUKMzCNUCtTYZWgs2AJnzjBzmuKnjMpaGmtmHXi1kWutbCFYqE+JXnxGi008zz6MNJm
5aY6D1ulbMknmrYUfKvvltbQ0ghVnNPfmU8D9z9AbKdO+HtP6mDqa+/dyiOkh5aLnAEtfZO0XPk/
eB/WXtlGZOODRHusngN5jI9yKJ2fsBzOdf/y3TfxAVAftsOiZqN+6kmymeNjOx+xi57o8L3N+iiG
0aO8id9gWoMoDFPq+MeptZW+l4N02dk4Y31EREjVoyhR4Q8ua02k+l5b3LtLPOOInN4soGVxe5PF
6xJsYrZ90kyhN7KzF0TuDj4thcE6bLKH1ZNxYbNoSQAa/yYb1ijSb3e6S2xruy+rvlaIcsJEZNOX
Ruyx29BcG3ZRRh/i4sG2yt6SufzkFPtDc4kY3BjMJYEH80crTj24KtJq9qvIwxjRUTELIe8wqtI5
FFNXmS1yFHrL/RwAHybSluviMck8LlgSMhsbAlruWymHxsljjdGzXF+phd1QDDH40bc7hERFw+Vi
a171K1DnnL0VOHkiJF34YDN0DlgseJE/Mfed2V7+0ljUvi2EwkP3iPnIVWzjqVm10T/QRLwhG+Ym
thDfHdyLtFyn6gNpR8H5CCfz6OyUBz8yjgJiMDhtgyFdQ5IgDwBDuEkf1TJXXY7JTYHh5d8Mz5KL
LUqCcspersICKiksCuKjR5hguWqz3D1xq4ulPiYsaYrzmr5eQVMjHIyqWFot1g7KenFiwY8zLg4l
akQ1sWWKBS7zEJyPGXyflGwAKh5XeqmfecXAN2rlEhjDkXs8/JlcIBY2C9I4law3BOPu4N4tS5MN
uiHfsfEm3DZo8+gGF++qzUSiYqC1j/Gmfk7bM2gMw3hjXhr0P3widaQ88jQ3F5+PP26ja5jRHSFb
1yqCh73qVewoMQhVyqQkzg2gmvIPh9G9/YP0KIWmc7/69Akh0wwkEG38vrnY+uvGwh0JDXzMUUZE
NXQ32ZHtXX7CDISGuZgy/+uiMBY9p+0NpZOZKEvxI8ld1X4kooUyD4FD1byez0ptaydlPKq0BLkl
+GYx/OFrJKubl9XoD0LXzuMxwKhGyIuDvaP/S24X/VllNAgcWBBDDppdDEGZ1sHqchSJqepRBsFk
7bpFDcAJuIhFt46TPIVMCYhOsZiyQgnmD8CV7fH/iIfXOza4Lw4GkNJgkPwqFyRT6ijKOpb6VzWB
GPRrPismQKTaTmavI+J0m4QLUp6jtR+Pnwk6L0ifljq8L+IXv3IYO+OR1iSIiN5KKhAJX4Ag+Kja
iiQFL9/yfWVBJPXLfFFgVXJVm/9wX8hBKkTMBZT8Dk1Z9pCt9oh8wiew/27zPAAhb3/90GpgPyTT
zBHKE/uHi8hhinaoXTbd6hw6/hReaKn6fxp7Jv6tX+ddJujZsI1wTGBe+aPodgMuNqU8f3Jq7sEe
3OeuKn+Wze/xvxYSovr3WAtPvW0LcJVbMEQ0HVEB08yOZXcLx0Cnn6rdNyDIIh7I9NU4mGQCvtxK
UCN+MGQbcoWIqFsKSQKstp/dcXe7Un3Pie4DxHone2YynGoIguz5DojY3W4RD7uZo8NlfvmDoLaE
obtamCIsWHr0sCYYUrOwe/QxFKZcDdBFOckyvKXP4VVDzZPng+QQ57hhxozGXtejpUBl5dWMG2R9
A22AjHHS4HKINVbI5XRKDm+kPMGzvKyndD9OE+0v0Xi+f5aauKcSlodU4NXH5rPKoJ/v3dUSvO+d
SPp0thej8BjvOnyVvafsmJBEjGyVTNNZfk94ThAzn+qCbKHud7eqsJsmLaa7+6qScfWbyxbHh4KM
8JtZWyLpRIqPwP1E21CzDl9pBg8zUMSTPFj44DpKM7f3Xpve3WKXZiaIKBJVgyrqPSd3N+8mw+qI
bcyXU5/Udo5ymkafO/AX1DnJfaP1RvgVFRrClVO8VcpoEle1+BwGdc83lEEp7A6SyE1Ax7s3JLmy
MOAgaVeJs1CzEu53G1YTm+cXz/yPAOA1/jDs3rGtGfjFoAZ9iJmBRjVWIBn20sp1Ky5FBEBd8cg7
lkpJcLzeUFfAlBZ70slirkTJpV9tNLMBU+GO5pjDLxtO6yXxq16NsaLkc0in8ViKEJKfCer7kdjP
hkaoJTrj1rX1+yhQid2cF5d4J1kHueJt5khNXeGm1uxILhM1CTlfVv9HJYwcb6M+jM9dp9bn59UW
XFFRwFvQAr0+G0WjXWqMUJ4H/bEL5493AltiyMdhj1eKjMNY9k6975Ab18O7cfdEDcFzHPzekRdJ
F7cZxhuhL8r1hYwOV0F68jNxS7P9IXdn8fHjF34pFS4fMTFKAtA0Z4PQL2NJAYaLUwz2NgP+vI/f
Ys7XZ552BGFu6AD29nYAUyhw+1mnHQajhustwRUlIUPty58SE++ramjs6hupeV3miBJXhH/gVxn/
yBd0a4JrrwzeOUNCqKi1d3bwGur+xLoNWK4JFluva+7h22eQlEHNKzgkTrJxvm64NuE+uGerRS7/
7W7XH2JHQGX7Iv7wD+3hb7cxHQbZsA0cusDToSw1YhHO41pq7DbGCs7ZJItOXraBbpBLARJiYzuo
5cMx9RbHbiH0BOTlyJ93gJ0sTNk7swfoqFRCQkHDwwC4D5pwBMaF/MA+fyl38ItQ/1H29VMxOe5C
Rndzd7ni2FA1BiOzED/Hr4XGJygLogyBPeu/ImnxwZU98g3y1XQUHlQl8qI36YytJrOTXrrkhiOB
I3/Dlf1EO6p+AdcqOzqYrxs3m9LDDZxnx7h0YwaNy6QhxviFdJIBIBizLfzJTmUB6zUKvyP1TKG8
5QdWp0EH4DG7Sx7Gcl0f6DoZX2qfzYeZpFAlBicyJ5AzJYHQdSt1gV4hX9WMt7zHSzgchgMld9Nc
XJldRlOwtnmGfr8HB9GT3TljylE+MMf4zSOoIR0DFrS7LPKQOtBhBSmkOd4WeEpUyc+8BiicVCES
uu0tWPccupDyaVREVhhpKAC8EFgBd4Pf0Wan7z5aflxYFSIWUPrZQ0ONIw+oeY/M5VMlR0BYZwVh
B57pB6B8oqp2Egm7RGpkEjBDpl5821fAGUdYsN05skBCTUI9nz+QavniMjiyUNuF2E5/gj/A1sVH
OBEtiLA9vz+PzeikkM4yTMR1vRYva7FKj5yMtxI/WRijM8EZKAbwCdIRjeDqDaO3v8IEHFYpBS9x
/Ljltk2DbkzO91UPoyGnu5XJ0arOFwZNqPd/UpSTjOqxRBTOB+buz5BaVJOP01xwVFFDE3Ui/Wae
qwR5ROJLsc4skGAS9zQjhqOmdtzm7Wq5ypMR7DWhjK3fz45DGbT4YMKJPERvYMuES4rk0DuwJddI
4RlQhidI38AH7ddeUS0+46QgiH9dkP8UcN0PSK2N6AnwRMiOKNYvyi6M4t2qdXxnGyvQEVDSv1/0
2B4vdBSN1DljbJAGRCF3Pp+8JCnZe+wxCX+3Wh2bAkONxacqLFX/59WxoEZKp6bjpAOdSxpeRJIX
oijPNcrFX+lP/aDqhpJ9ZcphGZ5nN48sKn9pCOgtwqRmwDHwcXauYkw0FLDepnrx8faoye+XHH0b
9jR4fo0C7jJ6j2krMR/EKn32iVh3FVhFI9UAsq+KAvbCXhjV56Noi/batmD5mTpV1r3d/aghCLZC
MD9FRmdAiaNpsrsud+R+pC+Cht6Jfoy4fe0DJH8i/n4rVKEEWFpFeD9tbvONdn18//l5l/pfdkWg
kSLXSxWXZEJZVPFRYF55S8VsXrZ65Ndxidg/A/5Rdh94TPN3dFV2B/BEABop8uHGQ8RdGZcLT1p4
Bs5amRpRzMqY6K60q0qzJFOwivvZlVPnR7lEf3E+S+W1eCBXOo8pauhbLz7xBdWb0JuRqNWgwolp
CL+YYAykcMSvRVhe6aUtjweNhweY/bqK8QR+mD1MU4W4DfSWqFPFrTwQAkIGbN/OROLT3qwaVt8F
nU6lEv9GmmcdA/qrydCeDZDThWEPxLZuj0XQ1hZU77rrV5tFjwcr4faepw4vSU2gnRVmIWhEqfFc
S6RPCk4/qFrVQCqufHJNhtS/T0tPqFR7fo3HJKBf+A9kLSkw47IPvhbzZj/fkMoCdYIjBUDMWY0J
svNZS0JAQVy67zrMtzX5AyOzvpOWEuu6MsVaJcr4oXHWjeD8p9etVBhUYWV07tgAMTXmxowyQJIQ
ahRcj24AQGifUfs045sk0j5Wa8gjfsInSsouiFJvo/hZbbtBf+8gz9YdUVZw184uPJ7n7Kq93Vlx
zWMY+ljrivnR+YSxsQOmQgwe0PEYt31+SU72Lv38hg/xQhAtxfO0Wtt3YE4E44rAeBa9XqycGoSz
JHbRyAex0XRe40ul7xwlW3D2raGxA2zc6VbYJmPP7J+zOAT1QNt/V03U4kmVUR3NdKBTy/3MyGKH
rBNMkGryjb/ctK5laBxesOwYNBzzEeEAgVI1hqtycaNN6CSof5+PY78uNJF2YJ/ujvFqczrgMQ6/
oPnNVlsk39BM3dWG2ARv1SaGTN6BC++z/FtOQPYhwozaqfYPVyPPWMjmUts0DGS0p2oV29Os/v1H
5ZFHhf/lcN6APHoWl8ZBE02TlaMhV9PqebWTWW39aLEmWkFIJR5LjWPacoL5gyhgFEGfMKNtoxCL
ZJy1cQHizuFMNPU8aFFuEXSnmHjIMglOvPnRBRQ0i3sLaApbHdjecW5uba2ftVma6JI+XXBaaBk5
WupqNmMlVwGGgHOyijWA1932Wg+OdS4hL/E95H07UE9DcoEzd6LDQAEO/aib2L7jNiHX3j2Emfgn
AMhpnvAqc0hVRXBq9wePl+pFPd8Xqfzv4KGjPZ7zL0veSSXrTpfEX7LmsiEPTJ/amqOHHCOIouGg
0vLhdRWXvSoS4TR9VcERO2MGmOL6TvRql/9nxOCQOxZHqipBqsvfMT1G0M+j8kPK1v3cLIzg/q29
2W/cfD2+C77R9GXNTJBpxGZ+cO51TrZc/YPmV4ePlz7OFOajtwzVAjujz4yQ6AmoPoW+KtU2jG+v
mrBDPwO8ZlLr6tkvct055t3xB+nLut8c9H/HH+WthfnFfMmAkgglvbi/GycEz6UZyea8lZ4HEcHV
JB8AX48hTSKH/IzIyoKK+zVmOnw4ur9i9E1URTIL5dIHJ6d3qvMbMZB7XIwVzmwKARuFHiC9mgoX
DHZy5YMoZNeeEfq6ROea2GzZdbeI4Pt1yOV37kc97YSGVrt3D/w7VUaC83u6QN6lvCjSflKuVx76
8QKWXoT927vf9JEGjBiZdFw2RpYZHO+WxrnvSVFIlJKm5jrapwQGHJrIxzj6xquWt6wPEvkZjiaD
48br2saG+McY1yN/S732B6FD7v9PrOjGGjHB0MhILbR5hTiOXXrM1UeYvTIdJNE2XbFrxCnYdQ4Q
P8WR8C1Dy8WEW8EGw4ryHAYdUzcTWtovMz7EJZYPjfMyWLFwoBoF05IQWnq4HKT7UcXH+LZeVzGC
xe84bttOeZYnqYjRAj5cdZXUcIpEulEvx7eQ1KnngY3GlfDPRiSft/5LbkyVxkZkv6597n6v0WKy
hL3hgkwEJMjFytXkUOxfZBBgJzPpZAqJ2/YMcOFPWB8S1iyjEeMswu8go0cGKl/SSDE7LG7tIpGm
znXG2QmVcfKDM0PX7en07RhLlcvcNus3/1C3yisD4O232M5vByVAWSjfMcKk3LdMzmgqPxqG6vp5
3c5FVSUmaYVNkm/Stwr9c1Sjx360rY6HiovtBPG2o+pLA4AJGaKi643Ru8yhhZKJH1rK5djSQfIo
s3uUCL8TOsDEwnU75oAiR6mtMyzyVPthi5qTN9L2MILFrt1vh3W9v1giiBDQarUWn7KtDTE6nwPX
DBDrDQ5ryDd2De/LF7DD2Lp/2+CyK+M9m7iP9Qul/Vspzq4dLA+UEM4dEeq/ahDPI9lrZs5msNkd
0iqYdHgNxJ81HAVyHM6i3WKaMLvsGKj/oY1G23HkTMlLjsNod2vd5i8r/W8H65f+WDVmEadxKLKH
EwjA3VP5VPg8q4m/NNeMJRu5q9TpjBGaSFni8XMp35vCidaOxG+S18Z//+2PCqtXo4hN7W5h36O2
sz1T8rmgOr/LCYwfneRybWHMsicqbu6NMF8X3RPK9xBGO42rh97J7cXHtr9MpIAIy66Qg8nRpbR9
pypdmw+3Zpjz+8Hc2N00C3xVxgKKxxzvAPmDc1C5nS4cmTzw1Qe54unySHsfsOGOLjfnyIGoJRVN
fUCZDRjC41kV6PkJpYr6TL35IsRyd/Tdr3qNfao+JdxSfrdW7VMUg07Iv+JXojT2p30FXddk7krh
o5cipcSnmtv9GeurDaQc4qp2k2xonLoBn/CktoFwT9wIUzt5LYun4T7gAr0YL+Y+yU0B7/lKxLS8
UfZ88GT8WXMIDMlWwk/MydJDRTkpkM7cc8j6xvIhwqCHYRyD5JDyGnf5DhPtFUbUrZ0sPxjJSX3s
xSa4gF9exLh9+Poc5vF0vUy3FLWc4mhf62uLdGK21jDXQfPg7u3yA9e3/hyqKbFk4vkQ52ALbijo
7QgYP1xOmjgYFGjnbrAqp1qBIT05LkCmI53UxHGZmk7ajlwg2Xd+7sm9NyeSday6Cl1afKn2tz0z
7AkXmuqDGV2mZzzI+vajM7PUKxPcqp5CxERg51nyLLJz3ks5vTAkyqy33u8ewKEOhwdwwACwm7BL
T+YSu+lAFh2xtimDcEb1vNkV+y59mtIQBMCgK265PbWirb70MmrZiTjCma6JlgwYY77EfVRn90c4
D7xE7MzoxvXvLpFA9T/VUHzouJ1t/aRodvKYiEdkqc08lJvUaVIISmkSm81cANOBfQox9KdMXaUw
AKTRjsPJ7zUS/NZJSYwSrgkQozSlXJhALd2CAsSyxuFUnHZ7VD8WyloOCRFxSZ//MdPW1004L4j5
bYEXMlK9tVJWzGSTpektdXL+oZHfie9HTV88Ly9I2RwrB+E5yZ8VZ3QCqxr7lHEouVqotvxfEU0e
G10b29KBlFbzlrWjf712HMSVBkRzlGJrHcy2TverUbxPEaiOMxAFnJ4BJ67HB5GjvOY3YiE2FyAo
J5VUTBqrSuhME+lxUnBxrmVrMGRmvtYJS6+FnQ8p3PAcghWGnYHmUWXR9x7LdCO2cCuQG6HYsfzZ
Fl+BlBAISRrTZvHMMWuFhOkO0bJHJb47pn0lQ1GMIZ/6JAzIVlKIVtDLCkxhKj6mvrUGkfjDXWGf
GumG1WQQ/Ky0BGaSVPlQzi8VlE2zVoz1peWQIWgHXyWHXsx1aZdSjIgvCGnH6nQBgWJ+djeOH7bo
KwREmYSqlaVtrQ+pnJhOjoA1/cbZ+6eNTnp3dfxtLcS8rB+evYP/LhNeQhJDSTpS/N+Uy0mQfse8
603glRdPVMcJIRnODOMvWkpl+KmOYCA6cRdD26VtbknAzp57oBfQwncgqrh02TQhw+ibEN55xr9c
UK1/9wc3KqbtFec74D9CjDR1oyiH0xQC6Nr2sDbCD9HRYt2OKYX76HyuG6HGmDA+so3aEHswQGhE
3VGOvBFJv3FzI+ZA5WYOyqGOaQSGSu54mWCzUR790F4PKoBple6IfmY9KJ4/omEhvpIJ5iqBrOzh
d+HURaF0L0BBAzVKhnTgMeGMiGkHdQgsd56j+Iys4i1QW2QPW4XZyfa3lIUWeVgu3rcSBA4Awcs3
fIaqOMzZ8Ptl8U7W8o2Xphe4ovPdIF4EI2fGr6b/EaJqmoTznpllDB1pQDXEz7h87DcMEVT2zL36
qi9gMwem2RP82tOFnhHohfevP/0ADjsVU12jp4lxKFTj6ddfBy3EXILlQZ6Vgq89bLyhzmjPs04Y
cw/8Pa4iuHb1WeuX5SFLUsQPd/L+TpFiMiQcVgwRfOiiE/VgqMjXayMb50jPdJSXyWfwDhJBKFEV
m92p3k7+Hc2k3vkCYWe9wiMZcC+xZLxrmZ/xcSoZW/z4QUgL2yGcqwvAe+WNnC0QXVU/PBvRzidP
dNfxQ4BVOADzjnmemMSG2NhTw6sb68g/BXUsRj7Nvz6207/BjHgldAwTLfGbr1y8DoMJszvlorDV
c2q56FjQqDjINz3uyA3yIpOkWp5MZQxyJqKHnh9T4lUapBVIXxkc3r3OWLq4sDb7f68/T8o7K3H1
2DBoIYNdp0yIzMwdAMfIHvsFdukRkci+tx4Uudx2BfQ5SY0U8q8/EO9LkRgkc+mhwO9BCJYUY1B4
DYkQ6VcYWRwnfXGMIevzyj6dRqkLP6EijTjjclfEwccLo0oOhR/zN9v1lA9XiE7I++SGn/AdUNAC
bTKNUINwe6dqCfb91Posf7m/5O8YIrsKZPWFwTKGC7hV/HgUsVuazuSyxnhtBTRCCsOeyD7KtHux
SJnw2sW87mUpG9hvqt1JfsosoqMJR166bEPqyVmVXjasolg5i527phsLzm0R8JEcwU+r8mmVvLaU
KMuTrMaN6sIQZ1QJBMdh6mI2Z5KjxCO794+izJgNo242N6vxOFanMHvXeWxx71T7tfvzBecHuLC/
5n+oSQ1jzHEU1+rO9RR02V8vR6tdrWeXu9v5ikKABxhvyb4qxelhyjxgc6IDaF+qidsln0cyJ9Wo
dQ1EPwkViE2GuvY8JN/PCQe498JDeWOkzQo55Vb0qXG7YnHJ+66oSk2nYrRXQ0JsThFM83NTEZfN
amNI0hRWkhntMhAo/BNa7TGpApgljVm9aq2tp7d0Xllls7/PHZwkMSFIFL9K9m6pOdcBRo05k9ll
IDh4n/tRDzHLVKpbLh4+mQJdTKzwXXbZDPhSoMPcOmLNATDCIDG0rXYcp/CJzBhC/qHk3Xc23Ib4
jkZ2EIa4cGBXy1dqnqbrdWHiynSucN1VY1SiTK026vnmCzjkrYlqaxYdAviW1dtm0qv0LhzIlZuH
piA5kDW8hj8X5/VKGBnnH5zDSvqCYTTMcHJUQ+cZNFjmCT5zivdRvgAOa4SvNS+HFIYRu6QwsOIR
L6WrEddmbmF7XF0iP3txaBSGv2y7N/SGfzQ5FB6OJf44rLkZBWXBIAedESYkLmF1oDLZPBbUjD7o
fhJ0msGyRBnoIiIEal2c/SNHbZgE38Pe09CudR+a/G1mj6TSIuvfJRCaCF30shuMtUid5w8zwiPY
EnwirdCLB2IZBeHBdXedXAwWzW57qaDV5mTLUPS+dKms2jWFFkvObi+j6a9L53w/thtsHWXzxB0j
dXuFkQaRMZ9JvrLAWjIzgs1nYu6CCxK05C5/0W/3i5rDt9xMNMwogZ66c4A3s5hA+6WNniq3K8sq
f1pKWddJQ+zV1TPRtQA5gqZfgxn5KynIOJ4CR7+jYIvGkrPS9OiDnQ5QakIg9cZl0S/QngRhcAB2
iw/1S+iSu7XtoRWLH5CYhEOhEP/HpSlIN854qIfAZQ98O4bohLkXJbq/RJIIJAH0ayuyQh3B3AqQ
88K0215tMwGRwUpai87Wrf9vDVY4Wku3qTP4HgyDCvvXzDa1Kd34QG1qtgsemS0eLsDNBzJDs+uh
BWVdO2bVI8mSVhS4wniqM8gbcpzgG788y3005LoAzQCis/JIdfBvdkLoFlNLMP7ksKsERzQnItmQ
fDnQ5e3tHBKBO72gr+PVS5d8D13C0d0iCkQgCfZubZdG7PO3Y9Wv30S98tJVUNfe+AZttVCF0HNQ
aXHJnSyWaAQ0jlWVdsM+pbBSS8bJyvsONJ11Fr9529jdmdtO7K2ywRayKK4Xv6LTdYSdgjFhnwgH
oCiVTv5Hn9AT9xHciXWw2Yxam3Rsu2w7cVyuQhL+1oWgyvsbbCdSW9KWsC/974zKJWLf8DgpochT
E7JcG2RZ59nXoBVQdCIdUKk+0jXqvSjIZ7gVnkTY4sX/0GLTSEBRRa+1E+m7yCbErh3g9b1BAg/p
OyZlzb30c85+9sv4LAv3tWAbaW1wlpFFy6mMCN7wKP6KOEwDGkB2V+1LrN1lF4i128LK+CMmSCkA
BVm4yUaMEGQpkxNxcVNhW0uguGcNPSlI661vLpnm/3a2/goVDappXI7r2O1Epjx8YBi0uSq2vdek
Z4Pb2cC3jx26IBV6K1LcrXyj0ZzoK5jFz+xBmVx+tbOhSlHJCMNZ2nBYl3lYzSXZbOcECklfypoO
SPzGQvSR9kD0I8xq04/Lx22VLfEhPYuevDAc6F2ZuKTA/fTrAp9cGUDjhPjsl0WCtkwyT7Qn93iB
zfxOMpzFIAgaNPQdRRIqv94XFWQNL3pkDBHqOveUyehpP/LhSQEpe13ZyFS6bhDXjdvBAPhbnYk9
3R10Tt+LtO3j+2aqfeZbkXDMAyTcAGg4Dyq4XhLwb6XZvMHzNHQs8qlTfLakBkfMwC1gNbZBElvq
oqC5DTEcspbjJDrnbuFq0yr+llhtT2gNPivmiv5pH3PEwACHPgl0LeDah9i5GafDsrY1DPhq1sUR
pHHCDrGrCyn+a/BlEamqRHujl0CTp1wFDW1olOZMQQ3IqCXntfFvBYKmjBAfkv+YChqZSY669pVs
casq8oEQk+XwGLBBzfUpMT+hKxX0Ysj7+8OF1miIdOMJFnR5ZyaS+KHWW29yRYvmfX7twNY9lAgk
4lIUbwP3RQ+re4rG1kcZvY4JCLYimp5k0bp/Hjrg+vpv7SR7A//Qy3TS3j+C1z/ae6VhoSY/gZCJ
24J+IQnXNsjr5tcV9RCwKJkx2RWVMMOe12N8emT8BS2ZyRAKYEGVevTy41tgJ8U0QtgFXruO6oum
cppHbM3TTsnpLdN7yEsivid9jFy8mEjxTeg4iVb41kcblfxZaDTwnbHxss5ZqZic2hfKyJRk/mS5
QoekHpBWCoZfSst6wrMasQAYFn456tJ665P4JoWS8TWfnc3+ZmRhHwS35SLHyc9WNjqUJJ52Ie10
21UL5ZCI4DiXfEyoJ851OM7CXhKUdCq8HWJ+s00Za3DHPiGe81IjX1i7MIzMd+7mTaGUuli+5dCo
pIOZjkMxmu02js1scBjRaazvjURnOCUP1XBThFutU9VjYRdUS8JCle9pl4zEpOpYVojcgAM4c01t
gJ4unHVvAbIqYoyKa8jXYEIWbJR4yafmnXdxBFzjf/cARVoUq/oYDXU+hjr+rfmwesOkBlZxDbbX
5KApaPQQJqv82wLd6xcDqqKR9PP2GlYKmlzvydg7bh/w+aeN1G0N9ue/9tXEWui5LU8NFlst4t7n
hjxQjWybgVnYNFpB7ax/rJPwwMHZb06XVsN0fwQbXVv2N3HliGHsr3Ds9ntV2vuY/6Cp3nmRHqQQ
+xGPS9L8Cutqw2QWChswuZC5bc9nhu9/PSj3yvB08SVF03XOoZtS8DDYuSRMnQPQh1msOigFZY5A
/K4g+ztoq+lhOahgq3MH9KR4fKo4b4SuX6RPg344ROM3HRf0VDpzd0L0L6ghBAVnVUpCRgFpoF/J
JJzrmTG4qSiyuUkfpcOBjfHtMbt2bENJelCmpBMl1byQGMPgxGoLdzVa3ekKWhcgmP6Bw3WK964J
9TIdJbTqbmUVsB2wzc6h5B/7qcmaq26+BFh7cI62It29KEFD8MmKPo4VfZA4Sx5B6UTg6Gx0F/u8
Qom+Akq6TUAcTaj9ogZ0x4LCj+xGTtqZN1Baum3mPgLMK0sEK5pEx55PI+byEHFerNp73XFL7m0H
I5mTR8zjQ3kk0OCm/ZwnA2hS52z9T10ZvUmu+qJxAepGmbWi2q/DDb7c2Ob2c3vP7pMG96IhDyrm
fBAdMsBzNQGnxlmlc9aT2S48p7KGv2+URCbzWFvwTLne29pwquQNUOL3HBTxpvacfZV5YltXWCsu
T1f0G3c5UGHK1PjDV6+TNMmdHe4qoH3XJEi/dviZvrxk/p/go0aQh4lnb+KRuD0gG/yvPf/3O0CW
hUzbeCfJ3m4X96T3jylLcWaQ61ANzZCegRNPxEFcnanO4Q6xaO+odqjV60U9As/WOiJQBthKb+KI
Eiz453xLFQ8Z6LZ1b2PQveTuAHPwYI1pApZANcJVgli9GzKu3/ioTxG09XTKKQ8w0w7cu8dW0d80
QrWo4i4M3CVyg8KMAF85wjrdMj9beKS2SSxarwq7L6Kh8p7Sc9XWmrGNS5UNXPYetmqz/kMAefKc
QK9gs9TY4jqVvs7E7x3Iocs34TjAzT6WJLFY98YtCCkGMEfQxC3mLRZmF5sQVQ7KY1vbgkQQj2Ax
ngGWSSZ5P3RMD3SzaaNlBY5cu0ZbVTDKBcbkW00zCRNDR0d0lYQyuCVRT53wE7ZIGTOOCX6OS3te
OfSb3RSbYq3ceQNRya77H5f/AGEQMvasHM8dD1u4vVnEXHPnjjONGa6K8S3no0kayYvCN/CQirbe
KRPHp6al+hZ+i/no+adfKr+g7pFa97T1IL6seyOeUMZ7gLSDf5WIjW9ILRTLR2i3Fz01Ei9PGRbF
U7oQdtmtpl4vtMaY2hR4TWYW7CDk1YMPei0WgSjjEzo3QpXqkw04i+ve4KMH5YQ5hCTyb6uV1/9O
2zQAKeNQMPa2iDeGHydO0hzaXCWSj3tQ9uyqVmCs0ovDGmrliaF5y4B3COTCsMBZC3JPs4Ry4XgS
WhD1LcB9fN+GxtvR1rTM5MGxAtD1hL9rTVn7Vn3qLL+6IQ9kY+uBcFLoMJPeSzOz+TbE14QgicEp
MLbh+aEl36mwS4/B8fTj98qDZpk3Sb1/MO5ITtYvzKQ2SUdYQqbz3x29Bwly0yrmiyyYp4RmiTF0
URPpDVsVwKb2YmddlMADQb3dXSgdShtHrDWcdUnz+JUv9OiM+GzbIgApIZ/2kqsf4qFFC6ai4xL7
QsvjuElaaordHlNuBpgeyKE7hHruZKkAkVlXB53shkeDliS7kFU0lPnWuaK3tAoNVej6vQQy9D+O
HmvYcTzdglcA+y0LhngPDysnlLJ5O9JRePGIzqaqTfPD5wGmzeYyo2yYK2Dpwp2i0tKEeO1dRTQP
/RB/pQrGtCyVBrpf6M5nfXj/5U9lEwXkprqYalX2c49bWwIiq0fBn7c7qRT+3/98ftnvzNOjzrpN
qaZBiFvKYOoqEm0a4tmjMO1sHnzIBIYdhj6DTyO8/Ey9OE6uvDnTTQNKXGGI2DuPYfjB6i5ujZEk
brPajLnddxuh9srWUQgv20t/TpDkarId26eh3uDJtj/hWL59S4kNS7wdM/GrWayMeAA8hs+H22yg
E83DdE65uyu33vBhtcY5Oz6VG5Ji1N87IxHykCiGwK7t77PIqaUnZAg/Pz2tHM0YDyug7LiJjpL/
bXgVLnBZKu81xi6ReB3enfvB8YD8XUi7zlmpjX+hlr+MMuLXlEh7qPckdFirzNl/zLVO7yTOy6Q2
ZtOyMulS8avdBwW+h0PXeM/VoPENMoOfRqYy2ts9HQEtOO3D+psvL5WTr0HtYFBKtQKDxnptVTSa
QJJN93X1rSDrdIKFfxr2orc4QDQ6DqfnlhyuJwMJhtayx8BxyhKXjS+1qfSluCa78FjUlkaydaXy
YV25d3s2wyvuAVkbZbuhVp4jrCafSB4Ts+Kuhzy1Xa8/HG/KPp9deFIGnIOn5xJUcrjVONJ1z4Du
Mp0nBnQtW66vjmvgf6Dyn5OZCaG4mBzhAuOFsXt40BVl/spTCtf5myXNMR7aXnik0ITyTsv2Fncg
ORkBBMDOPAuSLPb4A35/H8E7zU1vFj8xb9mZlHYZEGJbFJwl58fq4tBD+V1CdVLHStXg0xXwupc4
KTdeD2fx0mJl+m4mNeSmR2+AGu1YshZ/pUf2g55oZFp5QgrNN0RwoCKiW3QvcIcgyB2QHOQctJ08
swPdSaMJ6MCnJTfe29tPfjcOUpmhkuloikejHQmtw96jCo7e3+RTAV4Xb6xDBs4lzRpQZh6otCW0
89KaXDyhfAO5Qc0PQLgFYhmQCRidAR4PBuCHcDdkVh8j4Vu3EHYO1rzHChDP9FpYAC7hAbNW32bx
fUDpFO7Ij2mmmUanoQMolixb8SC9gZlobMy0ArCwuLUEfvbWbVZbMYkE58dW1KDiDXksl88H6lT8
CsVrAh+ryUqaUCKec7v8Oc3Z/0udZyDUvKjmE7A7qzuCOBqelyYWPn5+mWdtS1YTMIux74bor+xp
MiBVNqSApy14m2l1diEXXMx3eGPH1Yx3esvHzg/jHSoFtJ+GudJNu35A6uCO9f8d/8SIksCmqoXV
LFBujg+ozn1YrZBUszoTWr8YijFJq+qfI1JbogxDjL+C/TO1f6FUqX5m1K/mNFQOLIm/eP0YMXU8
EwRsv0BpmBVEf0rZ+omOREUYlk2TtLs2n8Adp/Qqtgjc/AAU+37AViCbLoRvgYwJTZrCF6FI1Fba
sXvXuW0Zxzpv0r5tiQNeFP07JifhzUCp8wSFkhd+Mv57Nolk/1k7C1CtbE801OUEhER2mrl8QO4w
pWavcy4hEjQGfnZP/wWHE4YUoIebgO3iXhMSQH9EkHI3XGFMiYUc0IEHw29Uooxg2aJwbPGEqI/g
bs1ZeIHnokUbUQmwyFT9QzoAEvKB8z6y+GQBfTLXf3CyPEVNyVp1+lo/7R9D3HWgnNtqjnZSbvVT
DmY/bkGJeAlfJAQDYTyxh0DseKplaEdBoOYl7nMPMfygpbphQvj1QzBZym7HLxi+/IXLS/frmjha
65NAT4AO4NNo2qZSIupH+2cskSF774EH1LS69cKoSyThMeUKpWa293oyyNMNrHEMijZ/ppuN3XT8
RtvQHdm3J+bOx1DWewfRmu8rnYjEibnEZb9qXgIqSTmxCNQ91FToTLrVYS2a7mVAlA05RqF8MyYG
rpZrxbTTJlJaY3nHAtN/Q3iSxt8+UJjtbLaypsbZCABvSrDP6zVrZbh3qOidWjURo5S7HIBabgy1
QQ0foZstDFPhosY5AigfWO+foyum6BTrdOLHWGhXxRvTEw236Wl4vw7zI/+UpPYawnvwz7xcBnD6
FavkgEuUeyoYYIw9DYDq+iMi/ZlP3G3xP+sNq+4vMJoEKNsbOoJyqeBWgfHX9tzgAbu9nhxDFWbw
5v9C1Lth26BZJmYkY+YIODQR9ebsokKm/+ccUMOoSLTTuBLXUH01VWKadtTafPbj/5JgDPd3dgpO
5BI775pFXrCYpGgaCv+D/y3S959UHWyebP3sTSDXtvM6mNWSoT+ilSnr+IfUQhkVMgOpQnfhQ+LU
iKXP14EdDcu995SdNbA3ZjHTnaxE5Hnm9gb4RM/7Ctstl8jOSCUNY2rJv9f3pvOnWV4XqcGNSqqh
tpYT2Hw9ePF/jBjbgs8b81EYpCrozBLUJ+RQakz1jmpGvf/Pydhzo6UsvqIqB+6aSbdfZDxVlHsh
eIJj5I8+uQJuzg3iBvpnxbWQRWxeI8WUpspTktP/1AnEqMgWW0Gw7SWVJDgeoxZxzTDqYSpZqyni
yIXlyEUwns4K0zJ4bprbYUPoyYDwK95poATEy3Wh5D5/qmgSk/zF6qC7gjVxJCv0nvveH/gk2bFB
2DhTkNiMWpT5u1O5L6QjY1h9wLGpryW+CyLG4yFbcwGFaEaH6y7NcUxvXVpdFDSOrZd4rPyxOT6i
0A37+ojfwu1PIgrJgile4OBLFxyytOiViWbFE4tT7kk7Up7U6Au6Yy4Q/vCI77pwPLruVLDsbg9l
809McDJj6cLqdYJKk/tKGw1Mwf5OUbJ/OxFvF8cSUWITl+6HUfYKSW4AntJpbh2C5E1M9s0DsSeI
YAKYcvNcT9Qx3NTlB04HgUz1+6GF4FJUO5+pwwgrqSQEp9UVZ7BrfpOxOPePQWfFaLVQBqBqVvw9
Zdv0VF5K8VJp3UGCFTGy8r3nAerj2RvdlXFX+VgW77HS9E52RwHIzRZWXloFkFTzegHG2nSvWZiU
1AbnuGsgwdhFi69PomGtqYuTKErKNTi5xPdjXVVyAd+3sXkvBE/d0ulkCC9jaflNaXd/8Z+zH1c8
A4DzKv0p5DDOcI/TQsgYHpdlZdZ8S1G4TLJN+okWvjRGMwOY2GCFLAv0j5vuqofHgra10VdHqcF2
I2cdMKn/VVhIgG1qVFH70fTmwGEM6ZWT7ehx1ZxlsNcNUPUZ2psWyKmN6wvhv8UoLSjdnib4I+u+
GDjB+ochOHr/Ez4YXBsLZeh8xmAarmiBZj49hHjdKb/pM/PTClF9AbsT67B/o95Dou+oEz+UgqDz
wHErbNtnrZTo1l0M/892HjL6Ls2Jjz2EVuez0KAS/sHBvQSc02QA7zaXytACaTBzXqsvUl/eVm6K
A91T/kPDhAlQAU7ZQf79yKSyxdG+FTGBD2GozNxyIYHOZ0kLqW9ccLcDJlkoCSwYifMhNAbTAO3l
IMRqE2cN/uH/pORyihxw3P7q91e0WVnI8s5MPRX1eQzOlh8XixPxEsq+ovDMGD9b5j+AqSmvDeSZ
GQ0L0xEUlNLE232o/8WYHZPuG9eyFIPhpkm2THgJ8LXcHOfmUkA2A6VBmRoqLKjUDEe6LediiZVU
IlW8iSBKxTZOfc9FfylRsX4iaI4NW8MHJ9SRVchmG86fTVFu+ij7CpVhEaT91SGLBF4WELY1dnoJ
LG7q9GkuyszRi0xarA3bwKt8/evHLNK4W3mDRec9RyNDgfu977M2XYD6ce5Mwc15XZYfddmIMEkE
S9EhCfulPJXmH4uldI+qpQcFBm0krJU7pLVqKZfIxJsFcqRagSeFoUVyg/xb9uohnctpKChfvV69
0KYD/UZmxSf6s5REJaDvIAWUWUTAOn7Wr3Zm89dPbU9LLYwYTgV+KWQYSlKGZTSITC5kU20YHioa
+tDkQWwBitqag7doi7s/kxCOwwb9MpjGcZdHqVrWEHLoXJ5veBWHwnvDYJ5F7Rivt7SvJIKvLHqv
CGI0eydlREYY8sDS7v2sGFNwBrzwxeHPr6G67ExFixIknDLdPrZAURho5KEAFlEm1ilT5qZ4H6UD
qdR3zUAanbuB4ypS8LfrC+RuAi6e5V7b4d2hG83pOFd78y6sf934VbIirJvlF+KUu0ihd/ZP7Xbq
8wwi0za59cSOTQmvVD4X2dOYVh/+wCxI6uhdK4VlNhOou5/GfuiahvktKjQIr0JbOZKepstmZdEp
3ScXHySTNMEw8MRbv1m7JVJgbxtdgDUAvrv38qO7uQGsBG3u1tlGTAdQoaJU5U6b8abxYPJD+Kak
3SA/vrtdg5ve0Mts2Nlk18MLQ/s+w8VFUwLyuHjBSl1acuyZhtBmuBmV55AGkIr5Kh34VhBgyOC9
Q34aPJSp6ST+l4qDTIeq2S9aR68kK7buuZDl9hNyV3vxoVL50rriBm0vQ2aTL2BRs0xNY75V2WTf
EmC3KaEtUawQFJDnFbUn8/r9DD7yGgG+I/QXFikyzL4k4lSXLJgJML7k2yyAYOcwFrOA5DzSJ0Wg
9G5C9xzSQo5/CYKJjVHcfczP2fsDtBmDhYjAh8KbtBbJ1fJCEH1osGi8zeT7/BxsnnI5q9KG4km4
uZ8rG/yix1dc2t/v7i4sMEHP3K8z2ggV15LlH1AZLsiPjZYXtDt79S5WLbXtN6Vob/OOQ+gkd1p0
FtwhmebGYeiTkEXRVDET+0lL32IjYBrklxM4WxbanT+fL8RDX8yucwrJQY5OR7K2rIAKoSu6piZp
Tx01qrWzTFBmbVpS+5rjuQpR6kmHhny8w97MwVZQBUzBxGkC02X4b9xHtQOWtGO/WpU5kEVtz5tt
yZw11fce85ZKJpvGxBZ2FMt6lSK2yyIXCged80v7o+psJCNCFzg8C9KAiQbge0StOeWurBesxbO4
HSCpmw1QUb9BvGAwFHPeLCSJFAP/C75O0dsRTH3jy8wQlLpKh4AlaQ20EYRZ52ceQUphaetegEBg
UZx1ONSUNPr9u3cY91QU8T5zaiQiwxgj88Tuu3FbmnkteZvNokiyHAbp39OKKyB36HRKWmf24gHO
PtKZKfek5b4IFR26/ix3iY/vVSIxszb7WJ8LYREaPJG51dc9iBTqGyoFm3Gz1Xf8U/C4zLPNBicu
tL5NA9cF/iPiHsvN4L+vtvdxDsKchmmez0l974dSOhKusEMD9pvnHUGvyyHC8QAVbdK1/s2tRuVV
3PJq7jEG6bG65DfzDFGoCYkEBvgXvW7hx+nbEEx22APkELObutGoiCa9wnnOzPi84LyrXfaHVXHK
lFTW7f1F/++BjXG6cmPTFdQdy2PPK+E/xDacds1F30QORTPCUDf29zRXCqiA+pq/pSZUlUbgzv1p
ndKcSUKp5DsYSsTNlXh2r1TsIq/rLoWiOl8AKUimvK2ObfSqQYUu2TjWmOYu9psRMeYByadLTL53
o//rn2W+2mVqfTtsRUFL1r8S2q/PX3LA5yQ2rOMUnAMO8Fxq0T+/A8pGETWMk/k/UfYzB01oYHWg
o7FFkwMEZ7wZ4nlyfdm6UVy3TEG18sD64pRVx5vtvxebNq2Nt3JmJ6d3XLHX0OL7qf/pccxK70nl
YwvEN+uqjyY2qswxSW0Z3fl8mPo0nV25V1bHV0BMdTWdzH8weeNVa34XxUm44G8JA7TcB6hes29d
uLShZpV3/IlF5n/NU4vEcZBYI1n1S15CjhZ6lSvS2ihnYzarsBlZCwxuP1ufyzbv6xx4euiysoOh
MiVkpotdNpFBccDpbTrkvtPfG/PKL8kxV8T0qK8s7uSkHaHeXi3o8BdeCW6KeT/W2+a+eVBuXBW0
zwaOHGsG1XR6OtkudT5IgjHOIwoX9pJvDnWpURY9a4dju73QSH3FWzry+FSTmfwJmBOeaeNVi6cj
ZgE9EWTEP3CnazJ6/ZrKIuoOXb5UiBiBaEk4fjJErs2t6fXCkF412Ys8IXtcnVL03sj/ZYjvOW8K
mqAwxZqZ+SYT60NMAPHJA8AIyrseVkQ3CKLiwPiV0VxkCtPg45uEFN+2OKdsd0gmc+WOCWwf8qsY
2+LfRmWCwnFx1Yajd7pddlkaEnWkp135JCqn8nNA79U2+FXKaLFCPL4Oo0yDhvwy4HCLmqaR/FE0
Gzur1/5662stMbANmlCYd2+px6oUmKCuwniomB8O6ag2OQPUvZuFbCAyd7kcdk5BZV7Nw8oWcyNj
WMxxtNNagG+OVG31/+RrBYzJCQYQWvFTo38RZOJ7iLBZ5+TvYlRVNuHpug93ApVm9kHL/j+xBdJy
mnZUeA5IGtwb1TPRVs6oK3lz6TIpf2HH7ijLX737L7mK2j/DokleTgWZmyhxgX6gquoqfWuX6P6v
rnWU2WtKix3MfcADudChsg3DYZfUDcqDFwML+1Fv3aedMY4HDT0pCYeGR3cgc33zeYa6jFmQg2fw
TD1emtitgqDYKPV2gYZbrkR16oytUUILAwjGolDyjQXGD0QtPjjq5E78EfjvQKzl8yI6qtJpiBOM
OFAhkEs5OfYakaYQzLEtMStLSfAre0+j/x4SALRcY8ZFmoJMgPaE7DLlguvLr+tqD3BQqRH2ekK3
u3GosB8hbpj5iOk1HD/a4DjosZxBP7l+pL2ageTiG7l5Y0nWs2762sUz+A/pEXdiwJMMMHA6Cska
W/kFWSq3bUolQpUtYV23chBWM0n2WIHG0B9tmrAtuoT0Df2A434L4pB5MeGneGrN2UzzrLetfbnP
WXSosyh+6Plk/FhtEB5s2R9aqGDnbv0nOoDfLmNMOwIYvJFTcb7QwOoYYBTG5SVDemjdi1Juvroc
+7dOso/LSXzyo2iBRf7V1q3HkTbpKsj40Jht4WqQm6eew4oCcYiIX6lC+JrVLd4kdMNaiLeqZVHr
W9tYNtvNMI0ZKud1qfNOkwulJ9+aVzY4/S2Al81X/paMT/+ZJXaXolCeXreXuaW6zNzTCS4wn8eF
QxD5CuHGIHOltPPqt9STLz4NC/u6HVTPsN203/cYgEGAACfA+micosaNdeVDtbO+f/Bivvtrvrfv
d7YauUGN5JAwhJP3BlKYoUIt5djZA2PtA7Nax+yrRzp0D9aVdkzjbmXqnrIdo+c1cRmQqUlH0IAS
/0KtlIBsPy9IJkLzHYmIafC9+qMy+y5W+Z6wq7JIi1ImVmIJizVvy8130I+yUecr3AdLXIBrBtWv
KTuXaNZPuln9MAzL9UCYueSiwfFp/l2ahgnlEI2c7bqYiJW0TXCtyU/kJ6bfsWa1F32+uj6VmcJo
0siNd7buaCG9egXJ0kwILnSX+VxjnG5a4MNkYofQ+A9EtV9BLIG9eW/alYh/5gzkigFcoYv0ZP/6
mcABAEq09oJMTUNlSeGveEphsluQH01s/xX82Q4Dw3MKoR9OLExMbfe70+D19pTmKUUFAO+2Py1F
vN5B4qkkSExStdJPa5YxeiFTulJtB40jVTprcXdpSL56f2v02rdP23oviBE7qVQoKtT/n1us1KL/
qIYYX1BfsprUdvwzSl6Yb1ibPxBqmSbxGsPZp49nb4Q89CRfzGSYywIHzvd0iffK2sWGrzwio1Ax
43RWc4RXTn/Uk27Bh8vHHPlOjbl2ejNsYFbhy+MILZ6jrG0tmuZynsDgW2UQ6aQP8YttjJYLelqc
+zl9lgzpZMSSTD6IEf8rJvvKV2cdEuayX03GW2VIk5axmMnNuhjCnl2u0K+bjxR8QyEY8Wq1FgLB
5dTDHgrSwbRTHkjnHXDDltWBbC/6KkQkvh/Gv2qlNGsfaWrhc1RrwWPkb5jPL8cY3qyHm8YcKQ49
kidHdy4xRtodwqSOugSrAIoDMZOSNBTOkOMxXPQx0dqNa/891dPALkmaJKfBuw+Y1N5Z0aMf9Q4S
UkoWeHARZx8IFB5CvvuSc6MZM9Td/Gu8qe8ALU0M2zEGb/qqUrTzAQL8Y1LUgT4fTvPWcj8t85tW
krE2c9BqiDgFOevus2hXZQiHXInZuOvRu5F+1ZDfx0yImyFpDDvaumgvX2YO++o2uo1y3w/fXUAU
9zNSannS4C88J7rQzXLWQS8gsTQse6o681luODhOJhsVHuXLPkrNE0RcGYYeiGSv4ZB4uCBquB3H
eQfvvW1gUjm7dtOnoEv/cTZq9Pzy10nqk7qtKF9/5Ag9JGSRHW0fJUvxccnNgMJ6gudM2G797Pca
SaQQIeemPZifP6hd+CDRp8soEhPDu9DWUj3fPc2heFnys4/UjjyR/GHnN+3Na7wnwYAU9PeooJ9d
fAE+QoxIUcbITMUUx2l1Na6fQ7YokrRLfZp7dZ22VWxydIJJO/TkLvH5IVaIR9venlpiSAe/vFX3
gR5RUEHYmOeEet99lAgAOYfXwBYysnrtqRb2jSUR3QQxY+U6f5UHufTdgugmkEvxTWrC6UVHdNJ/
SOfuqO0ovWfQdoXAWSlyT7KNU4qcwQ7PNThDIhbPj4rMqfl98mpdui0QVHUEGUoUzpAnfx2VlNjS
y0QXmIub69ZqUGRrfXliUISDWoIbh5d3TukqzGDyg5D7FDQ4zQm2Ye1IYmkTAlrJbHuEpHW5Qo5A
T3abnSX34OJB7WLIQMCbImoXP+2wHrnw/9mk8tm/Hl3JpHpaHy2+CkLt6t6pj39vSK4U4SSR7icL
atJkOg7Yju4VOoitteY9bnc2qXtWPf1H6levpqkBP1KC5R3aAYtZr/B7WTgh7/+HloSw9YPK8Frk
wBQKMOmFxzMyyYLRa7mJ15DVt4k7qn14i/AnnZs+n1AxdQ2TnrtZqB5eFZlWFY8TIierc79ubjZV
775OrEzCUKNf2NeFZRZquTKVnYAeuK4qtltTXPrnZgkxzhHDNVQwcrdc7iQ4H65vtJCjJpF1NsYH
QJExi5EJerPgHxWS7S+8EQtgOpQ3dnPYEYe7dXHB0pK4b1Ln/gMl5xJa0wysYiIjppS/fFqcXRe4
wdU9mSH00Yx4oToSyzgSL7ZD1EN6Qucffpq5puJR9HptSP+szWrPerUL85vLXGfAxjjkRAALsfxL
1T15HKziVZYQIbFt4YxAHQw441SHkAbPecUHxALDkhhGhtu85VtKo42Z9ooK0YQqfl2fs5a2zjE2
NxaeGBs3mVQ44Y/tFl/x7zD4qS7Ny7gXHtJFoF9xGp+cQpUf7SikoVa5e1yN2JOkvMIV5vpCfMDz
de/WZapvyVxBqqa7FbTITT8om6kA/D5/q21OblnQLgtIEI7hH8VP0OUeA652af57H1T8Nzuc951J
sxoKegxmZyHxNDUh6p8CaJlUznCkMkD/Zv0KzCEzf913bCvY88Z1iHemlqCtdYgiZ1MPrSto4zaM
qWPExwNErY2YadOiamM7k+z6ifrOhoLqj/F149M8g7ddbW/J4QDBmUTS8bF/tOKxsQgHd/s3jSBI
LV1UeaQ4xZnE11WVXS3DYaUwZovGkex+3cBnZDXOqEFOahN+uonbSSWbvwDOxtoKRDi5uY6AnGv/
TbK6AotWTXSB2gJqCB05A8U6BYuHFWVf/O/ZVCPf75K6+VuQu6ZrSJ2J2s8FrnjQVvVr8zYVdWjH
Pe7SWJot8AlFxTyR0HEv4xfdrq3sfjQTCA1t/YOXAKi/yGCkcP+0ZqHHUUiX/pGSSL51Oeq6ap5P
ugW9qhQhOofgJfx6fUZrd3pH4z0pvPFvMzD7WlMwEz/rKij2NjzBbYcgxGUsRg1eJIzYWAlsrlD9
ZrmDM4iwQ9wjnUPYsDVs7oH1i4BALtL3aUVJ+6uXfSv8dY8gkaS5BIDMk1+YJ4XzUGMZSo83XS8a
F0xhuqpdRxisDptJfLYQ2UcJ0zn4IJGH5ryYAFVRTXNT6/HQsg6papKBRuBjkb6JukQbZ/7PBqmJ
WmYIw2V9pB1gJMeKrXWuV2Q3kdJ4r240mCG8Gy/GZO1U7jgxjJ5Pd9MZ/BQehfX72epVqOfGMRhw
gOV7tGcOkOsSUdaPJRJCDG6ZkvJQg7zYMu4gaL191J8n4DPYKJfQevwCv1FdZzsDDlVfGhtIfacn
BfZLwyyw8PzE9iwRG9E5CxQ4C9yPohBbul+0evoEh1wQ4qV87X+HT3z/EtkdU4vlOJkfxYeWFIqG
40qUB667ycKOEII83J6EVollKtXufdb58aN+MU45keyBbdnAdWKYA9osfkpYfHNi/XvpxqcPVAhn
Jr5B2L5deuqD3kE23mNq0nhNRe6t1qwQpnHgKnpQCCFtnqNyoAqPBLbFquMccOfhaDWYf2sXxOy/
Z4vVxGg7lOCh8hg6rSTXRBCtQcgydudUAbtwaRRULuJCQkNNMrErHhE2nHtZVWvyDBRrBPHTyOfW
vVdxvPc7gz3L52b5tF0WcUlNAQTC2gVtRi7HwdO1hFUXGanhydjkUIW1uJMqsAyP1iLbnZWxPQop
uqfxxp9wh09CMaQkgvtDHym54fYKCzi8LRkiLxbFqDODKhEki+pfeGgx/Tj++DaMN7hU2v0FSoDO
xBQ/z6E2lBpN3LgJOsV9jxNMZfwEmX0JFo2Po0Lt7MwUB8KFsw3uf9GDgj2Zf5CjLAVmlW63upah
wOiHZKiQF5Vp9JGS9p8kPvGeJLRtE/f8nAxbp54VtvjcKH0CdRApp99h8yfjQhQnEDGHmYggW04Z
tQDuFa8/TZmsw7LqQlQLpXCgiyHIy2rEAOobgKq+bsZSrEbd/ibyVzJ1W3hGP8kMorAAQL0WqTNm
g6Miura9wl+0WUBn+ldkx9Gxh4JaQafakQmlIHv/z/aQWR9PB/RDUOQJdC2vcmGbNUeM/l7eJI7s
NySO4SfCYcLvRaNT9kMIsWSeAuZXZiEL9N6haP1whQd+ZDzlKcvFZLgoJbm+0Cs5qcNqsyoHGMuj
0xbOkf2S+xpfXsBgXBt/0K/HMmGmou675JC9TffNyT6rf9X5RXx743xOga6186fAocjTfx6xagjM
8Kwyu6Pl12g8Vhk6ROKbrST4lxMhCoISNTf2f80Hcez4e8fkbC/DPY6T9L5Oe+sp78jFarhvj0ec
nKa8MC2b9qtnVt30tSwHhgnGOp7JHkAzJWhJMtULPyVA65PSX8n7cqWHtNYTs+506iP5xIFBnbTf
Rnji8WvUXF/reHQiF2E8b1Yaqpf9amUilXXWqnTL9ix8dSlAfUiEKX6rljKb98TyqPSTpIufzso2
7p6BCSQO+Od1ET8tZZ6W6q0pkji4K/g2CCVqTjeZHcpC0A7O1GiptWbVguFbpcbyq6vYOsBIP3gd
od8QBi6t6orBr3tdei68zxp1nnRFuabDKT+9FQCkdc5gotVhSRfjq/j7IuzM/4FXoyshykCLOOgC
JmEuz8vRxsghTW5edrqy1SKTDlutmfgR5tKHBcG5xhnxMxVBbRKNeQtac90Euq8tqNzOPiBDw+nf
64EiJHHsC+EY3dVgLGrBIBHLMllmSwzlA1Uek6C8yWEo23FlAZmhD7dRFDLQSccmQxd8uKK/YDjV
QZPJlUqEc88nbD4srpi5XvhqLAC4KQKYcZk3DikBdYCFj8u/2BsIq2N9tBogQlbtegkL558lF7/T
2Rdwg13x2KuTFsNUuQGRDqbu0r9XdjSPTJHPEe0Vy9SmS33HRnFqu6/DaPRqf8QoJrFC7G0oQoEw
ZpW2c3NEOyF7OKOS5tv9+YNDZrxVAIBTUeI2GASu1vRn1dv1Yzh81IbCSuv/k0q9HvFEqRqjVyCt
s27HqPCSA7VKgsr/Mk8WlWMdAytsYvqSFcbig53P0ulW75n/UK++WUE3lQbZ52H+BWRlLZ/n2YOK
TPEokYmrbVCImGZb93vhm3J61hxu2WqTe5XajgzZVv3DFhd+b2b2X0mlGxZciBm4X0EeLhrSD4Aw
dJYr8mMgHgm3cjRf7bnM+rYtsDNAirxYGsIOvI26E9+WWHb9/65Jka1O5I3HwD5YkIJ1jbay4Oc6
IQzbhZZqlgy8/395RXvJrCIouQGS2/ebedIvLyP/RTFKph31+d8efIWXeuLD7M0kxu92WnVlaxkZ
H7xUaYb3SeZ/qCVWe6AKKzMNeqEBqv0lnWd/Y0b7UuA1izHAONtnroa1NMY/pTgIEt2dIdryoya1
RhRIk3R1O0LYZ+RNOICFZleG96sQY3n2Z9le8aA2lXCJWLUau/V4Suo3IaMZSADoEGGUjVkaTlEH
KhW21E10e7Gog/kTIWJI/T+VoRocSxJfNxMAyyAFFZpnLHYRVFBXmdBBLGhCR6CCYaH40kU1KjzF
beni5I4n0Qidv/00phPICykiVVA3qTEjbexZsDd9ucT02Tahfh8VjPJKSWrPgVDCEWjWNrk/0RKK
D7UOfZIfNxn+MDxjxJpnqhwOJPU8UAZJdt+nJsCZSwAkSe4MSfjaBBF1RXtOGoLZ5WMUbzLGurEZ
OugaW02yE3iqsSVQrmxx3XxpfSRZ64Bolmd2awz3vJ34Xz34LLLktDzcenUGgI3xjFpyeaYVb9qx
n8fTP/eul6ynumQV+XHIC4x2ofEJWQYuDmpB2giQ6juCNykZGd/dNl7ik9Fjxv3LnqMMmglgm0Ms
Uy+qDpOfhV9dJBvndW6NSK6abxias3aWYkKeEMb2CDM9YXkrnUXzaM5giou7wxYUYksb7fHpAhRI
zzFgBlIT4RqzrrwnIiEUYcvzGADWFHr1MDhHa2FV9EdlFX/E4+lRSN9yYdvsvH6jbP7IT6fzQwB9
oz5du2J5hB+xNDJCiLtZsSJZ2I/v1QSNErm/Byz77KkBzTrWa0V0SV6N9lDDgdYX6QJvt7BWle7n
6fTwYKfcglK5CBCmVBKJde+hEX10ktlD+AWPNF/XV/OlARC3EK0hjlP+NjNHvSOz2Pa30gNBFjEF
7DFjxXbODCkSDNnu/YVB/39qLFiH0MF0wwyJGRZG7oiYxFke55g+r3oqmYeZrI5Is/NQOjPBf+pz
0Ru7UvzTRwh4It5n0+MssIKA5LgJ8lwM+YBAK/JpaAgtxeh8BRYhUzN3vGhCcQOOWokP5TH9Zmrt
Fp9v5BdXlMNqVlEh/X+Hh6jOEyEUmw5HiXtwZefZ90xu4Ub42VgSovrTCyivxqkZzsqYyZ3SszS8
cOE8FYh/LHKBsI6/+myhwqBcSSpkItK2B31POyJO0gYJkZU2DagonrtQOK+/CcUjnq2AYnk2IUyZ
/DL+L1ye8/XiIMqIJ+Eg5TQW1ytErIYkfV4zw9nQUHUKHe29Ssx/ePKx973wNwn34TcSpMIKRVxH
cK9nOZAQF2vmXF2oD74/V+njMkAFc3LxtUVYm4oIxv8UhJEbwJSLiVOTWAWR5vuUWXg0S5haKN88
SZVrF/QufTH3tlMgFDHmhCdB/InRP9oasgHmN1U0XmdvESsmryODKtfIh9essQr9dlie4sDnV+vs
HwDTlr1o/pqGbNVQrhpx761NAzdHGKdkxQymf+GmVhKh8B9e+rJDK8VFxuCZ5c9minu53Nw9NLYS
Rnyh7yi9LxnYBVL4qvcctQk9Bcx0DAYwfmuZ1aTCBfJfZcE3tZpGT9pM6bnL+GDLym+HfBeAtJRs
KxOjuR/zfOfRcl8dKtLHRgedEd7l8cwipw/Ca/aeSpoDb85vJDrP1d2XlvyYw8kuHeH8jA3S6NJD
lc9mC/kuaqXJrzM9vw2TV2txY7TgFu5cRcbPtvICoIzGRgnV9lbjBqNkxbZ9C4vwnB/4sU9t1A8J
BGQblnZZCJcyOmSdeT2Mmto1RLct10NeVPlheu6GWUXkI0rd38DlQc670vSxID9wuyTOAMOknzuk
4GJC3X56inCQD3Q4GdZBUk/kn+5OL5/52nIBQWCo/ulM4hbcTmXyutzp7GZp4UV0i1ugmpdzmZnV
uYpXf+MJ1SANGUFVvVB2EovaJUq/1QONAFNBjDsVH+Jrjzirh3LSl2aiW5XqytC6g65EpUoDTSzV
mNdQHM8X/J2cfGIMRtRTSe2sp2MlKOGtrAVrIqMRvytFafUdB2ZO8I2vIRTmXNk0WXAWG4U7JThT
G24qK83mTbWoaVdlyWwNe8OESLIx7LFVRgYYPQOH7e1EzXdHbTBuZNm03Alcahj6OfoETJPNc9ZB
UZgoqOAimeTHQddLhCYoVQgRbE4KMhaZ6i+JUFuQnvdj1m8jcDviDRmaxyQ2jrxjxLpHMMMZhNLv
w5YAPaMHyjg+8px3cFQfWOFrPVQ1AepwiHirgWViFFkE/27Eu879PYwELMoyuRZslcUurs9OJ48A
qiYC/RjdL1oAsoD/svPkiHGPYQk4Xus8Nowmvi1h6lNukMsV+NTmgmrMuP+8n5l2EIFCq2Q8Uh18
ZvibHOEawYCDtsFQ+FQW/Z3TWmIsjlD38SwuhepEEHcdMt/uIVUP/hN4rGKVpdpm/RvqjWJejbs4
PAWwyTJ0AFvUYhUjbnamlyxxdcYvli8AJxzgrbsMETtc53UF8yDi1DwY5SWw+nZE06aMB9FVHwwZ
FjcCQSwhi3crt7/9eftORCfXGuRCND/Jaiq/KRRUUflXTalKuJjhYhn6ssHct12x3sc/f7RejG1w
HvOjGthFrM0+PGkqG5orr4IeYmRXEWUQ/TN7Ju2FPN6Y/uXWq/8Cl3NcSB6TEhzc6JKx5BmDcM6m
+1ANGIU5XhwAJCBqDpkLerAkbwSWIeKWGhDhR79VUy1o5E94XUufZxEN3ZxEyqeG9jXSINdOUZn1
zk3DtK2YdOEhxCyMoJ4cLtgGJoCCuNs3crlF0FdCwcC3So7nl3dAoJyDmssiQuruMwcSb/DjDRMJ
C7N6eiU2XNMnvFtyOg/MHpQk2BKJ1kA+EXSvEZJsKA1u9cxpJjROCrRcLDADrgNUlLVlLvklp9Y3
J7SiWBfHUQg/zNR61krj1WdmBsUrGRsK5+8cV0UTS3ikDBayPz/GuFjaQ783oAR4BtdxyNJciAHC
jHpkRYoK8engN20hTX6goM2gaBLEwEkEvuJikhGAMd6o3eJayVVTso6XbGeU22+EWK39NhJCXJ+X
Dus5Lj1XFcx5JLd7DtylEjpK6fkujruCQmFs8wbYFzpMqAPfY8S18fKPmbiWm6xG+mkH2jDWwxxs
8kD3owUbnYb6GH8kP6q8AOo0PCw7or3VY7rQCloKIG3SUo0cJoJlOSX7/qbaQJ2Im01CvJXoQEWf
4DWazcoZyxcjzqisGOxsEKsz4M7Zita57DJ558++vrXpw2Ajb1rGoBKNltzfolrxO0aPdb+pS8Tp
bGl8a+GKDgkJTDQVgrWmG4D9/5TGS0xB7vqvvDX7arCal8OC1mNaamuZpjPSOGCvbdFIkxc+i6Dq
Jmwqr4YqjOW+Bl1alPYhl6BQEvsol85/7FWgB9at+DjufZ+Vtsnda4JQUG8hDZgiu0wPobrpLD7l
f4cGNQuC+oU/7EiHIJDklSj447l8tWLMjQpd/9/pXlEtN25CkvbQo9VnrjDKydCmKzH9oOKiJF5j
zcIoT4KJoj7yWKT8qHmtl14M7Tx2e1nck/bNFKf9ddzx9GjvNN24Q0/C/TVHJQ/Qarbj/wFrV7Oj
TSlLMMYIOMyiAgdZuitS0JksYjBBtH1Qd6WEceV9V+BR7MPdLsjdQsW+i0s6XWhEwyvqrkUwRMUS
4zOXULmHqMiNU1LX+SskYboLO0IyJm8FBV6v7qtvdBSd3A0rCaoRcPTRyFAGPmHnuTM24GyTsG+y
KM6+xzqeqR/vTy4qKFr0+D/AYKq3CoIzYGiEX7BajasEHiUWH1iEL+ZePI3A6zz0GjdMKzGbnPpE
tyQ0sJEVG88m0fiCqlUXKvOWkQ5SnSCLp3Uf2v8jt+kyFEAP5y4rTUlEFz/cJTIo3JxxM0B+/Tgz
lfuevG/DmozQ0B+ro9qbEviO4ifU/6snglQQlF7CAGOFy3qiDYZcvAUSNrrSy2VUFWN40TSOsvBF
8cuxuJcUdcIDtGZMhlEkyiEAbDXwF8S5c0U8OlHp/hY+nzPRhEtrykdY+5p3+liLDoDeHy/uuig0
UOE307J4rGu5h1uADGKYBCM/C6WvHfvPkUCGLqNFyHisKtl5FX8FVZ6x/VhFAiki6k2GFeZSFkjW
D+ZRtn5DwUOOXX0FJpSUQ9GG01gRt/VpULLFzF2ZHsl/S9lTcj4Y6bxU+SXPGx8T+rag6SFYpxgC
IQGBzMcLE8mTtKJw2OQ1FbnlS/lit7A3pScCMYcs/Z2x2suIGA6Z6PVtniCABIoWLS0vyXevven5
uWVtmiEioot75m9ZAsoR4fwBdYd+kYs0IccgVdKRcwhM12sg8j3rsb/DDKdwad0/xllDQ6oRnrtk
BxcAPbJwQ2h6O/QMMiKpwyvKhTnS7SVn5MpUzNRZv4aBbppzuCwmaUXrS0HV4pEeQ/JdT/kKOYSQ
rLEoDbiXIA//fLgpTkazJS3eTHPAWhU4iV8sOTZ0CUCjiFD2n/AvcBIgSX57s6EHhQFoswnQZQ4j
ePlaa1jOCmHhVaZX2D1TCGHY7mg04lHKJ6/R9v/5VBZL9ea5qPsy7Ph0Lzn8PD+UgWWpAeeeK7Sk
FS3DmdGgb2SkCGcH1fomOkWDA2m4AKsMXcuAYXuGZWDCH/HEtNzroS/Uy8GiLNQtM+ZNjNoJUF1i
yNSlQA7yuxz8VYUrlAIMnwzLO9JiiNaaAPgH1TqPrurjYb8wAZNNIKZ0fGzoSen88uS5JTeCJ7KS
j3iZL8sIc546z9Rwpo5gJyBhWSCT3zjYaCMz6ToxnSO+vUnQo4X5Tq1/6kss/twn7PFSxmiNh63C
fVAQSG3OX5De2na9r2TME9RAmTd+/LIoYFFgjSUNH6wOdhlUqs3LdxntSPRhChGUz6nwKwjmARlY
tmy2zMC8zNZBTROp1dXy/bUcaharHxgNRAKuZNpAF1O2lSHVi5fdip9SP6Mxfd2GvtqHvaS+j7U4
H5rpiF1ozH076cQqfoWun1rIdv+jVvgarK9kTzXsQ+c/UuM8Ozt/sFSjMD79XqCnt9A1SLnIXLBJ
ufjfG598XmltyhOU8D6xWeFxNpAzMiVEfq4IK2T7d7JbO/sNg24k9Rpb+I6PULoEkTAWe2tEHurK
taKuzZhxBMeaTwg+MHc+oLPchpvBO6C8SRqTDaxFriR9IFXvUf0ccnx1fWcWMoN/r5DkamAW24BS
SJXPC6h/uj5DMlPqHk1jeDLakAh8Ub1PKYBxk+Uk2uQ575WDFqoPMaG7ELsyFAUFvn1Ai5ldCOCa
eqdgFLMK7KnXUN8TblZsCoyOFkCjDPpO38HpoLYGGBRqukQbGSDD7DVGe4eUX3yV3x47YpDuLFBc
TUWQQvJQqowTfFnDLtACkPX+NmXVR/eXaGPhgIyNUPI8xD/hU7FpC3xJsrQ0BRU2V356GvIlY4Qt
zuSr5ai2szdhtsURMhA2xgEc/GQwB/AmETz6B2z9YuNlunmYTFMF6UjXOZgqDkOQU4EtWwweHbgI
2aPBwosTj1e0OIiFcnVLaESSLz9P3QdHdB6pfcFrIs4l2KiN0Az4MIR+VS7CiivZI9AJGub8Hf4b
4A/vKrnBrnO4prtL/uNVqSH5yfIbb72JdX0gt9kl5cS0qa4I99zo5z9ZmSnpQiFKZfHrUXul72li
BMRfWGeAUj1s6uZNeHvoGDAUVE2dvZbr7ftXKSKhLFhL8q9Ao5gAHFqwu37MXf3IkN5aELo4aj8H
eY4I0H9Yi/jcBlALsgN4RIa+YnZ3JnwAUi0GqfyS0NacC4GcRU3OOqwK8dt5beFoMZh6bKPXjiGD
zOqYjdOdUSUV/MEpfnDJG3cPdqiJLnR7o6XT1vGKFyfZTo8H3bnpcNXxUaoG3CaJrzGcntxlTnhv
MIUh+G2WN0+lWBm42ydluc3wqoLHCBjLeSHMrgsguUOfgUOAvfCdz6Yqvb7hh5xXRSAfm+n2W/+f
JuzmJjpaVgU/S77MZdtLMEWSfI0Fybje5szUmcb4AfJijQtSF29kADO0OBpILsdT9IwuCH2nScol
KdYnpMROKY4DYAOZ/OZI77oCt2KD8+NgXMZxx3OiDJBJX/713/OkRduXo77SlRJ4+jpUzx333mAI
mqnSBkjs62/Q0qTk8zbXPPx6NOaqhKZFvAFlofjfH6qCf3Xgm15qaoQim1hOue+MVrRncxnRWBog
X8AzHPpod7bFEzvip7nd7T9rj6eVvwQAxO0JC01qaebOb986j6G/QuOMT7k4gyZES+Ah0uBTWcgR
2v0OaxNONIycET7Tz/hxLZYGno//9AlYfJiq2bsNmz4i2zKI119H9CVmgSq19qM2sXcpd72StCaf
kHngiuFYhqW6JnvPRqT0h5vkHWMb6xuENG2rmJf5aVFXOb0KmEaVofBoj75aBZmhp//kEZlVFKma
pImIE34rhRv52+yxd8cVFXyN7Yd65KJEi8WvNP+42JvYydsnfM0zXPM5TOYxTFilGMkiFg2+Khs/
haV8M/cM9S4UTw9r0u8Cjr4UYN7xjvg6Eyfk7CjBO63SCIVe03sW1TpCOstf7rZZyouPOAuYyUgK
mco90ZNqnO3DvrLgEzB6nKv4rDpjaqraF20vD4ZxSfKV2MdhOI5QZGg6tlojclyvdKFvTJnfbsLP
Eh78NaFM0Mur/AjcHWD1P/fOm34LgkeO6ofmeWJsE95AxiSjV6epsCYm83Esiq2FrRXOwJSfm8Zf
0fFS3lrFUjXsru2D37N1ftvI4aicGCzHUFo3g2vPae4lMGAAsgZ9vIqsH8iAj0Hr+wd1lrNHjS7n
O6J7shK3GYs1Fp+45x9nS7D1FZcOO4+vaA45CzDGeO/9GgyvQUvJtqqsFwdleqevpaCDkx091Gvr
M8iaaJW7UIwW655SDxfONkjdNNoKXEE4neSmbFa+TC0zbVsYuti2hAVvM9oO2JZr9t+qSRnOry1x
eOyRJkz070PFbK2oEYErin7VipNt3DMyXrCavApW8DucY16P6/JdviPGy/zjBNn9yY+q/MNQddfS
GSBI/6P+q1X5ZIcAMMcyi/qN3X5x240sRc6UQWiBWE3IbxFBrX4DlA4ghJu5pqY58GtjJlmGhoLZ
HlT9BA5WJ31F5VlL06n5tpAN1aGOSQ3kF9YDvuTA25atyIiQaGlW3ejR6r/neG7oFajIiGoy03ix
NaVK+3FDdzvbqyWlAEt5/MkFqZipVSh4L8UGaQ0dGAQTiYMNSTxLN5xCrDU1ngx4hYZ2Lo5O5N3d
wOK5+3v8hwRDCefe01pFb/i3QKamsv2wb80fLQhcaUmzGMRIiAwwn45WussXh06IbWESNxzUbn+w
+SP5WS5RQbWh2QzN3Ep7PA6HZ6aN497IAicHCpTWzZ/g7SbJ4z4OsIRqDma191T5IoVorEN8jrj/
A2AFgjO3ZGyNFDpokQETp91jX6iLPXhr3sAOrwxRpI8LwXdTFqHRrfW9q3bBAo1egAum8SNZl2Jl
J+vDQ2VWY0jV4DllaezfVYxVDeNMRdc3pfMQ2XlIedLUZGghDWG1GrikibvAfPc9WECERNu7BqUO
W8lTPLr5GjEyjLM1/S+N8dKaLlX5HB7oLDJ5BLpd2aG+9uQbot3sbo140OPwoCKumHLIP13RPp/8
yJpJ3REkcSMLWnRez9nK+IT2SFBOFmQQU/bh/y9avKwVZgrhKKp79Km/KxYiB/Cbeu2m0VXD9Os1
nL+N0GbejNBrnZQejrm7osfhw2vz+pVmc4+UPPyl8ZZ5bFW2UG8ifyx0udDqNajER3g5Auim2u56
EoAOejH66yOnVsyb9ILOeGK4n/t+46Q0W7OfHmKFf1Spu4f5GvUt+bBJry9+1vDYuYp8PQ2rTov/
pFZMgQHih2gaMzKD/iYHya3RQpNeDOysvkP1H3fab8Vs2E3xs5h2NZc7pHHpcnB4k7L5nsaRugO9
GhAcoZw2AiDfWMrs0Y0RVfMdHHjSNRBJES5HJ1HvzqfsDoCx2V4+p64oimlxEb7hrWJ3TloOyI2k
y5R1r0WSCVtc5SknZN45YLNGXGp3+tF/myX4lwAfgDB7a5mj/82C6JZZDuA0Bq8KA5wjLpmtgRtD
gvVn4nc9o4dnI9mFHcZX8kZkoZLaMJZy16wCC4/uKrJvovorzx6wVH07EBxxGy+PbfdTatEEeFx9
fuqViWST14zaEU1pOnGyzii9wowEsbB0vf1vk/bAbcDCP3i05IbX7eWyIFYaQp+voxwDjJn7J0N7
vdYpgZqWh4vSIrb0AV6BtXyWiyVTHjV6oQq6IhLeqa/MrflykNyFBw6XZUDfF/MIJ+bGY8+xAFBZ
EpOtANi+vsx/myOziuHrpoY6Wbcnk5YI1lPYcaKHFLCZOcj1pHSZGsugkYCgH2zIUbOKp9G13stq
Nx6hG27RXq+3jc83Mp04lxADhBouluqTZhQROWrxsE+XQJ5l5oEWksAWyNEXDn+xwvJMLyTassdV
ZcPNhU+//U4Z/x1lrCL+OUPQ+AKLk4XLBswjFX6G5TtW/9fSyJbdkUtX98I63W1IaHq6AWSsZQ3G
c/25GO6iLaTDGdzonDULLkMgMGg1J81KbhiYTrMaJb/AzhQtDidH0ozuGBPlCLANsCWbgXI2CMOz
KVppP/1ipbKsy8B0hwR0epBul+IYqJTjQ4c1YN9hlS04I4ja6tYQbQr42L1QHY54CpUdpWUw/kpR
A+hp1B4FEIfA/OuQdP6v3eGwtcmu8IIZS42FpTLRBxRct1aSLtsTLVgJhAtwQEQ04ve49R5G40Fn
YzEUhSv/bkPTHLplBb1VbLvwZtIX6kU9g4Q8lF95EnL8/e8TSzICuKL1b8xWxmKkPgn5N6ae82Cs
qJeycZWIxbPDqBY32rA1YIslzMqxlo1b6a4GdR1w4YPCxNRUetsVVEJ9Ln4kfyCqqPPlD3vqMO6a
e1q0ozuznqJun1Wr9vA27MYPpb/6j0/foHv7tf7VNpJUsXyVR4bqydwab3avtQh3Dfj1WmOA2x+v
Kx4SocrkfrXcVGOZiKknXYlPMcwLGVzDiUWCqIW3fK32c8YXN3KJwNsPMPXV8ItMVtbk91LWC+oh
Gpdj6g86qXJz5LPi8YePpADbmMtA2jWBpuRmep2IprC0Sb4i0ZrvlitnLxDAGNq8LNriHdCKB+N7
mLiC/p4spS4RXGQ4B99jRyD84395LFFyFPQ7uCbH+cFbJJSLTjGuaRrRnxbJt+3+evH77LNPkQLu
p7a+dSWSC3cWvM1dFH/HGyIRM0GuLYLjgx/xrxc0gMWdgiDXTQzfZHjFrgMR5nEB6KBPCT9vzcfI
HzjDsd5B8Oj61+NkYC64GSBMYaG6Fqzwobtbwee0DqKODrsniIgQXPWNF8TxRcgM1VekA+g70btM
AmyJDQjbC07e/+rcVZls9nrlxgixu2P8tvgk1jq8iZkq98g3rQFRTr5+rl7WbeI6hLxRZPELVInV
0FU1VZIAV/NSAbly1wkFhDg+K0rKhcCTfFIHyky0r4Nm8fgSYB/4eN715yyitgHERh6AFvHu7ON2
qixZsFRe18nkqNVmHLNUlieuGJDHA27h1/GtOr383RjnJmD4QCNtnfVL+ajtLvXaAKBIPxXll8wj
tJPZGYW/FGIrtm34eefnwIDOEZYaMbt9sVhUiPggM0wBIBxWkaUf66vQi0xzf1eo///YdPKyQ1hK
mRmwXmD+bauPC809L7HtUSueCJ0ZJwLTyVpl6SYVI5iOAjZcFi05IH7YmgvpqhTGqzu3HK0febfn
cbgqkYAMNURPiRf+CuS7CV3ecbvhcusu5MThaZ1vL68dPA59MZGLM/rW9R6fn656yqbw2UFjbb6/
4IoHBMZFWaBWK0KpIkEyoq8qMRSYps41wW+HAd9PvA2lJ6sNO2VUdJ9xJneudN/Hf1Wezp9/gK9O
aCedFPSgkcXFHSxVDM5hDVMoM2Uv0loqa9pNtGlaec3Sou2K4a/G5uPiozEzKOtNjHPWFa+DpKaW
kQ07DJv2v9Ry22iBL7x9ss0yuIFYtjibu/qdCXHyyGlkO1BoS/XW1BEo/f/8fQJC/WKm88DVR1ki
omY0k7OAeIOISv2PyMFdAbrLHhMNVzdzmb6/v//YoTmUkHw/Udz/nZncPAvW7MmYjKwdgGRxqEly
DnwdkNo3ftcueO36r4s+qTAO2p9visKEa99wt0+zhh4WotGGG/7sJF+1vkxcqTrMywPgwUzxi2nk
LBAVutMY6r7/QOvw0Bs5iCxniwJGWd6EWaEQ2Stg42vFrzk4jX3vIKqDRRSRFCTdck2gOc1xhugB
zyKNPGIB8ZGu+UzeKm3xkyM76os6V9h72KbRaD3Zyhs1ihQFOL5BV5amLuE2UjAxYhS9DUHtITDr
KGZm0lnC4XcfeE7aYj5UuiXY7fdqF4WvJ2E1m3dOYaBE2f+rfZI2CvhSdTCfOgWcGE4ACmdho/KC
YpScGi/ENK1OXW7mH2po7Pep2UzgEadNevkGMaZ4grG6aJd7kbsdQhzy/UyZ2Y22LxXeSSwP+QPL
NxqCPwoBHcQ5Ec+WBGWUgoOWYwtsP6GkCNBoAtPR68/uGKZ0A/Q6YCJCfS8bsmSKAF6+Vso8LD1k
HWvhmC4XyY0tIJe7CtVNt9O8DwsInTkJOcRnOUT4XzIiL0mrSALe3BAD3QK4iVSoK5hZev2i0Q0T
7mfZZylu+Q30gnA0YcK4yj55tnYtzWF+q2tuqcjSeEvHpIbBITA58Mh6IWWRBIEDyH/BLDYCL0Av
llwtEmy+myBVd69ufP+aVwXA0VtNpfM6TTrFN6OknjrFhjCAgL92LbMcc8BLIIWu4rTbJP3vKzuz
mGYlujevKJfGR5mfurs2bmgOeKWOBe9QV/CodhAIHCZIyBhQwg1dZ9ZBeMDwVKF2JEy8BOPP1iY+
c5vJ+FI1L95iDMZRffexFDYf+CH5Bd9y+yXlYDYWvUPp5s5o6uN8+XrC3sx10+6kbUJAFsCHhKuc
aBpai8zFEKbMKp0jCmMIr2XtJ4yJ/49AOWP/5sZ4XeAVaMJCaFTCctKIOpGlHj8l3JMDrcuyTunC
Ab4gdSjy6ap5pYCqVNTGNYrMWMtp8YnJmvNj6wVRhdG+w9rNczlFJs+vY8AV+HSo5Tfd5ARqF4+W
cqRYLTvXzeemwMqK2qwG+4kW3IptqOZpkZlayxVd+yAi6czNhz9w/S5cQfsowgHryPLxQJa+EAdR
GL2YCdWCObnJ1wGE5nYxheNnJwS9Pege0iIPQfd7Pjcuvu75KUUxZG4IuDzgfiMFFraVrNEp+IO9
zsx9pdnRVTNaRL2UzhIxTYuUdLQ7Dz8oLy1Lje0fUAFZsj9a/amgmbcawUaRYhot2LFFcJrYKjvn
PfpBisc4++zrxxZqTV5cuDIDc9OnTa0Q+cawCw7qbK1kskidxiMOERTO8ohkpHvDsbZlEZuoxr6/
Lu5bAQgdqPGV2zZPTOojZab3zJL8oh7tnIK/SIAN+WnPM0qvu6jrLsx0URxJyhn2Tm1ywlUNEq0r
b2cs/ybUAIz85Zgj0URbOe8aC2HVpivaqUbxX95sG2Rn2zfEMmFw1hjzMJWqfx2fHDyBvGccoDU1
p499lYboiGT8S5aiurBJ/yGuNf/U7xFPdwCFH/uVlg/LEqQj9PclAYAoyuFppnk4ntEEUpxqq0CC
9ZQ4PBrXpH7/W5NZlvzGIIxyifXs0T9hWPDqNCWYti9v/A6LeiaQQSoK4c42tGFRDpzLBRYfVzUg
nDriWSzVf7nolSaeQqGQF2JDjslV8QZ6Z0GRZMohWh8LITh1X6/FEZxqV7Q1jfqR12cDJ5zhFWz3
cUjlsp2YKB6YQ+bOMX22utmZ2B13zX2z/mNOD7itlQAE6AqyBTQ5UCYTMfrklJJ+zwqgHkyMB0eu
4M4jA5jV0FLtzBxLVaKmgaNeejlIoPAaywhZ+r2hHJe/Os43m+uHt61R/jUJHJkAo7hszQ8HEGFL
itPK9fUR+htnvlFJy55Tb0MEdJQAWgYxamhn3a0eN7DM6yp1r3/mXclquN5eygcgyYmnakImxpVw
jc8h+WP/JPR6SRgkL13fTv0VvrKda+eHqdicxVQJdlHEBXEO9LvKWoMZCfXr1b+nFq+BSmSLBvJq
NDVX4EAI2Bo7wvQZk02+hAfxYevydN+ZRPm5XgULWRuEC/lKNSpm4hMTuY8CsNi8XJ9E01bLmCKK
reGqYsOMH5OSpLFmmZOA1wfhSYrZfgtdwi7WbIvKnckwARJ2sZOC7ejSCNAGTqbgleioRQgVfmIX
T+SqMUf4M2YKCU+fKSonQvRDJPRQZv3GpdDjs939ycLTboXP+2mIeih8XrHRvRXU2BjhpB61kTCQ
IrWxDiiEod+HNvguwnC2KdGKILELFN8kOedhwUQUR9KybS4FExvQMwREqGNR+xOuDQM8TvBrpzM7
/U3dJC+lJr2Us7Kv2ciEMknneUP1jAu0ADHadXBq5h+ANG7vlgknLwpEZ+olcpploEtNF+LDyIKr
zHsnSxW8+xpKHxMcQ3jx+7+yzKO3Q6TpYjii/tRif/WzUjbuMwtm6oo4bGhRrm7CRlkHlKLlKcR6
TDUWmN83LB2AnaeGhof5yt+gDxXnx2az5VaceC56SY8iCE2iQTnE8YcuL4ZRv8TFfsJZtl8QXt+C
uToVw+HwqIx4YhMxXs4/50+/Tw+DQEm4abzFCbCl1govgtfk/q2XNTc/UHS62CEmZ7U31bJxbIHr
eDMCxB8X03ddjWUDfKIKu9YmBrtN39+h9XEfPPD9Upuqta6ja5M7HvdDD6hgRe0PrekqveOfI/Mc
DYEFFj/eF/NTAIHD1mZViwE0arF+aUPByI2Peeywm9obX9XbFypJn5mmXCTYyU+9fIpwf3m4nywm
BpZ/enbnT8varXxBkL41lD/CaUC0jgIJ56J161faGEV9kRIljdQUqmKPeMBcEFIVXvJ21vkyEqIL
AzbaHD6TuinrhKymH1u77CoF7WT2O5uLAegY4IXqmUV3lmWltjZfoSN2QnZmu+odeYX2EoiAU/ww
Vyacht6f67waKXlq1ct0A5yQyT9jPtWZzaT/smIUekANJKWi5U+6E28JSkkA2Z+wxOuYfM3xeh9a
XG8mVW9gxiZOmrkdKAM58A2YNX4D3fNAN/DZ3qmjy5fW2teZGDhaV+S6O6kVJAVYaeBorDfbytxr
HT1swmkxzgygqMWlenVyIekIj+jrc2yJFEYHrVakTS5yzHjxwY9soNmgCEGV/a3fGiL0EP280/zC
f0YYZ4mR4R/y/Nfj5EiyCZ2RB65vWGMv/POeyGX3Je0+WdNJu1JsmZCA7KErZOGhjg4vumwTU23k
umYHjMMzGZhPWk1S8E+YJKoVf1BtjloI6suLBc7aCEbOKYJkro/FyaYHKSB/+skF8j3is8S1toue
FkrBEO9IOJ3hQIWgpdC1KQFSHV1F/mMMsHYmF5PdKPj7WNRR3RDF107TnDU5Ow74uF/x2GCITOv0
eVELDSPLgL/XMIYaUdCx//zJI6UhX4l1d7GjOhhXJGx0Y2I9DXVDIpZvNT3/B2IChq830VY3QhC3
o9DslsNiuWwr6DHm1NkVB4Z1/iOUiUqLpxt/RYGcj+/mkDsu1A40fTPHXK7b9AkkEMLgxf+BCSsK
1Kv0B/NTEgx1r5DOfjXqsHHhwb+AsBEzmU8rg86hSf6Etws6eF0b6OBce3QhbiGj2Ei/Lj2kBDii
53QxfcMDFqzrRjY8LgUQpgviP90/gX96U49lKMdnALSKqWzpQTWOdWPJLnNhPCJ9cuV5G9+fslRI
7BuAbKN4XWh5ZhWOnPO58g55XOP9HsO7ssFPNwPekzEcUQn4Jp2LxDor4CG95Nhq8OduqMRVB+As
duw9axtBO0JcsO1Chw6IMpRi+yareC7hdvHspsAchC58vd4jEqgyKcqHiy1+UVMtx6BgHCPcuwlh
+VgEl0t7txMEYBZklFyudT/fdc//CMrdA3xWSFPh0lspHWTJuwohe5qJNUVAqRpNpZGTkMlLeVoM
igNUipdwtXdRMBpUCjQ9UdnsJ07AUdobsAEYZni1htLszvAkPkHNICPjp6pZnsmXg6agyBDWteDW
yYZ9UqKsXHl/LuAX9SBsVystQfaQTLOZbyVtFIvDOtANf0hgu4rvp45x4zHM92UEE///Vb0ibTtX
qMHhWvOnT7LxgdNTjxgT9YeyifNukxUtNL7EM7+DwCwObZWgUnne3jUJXvVLNwqkQu3TSuokltvG
j72cF1INcqFX5MsJ7Dp6g44zvVEV8pghAdNOyvvw0KBtstOnY6Mo+NXQ36xjNOMopMFuHadNHq4K
3iQBGlH84Iz4RFRbDaP6l1NPBwLzEfNqHcjk5eZXnpbzZ69GaaRMczOONQ/aqcoZKVRrL7T8kk2h
PTp61u9U4MjxIQ110j3hrJV6Pm9Y8uZl3vUPpfDWmoeRsbCW+YPkA0Vt0kpviQl59Y5XAK85iwVB
DQMMAEtM0kgXbdBzABqm5XIs1xInSTAPg/r27Ui1OHD+PkYXHFFmBvlDxMA8GqokSRmCH9X8fp47
HJ/41MCcAjCM3gvclTq4lPotzN9CsJgXZ/DK9DQUZL89YtnOZPB5olgc4oig5B2gy8DgpW70XBT3
7caZZp2D94QHNweqUsx2ShQY3vM+oDPljd5/UfgBI0FSwKQVkLaHimUmrztu2lNxzMCnllKvwl6X
Ep064fWydDQCR743nP5bQgF0iQw4J99/T7FE78OEGjkwD944c1NCuOJITug72kcR2l4YGFxc2yEJ
RjwEWVWXAoGJGsXgcUqEpmbC0krhZxDsPOkNEi56LP1V2ZEUYdPWxv+/HrtjecAprmC6UyesZ/6H
HaCQ4vkyZv8cL2shtLg8mL0rFxTUfCoWygi/Tm+uJYF0T7Wqflo4KT07isn7sCCj6QHb6mf+XMpK
cwuHn/fxFLtxIs39NGI7MwQPcvOh0aJyb5YRsGX8mt42acsYbt9r88NsttWuHDkm/GN6PyUF8cAw
CpA1X09z44TiMxrOaHuNGuoKtyF3MD40e48BkRzAUqAFZUEkCQZHKnquF4k8q27Yx8QYYjtVr8OI
BfuIlkk/6D5FhLyQoyqHXgeU09Y97cowC7c7GXG/+QYQQvew+jcLeXJXv/38nf4agU5kBfFbDpv0
qnp7+7LXoZHoAgCSahf8sH6kBj3EB45ymb/zVNK5GbHRIPWqVbqVdzrXNri0pbGhh9cv/X6t1VX1
nnzTaWgVg63xfwlCgdoxwKxKbtLTqY6KDjw0LikWdVjz60T12t1SsYSLvE8XIsQEoD6fJvpIP/LQ
5qB+Zfh2c0WHtIUdfhcuQczf7S118l7fgZBxyszFL3Hj2wbVMPRpkEYcHs6r9uXvoqTH/mB7xSYU
fpCj0ULGO+jithK73FRdmi68/RoaWzuoCJsWsUosYnI+TWpiPDLyaABuHIAkcYDq1fEQQWoQgRnh
k1jNoHVZa8SY8eNudhZtSfTTb4w9uCBOshDNw1a2gWwsrWflpBQ48vUdYqEzDlMBJQTIiiZMU1HW
DcNRaAknEzi9bannRFdfqhFiiI3oWwuNnZMmLQgm6rrDLXipSU5OS0SXFWsT2jLAWtF0MOF6tj9g
MhwJ/LjPuSfRTODeJHDTSpebDwH3xJhkgv5yhW0uCNWqJmwut23xofLK/CT0KVxCElFE/LZ5jqsI
ggClvmDrLXMZvgTOEPphn5UI+aIK/37OfaOVkUV6WIfrssc8d7MsVqgpcObuIQAm+MEPe1hbZqri
Nx2YB0TztaPMjqn31PY+ZPGyXp4t1Waxabmndw2+Q4G+kajuWdcySDaEbTknKsqm/AoA5RXY4gvG
vEvqw0lszvKNUBrVoHYndifUUmonk63/V5ZZC7myjlpYS9LT24IbVQ6PBZbeo8eW+4ikPmd8P211
Aniz+ZQQtTOmEn9lmaijsFsj+Wt6oGUDbdJAGaP9vSzqU0othwDPB1nYSAdarz9fBWK/B4U898Ld
s3xWEXfHsBjH72wukaHDOhcQwRD7Lpg2HPfED4q3xbC6p1N/djGmCJ000SvvxCmnaEONKvCjJ1E6
I7W51Iq7aYOSoUGUX95T8nXIqt9iK+spJB6cZG06XZqB0H9VVkDciNayAX50AQQ17CFqKL/Ejcum
yASKgUBeOZ7Hni5EIsyJSYlMc/7ku5qljoG+df4CpFnQyYIV2QNX+a8IBcKH18uFrzUWkR1LU+JA
Kwma+xH2tXperA4VNgrNW7Mgp9GBy+oC3O0OjuOzK4v9CrdTrb6ywI119jSOs84p5ppnKaeLo7xs
SxeOCss4qsxlvLQ8D5xib0ylGr7XXNcb1pgfXqfgU35WtutJq2gbQ33gxeaDm6NtHgnX+TTCjNrQ
qXu8NjiSMgeWcD2u9E4n7fFK2l41gYAhfgr5P2XctUF11LLyxW+td7bz0KO5z2p7Xja3/BqDui7T
a37QCFB1SsoPZ6fdUzxa6RHyBjvnu14ypAV5VeQkk54SzNbtxmv2RcMIIupvQpIZHAXC+JXqHooa
wo3LWOG5pmskp2YZb5cMtqw9OF+sJoMTUNP6AElzthUBvwrvBamkhEWlIHH3FQsxuw+J79kNqUCH
JsjMBTB58loZyRUlYhp5oLKcvneG6DviB54zERvWJS4vrQr7pMvIWKDzDeB2q/LvzxCGkve9lXxR
heMiyJ8NL46L8EGxtx7IvZo4kWtiEIr+byvsrPMOLrimUgmQeyrefdRuY6+FizXrdpyAD8+NzyTV
tQvSusqWogCsKzffJ4Fdgq2OLr0gN7tGdmRhkOmVXMWzgi5+Fyv/GHoG28jgHnUovc6lhQ+H1nGc
5jF8Z54vASrHr5NFQ3+h3vmI+UHuK0SWeJKuvxef117XiKHn8rKTLO1jx23+o4gN5h8wk7fFTLEJ
oW5qrJh3YcRk6Ny4xGmC/oEH9oU0+9mOVH9iiHkxfk0uNQIcFdnCoupgsRjj43xcSBEMV+1HBn/U
ZRY2hF4+4rbNO8J7lfOIxQPiWAfthkFsRfasLEQoUpC2rNbfHegDuwcgbWaAIE6e5DWu57A9+YNB
UVGGRpoe/uay5vZKWQexj9KH0yP9h2sMGDzuncXNbQfZ33R8KzQ4Z2aGfGizIE92rbq7FFUIBVp1
Fbw2Tg0vdIW5fxXgwaOQ7hewBt14enB1Vjix3JRl8ijDH92S7PSad8pTrcmy2SD+o4Sn6gKNuS3J
4TqdVcaJ3NPbJDcfhZbWt5xfiUHq7JZ8/JQdZYIYZepOuWr38Gqp5j9bY5Q/75j/Y5lAml0yLsJl
B+Rtz5epaVSCm+6Y+e+YnatNuOv/7j9Spx9C8H8RIOsbA/x66WKKHD1BYiGrWpiDJl+PScyjOwWn
1exxAbZ7NLb5bWJ1fcDGoAmLBflgtr58DWdCh3F0WxqRpO412gT0PIotIIyD/MnopPBYdTXi+lfE
PQpQ1+bUHowAHjykmyycGFPC2+z8C2VFVm9nzfZVq5ZzUVWH4SOeu1/W1P4UY93GouoDE0XcSf+I
kAyggt710nVP0/dNZS1P62odZ3ISfHCoyWhD4vvhnFczdj+kYpp27UNvTCHd4nYvon6ZRMjU/20J
58rKzJo7zsKxpQg0TYOJoN5s5ULJUd54kZ594mRWD5GY+hV+ntEqWwAdpkAZ7m4gKUtTcIxUZjnY
/JakuNes0GyNIBOAS0kezLDxUTfwm/pEtniRYK9t1/W7go5qj+poOQf44GbfiDUkQoV6Mkhh1IWY
wvf9vA29xh6N7GYiTWAH01pPqHw5rJoq86+nSvjKC0y/6gY67pQxJwdgk/w/5ZhkwZFYiECM/Tur
Ixh45n+vaYuVo5rWp+Q3owZsqgO/BzcdUl37aTxzTH8BFpczZe/QrLxZMtCvYxUXirZImtfjR2dO
wrFxEnBZkfmfxzaMsiLFT3OpPj1+A2vf44dyExTKTtyGKJDoprVfq9fvSEKplRtgu05Yya/Txb5M
h/J151K6vcNnfHMGCl0U5NuvGaCNnUDJjO6RzZLF+KpNZPTEbQfRfbtNMXVOjKYJT2JnsQmwEUCq
d/cksCWHUAjZg8PFTcTwGelEFjVCeJkQHfgniavk4XYvSTt2AllOxmK34s6T+D9SijYmt5qPdYFt
xGWI6TVR33gSMLBFsC2NnsUcVhvys//V7i2hep3FQNO6M7XfJAI7J5f714dyJ6HWlTASkEWNceOZ
hJ4VntStUBFvpmvZnskMcirEuYyJx5UmgyenjbQlA+0zTX1M4bP4Be7sct50WFSf1DsmNjpxPeWZ
tIJCDP5SN1wxFAej7A0Zs6f3xnZfG7MPG5eoyl/lQd2PSAC32HPedAZi5dlsF2EQWsooc/YzW3tO
C1IKt66iG2rmAoN8IF/UgThp70Cczk11f/Fp/+0U6HvUTOBdHoYg2RRh8pgo9bC7k9Q03/dvDRJr
T7pIF1tx99pTBTV+aM3ip3KEZtyghllRZGDUfPW9GpNdMBiCY4ZpkzRV5lxO6BlWANmeDQooDrps
b5x/p7V/dpleVBwSGRg8z0AIXsegIZouDnuK1G2N0dgl6ep81ntNkOzJxxxglzISDISxTr4dZba1
WWjm6ho/2qbxJN/f+RLfSRItZFLuXjJXTNfWaZWEvtEipB7sktm7LORqZhiN8Ow89xi+efYRZmCK
8iQNr4/CsXojoUEV583ZIXYCIyxHNYKdqlVxya6UJa2ofp1hevBe6DsUsl6oOf19cuGv+LQvjViG
xyRqitmydsbLudLpqoGeaaog/xczDj4XxsXzWKrNVHD1wI1ZL/8vfwZB+ABvoffDezFWxBIlCgq/
e23aYSGYZE5tPeqoixmA4WkYgJ2Yh/9Kyu9S4cIf8VkA912ymvU6ufWG4qBkrPdVa+ktiN4d1Eh/
4oQp+ZBL53fIspRCCImrlaPRkbgwMTxbzpL1O2IwGk5y4TOBDA+LuI8DxGN6R+LyL9zTgNgEpErq
g6T/e/eBKUPzt/6b63TVwmHvgxlCKSYlp5iZwc6llwdLxLRj7YXOqpoSYXBpxvKKvsH/JNy+trmG
L1Zfy7CzPAtw//p8pXYdDF/2RqdfWQDFGW9lVxi1/fde64YRpVmlho3QF0lVTnxTmRyM9DOY5OLM
LeuI6w9MPcwfEIBqNk3ocE2hXLx4YCBlypAWv0wJDdHbIM3m8iMJ66gm4YA8NBOx3P6aS/9Y+ODC
wE18Ml2qnlt2+tIxVSBoOiTtppQpQJnQeueKvuF5yF2GF1MaUiL9nPLZ3UxIX43mTSK/xXX+JJR6
yP6bDNtpTIGoK68ghWL6NmozFXT6+Rdy5uCBl4mAUmBYz3Di5EyqdJVr0xYzik3CaEQ+TrghNLUS
opNEOTmytkuc3Rmyln9EMRxbKaSrblaFUYFlKaACsjJcFIoqEinMNC1V8+QQNdzV++/gUyXMiRO6
KHulNuwfFQwIlxQcdmz2PvLBGV2UVDfMybM/6EVXf/Tm1lGRKZE0u4x8w2ZQvbc3DDlFeYoxrlLz
Jn3SYhJ53soHHRm+gEyxW5/niyzj/Ot/3Vy9M55DD4tpADM9hzCDNhyRsoIspCATgN5nwVZDivQ8
D+eTGI66dd2YYW+moNKDUUdX9dAPY6LwYbVeQuhacEkd2Z4QhPidbFy0QunUN8Oaae2gEBhhEdVn
MFFaqtwd7hLrzWUyupCsbTl7X8g6pzXdZpooVi+3XTYdRObZMCwTug/B6VFUsYW9n6S052fuGUJt
skDY0Guhx1z9boES8kVNVRDbf1IYuCrIVI3go7oVyC+8Lnrdkp4+8ygPOqPTXIpmxF4NaHCD0g3h
X8+SFDsDq+ExZwscuJgcJY3Ywat2R8DMWYdLnZ1QDmQtNBKHBgqFOpOMpXmQEDbs/ISGDA3tmhfa
+Ta+kKsZzQbkO51zpCiHsZJe1XOi1SaKr/pQ1OU6eUvd5GaOoIAuIy2hKiv6Da8cUVbPIxlE3q/J
vkWFkRcCkqCiNqrm8PHwkM3S9fMpy9Mym/essnSQi0/uFPR0imduFwIXTemH6ibpjyA4WDQt700t
uYaRxSdpTfBoWvCRNELxxQ27Yrbj8evb04N3K95LUUZG0uCLuPQJ/ObyJM80Oo+pTDtxf2/ZN7Rr
pjeihsbRDn1ZvQjik6yZTkKkIpd3kaPCwYH0C9GEwgJLH6sQhSn5v0jzPF49ZkshUmbPMYl8P4f5
jAfrf3J1rbOuAxc0eJfN7hVSJZaWGXUbypG4Mq96jpndzc6ZqqrUg7i7UPcL7WJasp61DZaUpUbg
2+zI1sZDOPz7q6QQbVCZDs9wb0q2ub0rlXTI/RXhY7oGfSjPk+2rNRUGirYFd0KObrgYCNwC3HRm
yX56qwz9nuoLGKiqrOYvk3zDx29xVAcgPcXJXQAnid5EBdd+doJHUwN8OlKwPcqLXp+hftADbsW6
p3PNp7SjBS1KfBAK0Ms/8NULRIG+oMKuZg/5epEQpDLpS+tAfCmzawo7PTfynrgk4g+XBSsO41Ow
fw3euWIMe2Fc/I2fW9n20G/+m4kjKt3HWhxeqdkOCCoSKx1ak2MjeAJnznt2FB3eBONAyoE08fnu
JMAqMCA/K+ohjDgFtd7S8Y7muA+7SgPAIiqELPpTne9csSXgTXBZEjRB5AzSYMMXnMPimaLcO2/V
sUbVBh0E/aSzrCRen/oaxMf0DrAsFUxhDNt/xy6VkHNVqppBuNYSKyTr9/w8jjt5vjbaYrf/hi3Z
K6cOLh/sOARhJ9ylhLJM3Pembbb80h/swCq21GykvhSN2Ktd39Z2BH6YElFKUUCp7MnFwgJyAAlw
4knG/jdgwEMUZeAEpyhdhHV4ZKyRdks+z00p25UuKjY9FG8U5Jh7kTSzYiw8ThsZYMk+3xqEEvOD
pIyYOyBJKNX+bVKE5tZeFw0deqzp62mqQdzFmW7vyeUVNbWCMlT4YWZ2T41vmI6DvWDm7Z20l7P0
jL4rSSX1FA6ETB4Ds2g62RO2rYKkszJnYlXh5SAjl/2zu2t8JHYsZZBAZkreKH8HbXeG3oXn2mp+
bQZgsBp84yxvSqcSPjA/tQhJfQNHVgHJjkAZWF9p2aLNUP2KvpTRQCXcKSfhs/mQWfDweiIDgfoQ
akte4SFsXM9iwUXnNPJUaMEQJb1+zQIHG9tlJGuox0wpHIMiF1sH2MdL+9PR+h2vwNgz2GFkn94m
+T2eU9XIRHd4StR6Uo4LevtcqtyoLcbRLRifuYvVBqNQVMxdJefyVTdKN3fx6t7PTa8PR3gma9MN
yGaL78cRG+Yl1pwMPqAKTEgFubLLlq49Aa2L4d8vZlA8HCuivY08l8eTMWFv9aM8Z7+PFhLwIRSp
vdDIqwqEvdnTJCoCLBrU5maotLQXl7JSRWqbtERlPaxwEoZLcDI6R+VLACvB/9i374nzk/EF7irq
LKGRoR2ZW3M2e1qMGW9SQOzipfk3luIe9iEhxmdJx/zi4jeMYAdoiucYJq0mEqyRDWu1N5BMl5Ls
RTXTOjOMhuyr2I72oXgkPlq9dv3TEtTFDHIrZCMrQa7DscKKKTgz22yRiYTb5gn2IxOi3FFS3Vrb
f9zLGXhmwFv0xIBCTaGe+vwUyqFqPx9cU/GTCC5zfcjGqUza2kUG+/k33obn5Z0n6n5lQjV0RvnR
izzEhjJ8PB6mg9t9plyFR55zCQ9TX/f2+oq1CRJV9NeONR2Ca9Tio4w51J0tFPupPHcCQv88us+X
mGe0rgRINX+y3kO0ezvz6IVUfter9C/Xo5sPrVSMgKFHJbf6zfEvC/px2gRoedC8sxqEC4ynjRAz
ESVfaYs/U7Euo+bqy1XaB87ayMfNhuvXIcOIuuLILwOpIjoL8qShoFnOYXlDEFq4Ts3ZdUBFtT5T
8vVuPFSbTNXynOJ+Q9adjtuqDZH5A/+Hu7a6xGwWP5bSXwWADaml/zGi/JLE1V08KyGDQj4lZuXC
SbbY3cNHXUIMiKB65jGGEJsKzBj3gyAzT5ZQ5FTqQp07hemKhkeIGhUt4O/dqX84BmNLe5NoR09G
eZEkplr6KCRXVznwl8xaz3aUJKDD5kmt65Og1mMdSbRR+dkPBxbC68uyBkFx4d1E3gv+JdLyXGnH
Z/GZ6jgPjQ/qO8IKP1t81Au+7mYaiOn5UyxuIuKoQ4tKBPudyQdTl7P1XwuZUeh+HmqJU7iOxvLB
CytpV4nY9NjVNNAWl4rRczVmu40ZLQVhkel9bcfXgNND9R+WhHShM434hdJzusxd6ODWwzlyriDN
Kp37ht22MzYuO2/Rjo6nnyEv53sbM8fnqgjCUFkmLRSnfdJwahX7Tj7Q226dCNv5/VH1zxivypu6
Dc9JXcdDIXJRR5Y7n2m2rtgXGUMmSpE98TguwnCvRVFA+lHTttZHbyeK7/HgIdv/7z8inLMn7xpD
haRVGziIvtoKDATkejBAjKVU4PDwWSu42/hcEbdN+naXlo+itddglXWlOoVe3wnPJpOP+4Jo+da+
hFWoR91lJg0kLvPudlNTI29iktCbQjyus5iqbekWuH5nqwPSC5s2NXn2LXH7hv7bQKvX+Ci4IGNm
b4uhU9D3wa6cdH6pq8+Oanb/ONx1b2IP03HN46z0mW6BPdpbAdBie3MYDS8eigfx5F4rknVwd59b
JNvG/tHQg9F9v3Bh/KdoIcUsk1Kt1+7ZN0ndY/ycFQ2XFED0C8cGIPWWYDmBXC6u8wC78MMqUuaI
jk7goUjLbqRE2IvhGgqWhZ6IHWIOcfKNVNrJezx+X6fX0MZh5p+biYuJqgt2j6x/+kaaypCa+mY1
AiE+0Z5pGRZk7TefADU4g3MhLMo7ODlSxDGNeRwyCyI4GsPcGk2YhhXyd0NydhBu70H6plVCJADU
S9TQqFnhzsgX+fKgsAT2eOJ27VMlcGyEOFhiEmeOVLOZ86EY4iMmjVvwNFcM7IARodHHm8JOfTOt
sYPm0+BJhhs8nC7V70rOQ7GkCHGB4r2vcZQVCeOY1VNDYLPlHuflfb4+nC3AapHds/NGAc1jTGoi
xk4ukaIArG/NehSqyBortFiILAT/A8nBG2ft5gVYv5SrdZuYi91HOhjX29y+97f4i3ME3V46csCT
nRvo2/MMOSBo23uMvny6DO76iWvNwmjTyehmlsjfDEB5fULW48kDOXxtRLI7dCfgy53Qs6WIZrl8
i6DTl3G8pxSaRc5YS3vNI+9Ze6hp67Aow9u0uI8Oak1VYBhifS8M7Z6ODRTtODq1tbQj6Fi2sXqO
1WgAoP4q7IEvWO1ZpxD2DE0RPrS25PYfndf+r1Y6znPHRDTrZbBFhiZLfbPgPf1rDL6XptB0oF14
dXHIQGKIBdByFWUwrcqTPUj9qQGqi46pLQK8QKkwWB+2lU51U6eNL5lELXXhqZxbbJ6i4xwn74Tq
W4NOQQUhgCdO7GQN7AC2Usl5Ho8yASh1dmdgghnYRwR42RPFbqCMobx51qkq5Y4hmUnJoK9JGVVL
VL5s2mvufrCUp6rRQzucxCOwdQs9a77zAyAJwVVbgWvZGaTmNUeeb5lm6JFdNIZ+vCSyNU35HkVD
aYcoJkjklXf0Hf70eQKIIMDlNnxZig5IDDdJCZXCjGuNQ3peRXQ4mYsfmIeAHf2MFjbY9Ihlu/9O
DpgKz7lYNVxXQ5rYFFmQFtgipgcCIgpKKOEw4x3+2A8SzE1I5aWkC7Jjxs3ZkVslZa28DjSrJpbg
zY4Lc4ndafHvltWs76EMVqyqd6TvuLm+/8QSXB/lHD7/4Xj6jybopYQZPzyNNOFYqXSpdhjr3HU6
2kvGg+uJhU/1YQEEp7hIE1EP+OZ7G74opgr08f8Lxzgx2BnuP04sdoqoJiXxMYR+jZWCgvrh/apf
oif1qXKYe5XaFwLG1lMTJ0FdrnOk8vh2GFSF/Fw13zeQqtihenTSOuIn2Tb1G2y6xw8boiKj6COk
UGvpetlS34PjH+l4pPYX7QZY3Uu/27A9e5CYLoay7l2owwxHEQ9lzv5xUQ/SMAhCoIJnbOWI2xxY
JOy++Yk2MEEqOHjRJQLyAL27jxg+uO7rtJhYK1YTeRa0pJFOlWh3njdtkUPAqfAbLM43tfeu8Xys
p9t66jPs9yS5BETE1apFsBRCRu9EVp6PGm58tFMsf03U0f7szwyi+ddCPLFUGfuCBNan/06ugpiS
l28iR7kxuEk5/EsJ+D17P3jojCnaUDeoNAmi3CuXpToW5Yw7sOdlJZ4Kwmsau2IhB3ERUbxnkrYR
37qgzQ9CQboue+acVkXBjM/72ETVg2dv0X8O0tkXb+C5FWUqbuLuAC1jnXtEFUSPv/eSl3MdBqCN
nidWqd5ABW4eGIer+ovwXbSY+48Tg+rT5PFtlBU63jC7XNOPlZ/x4UuPEsj9mjzenyEVSfa8OjCp
SxSKJo/mbTLUulmD/AKQfyFNCVZPV4r9xfbmTKQMmHgkmOLnRAhVMtVdotoagOemUZ4CSK1RNhJd
BNxG4AQcDatTTg0RjJHqgZYs65LYws5uyy0EF5886rNtZbnvzGOeftp5izlORtrUNvaYPmhLv2/Z
kFkqCVC72+O7kEUYsII0a7nvF5LSeqVCTZ6GlsSr0ZSgrAplHNNLziAx8c5CYGhiVAMDti2En+nF
vDCPFb1Y4S47pgT8JMJT31F1T1lssC8FdnG44lil5SdDwTHEBfGNbqi4usZo5lAg2c65FpAe3wNq
OfVWcf28TPNDuIRHH8qay7Bf0arMV2BhAyZ+Q18r1eK3wwBo48G046jZyY1Qvjs3df1rYmeUqrIx
Uuxryk2EjCEyRIWE0kM+UgVG1V/G3lA7u8FSmpQ92u6dwLFcT0Do1KDsJvnWWc01SUBGJiOSi9rK
umW/b3/t/jRAD9W90NfigAvQNcK5RELVY9DQ/LrmDzoUQEBzI4FTtSCdW7+7cEjcB5gC6y1QSMZf
zomx+O0D2JmFEnmehch+nb9D23p7YA7aAUv8VSiTOaih7e/vGYuhSDoKUCRSsSslTKyDVLD/PyRO
4e4T9Ss8ZZS3bAPVIVMbW1LShChDlJy+4EkobggjQf2zGmBQOTX21mC0+m6EWGyTjgvL/PCGajHX
haB9Ags7qWH+YYfi4T5fVoCT31auhDiweYcho6fcUaU72+ZDANqPj5a0tw3L1ehb6U8WLfNZrrDq
E842byiUSudjFVxZ7qSKAH5fHYHmN0a9GTn8qJMsHsLCbYiRuIn3cKvHNf371rtE0Qdiay3vRhnQ
zJqXxR4/czsno2j0Q0tJoh+IojuaVTSynt5xgtLsjun1ZARXSgZCN80Dfxnw3NypCj22LrgPX5dW
ZaVZhUR/jEb3a5cFjQK9NChOrwny3MP5qlnBvH6GBTxC5xJjb2n4Pxvlsax+QVJrY6UOYa/hHcKs
8zfty/WX3d9+it5wNJjVflzYhgacbhAYyKfn8G5kNvtOuJ7+veyQeth/oMZu15OtItV2hmLXY1TU
EMJz0Gkg9Qy+nU6bFQ9RaLK/Wu+oneaVfQqpeFRTV4/+6Vl6RImNONk+M4jVd5dggOnRGGFIDElC
B/KpispJsEgmr9CjUi1OEoa9Ga1c8J2PIEq7DL+nZ7CaX5gs7mkjyH6iCvaM7/M4uhIRTt+gQlqD
dt4KaSPDqhh6Sk+e+OFxUddc8T8/dDZ3sOI/hYM2TBmE9FYBvnF6XIhBO0QS/ZbEeT3aA+0HIKzT
kIp8WZy2NVHCwGJl71ili9coMiweqJPGWReDiSzKz4/n/NFxDnnV7bO8cFQVhAderdPU7b/K49B2
DQIA2s5fmPc16BTJ/zNXwWxkopTGbNGmwReqKQhRkYE+hq+V7/lqeKDKUawsF+2cxkUtT02m0JQZ
2uNZKHE3l1FwWNqirBG3aaDkvM5pmA4hoSXJOLJmpoN1IHl9vUhihOH4ZmWt6RDOsX74Zn0DPqGq
wOeQHwUUODW6z1zmHOhB0WEQycuRvPGJkSCsC2V1XazosSOrWPGfaNeGy+Go2F+GFK3Di33oEjWf
c1SBLdzq5WcM850xsm6WMuk2C4kMSBllEJ4LyIPW0/YWuuc2RnJn180r+i7SrFCCRFtXJGR01ph8
cpyQs0IwjAw9wemAzVJKdG/hDxyelsE6aIufMZBi59Xhmg+vqPnKla0O0e9QO69yS91/wRLXZIUm
UPaCM/1K6iH6RHNMe2+vg2v17h2FpmwvRjLdW9ENGyBM+b1gL3GKcTaEGYh+OoboikP0JQNRW1ox
jZibEjqNKjr6uoGtz4ZX9jyt2QJWeTJph1uwZMPi2WWtSF6k79WJxFjsHLRCt17De61oGyLAYuaF
/sfqhRcFkCjmTvsh5CTJmQ9EKMko/lGYnfxZdxa7xxT4qUyJ9XSRSd9j/fHIWc1fBTV/VlFvprhg
n0jXzx0L3XNR3i/oYSDxC0bP8dWXwF6vOs6Rb5tQPtva5ANood7HfFvbO1RrRujlYo9uEpl0rDNH
GhRrL1eBdUhL3g4Rpgde75tX5i2aYia9OFrOSCTCzWI++zxBJ+89eQy1fyt22MbIYIlBoN+EZM3r
YsT686quBhK2SZSgtzF3EYkr094Eo7WDqODXMY3RSr6/K1uI1hcwMy13oEg5aD5Rj0YcoQ5jxl3k
PzWdVxpQyzuxn8HseflM7KmA1hVZgZltBkT6TGV6hsGth7XB2ZJZVO6cwk9wIBAc9wLbBEjRNvsf
Y80n/znHJUh2P5uX3Db2pI82b2hMwnAdnaoGH98PesBjSacm9nSKir8pFRESyzxiUYnWZZuCCzc+
bKVwbjf0JRem8hCiXoHpasqxGbhrchQGJ3gRjtHyequM126G0gP6uSKCC2xT+7eGjz6H2vxXDzKh
vKCHo24fkwbgs46uRBaMkKiMcgdIQrW5f06qCP7nGVd/luPcGH/ZdxBpgpVg12ywYBZ0wXmFzE8b
J/AUIuKQqeCmw3MHCePw13qIivj4twBLn5K5lbq+CulXmIRc2MHPr/6VvZR4+5+6LqzOI5WjD0w1
OnkkcgrC5QqKHs94cBJTuDtT80tSNzk2RF2sVxvrAHF5dHIeh1gXy3sJw30jQeZo1hjd11yT6dFT
Q8GlWh2IHSZJ9XjKP8rDjLAROQx51Ram0XGiLbvQme3bHQeHS1nZBVmhOhdn8J+xg5wStp2iWQck
vznRiFGgmo3uAWtXcH5ng3XJ66YU/5AXBfE2Paz2ZFEGSzkWG0fqdfbfwEb9zJ/JUSB2ksw7q6W9
OSHJfoI3VXBncbGTLJbadIYqqUTpW18hHV0HmyhYAWOeiE1ua89PLzaGk7K+0krd0EocOhL+wsyJ
11HBroXd4VrCfIwfruX7/NB64av2SOaQMnzJRL/BY4ZQrArTAgz8MrLkb1I2LQkILhMxBc+ZP+dK
4ZLdtDLlYpg7Oj7TWSDE+Zp1qTvaGcz+rEERM5r2DxAWfMbqd7HLqqqqGO1mn6SGqkUIIe5RcfLF
lMHm2UdHmF6EWKE0ghxP2cVRBnhshzx7tMguUWpaWyUD7nzUcOFdwlu4m6Yf527Wv3uIOcgSn9Q8
E25diaJN1m/F8KE/3RjjIFSS0ODFpQnvfvq9t5BO31Ygy/lsn3mF2TNpBwy6hdOaMMfv3jgMBLft
r1SiT9hJ5DG2FiLVL3M8GXZ6ySJbRmk5ucVTTMLJ3jXHdR6Vj5ZXkhq/oooej2dIz5Unz9hwtsOY
+uolr/PTPJNlTvl1GMt7p6QT2pyEQsTWxkf2cLi0US5Cbr7+gyAKkgXYS7dF656jjZI2Lfq5FpvX
zNYvIQSDf1ohHgQh+VcngsCjd4PHMMoOaAZEjJSzfeZWY1TU6CvVKHdzQR0DFbBpe4j67FpY3TpU
Di+8/Qey0MumTb63hWzaWJ4J9jVXVO7E6dqJA/TsoYzfeURV5kFQgiYIZmMp8ITVCCG0YRJD7HW9
wy96FIk6yAZW+6UfqKQV10X0Yeg9p5enlVSoeudgKiipCZqMJjvs5w+EwypuNnegO4LLyvmws7Ot
nv8/wgIReEKqo0y464ibRZcFv4aZeFjBaeSRo4YDcBqyZzS1o/JnO7HAJZ6kWjQ3P6BQCvoWRwgm
apNmhpq1e0k6H45WfbNu2XOP9Bjasp3ibfmO4Im4JAhOwB3qzK3t03PxvX2cxtR2c0rdtfRSEUws
d4q2Th/Y0JUNKuIFzxnvIFMNj7Yqrrj3uqynx3kVfGtXisDhs7djv+xDm5tPDG6dqrtuqyTT2WJQ
Pw1eSlSE9YDIjjkyvkqnqzQcF1YPXNM8wF1un03G7wBdxoSq3mlPHtUGsmyE4gxGqzeXe/pZ+rdM
AB2fcYOcwO6SbL1QzWvZWOYvYFDZLavcMwQaQhHpmONbpLq0QxJsj/0UoLgY7d28Vy1UfS3ysIzs
sNA0B1C+hxy2UECrd7Csg/zyPqQ/Vna5D/JWIljZMxQBdMgzj3PVrRtHkdxz+SEPOL572T0cFuKu
w0K6o8bRjG+esUu2idSvs2jer1monVbCnGqqJ6vIeUv0i6f0iaTVGgxDxU95dqFIpj2az7QZTjRw
2WSUCl3HHtNlZP44jUI20c6GpyqD0Az5KkGhad5DOTlCcSO/b0S3gEfRxNSnXP6c6K2af1LXLQ98
RIhgWjc6TGgPGTZYc07HTfqM3atUY5KkqcyDXDMXdhzmVn6ADb7bIZ36qPEGMz1E2CtnWmO6nhHr
y/4feNnSJMGqNkT+JAf5kbi63obCpGP5lCrPERciJTdTChCtNxa1aNHw5gDhwMH7O5UYyuloA+ME
C0xCxMzUEjS4LJMccwzPXEJMWdJZommWrXmJtSta9rrtYRWU2bsKHpMDYne+eoxMUdEqqKNdIeFJ
VvczIrH7cc4s8enoskHj72TJru1w3NvWVXwuaLpj+Ii1Wm0UWRdjMPLdeWvstjEniHlQWsj/I60t
GOTK2/VcfAyMBpV5zMWBMRaDZ68uTkJBjnuX3xiNA+DYvLT70Mj/9Teuwv+Fb2XtmQTJD7gSr0PO
pvaZiTUh33sfuEMCcdUAfWjqxVc4DtMM9OkCPqS+N0PmiJrtN4eRcaMzMmTREQHsTNoVS6MLlj6R
RJCLsqN5M1nM/tbWuet6UNXs7V08Wc4jrvXM2TOVcxwG4GJWF7C0q8FNL/xTDr3pU+JhnAGEnb4n
84coVxZa2bP0RalEOW3e+Ul4JvpQmIWg+TSV41KaNjzdOt627W0NNgpo4HTf175yDY+1EtKHPBjK
bbZwNWMMG0CGVsRJq4JERwSZfw50ew1P+Phsfc7vfDBXkvuS2RHbN3RpQIqqtiUxecHy/LYrQRuw
zIAt3WvbI4cZSLIbIbLU1LG7xfJ7Rl+7TD1qsLvU81QcUxFf8y073bSpye/OICQC8ZjVPNDDmwZx
J/G98OMOdLHnStkKKPYxAxLMbOZMqU9krSp4H/9kMpngEV7ZC8lFyyz9e6E26TgcdkWh2a6TjcDz
+rTIZFnHm31zanmeCAOt60AwakUaYMWXxYjRcs+mBZ5NGc3eDXBfDEfEgIUU2I14mQLsJ/E87fo+
WhIjRIWoyU145Umzxn4w6viSE1qkQwsfJNLStq1e5qKHCWBG/xSA8h/Mzi0VymPyUzsnJO+wOkzd
KLCLNVxFgg0w3mNgFJTeM5+n4sXuV2I7vXL3tWD/bSgio5QGaLD7FObqiDktzwP2xPeVULh2RPj2
aMYbJUAirTR5vzqdEdBol7T7jQ6seON6qsg3z+sjYEl6qOt6mdNy9iHxDftiXYWvnrIuKfNUbt+F
kXKfLzGCX2gfx9QvOKxs0dRPomLtgcPWc6ZiqlibICD97uKCO8UjIqomENqvxekb3BpVVQHOSttv
Vb7EmGSNgPqz10v3HbGVZ2CdWu1vF/1AY/ev2AneshSHqlX8N8amQ8uIH1vAn+p0uXJCxiTzUM7x
Y0X6wzFpL17ofJFgQ/YQ06W+RwV/Hr/UAtC6Y2LjyHDPPTqe+snNNFiSej3IqcYVOX71B46rmhdu
14xmnH08BN2Cjwq14jfInA0aSOTzqmMTS3Isuu5DMqORQVVNhXS1i8+SztRfdfBrDGDti/ygTS6u
ffFQWZABjsuWCmxBU8ODr9Hp/tNg0i03yroZWKwJik0yExkU6cR0aXQYzxvfKliglKOiIYJF042F
FqcYZwLMlS42KooGkKPsnVXYDxgMNeg38ftZP921N9L3h9VLallHoPzOKhPLjXs+FwWfymcztzc9
V+aC7W5azPckQbD9uzQeUBq17QBN97FdFQF6IpqYWxNYMlsli8SUbVNDNa4wvlaAwOztxWcmXfv0
eUCDWXr8yYIieS3wHXaaUvBkxRuglkr4XZW1nikC2CrZcviy2omEMiV5upmRiCORwI8vf0tK9X6p
hHuPLUZZWtXuGT8N8fIiVXOzzwOwQcPOGcTORGMk01VoTJozQAlwJMdyXzrdFfvxJ0X4SmAcPHvg
feBofxsclLxmFEsTMZlN5dIQ1RV4NFbMUzcM/cVdBRm8VLXNrImFIDi6O4HUeGHfVkjY5HWsqbwr
hzEl2RD70jPmjvrdRFVMiIJv601/XyfNJ9M1xrjXh5hOCjxR1jpt3RhZ09g/ejAU6cvyabJKDXYx
jxsdDwRk+FXfbv/Qn/Gq0PIInhVOMAWXMib4PGlb+V0mqxpogWcIpLfUXcHM8C6yxM4SgIWTDDw9
TzHhCjz0NvoO7K4jChJeiUXxTsfeVZ7XgGNdmpWxO9med6bMURwfcPKnSfR3P9PuBujjpEkDv3qu
+5T+YGOrRx7vUngEUwwoVFGt59ieWZ8dSiOHKE90N/NQWw4+2rETtToyAd0v8DAtc3pKipA3wnDM
LfO5khUDQn0BpjWC6+DfaToXjYz6XqFKLIlFUOrgrx0HmuDRMdag/T6JsVK8u+JDp5U3v5IQnRrQ
o6wWhFgeGvxVTxIgL6MlMN8jGHS7S5pWQzdnRPPZ3/mfAgfV9Ib5tQ9Wt4lWXFmjhiuFOnu0vUWo
4bnY0aujbNXUfb+QlLVQ/lp071dPAmhLZ9YWLFr+N5WqumsER0vIZwy830IpYWm7tYCRTPuSvzxL
ubknLC20wPir2bC/n+8zc3r+Z4sYUi9HkIwrrD1kjR4xKlQdrFQ5YVLotpoxlwNui1FUR+gvb0Le
QASKrQgklkgS3TstYhkOiZbpo9M2dEueQgC5XFu+mXVJgSfu/YOnW4Ax497ZsgafryH/a7k/KaCR
C3NGBfZgGlrWyXQ9veQ4bgvfwfez+7hQfCzftXaLD2iCVhrHCH7SFGu3QVzVBqk44hsM6+Y/OuN+
jTjvQ0iVE44E986Oybz4FbFWlKSdVela6w6d5yWN+vcyphjvLQ2MfudzrDbk3Hb/AaZUJ6Aak+2s
F+sTmtIXt+3UEpaK5Rl1HOuW9X4qIbm9mLwSmO3BYyD2LIiRxd7Jbgca0pYGiSQRdS2fm4O30pwc
lPT+obhTFNPmSD5UuOp0Z9ghuw67+fP+TlbdCpor5MxNN9Eq4ToiMusi4jQ5RLRMGiCmx8LWjRDf
tkrh5B+lQbkIpX1tazkf+0LEFG9YL7NJwQ78K1MJ7wD3hKNyUISVbia5JTUV6fq50kHWFvhqsDON
jFzs3mGVivW3XeuTX45wICJh+ItbBfPcQ7Sbylvh5Vy++TZ5Grd1QHNUmhiUqieRtvcyQxXOzpPu
Aq5Yb52ZFadxfbyPnN/a5OfYP+0DaSHaBBl/H3qTlQ82vOYBIGUmo7s+23I5W1XOJjHV0PSEXBzb
PddZWQjtoGNoFpHCucvwoFRxkkL0Fd6l6uG0xHeQEMzcloA9keNoD9HuGj1D6oCgBRY6doYvMJLR
bdxw+IVwr8PDDv1HPga++xtjswrFPj31+2z1qENCVF0v8P/HwR1f3OfvAf2Qo/8KbD4JfSlF7/Ui
lkwlLQ739D1EABLHGID8H0bumHuqR3dRAWookxmDLQKB3KpxJHlBPs8OlEQrdUTNsUJFZi0Q1Mvd
yEJGs9qGdG8FPau7OmOT0u65mV0sHrZ4/YCz5iRsirHA1Y3lt/ayGRUsM6wnF5THWRS44h9XukvE
4/rvz6AOxQ0SIFS+ZyXwzcoKhG+FBbNfdnRZNecVIZXDI+IWJTMyk1DwFwIFfnQNbnF5bdQw1KB3
6hKvBpoHFhhsNOcGSt0O71mRJkGFj91UvceE+wLxE/TttV/DrBl5YXrHK0SwHZopuIz4cNSsY0gO
ep0dQsC+ZnT5u+TjO2F0ffBtrnVlaet99U6rf0d4Rwsjc4zWKWn777p8S+7jMBLsKytjcqFQIBGi
A9WgvxSo+00fCsQ6foSClfOnXhJ+Zx6UBD0Y3R8uVn7e06Ay7ez7FFP9YWoIFE8bZq5Q91jwSnTt
x8PRLKHSnM9YNmyvSym/7BahXctdCoWV9WC7wqjBhV7RRJ/b7LbxmEzCjeyPsBJbmoS7blE0b2Fj
GhGKzUIjB6rqVlhvCV7LuD2bC5hM08mOagsxHVUPjuHPzDLmelgNFHtgxaZeF9ZWFP+Sw5sUs/Rq
KkPJUzoMEY4c4Q0llJ3znA/WUwNm7S2JYBapRa5fs8wFduO8a25XBEc3rDbdE9PhgD7AMRPf9jVg
s6L6QnFJNCwoRBa0DCO+97hENBbk6wrQE6SSKrgq0jMxTyw6jONBsmwCsvIJw01+M5ZhVaXDWrG3
DOV+6GC8NTdrJ5hUeWq47a67ziiBsDSPeHW7Kqs8skE08KLxBBYUZTDL5bcwzWtjB7clcotMrOd/
/+972P4dk3b5RabQcp7YVzt8AqYOBxh2Fg4p5E9j3y0jjy9k6W2NRlF4L8awiu4Gofzckq6pAx1w
20/8f3gZ+fGuAHWWdEynlpEr1vvkSXRiUlMjJAEC7V7bZ1ViVBLJh5olD3WT6KK69yju2dIF7eHs
sqF3Vns4/crz45RMQ+LKfo7odA6jKAsdk7tcXYuQCUfXDY3vpDPQafRwjX1IuzS1kEW6+rG9AAqA
2m1QhFXwtv3vQ5NmniXSKizAAybxY6jg3SrvZRfV2jOIXJYSGc3/k4xlbZVeQ+B2DNnbeFa87/h9
70vivnwWQHcsV7XnnBiYXhoth7xvfQYN+QhvjfN4VS8SaIgenQWSpLX3IKukH7QOfnjHyIBQxa5f
u4cnTDSOo/OAHvki7ml/uWL9pf3OU16CGWDqjIZuYzSGgW0AawBYqErHIf8smcO5/z9h9gm07nxq
fiDZOE6Ybr98crXBjZ/54gyhhZ4vfI6gky7snotim9FVNe/q22kDaLDtxfkvKar3FBH71hT7Qe9I
9yiL8ynuNkHl3BAOjFlfaZLVmSKeiiultwrQJXqjE91veRRFoTlVT+C0zJdR+YQP9lx+j0hlr/8I
e+Fws9B4CG5X1zbmOXB8+8bNI1uLS5BYXVUKvNnJvEoHuP4NZjt1U5m5HYb5It6NW3QmMAdzSQEn
RNOWqIojSwr6yYQL2bjUcde0NDsXn0MlsOn37V4BFiX7UQ+TifVLuH6vD8X+nho+th7N4hE76RD5
iNjtnl/WFJpSEmxdfHrnj/TCQvSX/jyluLdi8mSARAehYJY+tRg0ON2PjoXoToxdF1lUkjfbFKkB
zFQFs7lpjZ0wMMG44KshbnkNP0mzK5+o/O3xHmOxb1HVi6M0NuDa8+yA1yLkNNcOM1F2W0c6xpWm
n27QWxsclW2/Ngk7pPO5A5P0ljrFFXycYI2QoJQJd0ppDwccRMnTzz3zMV39QFyBdOBVai0DskFn
Yd2Ibgt2/KBoXuMosvlPobZrvQhAR1HJRxZuCBaP5SoZIbYGClS7KZe3gjQf1JBwPTUjZnGNyKQz
5sbQfsM8Obn/BB8Ky3eL4PN16uTyBZOu6+LBnu3jQ/DQYk3HSZQdlIybSgU00dUoDDwHr2zp7N2/
s1DDqgPj44e2TnqH6AW7TnYx5g+PEXLzp4Y3MaUnmQM5MprZtuGP2FB2mV8Cl6s7FwvoP9FiM3a9
lvs2R4cs95200OWruK3ttoNyVXVghl/rgbOI0Ifnb5xv5EMiZctDxM/aZKFbiLkSON27DHwwWrgo
tPe+D7tvhh4syrPnmgiYsHfTA7lZdiPXrXQQFl7WmylIl09uqZGa2vF4Zfp7lSpGvmswcZm/dGXI
CRqzwhIr+H1jR7P6+x+FucIEkefiwyhcYKCLEDBNzdt2ynHmgf77gcEd5TpPD/j6AjFHiO7WwvkQ
tlPRjOzTyYMeB4ghFQnVJ/eeW/vIWvWL/NL/yuKfDFrOBeLRuY0+Tlc1iEcNuO5hKQ2rufjL/hHc
5kzkBgQBj1Cnbuf9tlfGemE2wfk3ha5ED03bfUioJyWpvVnbSKv1JFbbmGmZin1FeBImcjyV/z0r
PuvElXWewIBx3VecMMxar07UP9ygj+KlsiVt2lUvE0j5z9JVAze2NaAylPbfxhDThXoa0kjbKWT/
bDdh0jGJZ05J+vaTUTOXZ9UQklejlpdcjeR8YwuhRh6ZwblQ8gjxzASevBA8XGj8iYHKhuNlDSUt
mQOWNW7BGK7FYj+ieZBYrsNaN67x4W0ddI/ZEcBThhUWxVSc+u4bqzgrcSwOdn8F8UU3ctli5xS8
aPn8sEVYLy87bW4eHQqo2HpDlwyKyp8Cq4N6tF6uQU7ofrNfkMfzYQB6D24uQ/JpLrVy/+z61ZS3
IG3zrV4jtqSTikfTEwyPEJEim0ORd9TT14d277Oz/B4geSicWMMr4UmkPC9Rgw/mMVPJxA5NU+fn
PhGqU8rOSIkuBmXWynU8LqVgOQqRJsWmd4kVV2QC2wc1k9Oz0dYwPczw+quWucLfITIIMBwleJ8/
cVRwElbgS7IsCziFXyJnglw8E+gwf2idmsU5Kw3fnQi25D0dhSufJ2Tlsrl8pySFwP2SdVQVb8Z7
uCy5qQjrqPl5TR/kdWuVEw8ir3iw4vbnKFJJJaC4GXVkfY6s/trPTfH+BmROveOHr7ExSukF+0bi
KBfST8BglshycLySAYTEqWdTmmj9W005W8horvzhxMFDoXhYEqwxWYDfCbVk6Oh+O7f2JLB9O2/s
AJU0oNgvLu1+0e5QFkDfFruIHaGkQUToqs6p7pVwXna5Y4vvSDYYQDNSgkiyPf/milnV/tHTDTv/
rciemP+hMLGk56t66N28CCw4Ews7aBsts7NBkVkyycZFHDnEwl2XQafr4jgZAxt5xjv0MqDDIBVx
uS/OwnJIM3DO+J4rraS5TJOleViU4S9eMC9nazf1JfRNmnKBoGoRX+l93XhIbFzpq+ElVh8cC9rM
c9hkK4Tjc1Ex8PyBS7NJD93hhmOLrDAZy2qkrBIjduyLJe2M8KA6ey2ZqgSq814+4DI8XPNSC1jl
kTKn1yacoXgFnNtwOnqewnubR9AoGO+QNr/w1QeFDZb6aiPDEx0Ewsf4SMqh0zQz+rao/arUN7WS
1WD26EJf2yY2aInbLzG8pkrr3I+vikAXO7BO27MtZK98Kya67DmYOvzF0qgSPuzS2w6tsnAk1pLV
n/iAbsEDcva8zFDwE0mntUMLpxkOvPcWXiCjm8ZNTpjRVrsExVRBxlLT6TtCNBjmsVSi8s3MH2qb
ocM/ZMTMMfLbKtDLtKpbRV11u3n2NqX9qox4oVybQVpN3dwyNUnvdiLG5G9qSfxHMzyGa0tLzc/V
nqiZO0pIjQh4Cjq9f74ZgiIOXCqlJjC9m0vVSG0lFTeGos+e4UkmdEWHjVufqci2qjo6za09DSAT
+iWUEkj05fpJz4FhYOhC3U3UTso7dhZL8H870uGz4EfF1+Mgo9U4OJxCUFeogNJpmXiN7DwxjfKc
QmLLwQcjHcAXpc9zKRITsubRUpmawfc/PbKKC6GS0vQGcuyYLhW6V4lQ5JsODqDkAqxs0i8SaSFU
BtRtJBMOv5KcEy3MHc/px5+7IHQ/P59g/PLiyufa+1RxWiVYprcRYBJvNunPOXpSlyoHsifK07WW
rect1EL9W3rvIV1STiN+h0XbBN/yC7pnfV1z9Gycdsd3MK9ZGqImsBvgo0Lj+TsHs5v6VHBZw0c7
DbfWwctAnFntlhKO/VLzKpL7RreL2AtAI1P6yWHP9qHCNjJDOtOr7/8O8ITkBbt/O1MIPJurV8zM
QinvKM6F9g6uxtHckfkULABCFJDdUfnmrYXF007TnIIrKfrndglD2kgK9yIk1WAsEnIE8swnaW95
Y5PmjjBlcVHrLYfcZa/99ID14jfWxOIQ+wuk5nhHH4N1WdiYIVK54biF9+v41GCrRcRTcjWebEtl
2T5q6SyvU3YwteGKp+yz4LMXAPhrw0BEpW73DcrWLQYY8flGtmZ7QIE8CEsK9xWFmTH0a3hW/aIh
W6HdU9v1uGLvog3c8D+SgB2OswJ+xrN5zGUwyAsvfQWEyYrJWmlBcZVBYmXu8n84gA8NopcTODrh
TNxWXQ6rDJ1DDI13r3T8EKdryl/F+Yw4s7SVlLBTtTp83L0sLgxHFDFsoTcyClv4rIUMEVwEd00q
N1dDyHQV35ZC7fc2vusww+WjHp2qOv6e3Y9nz3ZXLkazapCE1JyBHCc2EAGfYKr1DhUd2fGa2iOe
5yUSCmwuY7kYbnkMbonYQ8Wjc2EStLd5nhr0+h4TLhmO2iSznDUK5z9TCjn5FdwltDiE2wmC/Ah+
0QHse2fsohvhvEPKgO0/B1wGHjdzZ1T3TLZN0cnKg+Htf/0GLcO9KrGgbe/O5rSbPlxA/s0OVsL9
wIGykmhdZX4IIN0MMgS+4rTzGmllFo7MFN/W6QM+8Nz4+FlefaT85lnewyerTb1R/saVbNZ+UU4R
3v6uNGy+AVs0QxPwF5Tuo7NK0dTXpKBbwrZokxo7fl5ywJHGwPVRFiMdcDbdDwNmU9UJKR6oZR6t
zJpCP5neQIrxvtW5mjYXoQblyHvDfnS/9+0lkkFQ4k8sLivDHnrCb2aqslYH5MtCwslABjD2gNDj
3u6jGVgtICONcFFEVc1PUd0Pt7154VU40ZHjGucgA3HBI/+B3QdKBMjtOG247mC3iaAHCtG/spxa
QGQE+/OwoUwpYU2yQGi0hDLr1YAj9G3mNg+DDYS9I8d05vx/qu8drifaTQSGdVanyg4HSy0jMHEk
r02/COdGqaumeUvY0t9fsTMFq+y2DgZy5IiQjFJhCOsydOLFANyhQvdUa7eE0m4bCwdX+MsnBGkv
C8agmU5brlpdLgCDFgFUEjhwwfq1BQaLB/BSagK2WplK+lyHhvdkXo3ORKTtST5I8paq+GaEwRjQ
kdiHZefskR52GbTmA1/GOtXMdf0FekwGwqnR91Of+9kN70mPcnPtM1ikyOMB5MjeY8VJfbkQlD9a
d3Bt6j3E0UWNybBSPwLVKizn3xlxjT3FijuYMZv0cxAlmvQYRzWgTVk0KyOx1OQPPbc9ttVhDub1
WgXS6T8F5LVlttsIyvZ0kMWTt5igQHCN2WlduXlkgtiZm7dGEKXoXt420QBXYsV2S6LCGSvpwbMS
FmnWHThTUEG6KKeILlUc1HBhK1UngOAcLBbqY1o5WlEnUjtejJndL2W+ASU7KAxEUKyIAcC4Brzd
3AI9kIrS/zrT8irM+Y5eclRtioS38GPYvXphfNXb7I27Q/YQB4TNnwMZcPRmK51YMw/1mw62PWpM
NnrLxw/CmkVv3ZqmTtEo2gUHQDbaV0xD9BOP8dVimuwK34PK6D7QXCD1fXO7JyCUC0vPWnStcn6D
lA44XV7gHBrd4jUbBfD12O/khzaT4hTppvHEZuEfYfEI+MmRd3gq6laOwiTSRCKvAy47jHCvBSjK
W35hdLgZKBwGJER9IpBfOq0x+TAOKusyFUY7zimRmmUULXsC5F75splmBrbIgbFjo9Qsw0nuW/NE
Po1aEZcQ6fVwtsWVVXZBItJBF/PgFLSZiNY+BQvXTaFj/gtbmRQ8wXVfv2GFcXjZ86bJCXzPMiNL
X7PDwTg5adgNxpmWrUdp3T9lV9f4G52QULPea/vqHTvCmn9PEWx42PtZS40avD4BOiRKfd9hU35x
2Nf4AczzxSb4U6r8o1bEGF/VXzzaerhBs5jAPemTCYBYDgjmj9jVlyeEwyVUSk6E8Kg36biK0sXD
OdIZr8hwVkYZYwA9m3qDInDXlAVlSNdm6palx7wj56qx8N1rmo3Qb7l9zZg/98Ir97NKF2hC4X80
5EV2hx8Of/+r2jIwtvi7YMpP4lOaHoZm24LxODEmvbUuLkYLKaDIrikADVs1XWIXCdFzYO6W6nIY
ASow0S34haxJKcIOccgiZpbnVlM4ix2a3/Evg7BkY30TCnULK6fdWUsLvE9g91yg/VqtGeLRfcC4
QbSgBuOXa/tpByx+kMTwj06kl79xfFHOnbRaswMeRsZ41loOxo9AHiMgMOrIsfP7+Yi+mqHOHEyM
5IBopv7YLc4Lfadsy1UyLflFp8kF0cN+ZNrTZ3d18ZH8KMydEmdxaY7bawGaI4Bouq4JNnASy3fe
2Ms0OSouH1uqfhyDe3RrDMzqnBpEUFdMd7AhBj7sj+iK9hUznjnxn30ohiBWyfviVoJm1WAnZziw
px07zWrO38Pj8gZoHR6HBUAih+Hn/9OH7yXksuiKC4+3kHkmxIytGjb/HBSNCw7ZlLgiK2hExlwf
LiixBYTrjF5WPRU84hA2CK5RtZ2Gf48mNiWqzFxOxWuMdT3xlNn4Fpo9EXfatlm3trPfKhqK2KV5
ywn4isQgDnhByQnjloJkI0rV9LVw9SZJxDMRL4BgJmUxTSDwgKXzPeLchdWxToLtWFyEb2U3wCNW
D+5/kPuAxmicc6MStZu3dMvBD/Nj3+ApJXs+97RpMyo1UMLGCCDYd/JjfBerfLEUKlg5+n+Bwj2c
UGay8qQk3Z0yaoioCKMQPL1hlc9ytTJX1XHXlFdCyqU8FZ1yqpk+ZoNu1AbbbZgBZkpB0uCF+HtC
qIi+oBDCG4OLRGpamIXRLh7KmnbrS2Syq7csQbP6q8rhM7SExn5Yt9ufYGeC04eg59oC3KwUKOUV
bUuTL0abW4taOGu3tXUKzGLbfk4T/acFBqKE2WUwQMjYvUVE22MJZ4drdGMdbH8QJmsil1bZQo5M
e2skvp8y7R4jcmugPrM0JK9tFB/ldUGmSs7kufamjYjkHJF4S4BjB54Ej1YIr3eUGVsGbv5s1qI8
dnuwrlRBD1ZmiSnE3FRzr9R691wzYjTaIx+M2OSJFPL4B/oPQw/sDphKBbjbv7retljZ3Mwdoq4Z
qC7okmT6+qUWpdOiZ/omy+B1R5wdKau87ad7Yfltmucouf4qGRLyYZAuYbOFRhn6h60Uz6mY2EQh
PXqzLcGvQfyw7O+veKf2DbQjf3YbDLcFjdj5KxugM4SfAnLjd5yunjIpOJcFoUO7QSg1YNwNRaBA
gJuymUW4ZmKp4fgvDrsWdqDQmApsd4rBdeKVwsKDhj33x+oYJZULeHWGHN5t4acPS3BoCCWGpp6Z
1N7GsEQerijn7c0Lr+kYu1TfVZofGdBmz4oK5fMCXvSviwIH75LCpnWYwoMzyQdO6vr2VqncVo+F
QGAUzojqdcAKT/kT+oJm6pW+Qla4P8yVJZhEwW4qCcyTM2gjLrd/WETRo2l0lBgvUn5tK/sZS2tw
THwF9SeeQvMjuTsehtRl2aB7aJ7t5kJHv/xpOSk5ZUSfr0UDLoFnmLub5TfbXP2D4invWaQSAhLp
I0I5If7wCY8kpgldS7L0mRrUKFVnd54hRmlXKhegIAyRuyillZwyxZF59bRCfyMxcDIeB4GrgSTm
4E40/wYElQ105bqQyN2GM85cdfcnct5tNuSe4xrqMqhjyLEgN6CELJVQmRqnNXQUWi07cNfDux66
zOKcN5wZcdNow3Sfb4Oq+w2KBzmF15UMpOYFyLm1oORtX4VJtaFTEkrxBNMBggfI950Dg9vvonxo
6GNs7cwiQmOOYlqdXexG7Q3FsLvJms+VV40VBOSjbYILlZiEw4+I+SQmp2o72sIidmWL2e6PwAE6
pIZA4ZJFeAzfcT26q0Fp4nr9f2seN4Eq9h/IhL7SSIa8UcRr8hoWV2wcGQBU5FnspghwVf+XJxAg
HVYNt8z513DaJoQwqS+HP6P2NnL+F43xqX6fGR7Lw649sq4d8KTAZGESsgc/B8f+Nh9zcgYXYVGJ
QYTlX8seW7G/MJqEG122z5Zkwr+8nxM2Brq12ohY0R0+QPcJFrTYCx5sghdH5Sfg4YwQ/6RVP210
yU/XY7R93SlVkZugs4LLzxJwwTOd+VuFNPiGnIezPzyjLg8I7GTQzDvn2WNFjh9e0j5Zntt/Sg+A
nvgrqC4LAdwFm21pmjVU6mlMsDVxdZ1yWKUUEMdgp9DaLBK2MFvYG/u5MkZ3i22eHuuaf79sYnKx
fTJFVWkEWmOImfSMAfYWGlA9315sPWC5ipLximWQu+sCxXowm990unZI+9Ho0k9tnXbOCZsn59MB
uFgb7Q5j3Tou4v2Fbv6O/102KxVbt9AgqJOeuAs45I0uLk7rIfMyVpLkeC9My1wt4K5E3fQltiPG
vrktCWV89CxHrAG+bgTUDnbs+n3A8r1vsjt5+6kL0nfj++lMGlIqZfQtOIUJbVBA/l5tGt0K0cuj
aQT4RdJcimnRRwvaKJZZ2dY6ZU3j5lApn73r7ZEJl7d3DrePtY8mv5E+Rg64udIuGR6Rtr0KvAMz
hXnt5UVyZjUbOMpMSobwKk3K2rcqajwRqg0TlZ57E7YhBevCTfsrhpZ5l5NS7w8/G9UROKZgoJYc
gpRD2i7E1hdTllhwvibKDUpBZjoZn2kb56J57CNcr0vN0r4CmcfL1ccoFXEyB7KPCsUppdHhLyed
+HcqfGy3v8CmbdbNYzZKq187BYgRdyo7Dmu6tU0I7+DvupuMSb6FWGRzzKijTtay3U0X++OfXKTx
ZriWA6TBDVE2YsQQ/yGGoWKHj0vYvbgwoPGTvOfho6PtljHU/qQqha3fTqnqTl5JTRsdcgtVetW5
mzB4bZUutKt621IfpV9ciOmadUwHdRUVUXgEmp2XlRSKP0RPDEH10X/T9HUlSQWjDzBrBZz0Sur9
Fb5y8zokRpj2Co6ovDVE6eah2E07ifaqgjsTzweykz8E/tc9f7uOJBmb+u3n9DT3gM/Bm1vYMqRK
s5MLNPB3ZP/6KypyG1GTu107r0YvqIbkxJEbHwveK0PmtqvC6FtuINW5OnJ9Zjzt4X+uNLH8atlA
xViuDY3ePzll1Go1x9lNZt2rHqwlEpDnjFOw6OP/GllQHph9tTxw0p13WMLF7tRlCxIUG6jlzAs4
J3RCtASHHQiqcIQ9OTt2iMvCukMo6Immp3N2Xhm7yhl9QSbmWBAQ2vQM5K3HeC3cPXIGSPROtWBQ
Wfrl3a2eA9o4u0Xcv5mgLYtDRviXW7rS4vhlAJrVvdo8WdG8odRORPvquzPCGZwN80qLaRFlnilY
AzkXkxMoFvJj6hhFxfRNlaxdIONS/AxiYWb3YllprhFbtHQkRZOjZp3L+E+/lgV/McnLiazb+QQH
3g5DHa293I8VGijzuNhmjvOoAOI1Bo+GfxY+Uz3hMVzIjCj9at09/NFDv25RZYfP1ZlKBh6a8OU5
PjR6FSxXUX7oyiVZR1VOohaSQtI06/uFgiU+8OJBgcTtzQTKAXo11w46a5/K8QK/Jq6YQNea/ZNQ
ZdFXggkWMZ9ZKNHcTfI17kb5WDKcIWkuStuaYUrJG6EImshB31760YhLBpf6ZzVl6WsOJtCG1clS
8XncHuCXjtdOj0kwAbb5g23aaDh6Io6igo1NlguQAEYg0LiVBNrjedzUZVPZKdf3ftxD4QixPQs0
1hl9Mdsdl+eUZcTv5k6sh/ZOlXN345idsrVrPQ/2mS2fH0v00g25Tq9MGnvoL4IY45Nm5I8gplpW
YEngfueTvWRrArMZtk6+c/rGyXua41k7AWiUI2btVo94jT/P2krZl916M96xYyLYcySC9eIQ98xe
Z3Km7FLMoVpZQ0etVL9m/TxE52uBW+q3mQWb1eISU+6y50fKjFgkitrsHyIHiOgp2FNigRwiXiQw
iK38HM8EB2nWAZb07TguAOsIFnEM3HNRB0OaKQnkWtCMwl44g3+eMbdiUWrgdynWTivgTDxNP75v
Xcupw6JjA1OSoRUwlSKJd0YfTqF/SXtQ4eEO9Z4GmMhw2rrX24DUviaAXUBoQzNszHERIdprxGLW
1Jpyek9kQzH20HiGAcFE7OqECIKDgMjXZE/oDJIFYUcdngGlbIFNAK2buE5/jubC4L1ppkfLPIu7
Er8zLTBX768WrKhTf6Y51y5V69yDGA3RNiW16NnAxxjikldXj0nDrNCPVkIcBjGNk3twgH7OUqjG
g/4/I8sgLFatY6sCzvVTMHyLnkmv4LIUqi/U7naSlAzP7rY7C/ITCiqTOmSOv+O5Cdm9RIBowuJJ
R9NKtjfd0IUmPlJd2iTBVc52ZwhyRUfWkKNxOL7wqp8AAhZbctu5gOrRDXuhJxhopmp2zirybc2a
4oQUN3jJcgZ2OAEiG30UAinsOlqNlm1rQtGR4vl8AXbjx9wlMMXcqW4vR4Y18y+75R3uv2U13eCp
bhPs/pmp8RDfp6Ya2redQc3Ro3Iq+BP5zSgxmi2ricGRm24Nvs3i20deJ1RMypHB2w0WMXXwUxyx
tUyjt4AlH/15OOo2X63VzKrp+J2U3Yv2VPPrG8+nHeT1QrkEtqe/vQygCIKZFHWLpp4VfLpwk0hR
5vLr8Tco+uoPkUyAHiYwhMz8A7tLV6DU1JfaEMYSWCEOhWFuBOMGHd6Gg7W5PRnauD1//iFg3FEC
yoVIPSMiRNR6dOlKKKjDkApAnIa2eT8ITv9uDn58Sg64+qtifHZR6AHZyWS6E9CVvM1RZO4RYnjJ
XDgXXNymuKL+ekRrYAxuLHZtzuk9tHHmUbOZwC4D7DLKL2GDl2JbibOp/px3JzZN7HlNFyGyWen9
1yKiwnSjHy+3SNJt1+TIN3qacpYyC6iorU9R0Il1hZPsjluxt77OiEI+6yTj8rfT4J8u5AWxNU+w
/Qb3xXVy872pLubWeC+EHekNu9zyXVMQAm6XuE67xw4SuT72X00t0Cl99daXvIVvkfDPriat6Wyn
44HxKq2PMLto9HwR2G4qGEZu+9TZzVUC8fp1UrL9a1SZFpyJUt9ogbKZpMDlwtj1bMn4QS7rUZOw
gPJCLoMfbUrOUj5v6C1jvDUyg8lLGW4a+eOEq3QR5r6vwLBuGrXmBUMe3C/+0FSCWBvFUrevU0lX
V+rRHzKG2gO6nh62dWYuZDQNHHFp5G8pXVrjm6H46gAU6QM7ZGt2bcmEZGgwr7d47ZTHoSE+Gv/S
+/2Q1TVRmZ3thVcTxr7HFTe6S0H/ZL138ula2Uc/OTTSNl2uBkfxn0jlviIDshYoEpKXrvoo35O+
GGELj5in+eZe1FgBbg/loIYnNsV72yK3Qpm2iPJQ5x5uTttRmaLS/tKi4dL/iNpU+lYiDNa0rX3s
dBs/OFyfI75JcmwQ0I7w7J4baYptTR4sY/42SaQK5/0s8naSZkw9jMYH27pJsY8nStDvpidn6Vp7
MLAGTNL7OUFUlwSQ75meHIhOb8stZ/elShloZ9O3HZFONjk6EwFx7Fpipd4rMFgNLUWit05nFWAd
fKFPuhMnxVbfHN9CgcrkijXp2xXINp3s+NrZbJ4yx0W8A46n8Tnl2S4AKBFzNDRvYqHtqhBHjiVR
N6RfWgzJcJ1IDEBqnGlYrHbOh9+AgFbKlAPa3v1BGpk0bogO/iyo4Gn8jviTnKAdaRRGJYcTiY4i
s3cpw4asR9ZBDeQtZSqsCWqANjHOrY3kp8PHugLL3Z07jihABX8MJIAQedkx9l0Lh7LaI6kQIP/L
0ym2aqMNN4SQjxovn3+ZB3oPBAJvJjjdlRIwnJZRfvaXEcYE9/K49mQ2dFgP3LExO5Ou0x+W0aLx
HJnOq34MlojnJ3IlxvagcSG1w+ZHdazy+fTNh5wlCCOfIA0USOB9d5jCO+ZhsuILZ6OLmXtzkGEy
Fii/IATn+XS5f1JVAX2JgB+JBhhxLdsoPx1z18IXSzG5AYbU6zY1Hre5iwAxGogj8mlt9LM4U3z5
I3LCM0fImbzcDuZyRfdNhE86FOa9uwhJnYLv2gKFPP+X/nor/Pnk5boTH9AIJgSsTC6fM5a2WMAl
kWbcKVyN5ByAk5iSEUBzTDResP/yw2rAXy4myW75PbMbTIz06+F28C4PKprpoiGidfxOGyre5hCN
ILjsP3q6V+Cei/bRuqMKuZiJOnXnBmrrvGhEPxyGe/3Ouelb3261RF6LLAPCPgec/OGF8td2ohtt
dqBVu3kafAun46360zzxTaAjrcgXEoIZR/O0jR+RtyR46qmliuA/eXA2i67BnC1SwQtwV6pqRMG1
9+EdVovKTGzUJNX9tUJtEYfaq9oBcwEzu5nsDoopbQiVKz6qvm8MTt1d+LS1o5QlzGkKsoEsEWYN
yh6xvLt8oH5pQToetp0gbzNfiwCcX0xRIFggTCQ4iFhvRmp7E3+mkgvpYmDurM+a6yy/uxLfOR/g
2povcSOIDwMLompDya32t0WCkxD8NkLpcgmAWYz601PLjXgWQAT0TXZypC8RHtsUz/apYdgRuZtV
q91m71cq9y9wNGNhuLWBmw74UgVsGaQJVSKa+ONZjr4EY9RHkymW02IMYO/M5BP8mcLQ8QHYGkRR
gDTHAD0gkB2KmCr2rmBWFtYn/+JmXZucd/IifAmKWGKbuSr7U1lf3VmFvbSQueMs8ltKITGm4OGs
U6WFVX+4s/UwGEzpBvj9OlIg9yfkuJBZ6hRHbAom1RccDmkGGiafe6pts6AuUojdSk6bec5CDSyZ
AWvOFlVNC6fSiVRwhREhvfdOCCCM7d8YutCIro2UAcQ+kLlA/h6a4Ec1NWNsvfW7T4SrG5LgGcfN
ko0vEqjGr/yBEbj+uwDmV7ffoYO/R/NxE5tWBsjUU4iyu1lZ67MXVC3vr8FFKobFmXI+9OthiP68
ltmJ56YwYhBtZ8epCx0HiYU5FEIYwIB+PgFHUh4jHHC4IKlKEOYkq0VVVvebj3LGgd1Dc+ogHyEj
gQENiNfDS3o3N3UGT5QJSgo6iV3Vj6u/TmAotu9qjAyyNK3OonrHCwSK0j6SPE5ffqcByZv6qJJb
o+T4EQJqFFspHtignqcGb5XZtPJbQNKFioZBBm1QwzEzOgh8Q8GcWtNnucWCXW0Ov0i1CazP0fnh
Khd8ClUV743TUoJNM6dVJ055UCyxN9eQJJbxrBu5n+zhOXqc51ydTBigsCTWtD9rMfDwfvZzwzQM
xpfy11i4F66zLpuhoqExoGLii9JH1s2j0zLHit6YX9mBIbrXMdmI3bDCxAovBicrJz/L1Fu0RhuR
hQjsZFpTEuDMW/E16rQ//LiqBlu1gEV4nP0032MZS/waWax9XWzhL8t+JspCn74tJe2xxVjp65RE
4d04soRZXNyPp3E2e4Hexbw/GxVP5nuAoQY+B7aXHSDWuFwyMSBa4RHS7wbw9q15Q4yH2tGVYD6Z
CnZ/LZ6SAVXBCGWf8Mc+LdJzUwJ1slvNc2Na9vsHT3PsUHPgqv159c3WlAQ/58MuT1eDz/ShYTMH
MvHtVAgwir36mk8VNB5VbSOxHiG26a+25iuhCMauODolh1pdDz2DBSkJOJxsehwDVSQ59g+fKyte
q6NT2CaiooSUwI3vOG0znuRf15FBviawvBELLR1EUYmVWZJnSVJXxsmAssXHzAPNkYQeVVbYTADx
YuB8g3nSh/6MFlG7l+Z5MxjmMhAmq7LQ1JVMNQ6fKRQE9iKJB3mlkvvBnJc0BaD/r1x6Q5xEaIpa
O45M1H5TeqDB30ll903QImbLQC1X9zJ7laBcNWIgZUmMayjjQCHWN088qjYGZUc4vghfCvwxE0Ci
/nWXMCxExh5+pd4vqYUeIWGaJxUsGpP4KUoJXj5qUGVBgO2dcQla9aSECzdktqZQCsEfAB3l5cmV
zOplpRdl+d3huWddJqgseyNUYhg1lNf8ic6AUoRsaoHszc4vf0uf9DVcDWUY5jl1/AZGFmAUqZfy
l5aWetGULOgA8bmP1ikV683DB6qZaMQoDhNO2yFLTwuaFVC9k/rOiXZQ367GtPF4iffwc2joWv9G
DMjgPvM9dyled3s5DTULC5Wi6VtW+ltI4DzcCBTnTYWVY7oRYOIHrgedbzSzFURtbeYloC8/9ek9
Aad/Rg9cy9Nwi/MPXJte9gjlwAXUy0dErqzihwk05OC+NGJU5CUaBMhzQ0bhZ1hzKF3mcQYKocVj
j9D1Yu7FVquXgQNhUI1UEUxWy8shaV/jHJtpfuNLeq7b7KO0tT97QnghsWbW+6lcbiSne9gUooe7
4lF61fxkyDjRaJF+ZBLy/jCc4/PM64qBHmEQ5C5D5j+7g8e3qg39aTCn3zRDgnXlD56psfXqgD+h
8ptmI8G9E4TVobIYzTbTg12DrhO8nXsZXASDa/48O/52/IIDmw3OnIyWFAZM+31UvqYS7RHp1MKW
FCV1v/yYYSm2eOvym04gpJR1BGhiAYPnh9h1H9yzGJyDIfQP8pZzU8SAevH8GE18vNw4RrhTFMik
k4GEXnoSDrkQn8QunI0qqJaspCRaGB+IG840J70Aqz3Lb4bfOZJv9BU/nbFan0SRqnQ6SwmXfzGp
zaypZwAJU3/a7JDFH6jXzoiIIddyNiWBT7snk/sUD71WmVHO6jYM4NGl/0Tgnu4cySMWwbCAjqUJ
172Q1CcWUpZN/U+UgE65uX/FwylPEPsD3qv8OGn6mrzYn6mW+7y9nbbif6IshCrFYEdjJ3RSgcXw
WOM5D6wi+RMov+RtWpOn6Z2feq2Io8sSG9UVPoQ9O6VgXnFcJDQkdsH+gQkzEIUS6r8cEmrIwn6n
IP2iMF45qOBBbLRz8bGTpLffi9Cd3hcrO22Tto5ORpU4YMoic10AzFhZZw3o9DlDudre6RiKuEwT
CxS5lCNBeInFNIfhECSFww2p1ebJIKTcF0yzjT7cwr8eBx/IvpUM5PT/IH/wzxDjrmJtjq1kogED
O/iuyliKvgxfWw649d4VpCRFEvlZ5yGObYhIr7lDuO8fURSsy+RmzL9IfSMgo5DBTwq1GpjTpfHl
AmSYju5Cn5uGHIHLwkfYv1kbSGrv4E+xbUOLZ18dk2Ki0LSvea6ovG4yLbYDcalf03/2qwTfhcbl
NTocvgSjKbZmBSgkhLcfDC9CViNkKxOlAZXw8klkto/OAn0WKePhsN7xutdyBbsYPo/xJI/JgoOQ
mQHFV03j5T/R649XvRyGsIPbsy1fmh9ojeKIvswxWNEPD+Ys4kjrXaLCi4MaW5NjqqnmF/C3Q1lF
y1W64qv1eK1Cu8KS9bJacGJtVcbT+mDdQ9U223rbDKot9Dty5l+Nq4P72ptC3T0rwt9OZfbr9Muv
3mu+ytpw9FfneRb9yoxAlMvuqzxX/TIJyGQfu1qawRg7Xh6kA378pQEqRb0sY6HokX/totFr4G9G
41w3wyepFBKnW8xDEWDq/ZOjSmQKT8c/sqToYWXAnWo3MC6J8Ncm0589jcI80SppwMUer33htycq
URoXB8Q7i0nqA8mZP+Gyvn/OOm2TJiL4lJkbcI3LHd4114tvLB8vPHt8ug00wNgF2JU9Bue6r0pY
3MXInFw+YK4zKYYefDqy9I2v38A4vGMMoKBcHN2e6qw6ma1C0LqJv+LVrOlpTNfc0JvZUUphXFnd
RtEsRDQ0YfZRRRtBNw71aAfrZsJWyo6xgkkqZi9zPh6arWnSjybgMsLB3JawfVGMFC1Sxc/VzR6L
ZNHIoxdvOY4P2SLRcVKdATcd/5ytBmctnJMJw0B42uZwoynudTEWlHXyTLtUpw8GFo82s9pP1iGD
wQMD3kaXtbshp5QYAFd59mv5XNVUtkfwwdmA7KMnaZcNN3mONmUX+s/UQ9Tepm0KZlctAuJfc5mp
6EBdkfSPqNt+1OATiVgI+ckX+tQKcea1bvGLYhe7EKlP5XsHxrYbj49fBqiDIpMEr92ZEH+949AS
burAguSY2AE627MNYIPTMSNQu9nesHLUdTgC+H7l9ZKgm9gL3Joy/PYguhzX99YQO3k6/i+9e6xx
TWVh5gEhi9i8B2HDsW2uBGFwFcX2xuZP8fAyLFMnhDQEGRhXIJ7Pa8t3r5teajjDeWSCaYZ8ZZwP
tUzz9Q8L3M2iN0Kv932LGp1rrib1aDWp1+1kY4OK9Q2EEiISwKemMgWHnMNyoNoouZlTESCGF/gX
DDLynjOmBvOpP+aTz9u6AEMwIrbV3lg60tpU3tGBkiFnlgy0+8E62TVSC6EMZdvNVTAiITsih+I4
wcINaYOTAaLFnKodTEG2Xr2g7OnzQMgehWX1zT85gD18jRsFjdgQzcCnkb/Mu47au2MTGCW/zNmv
UXvJHdZsd8z72CBTusPGy+9GYDgCZ0/X8gerhkaqKycysjLI1gCbB7bkat60Kd2OrXdz4SmY3NKs
vI5yicf6PFvR6F0g/EC23MqtMEg5Lo48L/meMeS6+oqb1LyZjTENVe2N54oui9AvMEK2tvhL9CpV
I2EqrLSsB78Ept9Nla+yPJo9r52PmwlxskXaVg5rxWrmzZr2y1/BcDAAw9Scj7q66o3TS18dItQ/
Ej/Cm3OyXwmMd+kWhNrEjdyLzqzbQPw7epy2TUYeg57Q2E5bo2GgsRHUBa2d3Lb7yDZnpeIpwlC0
jhtvrbPzBygZtmeqKi3dTXThGTSqvAoPAd0KUccRVdj1uXlxLUChQu5X9Q+A8dMvmuZDgEwjf+PQ
xapNjuwXw8ghUeyvAp/ddWz/30x9VdXBa80HjYIRdgt03FoXTHSmPN17HN1hmQnzcjpPC6EkyaH0
RgNDuDJhAN4O9xyWbomIyCZ1Lp7bvQLiNNvffSKTLjBreDIv0crvox70fm4mc09MZ6UtgTI8KkQd
p8nXKTTYOXiaHMlAZS9geXoP/2uRcCLQSgpcW4sTqRwfIFKZ4SPvFHodDhKHJXeU6Dizzq5jN3z3
kxgeUFSswLBn8RnlYHNx2BF2R6Fgdan8fnZacofYF/o0IHsyNHyLnxHZmou0kMpY1jQ25InaakEp
wbs9INGQNM0RRnfllqEpf5xn1szbfMU66PPGhaTSNtcOin0maPd7ogCxKVInEi53LalEif68DhzJ
N2N30OtIlBHoAWaYAAy2kPZNj7lOGA1+gFhYap3ztjy9AUUB32nUVaan1zNBHPusn+iVKiA6bYIB
VqiQOqtk+B0/Qm4gdNH6Cq2FT/AbZu5kIe9uIuj7J8lAmNDusYKdGCxaZTsZmUeVIa+SG1JmSnvg
c0t21ZJGLdpzHXdU2YGlU0gb60Z2uLC+zWepOHwipHndggSTNLzXXFWIDzqJSUWa5HEuV1/vrs0e
CsSQ5XNpP53ja4GfkFczuM01YrxMdxB2IZRr4LFPL1yif5qDNp38BzjtH9NgN6swGDvfXGC6NmFp
5mU6W5yhGma9kDYT2UD+UixR085s+0qNbvY+TMOk9GEe5MtIH8Wsq2/s/xKg+bkOYNZu263Moyk1
ShwxKdQPuoE/tQM4OjqAh9yd5bV1JUKyuxtwIRTHmPbf4OtKv2O9qqg1Fd8f048mnYEolF6Y4YW3
mwn1pmcJrUxkVU9ruowrDR0ZnM+ldrLapcDQghKm2iPLm9x834WTdZnRHsH5Up8aeLPcwzOpGwlc
BtmTobDUY/i6yXuW413my/VTT1ors/lTUQbeXAojcHx/2+y4l5S1Q8Hx/+Ed3Y0WzHyEXUpeLjkY
9VwgwOWKQOvCWQg1Lt5pyWU4JW68uZcllW6LD9Q3WkTR6e4so6QxaSR8OGRnnTVVsAdcJuyZWGDd
Ah1KwJ1hqB0KGiUhybEDrHV6QUgVjC3ZvpvmYJCXsd6NfskVUOTHFX+Pau/T06Qw8BLM5M0NjZQx
xC72sNyi4fJSfEqsOJNoPqKpP0wVqjYNscQyymAgXaj4G/E0dfaI28trE47HSYvHxlhj19MiLu1m
j5F1Oa2oeNyXbtO3TZF48INLJNdeaHyxj2hUuJWbSJnUM+cu/mbsC+qGKNw2NO6XNL9dlyIHoOma
ZhyyQnYV9xemoaukyyfFtEJW0YlLu3y+cdabQYcArxJx23OZRI/EFrb1gmEQoy1FQ1Hh56Or81b5
ppP9qUPerbxmpWD33kDnFbrgy6TdqskYMFo5LWI5aK4LmdqSnb3tFNZJSwr25u6WIw1xRnslNjpQ
gzfr+F8NrC3BVuNvy89lvE+EY38L1vWALv7eOiApVj59QzSEWlcTuukDrkG3h/fUSRPZ1PdOcsC9
ALZG92efE95OJL7GEW130O4GeFb41umxyxT21lBGqphzc5HB8izkKJwrbCLVRFoZk+GWnH8wiA8A
K2MPZmYo+bAAsjORdiMuu8rdX0+cfNEuJ9UBrJDKspcCjm2exe37nRmjNCyq1vE4Nin3w+qebcM3
NOiN7MsTDU12ybCs1ojcw8VkJhOUBrPzlw1DBHVz2YEXIkUPl3grEL7mV1n25AYrRZ/zmxmyJSIk
0miVeeFUHEcoWwq4dOpTC+n3pwiCglc6xq+AJjz39duWOXdBWpUoIAtSA7okxYwRf+Pfyo2hcIC0
UpHG7Lfj8URKd9oJk5clQSOy9dQVtnB5vTvU4QLgw0VzMpHJAwYXfAKXwc1O4dYmrSbFvtiXJVzo
FN/w7vzt5aMkmEXjjLHyMWUxdKV0OC5kkpy5xz1yLGgll1zemuORzV3OckQ7z6jLsfQkO1t1wvvv
jVu+rFU2Gyw+Wl8OC4nFvo3g3dgIKT0kE0dbvI8748NFBjhpnjlJ3VZvLY3rc0unIONxMnB14oUx
HF1/QXsvhbBAYTnm6CMRiPEJgG3OQI/xvBgYhXe+5qIWfgyLUqMJJwgzKMjw4/0Ls8WyhKXN8Heq
cHY7CGKa/ylc7Zu8RcOBUsHFBTZJ1SI4TZRwZroQ7jiRGhSwKFxhbWyXdaInwVvJiw088YDnHK+e
t42uoyeBEq0EfwvzYVeJcp6h2KxOuOC3+N/YEfTXzJS9p0tqrj5FwFzucaN2G93bLqUle7oitxMV
utkmv/3I1+d3xaGqdEw/aRd9VJn16Q02MTHfr6vphX9/wTbDtuURKkcb8/L1pgTj0gd+ZPGUUl4j
D8svN79ikiZmTlFkkLZfr0I4ltqPDc6dzPOooh59DB+3irENnfn54EKqPqby+817OpCVIbGaSQDv
L0HEFr4IwTbo9GJ8yKk4Dk8167AAV+2cyJw4hM6MMcP+sKOjgVwd9tUoWJd+h4JuwCfzhpLvMVXR
V1Hei1AwifZjkPWM7inukVrW0BDfFhR63tbGZcRll9AX1E6FoVwy79b0L0Lxc5+OPu7AYO5DGp/l
JYTGjqbnlh/z/5KqADgMftZRlXbTF7azt1E4oCQMPjzgYkg9WHv5a8irrD5WFwATafd0c5qprjCp
CZjaIWDhW2L3+HDWo3ePQk4SXvL4OEZSZ/theMSkLi4S0/ekDnI1VjQGF95adJeb8236vJZLSz9k
QBDKv9oH/5/IufQaWvyRifcLZxnczSeRVWncsmvfX9kDi6aDjkBy2O+4F4gFg3lkVJksmakWhN2i
WsQQb6K/A8iBNUYUWThhZcDwKrIZd37YdiXrJajlhCAwgQwWhgEqv+SrEjJZwhjGz9AAXEKFgua/
ImP6Z6vpDbH/Cd/Q7tipeEnj0XRDXMbWledkDbF4cBiEAPZCWSTtns/bEIjY/nxhmyS2E3o9NUs5
FSwrR73VNm1pSUTZacFaJ85bwBcrYtKN4k+lS5KaAX4k0fV7NAogByofMHN+wKW0TL7dhPOQsm0s
4GFesErbnvcBAcUimbQGZt+NUdPaDezgkBjVbuTFZUaRZl9l6rqYW157FAyVSZe6Lgwfqi02pi80
C6iWzCYxgtq+aimYRVSGK6CtrEnjNBBW9uA7Gd5EfH0cwGQkarZdzr50xA/TdAWZcQ92mCML0FX9
C1jK56/4dq82buC10X5lo8hLZmE5kdkcvka58GS3mYF4HC33qq0jtBJjuF19iv1biSdXhr3PDWAP
CAsfOAFYij/zj0RjtDqG2i0cm6oHT61u1Oyplbn4mpMDcmdRIZhkZygRj8f92syAOZfVCJSd+UME
qTIDfFHxth+ZicJejhbHxIiI78iccKgGBBxveD0BhJnA39FFEU5j81J2/q9i8AzWQzyYiMBBJLqN
SErOEmIxbx/ivj7/xiaGSMR9vAQQP6crs/5sD+tER8qqooCQah3fJ0QBOFvyWE7Sb3AjlnXXFJ+o
bTjJEKhbipRqrNqGrKdUi5DcLUrJpUpZpK/G6niPOjUbayQqUqA5dHJsGtxtBV0HiAuGG7+RiirY
kqUKlr/fGv0OPF10rOzCKTMPCb1v3/ViFIHRczUur2HyyOc+KDUFiA8hG5bFdHyQnYPczjisAy35
jRQuMvBzHLBrLUmJy3LMu5InscDKtj0Gh0EE+QXq1gerpyYcQa9v7yVKjQppytkGqQwGdAvigiyR
+gth3ajJ/QM3MA0E9XTPtLeykaa/Xw2Oasl4bCulx1UVVN3cAP0z2HAewAfPTe2rNXoDkfLBhbCN
YJ/fZUBRfdJsp0lNs7P8PRKZO74siKSUxsX/p+4Rl4eD9JTslJU3c9p7Yno0VA8dMwOFyW9C1OdA
qHzRtT+oFS/MvXywK9musK19HtJbp+ILtqQ4rontV71IgOZjI9DR6Ne1VDru1lM2yZAOgqEZqmbF
9w1XyI3XwM90kFBqZcg4fo7nYwPCE96wQvQ/BQVKlv7NKvLpGVl79M7GydPjl1+H9ZgDrN88SqqO
MUUuppIjmiaKTgbEXvUmIVvK76IlFzURu5v1OC9yrUV/5yyywaTAwvWSzpSrIitwVyJRishZvNO9
ZUgODVey0n79ldXIkYcU/mF1Rkp9PWwNJpOWH1dqVGdPNebOwqof7u5WbmaYP5PDazH+nOdiHNS5
J8gtnhwphGF+P4L5M4I1pumFnJnF7UerYU6U67GI9dzefHXggqBsplc3EgdqymWPhtHAbYcbFhJg
Erh/+A67EXJjKveiWG7VGrSclOwNDdAHOzFDnvqo2oOn3/GrIq6Mh7h038eyd7yzCCYi5nibBPBK
DQhxZ4MghL61nyij7e3ZkPsvTS6LG5sAMTLUrsq88/RZHgfh4IoUksmMexKG4V7NMdQ0KxLclkhg
BfUAm+pDwgN1NuFKWh/OuFAxrkYI8R3iFO5hO7TwDK2oG1TiDuK+LeM91183XQkG5SQeaMcj/x2b
mMFsuvfXdi+9z91dksCGZEg5D6mWYEfFKk3uXXegRwPAzRXp60rz+DVrD9yIaBCuLFY2T8Kp9RzA
baplzhMuSmIgd9n7feLwnSd1xvK7M3l3CESgIVLPRevdvZD1DGBOW6f04gEImnLV5o+hZeoV8NRV
N510pzaNPoW7MsTZWXr6jsvCrrCSIAqC/uzHufaE6NqJJ/RNBJ4IeUIxxzSdLgX6Pxhd4VCgOlsf
rpsqyxcyT/5vvAbeKkcXErMLuAsugE+ouC16Xi6Uij8TQzThpyKM5SLdQOz1B3Xno31D0/YMbqTn
y8j3tKHBPhpjjoRNqmvFaIL2pP8tdeX58tYjSyqTKNHYlgQyfS109eSWUkRQy7qm1X3DPcpVC7lt
H3SZTifzgLuY7LsdUhSWPpOb4nPsQFKEkDTbxkoTL46jwkgr8nkaD9UFjbIUl5uFAkJcLoLg/n7t
MmVPJ/YTn3vSqR2v+XLmoHnQcd70gO2OnJWf2gspU1Yjj9roDr1NrH7zYmpq7CIf6LcG7GADU+KA
mFIox5cLrOJpBavQcA/fD/topPhTWt/xqwd5bKBdlsVCKwVlQLc8AG1m+cEQVYYnJQ1vtP2QspXS
yCdmYD0oiWM1s4C1IyrXb/cDbRE8nTYoA+NPZIe9He9PkWOE7bU54VDwrQeH/HnXUo0vY8PPxJY8
9CQdEZHLRVoHzf6TYM7B3oTNHURPiTDA7bhP5R1FQgYxNVn3y1kAOr+couHgVB6SISq4Jt2/9QaH
u9K3bS7ia9TQ5PFSFdeARY1AlmvVV/65v2V+SFb+5BcaM30hmcjG9iANLKhAivfLtXQLSVwBcEYj
hsNWGUGgB9jtCfnKeprzD9KhHumyiVFwLyA7iBiRWkahoTAP8KtLsIn+WDPfackg4f93hUalq7Pt
povqcPpSOspqUtqZxe9IBUdTOQtKcn1cyJ1ZsMcVDcfWD5kQRE9zVsPEETbzAki3p2QTiCNLsymU
l1B5n72P+prNzbalqFvOuRwxhPwKsrF+vqjeVEP1nxCGBOFO1I5+tXN2zA6YqR7IlsgBsfzxdG+D
6945vbjw3811/G+m5n3NVGv+Xb3q2uSgVKM3eZCPpj3D8jKYHGScWoX9KL24JqBUH2Z2cF8zFMD0
5jQ9q4wkSiIhxK8hns9CSZy92TS1gzRnwIuKqktukpLfkRu/TLdOSV4MZzrLZ3Pd6JLg9j7C9GN4
cEY7o84xsJSXvLVkFnQeOMneFa7pWQWaH2/zGXjbG2Lu8yr802VaosA/yq1CoOOckJi20WiAOuEN
FQiTMEuZ9+VUZW/Bnbns4BHMfAXpQikSvxf47asCOHo5V/9IAW0yOD25XMdEqVGlHlr9n0zQJ3+K
9ax5Lviym0zn0GXx/YlYHX3+f4ocCGp9GrS2Vuw/p9lpvGwRm7ktgaSBeXw8yqJBBjZGGNpvuOWX
4ZLI/EHKtyAdizBZIx4PVvL3kqqnQpt2t8J7j6MyDASsaASsAsWxy/JPZQQHsfhDO05UoOetCvpr
xziF6ti9yjgTZROVGsAcJmdYzU3Kj0SbStRq3Hy/GF6/wx/SpJLO+27t/cjAf/hHB+8+kky7RDI1
Tgy8TFU35HhEtY3M1TC4RprTu1CY/9g3A4ZRqIM8TLLemqJlchHYgODsUshYfP9hDBaqtmvycZys
sISh+IfcN0RTy756/UpH2LNIXJlF68hFiPNtwxayfNy4Hn/S00NWUrg3XlIjlm+dRK+QvsJ9I86U
01FOE0h+WcQi/FU4gbYRVUM1xakQ0hzIooIwhaBr00xVpqR/1h2AcbAHhDxv7vYLYOLAplCtTKcD
5cwRpwenb7It17ArlU8FrwF+io1vyBwlTJR0FybCeLvYjBbDtbN3FWK91BhpYBAugf/BJ3oOgUD5
TkrdocoNROgaxwIp4Vw2mrVfC0dONJuMzTczNax3hKeEWuVuAS9pTFnT+TLeznAXu231xdb0Cv6B
uz/CU77EcYGBD9WMCeNxJXftPjxTAwyTLTVgY0YeTLfwJ3PsteHSJh1Rn83BSnG+T125ARilriZT
+OzVM1yiu/1lfrmu9HYTY6PqrKAgIke0/h6X5hd+uko61mKjCstG2PetmGnT1YiWRNcf3y4Z4al0
B+e/4pLHCccJiAxbemq3La1d52xhaHYt3/n2urTPva3rTOQaV2XkEB3g/ZiUlpUD7GOwKwDrtO+K
Y6eZ0BHB1XZk3pkKl33cKrt6HxPNPn5hZ8wjbbBOi12jbQiqkAP2Iw14BjvoYM8+Eec224hiX7be
X6fWBpssrL9LsI+tpZeOQA8KhMt+Oe0aJ8kCEW4fVUoV2YE7UDGDTSghIMPAV14JBZBI3uLBXk6t
sSm1xPTFQYjnH7qNvrwsOLEj+eKK4s0/BG4i6VTjrKmbZ+f60T/ktTQsVOPq1DvSZBhGFIDQqQhT
81DZuWNFZrJDUMRZjmHDRY/y1YJyo2TZ3mzDOAwkzJycHpFwaQRUVGy04GHop2tt8Rh9Qzm3MD6r
ZaY3qq+3GwUZS/hmdMwUf43G61lULgrj7wDv9EkJi/tpbKT9ndcySEjbXiDiK+XJtevpMnw5oxG4
Bq/Wa/0LBH/mev4a3Q5xgqfL2LykVvb6zTfKwFQGCpipb11oowTUttdJklq++SlfM8CineLBdIFM
mxRFS0qVkMkXUD2aPJrmD92bm5PLKrugThIJe/YDlsEIf82cWg02BxBqn3D4my88YT2njR6f/aHZ
C2jbtYwbwjA+6H1GEp8as5tCp6XTVvE14hn0aBsaopWL/S/buAjQPipKj3JTJQmNtFgHAsNkxrEm
mAnX0+6JTgI9pIeh4ASPG85O9grU4xr8spFnIfU2lN/qJPwFirY0TsACu5BoxeFpF+xHx5TW251V
mRRVChwc5/M1wHMH9/wDxo3+sSByaI1gLGJl3Irdlu94Wm1xhw2AUZLWMJj5kNRdwarP5RY/eU1j
05n/KP+uM9ZeEwEjoxdQVyb+YKV7wAcydEfE9ieVtDjco3Kqhp+j0aSSZopdyEShoi0e2VN1ufZD
/UHAoxqO7BUj/tYJ7XSTMyWjFygEKajP+MwMxFeIzLwzB9TEdWwJ0CDr+LvqYfqcHqBwzOWMure1
PyYBAQQ+EMIY0HflM3BTs4unzp86xb+uXlsGUTptHml7OZAue1gY3PYyBk+o7Uv7Ck+SG6KK1zT/
zqnY2EJHqShIBAz6c/zQP+SFF7lZOpnDk1LC9GI0lYN26da4w/VxXGic/9x/D3hAuGnKLI3GdVZR
M/7qhZirZcvgoziJCFBIoyDaNfaz0w/OfjL+2vYqZ9POZsSVNbxZAtESzNbVAe9khCVU5B8wfbXe
uKqZJ+xeqIWQ8TnKtuMIwAOR9pDr2hieQSBhnnplu7kTpbGGm8xmFmkuqDqg4tYGEhkIIi34FpU4
kmGKeHBwAWreR650RnBa2h506Y1v2Ov+m7AMTBM/U92q4y8KkglYDBdF6vz/mVwwrIDUMgBRng3o
1RrJo5nB7drtvfg8VezJcddyVBU1nfKoyLa86MYBzg7N2lea/shMCfqTAia9jsUwK5zOgQpzeyCY
Ld1NjFbAITZkQ+5r+DKrsypQJgK/0GmHdaRvz0ZYb/T4efBdvKk9QhPJzqmjmQIhyaTHH8R/tjl4
tIQVVrr0WuxRtJbkQf2et8/OMr0AFdVHpAPoiVc3tSpphuFyHcU9AMsS2E+S8yVWATN0SScuLn7L
PHJ0vwHfqqeal8oN/S/f+HbD1QPZoTR0dYqV2e0ut+hxkLOq7DPsmJGeFa8Srr2k3zUH9rxkTrxh
mOvbdyg8aKrvBkpOby5MrIatiu0o3tgZgS5E3vUaYYTG1PhBbJXE855lottr17KkSgGx8qsPVW6k
nfInlnjGUc8htqGxby/PgdAEDNal5yzqnKLWxNImZJkEWmdV0UsyQteR0QpWQVAi6igiuIvzSLBa
u+5uqK8D8Kcx2yG+flTzLq3B9EpSndbD6B3kWAPJ0Q0ITJhXzDzhd0yNN4efRU5F5rxxA0KVepmF
h8pO2oLX2OfczeYBYf0aof4OcxfJi8emD4VhROW4jHrbkoC6523iKwHcqT+WYe00My5RU4/58iF9
14JaJZcN3opki9aRLhLBEbK1+gzfTc20gBeohMq8CF12l5P6aFLumfJiL83Wn3H33fOpP3NUEYWw
sdQVTz8C7TJGA0NeVaa+avgG2ROacdpqYd4szXO+Hg7oQxb/1VJRMPbQBbyPyhPvj3jUKzSUBHey
1wj4cYrf4BcyEgar7LWYIPhXK1kc6xSh3usQkUgtseL3KpT3gBqHl7jzkKsPGrYmTGBftW3vM998
5ofWATS9gagtvfo0N9o4j8SiFKyQbvPS5FLdNJkEQ0mkw+lXqG051WAbWMWAeeYViZIITDDRyAEr
GUhMfD+lBHpCngnm9lCS/TbJzEUiMxMZiSe8Ij84SGoxjklWuQP5mYQpxEPLIp2BBSqjn5cYZOsg
r+o/jcdtocmDovf6JHPgtM68S+6+Sn9aqQI6Y55SgyNGzARv471C4clIVjzTI/0rdIJHLmUxGoOU
goLxfVrIQn7+/SVs+QeEt355zh1O/xzQFYkcTYRiskq/PKTuM2hJi2GqavCexhZerVMRlTfjw0zx
Xh72uRdfHDIUubtSszAbNbp+k8i32azb2xmHav0UuO/CytyzUlJnpAiBynBwg3/c5nHpBPCMrgAM
KuX10JsgYHFGOPqF716QNdTjsSsMbwbNWrJvRriwKAq95eUAUxdSb3u2s4W3bf8VMkeXERx0SwuR
q/Tx3jT9PM42SVc0IdHjOORcdOKD1Pvl4Zed/GadzFTUslKhshSTSa2LP74APvKIXMSSklUWjX7Q
hkYW9o7jdcCVRohHbRTTnIHBGvIa/IiaBlbsh0duO+rZN+dIOBWEOtew/1V1TlS8q1ilwLKFmBOo
fie3yEu2dwMry/MJuMxyHYZPP6p3s0gHK76U+UPneOsmVJU7UFfYQFL2xLENIxqxZwttGyi8Q8No
UyGo4s2tpUIeu1d47U5tJjuNl7LiGtxyF3V2PZkAsPHB4LrFuEnDeUWvGVyl7yi1gfk56SwC22GN
ULFsvUwG2ULdxLR1rFfH7qkf8xnCj5XsmUqN2S1SiN30sYe1Fus7iOk6yl7O5Hj5/xktwsxWdfES
r7L4d7NNRzbFOuWQrsTk0Z9Tnc85jBPH2PvejP/zcWFDs5U4G9WCLZRQ9BN2suAX8gEVyo0srGdd
fyIOTmnpVxwu2LqRAlk5dREcLNs8F6piwTfXtUPZCfl+KIMZ3Sd+itczrMW0JNcoYfLVbGn4BPd9
EkqWVZD2EuagPgqPgMeG5wUmLfSuRGHE2TqseZP3PptTbjvI7U19AXdZ0RKVbm5I/QMoUvDZjeIT
b0PSEiBLA3SYKm2JRmKm0lK9awIdkt2v45FDiAhX3/KJVIS6CKt2VLjZR7/mUtCs4RBjNrOUqrDK
gVIVwGfO6YV+DPFhJ+Qa/rh4MT+mxSs+v9/CzuOvL4Hqh8xYs80k+PVuGZNEoPMtRzV9V/xvKMaN
k7yBbBko/r6rsvbSw1vhAh3QATHbasxJeBqwOVIJ60+zj47CuntQ8++NjJlNMECyT1bvdx6vHUf3
rjvkv/CDgR7NbMj1EqkAfWF/R236PYiCpBUns3ud80q2Xlj0SSq0jhjiLca2xtz3K0ftxBnNcXKE
+nRoYqH4YHh258xI/cVy9X2J9kQ9CXlqyZxp4q4IO8oStH3MRP7imD87mWk6x95/kP0ipK5UlNo6
i4JUHeavkUXlqjCfthgAQGB2RG59Jx4XoVtbJisHkYb3bXWOdHk3XOmzpBbQxB7bbvAFISpJOALT
sQvDMXIu7obe4T1Hw6t5CNnkvfR6LNqexFfG3aMPmz0GVaTnP7VChTdJa2FrSElqZoCZBFUyeJuj
Shft4gqGXHYVS1VdtHT0MwQum6itPOfftzIa69M3J1kHpDEXjMXV+yHxCQgKHXXkVqPoK9SG9V+J
LTYv8YD1INsI6MwZhKUoHGYCD7GItvTxYa+P8QNy0UGGAOEEuwT9u3zYgK7dvAJ1vox5A5xLKzsJ
3oSTkuCSQkhYsC72HJYAzXzu0GrugDaWRQxqx+hmOH1N9v5DrWYHGDnKi5hemtnD3dwpUMTdCe1j
qsw9MN42yRTDrEWC2E8YxDiba+v95NYV1XzkSw0rRFb8ZDBzZlGKJz7AdEgRVdXIYQvpawKGozg+
SRLM7+K1QrnEEsHd+MIIfgp14nov8CGqB8w2fF7h3eyUti5r9JuNWcQAVF3S8ZcBxx4VzXfVOq4B
IVNdhz1deHXOYIPiyber89zycly2LWVHmyaxquzIzDM70bSaOCpTh7+yAdY7QF2neLYIOL1MuVuf
w/0mTMqW+0Ga3rmZWtU6aTLa6kOhYRfduIvouX/jqrYQCxKXwn1mIiBCUmWReqQtBwa3G9x1stZu
4CJ1OWEDn76i6TcawW6guZHbmc+0UEWWPdvXnfEkDnWUB5+LP9O03JU0cS8JoVJNnJW1672VVUGG
Z2nmMsx6ODGNAs3MMBywOzc8mQN3KbD7Z2K0IpnfEvMkvqLoZT30gQUzDQGvg1Dlf012iYEUxKs0
QNebBCvEW4RgvYo5iMr5ZCyh/NlZ7GeBddB54nA1dzsxIuqiRjsNBoXMggxKmQbAmfcB+cY4cUoB
CwVzjaZPJF3EfjWfV7N4NcIkPjgzqEMHVgofcUT7jsnL3ozr+L7WrSIKGP9ElAwhOmH4kai92SUW
6nCeh7En+2JqhVseMWPBzhnj33qr/1f+pnettL0yeHqzNgOHS5ZTFMdUCFtC67O9ooyc/JGcdEAL
542Hk7Iz+L4U0/BI78Gcz/hmQGJrC7SNrlMgSJxYGpgRKCuusWPprbARje/+6zHs/Wiq9xti3XGb
amLPZONOZTJGuhzYOq5tJM/bc0mtP51gPpLc8PKCZlJ1Wrm8UXyyfWW1UidVqJzrtTvQ17K/umOA
vWE7iyZ76LRQhjz3F+u40iTVY0IFCz0JyFs89KGxgNe1CWSbhfzJE2w9WpVwMQFPxo803ukegMsi
JJGWnhEOJFO5o0TFExEDxSXzk9pBIhCWpDgoWuWFX/RWV790PqkJ0QXU0uNlCKyODw0RGtC05ZNP
iTbaaWbIVi6mt6z8IWbfhettnZl53YYtIHfdsfGAYmggIXGzSBD/n8Cdy8rUdoZ0qsR0qiTcCXcK
ATkC4Dl6QGQt+u55YEKjtMVKGe/IBxsuYwAz5v7AkeLQTQ0QMZEbZO6k+2SAaoKqFHr6nQWSwZ3f
BMhTiJ3grO3Zocn71lxi71yq8csDhLP3cCq02/QQf0A78+/76xXHv1AVuhaptGvzUVYqZ2LuBXFP
6iKsQL2n+4iceHDcYhq4YVRq/rSnRJ7VU2B/+XKzuQYAQ13rqyGqzhsQKx8I4MbVzjMr3YIyIoid
00N3s9dn6VKK97QHqBMkJU4X9ECaxqUWuxM6OUBuDQ1OmicY2T63rB+1Jo1d8//NLbloGKTbZCWE
pVITufqSsNxSwrkD5jxq9+I7K9vQDd4kkZP4jrlmzgmY7VLckWFegHgXMIEQ39YwXRFp8l14VC64
hx3YRTZnJfKRb4hWrhUQQkIic1NbwmVT4TxNckG4eps3+scK4s4MnITczJ6v36RAzzzPL/7zBFRD
peY30B/BW/CvAZYz25Fv8WgD+nFnfaLf215gUrCkHWwLZ4D2To5bu72ymMjIO5o1Ccn25ZYVluKj
tIdkFRUjxbYGyMAjQUijmXA7SHq/GrleN4eGeyl7UN50+6shq/jvTBE1t2sfmEBRIQyQZwn2phrf
PwEnCjZLK0pZi/ZhcoRrq1bRyaZzHLgNuTx0WJnMRBLaR9tiNDe8UJuNo+DWukfaglG4VBgjOZA+
yio04P4QMzNDKZHgri5c+V58s3FFlNWQyUb/zyBgSjQRE7C3yk+9ko+5krQ82OAKukCICpSxTWhe
Hfpf0zlbV+5co76jUmYeM3gcPzI42kJSWeIE+nNR+dnlz4hHCPkIJApzmf2SpjK0QBF/74xcb5B1
NDiOJDcPB4+QuIOGh97RgoLxPH4/la+rFfTplpiX1C9Qc0o57xugUp/KyKtdPQYKA4XZaNvqiQi3
zXgLFUHdnn7JWWxzVUL2ZnfIYn/Mwx69gclXKuLX7X65r04h7iEAM0oEzEYd2RqOgPlOst7y6te7
/XfQ9pqEGrAQg6FjPRoO88QtS4sNy0RNIHPHG++MJXdRDYU2mLrVuLUREr+ag9y7r9a04QzuRdYV
RbdbfeODVqnlzKN5/3Do60rOXaR16X9BgxAfVCE/mVOG4irwcUQ52GcIL/S10y0gvHLyq1V7irol
onYe5aPzvCnwHBEZI6OFxTU0B/VxYLlwKlun47gEdT1F/cIqlyqtGQWlwMAUONE2+tXmTwYmGaqC
a1Slx8Ix8fv2fRB6lx9lArlICtMnWxIfv445jtqb0KHc5gLAtsBym/oNuYkPMy/762GUD/qm39hD
ZFoDXZhJUNlsaQpDtL+NarY04xP+LuNwIqwrDL1zNXAWU6SYasXA3T2uTlVVSdpBO4xdfs/Q0gXH
rgJfn4PS5dgL0fh4t0nTuyIJ9gheNlI5+doOBVtwlRxUAWjvoOHzSQOW0fEXNaHYBEmOJ+F+5ope
Xd4X26/N9uQBh7Fedsy+aBxFsbofpqxt504eWxhOv2ErGBs+gp1k3Oi5VDtnliv1dL2kLV0ozyg2
9Ou2QOWqtcUyOTWjo+zG99yE+fRBQZZLMdjFynLqqWkojiX81zMUa7v/XY9QaRaeZbWLb1L1+Q1C
2qfgZnzidjDmZH4MMu1C4eCUXmeYzJfKQnA+f/Jn97+0flI9zxqrFsBv3C4xVsAaT7fttfQ17T6k
/aenrgVYwW36Sz0Z79TC9nwOjgsF//YwrJm8p8ki2J/4GeLt0MonmYtAjcKgwEJT15PUcSKWopyO
DKarsgZmqvufcg63Eao2qCYODvM9vCLdheg9w2nvYdXUDXi9m7KO6URW7DVMK8uUAWgypRny4BKo
l9UpGBQ1RC2hhAvJwTJR0J2xYU8hIHV5o6RCUHd+MZHHv6qsZjZSPtxM3KlGJDSBjagaB66LRwPo
0mmBZXG+iwObS0JjV+lTq0yZhGzG5Y7bGy5iitIVTRGTH/rTYIjYvMer4xWIQ1G59QQ5NvX6fP8b
3RsxpeZ37sCr0MkzX3q/5Ryq6CqhU7rhzYfq4lUuszxIcWgAcHjXpWqhF06Wd9RXtrfxsHbzawBu
XdFL7j8tquQtgnN0GjSYv5WmXDpPaeDVj7ujs56kvRjKSNNaqlIxY00ah65gBFZufKbisCg/qYXn
vKAUbYdP9EYO45TxGOomrqdd5IYMRhLqKDumsL0+CZ7oT7dlNL8/KIvDckmJNPwYeCxPgTO7SnfH
4xJ7d2CatLWE8/Xgza+vzwFdoIEiHPPkXaGqt5O/X8WAwzzDdfsUXYAF98z0gXzDvKS8TptlxIvn
XxKiMpwF3WTeAqs/qJUT7lTTXAYX7sC/1+XtMNH57FJbF5u/KUA/3dt40pl6uHKrenXPnbH/g2bP
qiqNl1dSBRxTRbNFAcjo9XcJ7TQ5IbvGjzBAUbhXF/vUQAND5tSNbtb4jhcoPp72HBZtoDmCes4L
shw7n8V89CoHxY7cTmAPLQnh9e7vDYEQS/izq0qdhSyM9ZpBhUTcopVuB/AYosPxRFikCK9sQ9Fs
EVOOCdUcmnNAyFpYXtaGaZsKE2qBM8bxg1dCjZLeiX8LpqFwd/sBrpSvq68oD+T/G1rrtDGfRtTl
4QcXjdjyNPAQb27Zi3Bzxn2FbG0gy7QfkF0/UpU8KBIz9V8Zeocp5tyWvu5TAEPZ0XBt+j3BXmsa
ghNnFMtqrjkTxv2g8CKpUe4ycrXZ39ak3MkL72HnVTMCo2lvIQ/LxOsxu1MNkrhj1rb3l9BAb8Ah
oAjCdpTigpPBQJEwq/vqT8CdcOIoVTaah1LIp+m4Wc4IpoEafa9Vdlb0tki3n6DxDwcfZluB8HB2
/+n//DbuHWBLQk6v5tex41s0OB9bOENqyvbwp7YI3tN2LkANRrcFEzoxxl4cnV45sNkpOL1yEnfb
sLzBlJnUY10DHo4RnW/S7f7JoOflSVHB0ecDiZo/IJVJWo1DR753tALVuao73WAQFQ24QvqCn7Fk
QiuMTQq04e4irWg43YY44Yb5WOrtmDvzokPX9RMfUHzL5xO9cx5UF+yEnL6AelvovhpkKtzGulJT
EXoKDhBgT2WPSQpZO3WpyNMAx43GA0SWLc2HGlTPdR3nRKNh3wAMkwtkZnXdSI0uVY58istniQQA
QbSybV10B+Ptgye773H7E9YPlpBZXyJ/NOGaet2OQWYGkyj8FxMcygGdcEx4LM9bcD3HpLmNUOR+
A/bFkudQuRrxiy/HWc81PEmauIxARHk7asbierPzBvydKC4TB9wWhx9SK3XcNc/fljGr5InDs364
fJw0uwuV9uCZ6nP645DwFJVbV9vZAzkDIH8cXhxkVSHH0xoxCPhNcSt8HIVOT5QIfa21xXThWTci
442ufDioq5OGyIOJFwHOiXx9MsXdWrJIrj/Y9EMFRw7hW7LqbNvfteymiSbY4k+CXl4PMFwmMEWP
UCVV0/jKFWEuVl1eDUcq1zOs0nljVjEBRZnKRccPYJkpJzdYp6hYN0eH7W+uSqpAxOTm3EPOy1Dd
9Oy821TmTviHZ+uQ6s2ikCBNlZaMP4FnyRUg1COx3LEsTPmvzCpfi/aDGBEDfElm4G9zIUfrZ3If
RH5yYm/uoeHQhAZZL8/6HreRutDgtvEIpKe2YARpDs1xYLrg145mHQrVua8vTcypLvlvHz/NsGaQ
1pFgkrx9ksQ8FEd3fuNHQs8UtIDnrHH2B9d7422U9Njcy9rku/TpCg6vODC/Dn3zzTCA1uvsYUdv
eeyD61+TF7EObecsDQLMO94bxbhyRS3nCAg4kPoCoaah4EpsKe/rrLXExpC40hCH4V6u1v7V/W2w
7hicvAid/lmXQ8lKXBgI2BynW9in9ozRl4VPd/VZLyrn2Nv1oSKeut9OqwvZtVXDTErmVBf48UhV
zaeN6sRYeOKB2Jfj//GloGh3NmLncH4gI9RJLm3MwENnsz8EuMNSVGoGsiJrrxGqrUyy7EtC70nT
WB7LRNnhw2aExO4FSnbaoAPI0uXK7HKE4Dx71gzZeA1kF/KoQpsJKoANEqP97JCBhMX2pJYsxXh6
/xPTjZChmVeGuU9AdMkTBi9Wk4WeDFiPz+V6M6wymY3/YWJmepYlPbYNs7cvwldpuO6+GB2cjcPP
HYIxdz508hBNa+9VA7MpGYCjwxX3BFVUUygtFRG20A3TI6NAuNVaT6KJLIChlOS4PtUIqc4lmUjb
vsY9McYm33yaq6BNeQCR3vz4naSAAZ4jRYaydwoacj3jXGOQsDXnjCLMjvYPj0tOgMYE7yQUj+/P
A2YqmHJ6YNk5LKAzgDFQ5so/KSUcIwo1/NG7UEysYxDE6QUncueAKQ8/r9HOEBaqXqMA4WTWLxM8
VrWbDyRs0wtqMLx73vZwI5wDaZklIneuYNQQZO+kOLPTnaCSAThmjuefY0uE8rro/k9mMKBVS5II
izbdcApkPBIbNWf0J5q1wvPrk4woIuLiF3sljQTF8UvisCZgM6w0ZTAmwKWTOvZ7DneMXh8mguTF
k036a07g2YviCoaz3vqnqX0eIkKswRaFzTuZtD/W9OUrXE7LvZhC6PYPIhUN2HF0mg5ogBVNFgVQ
DikorYeJkB/UkRyipkoB2BzRRM61SWyoEttDtmwNj3zFJzZ1n5UMNt4VvjouCT4eWunqSwo2x/u3
9gPF2tZTzAQFWdERxyo1XGg+Yes8043/irf1Z3MyQzfURItwf3ltDznXbNx3ic0cBclDpJ3OiLQ9
QjnH1PGqpQTbXI+BroPDCEDe57pCSSBIP0rf8g86D3RTCohknD+PTSj2UWGLYvcQU+AgRDjqO3Ub
/xikAMg46eoAGGWIELiHDj9KhLczb0ZUWu3UYKl/nV7DeSGmcXt8LcUHkZrncRA9b/c1MEEM6V1I
r1CpcH8AW/Rk0ZSLunULhEvFAUkbImhrdvk9p7Mkz00hBwwf9W8v1ZZcf7NPMmaPRud0xSV1luTb
6oiWK7PAGQ1dORhdP9oaTIkUuJ5dwHTtr7UZu9HXrnfSMq3zZ98O3xKTSxPk2MZpwW852TuZ5RuW
+znURe5HpRRrP426Ih43jA3+fk8aoSNvae5GrGDUFLqi8DBUz7Mlh/5Gu8EO/wnewa2koh7jRzSo
6QnGk4X79l2eL9Ons5FQirc1LtoVcLlGbDMA5dhuOFARO/T+gdbGEqOt7wwmdA0OUhvtHmAvW1qT
+Lw3pdfByRNOgEvVM9PKHQ0G6ETwpVDmIaHG8VS616J3e+Om2qhkXFgh8cl6P15M1WKeI9ennmsa
QJrLiTFblLYi2RuzL4lQDMwRue+YEZqR9ce6j6ODie9ixWdN4EbZgiScMVzaT35+/nnDGRBSWOVn
AAmZlWALC3e/8hN904u9BDxh1IeX80y6vhXOo38HqVyl/r82ZuUw36y58n5PH0RDGP5O2UN9tLgl
Np5L2teE/fNNLO8v2cwOvaHRfmegjSfA/PYP+3A02HTDwBJBDaRujGtE5ndGKjhCEd+j+ET2AYB3
bs9KB3RVliegdGd6td9drkqBjt5qpy4PEhJIkcip2HqKOklv1Q2sD3gvNj4ETdiIZtAeQlBlBzhR
AM58dusTGqEO1Y1XXG8179xw8A1i5y8eoyUIYwl2ZaF36NMCDpANVnp9DG39V0RDd7eS52zwm00B
NrhpJDsIdozxWUhCQcynEmQDgf2B0KNVltrl4ipIca4H5t18PrTg/OSmF+8ERnW5RBWENfXCqJKe
y5CB47ykgTtwEMJidGiv8LGW32YUyixyUtdit1zefzqjxD24P1VOL2VzwkDvpkZt8qAVt0KnRs8z
xA8jelqx2hp8RrcZ0M8nLMuTx8Kd4feIel2WKL7jeqpZh5el8uT4Zd/QuSrSWD9GdwlSu/q6Tnni
XpdKIHvM2wZ8wQpYnFpA7HDeP8oMTDiv/1kNC22HSe2SuPCwhGN0uz+Bi/2YdZNAlxsENeyil6AJ
FHRe285KtRB6KEOucqv2Sx4Na4cg3kBgqnSdWJEUDTdu75KrcQXK1ogjaaLwXtMHNJ+0vgWn1D3P
lGBYR3/ZFeVoCFow04Kk5ugIG8jc4uXjuj57d5gCzdq+o1GgcSyhV2jVqzsaZdb7uLVfqxGW0+s/
/w4BO+RKpHj4szSU+eQtGHE2b+Vwn9hIgl8QW0387univK6xDVIGnHHQBEhH1UeZvPvP3iCsQ5cW
fPtHV/cOdHIrgOH/FYTxFu3HAzt+vYxrGiRR89cQisQ6/a0kJN09c8iky2BV5Lu7SORhqasGAJ84
qNa1r5MsNz8jtOxzT8SJ5gNKI2Ybt3y/IkArI3BttHVRueJmZ28EUOJNftZQbB0jIk8MUE/fXbmb
dDKeOCvzFCT/TwyzwQtfZVD70MCQoHEJyCmZ8uRHc9rS3dTqvW0F0J3DOFWtzapjcyPZlUIHL831
Y8pXH4G5tTBjBCzhy1RhXeydUFfSOX8taNP1qltD/rqgUtXFkxNNH+ABxtAanAehnwveiC7HEEPA
vwXZhc1VFyVJdtFLrKVBlTXCwCFVB7WlQxczADBPO1SE/KSiWYkut7fbv1UMXpvD4WeJpfXKgUps
gahfopSntJRLecJgjOsE5br7UF0fFIBAqWF37ITFvhQatWDU3k9PnnI60W30Jjjz/kDItzipuKK+
NiSlC+cs7tMX1sNyDemMdZ9etQEF3EMVkrrn9a9Di7/RvEqsqJ71G3C/XsAz9Ts83gOaTPucbnZx
IXVBkuSgZk6D84O9GJDQE7d3Zt9uNljE0Lx0t8p0LmEc6tLqe/vgAJJVDkm2dxBv1+ps4LBZse8o
Va+45kug1dj6Dge0cSbolEgWt7MixtLDBmAYEi0NJVEZ3Y96snxgyNOTLar/CWboZBjAFaQ+bn5z
u7+WoBrbcx7yjXK0QJy8ih4xl6gnD0ttEI8k3LJCvM//Un69th1a24BBZZafFscS1wNdIK1ruX+m
Rq844h26nbN3pp+tYGamsi68vZk0+T7LO4BaRoD9Art0hWHCVeBVHJ3yYE4DJw5kriHdv1X0IBF1
VzXGFG0Za2mZFqETuSXXccszYAbwbGgKk4EiT552QaHvlcX7H5sHm8rq21htP3DS8pmAqie+Bke4
Wa5zKfU+2Shw+HubSCoeWDGJC0onWyKH8wIQp5gDwpgVoe0jQtXFzQF1hrPz0w8ppm/86cdHlLyC
1XSKaQqoCDvmFDWraiWYCd4x8eov+Oin+xBq/CgwCJX3iannPpQLvLmGuAnhaGDuAJcBO4Je3yh5
wNl7NerWkWolGH30qIPUC18dOk90GPOgUMQhx3cZpSgu1lCkvB8leuQVkyIfqVD40Lbi62u/RNFS
KJ+nJCGqC3fGlxhLKKueK9DNpa+0xycILVBWOqusOrCIpvrGsnguC5IXpEQu3z1EpqLjfL7Nfblu
BU+F4CTOSYK5y0WWVmQmVR/mSEX+hyCzEGLT6v16rLise4ApCXoouHUcYrUPMpLnReTNUJ8YuwgU
u+NVXuaPa9XLNIvElViK4qoKuW51KOedtDr7XZKBnbNroozKwX8NfVotVqHO/c4WbrdQJhFDTFa5
qxVC4Gzeg43lnXhjDtdnYfCJM6VSvrkglUflRnZCCKGz6AKbGR9/WhvlJU/tyJih98wht7o1Q59e
qlqG2EmgQvUfOLjulZcj+6bLoGMvfJSTDWdaK1PuFvdZLXeeWyC93eIsmRk25F/gQFRw8g/tNLoF
I/xvSEE6Zyvt6oylQa2w7xnnzUOxdcmFwocLer/cPcb6FB+3gLz8b8OzL/tiaMfhQQ6FpGxew02j
wc0UhdVQOUOy/N0sjNnNkyEoy6HTEUl39GLTfyaFg9dmoPr/cIf1rr1Vl7pph7jiJ9qkDkvmfCis
IqZfOtbSNFwQRcXkiASLqQ1Md7QSBTlNfng29la9fEPPkX/uCpA+AkjuP1p4PJ/ntjO93YJgZtRf
bZNO+9O/jqmto8MfxAhzPNWYZ5SvdLc5BjDIis0UC/vtW1xrmPcHqcbXSU+Fa+xAkYTZsyfYrhUe
nPABmxf64hZjVWijXzMjbo/R1+vIiXvC+B3j50KWS8uIQa9ddDWQ3H/IC7B3CPglLx7D+Y3EBCr7
dRW+m+4fMxQW1iOmWXtmDPfYIVxpRsPo6t7spNbwJZNIqFNKJTOMrH3bK9ky3EIyb43UEFtdHZsH
CkRvrbrInIXVmnBGFzcw5JYO4aDjLI1UwZmG769FBOK6ZnwkxSWe7QvdCqLYuhE+Wk9E1tG3c5HZ
hyGiDhdRheYEcIYKUWoRB7a1FGc7t1INTbqXsT8QWRIOJgY5Fc2Z99/NjXwFI47lHV0eoSQ7Va2m
bwudiPX6/PkHN/9fcOQpXWJOhVUM8yBVmrv+T2KzWKskYB0Xy9R1Uq7EpCCLyKfddcAV8zFqQend
Ba7izFc0tnPFo1t2SFa/zfeVBpSbX7spjgOCE+74TbO11ozbXTZfRQlWPg++omHxQ6hZJGyfMl9V
dxpefEb5glx9IsHR6Rsx0mVXn0nUTpwBQOkvsgDkSH0ehHH0PG/PNi2nBL84FdhqLjJXx2X5SWnq
oLErihs5uirJ0fU7Mpcq3Q4j2PlOuHS5BD+/eFcayOQkDtJK7/WknQpXxB/X+OKyoj0ftqZmhgyy
3FxFj+Rx+32YsD716fdIryR7ZcUUrnL9Z+b0J71FlHsuvGi7zKlnb/kvrtg0HbXB+MOgbxjmQ6X0
O2p/so6p6PFCSLgAVmPB8Wpuch1w76ZAvkQZtp8PNIAhanZ0iy7d9zM3HJJEBcxUIsLDYVQVvUZk
naxbjV6bBjoB4k6PQb3LieO1lYquR/kIGUieixRA9elGhkIt06/cmks5SuvHdrnRVPigqW3dUoxM
qOTa1NdDhF8RPU1wPV2tzwb7Hmy8k24/q70ZXzaqf1n5JKc8JSpxFzDIuovokWkIrdXz/qfjfq1t
0f1bdsHQfh/oTvoJEYpScdwGPKT7il40uHXugY2b4yEMYUA8RMhW9DCTxIh6nWOBiiWqae0Thr51
KBvV0+QvqwbhC7zysoXXmV39CmGoXu0Z7QyHcnzSgqn7o4GnlfPxChSJuypgZO4GVDlBdmN1/Tar
/hLcatrkequl5YWiKhalhlSKW9e47hqfH+ON1PbvFPfgHxB8V7JD7onRwgu4uWLsKoOCKgfirDh3
DSLP2xmd6y8jG83WXfNRpJ/YDeVChdIif0uc3cM0UxM0wQ2ftK95hI9W9LLZuR9OsimpZNl5vlSQ
l1SBS2Hne224eT8E9mrsZHEOHPrws8jET6XNln6sZLC841/MaUJ5xP+my3DxKKBiEOT8LS5K/2iO
jMSFxy8kpPaLUVHjMCEAk0Jp2uogeqIJIYGFJ+s0Y5WL9JIKPvBPlGyMskcRSI0ITiuUOG/BlhY2
sk5vUn1w9BtswCIRZbzfVRj5R3clHmNBuy4d4wPNQoM6QWMsLMSJgEMeqUem41yLBkyUwDj2YCUi
53QuqgakkmYtz+YlyO7aTiOhyhDthNVeCl2m43B6BBr0PZsKjAXMIUuxzl4AjdpEC5EtLME9/9PP
kFyUWet2HhwZB0wvoeIRtAKMhHJ8ML8m5dbvz3W9WCkj56ks5q8sQAs9vJLZgMV0H6NBKGqFBeTA
6fwDapboRd6Es0kGlH8Wmn2AjSwu+FW1Tu4Ew8Gj8lilSuvNogULUD0UUMz0I70egJhbdenMV25r
onmxRwzs3d0vcnljQNWzT5+FOwf+XiojyBIpUmOex6jwCbo496+lyk0L/unRPl7D6juauMngqAtW
mo4TiGUh1O7Z5kYykOOkSgNbXe8spcgNA8xhHDC6NT1FvhNbRohJJOuiw7l3lX+GYWkxu+YuUQmG
f/uwy8fdbzagqIw8GPudob4Qpx5axDdJKGt7Bn/IDlDC5ah9NMMqu9KjpQXutSgMx8CkhFxQGcU9
cElBWTbSDJVknaGcUThsw7UYlFEV/BvmQtneHKddTXwXV6c85C5g0ht4mwFB/AVIJgbiJwWGgErF
NgWcsrLs1uWdMT0AskIpTLDnze21W/1o240P9ChbA0QSHpwxFoOZ0Gi7NP/pfmL1jKfdUyFp+Ima
Ej5mIPAVUrkQd+zU6+sWEi2dlBH+sBttr/iJWh3uHBgk7EVz6LMm0f9C/TOkF2LANruxC7b3qGo5
Ce6U/K06P31GPD6H3oH0F7qx4BbUnnqdrshlxg5scnGCL3qxgYBYqVLBZFCRMh7GwtPpoWeVTQjM
0p80+PospZkoSbUDQm5sgisDN7hXph1u5DHaMTPDgtk5LZvkqozBVNEEmlXaC27hflwOBo4Wm0Pt
fe4469KOaHa4YRs9ap9HhstZ64QWMFt2sh7vHmL5YxlB17//b4jwq6sKRjC5b732bicuoKPstK6x
rKuXUIiWCZ7kjay0NCoYQtIjYwwukI6oA4MaRLOVAl2y+EgKTaFL6H+G1r1vNdJy0KpYjVz6zA/L
YdD9V7+akH8UZGfZ++i/fjtVzJ3pH64AUwr168aQcSEn4gGNumPJSgFJpxcuYC//zYIhqgaG5/BL
PzBoeN/5Wo/Mnn5MFECJpme3TK/TqZQkSTc2+GhSGtLvnhArUujuXD/it28ew5SZ/CLCoTDBG1UH
RBC+2sKyvkaaHiJULfqZ/cP8oF8J6ihOzc7BfRybIncGPB0h21wisvRaaH8c8sfUyguLthBoOhZi
0oz2djQS6wjvn8jl8dqxu/w32xWBS71g8ZHa+R6DuQ4FW1uU853BNfi2m5fGccMWg10VAQOMSVQy
V8nIsP8gvnXWeCowEz0Mnj/WTzG4helXwAoxN0lT3TJPcaIsG+9xITCHJ6r9z9xT3snWhp4jBvS+
7B/Nzddb0JKJw4av6z42lePTJ21vzuSCHi4gJv31plnosu3K60pQbya6oMdsr20KAI3jH64kvoS5
cQGeOP4qUlGSRl1NugFbzYUoeq8WwhlDv7VdzQjC6Jijy/U9v/tz2TYy0JJmXvmbrtpmSUuCXKF7
M0k4oYFW8PToWbu/Uc1oKB+K2cSycCQ3urEeiHr6in/+pEFye7kNbd1Jwp50G4RNeVK3ptaFDoV3
+CQxadb+cLtcoNM4vuEngnqYszc9CNchtFyLg7A44rMyK7t2/dnSjUup3TWKG+dhf8gAkzZwycP7
cQXq9KVEf/DyrwIYAnHGa69e6VHsqS9hnAk6kqlfxMurPT+oGICl2qkBsHQG7U8fBZPl6YqpRI5l
pROl7bSNcLvWq238Y2+1buT1UUsXbGJHEKWCcBm/yW1/yPm0TlAfPwvYCHST2Y2WTy3itENDtng/
/4fzWOuiEKMI9xJ/nrMubI2IUUFS06I3fSbLAxafJirtmfxxYvXEVnKk1NRKsAkhc04VbwVfWVs4
L5j3udgbDPgs3xsbg43t7GIqHUcGbK+oc5b1PM5AGDaYPseSCfbpvACkTxy4bj8AJUImrt3qfqp+
c/HM7+sg2/fLn42y4XHc4vWvEXlwXsdcOvbTbY6PcVzOnr7/vs8tH18vTf18QH84j1G6zZNR2bn3
eW+TaP1x9hyNzXvS7+A36qlAHRY89MDhDPnGj0aO6ke/FsrQu/FlPANkfAlwmQ7FQnoekevEKJ5b
IbXB5tMVjZvAaM0lM+74nMRnPgiunlI0huplU7puxsSegelvhlCx2t6t+8WM0/xpbu/o1TFHPsXb
vpGM83KC38fv6YAaJGYZOUxlkEk+yqNE0evZuexwVupSaBPU9+L2+tUAIi1glQQslCb4RApNLJGK
oljOWHzUhGTimFyr48mJfC1/UXHu0/YVkIUAkvakLY1HaGVEza6oWsbP0B18bvLLQ4Ro8dBtkuii
Q8r0P3cUkpDWY5AgGrjHBwV+oGFYGZBb64LeV92FKSRmvhlbng3Z5nIeTPokKzcp45quEWFhw9DT
lFEKQhNu0s/abdEndvh1id0W+IPA2HMhwUeOBmXKsEq0jeXoGUd0aRuAxKgi3AoBY0myCLcTkVHe
YHYJ1bVJsLMgwGw419rkhUfpMIPH+EnPaINm5mHnKewxMKUBx93y0BHZkHUeOeKIWy11mevmsuvg
CSP91OFrN7I0AL3/aeF876UYwnICUPOLsnUrQxuLWj5n/ZcJqlH1mMEJL0DjySIwJEFhcm0uhiJK
d5YxGPF0GdPlZX4/euzTvw3vx+3YssgnYtzwhqjbZl/GYfJHHrKMtg+0ACXjDDhFYlIojU5g+xGy
5AUIhpTIYPTCrBtBvR5OfkGAyL6sWV9CoZ6aafDXQa+r5PXa4IgpRfVDi30H5hqhHNeoLrXSjTEJ
ichWR6CfWXjRARrJgV6VhnmqIPgrNfowC7thUFAXHBHndkWSFHvj05J2qGAEdetEB9zUu9u65IhI
haKBd7kzOiYEIRkZlK+mhCsy0hhL0h9HLvf+iuV5FHbyI8aV4vPUwq6VmmuPF+IYeosnAyzHFYcU
R4G9jIsM8fe4cZ+MRsokHqxvFjZ/LvIrOU+J2n+pTCL0ouSe1BMeiLRuX11SoySF4dNuBFotVxcb
0LrCcFJmv/vEl2qWWOCocTZ9D1bn7vwAaEdvQRO3dyE8BcBZg9bCErtamosNDfgPLDPJOuC8sxEh
ROg0tzDL1cOvRvJNr/1A0A0VVaF2hv9t7CjD3o2+Ff4DzERttfPAEV0zEe+z6lzfylI/nXYOsZyK
mTALNA+spJcMuMBhw5GNE4Xu54y3GwkvpbSpOqHyvYoF2Rku7gblHxaH1RTVdG22ns3dsE9nmSPG
dUVOJln08xgnAzVl1X7B2rOJvF2Rvo3l0Nj4H5g8kEukYWlu7OfV5z7X1oiOEjo5KfClh+z4BQDW
fDnGtpF1IXszAyR6uMp1hVo8PNZcg5aAImr2mY/oIEA8nGL1NKfoMfUPK0J1+KARAm3c4ER48kes
LoVyAngGEhQMievssoywBxuYLnx6BgD6h/KCDvgBlW9yl0mS133TEeEhqsp/w5V6BuDy2KkjqUFs
SJwpv1dxKbEVglkYrMzdBisIAMcbPQrKEHZbfvUjA7eLVkvDiHRuxRMKgNcsnWn8XplNzwAMJ3RV
y5iE3kj1/WwtDnvKyZQxPpAxU0p6PhwP0oRhr1G6klHmyPmicdXOfJLR1KBqEp2qbCB+dnlKni5a
T31Nygdavnhw1048DgWmSPz6+JsFMXzimYO7bhkttvjz+Tr6c2d/0d/yPLtMuxOrnkb+LCWcudxf
eHJu3O3ofUz1b2ftTaRvNjLDNonIN5RHyrPfCUoynumQZ5DpX459Jj0x6vVPmoP0/RzKDt6cHTnj
C0jIb27raxo+HrQVZZG+vsM3TZe6TZozJi5a/TiQOrix3qJH65+oWxSdmG40lLPzyTX4NErMB36R
kZdy/y44lp0YcvrIboske0wVg2wt/wN6qRod2tgD6IOtd61pXSlbYScTjO38XlTqVXKWnD0v0OsH
XcmbbhpV3cpuzI55E7cYM6Z5fFCC0/1UTrvqdk1Wv4gDKlL0S9AGAmCeVpgr+/UP7XhYkWuIdc+Q
mOqOZHfAwQgEYqCcE+6CQUZ8JgSkfaXxjCMwYGFEQK21KZW7KcrjN34AjtMLAQM5rZNyUyrrvvKm
v8PfZ1k5M0mvU5tPKxQJni5Roae3axx2EJ0HdZphKux9tXDCU6pJ3+BkqwNOQTQj32cY8dsQN8bW
pcOAgQsEXU44HWnnbAbOZe6sMZDXWg9ytdVdtOw+CAczkYCGJfenXQE7ejPOvH8XNUe4IP4nqCfY
xTYqItjPRDu7XQNlc6q6Cgn4U4E5vVijn8qklpG8o+hIIKumh4yJk4VdP3P+mUIC0uqBHEMXpSa7
lDUEYfxZ6KqIEykI9RuWek5wiQ8DSfbVfCH3dbLw7M7B2sm2HabA/cIrcWO7dFYnEA1cC+EVE4mc
Ub/EdDoyEyCAp40/WRrkGSme2a8wvoLCGmtTtsFajbT8aTNKhZFBOhJdCMuRjDOb0VY4b5wZef+j
1jZdxaRLkY0dHM4lC/DNDAc1Use2IrMHnMSHgr/mKw7PG47rZYcxtq+7mxwqPPP4E1z53seWxMsg
3+9tYsCmWj3k/finNio+3kzrGOz0vCsP9BvVy7zBkYLYiARug/x+2cxxzzcoB3MSFSlnAzbOLJfY
KYUn2w1LBy6Kn5BB62sDyEwp4ggK2yC77Vp0YhiYY90c1r+840fJQcbETc63e4Sdf7D/AXfyOEi9
XL4fcXwCQ8x+0O5+wcyNWd9rHaVwkT0wDaicCF5vKOyqh7ChC+C8pQHthi6dRcgvrezQb3frL8Tp
z3NqefsDBCB+enzcisKW5Lcw2LZ5lExTv6seZ3cIaPYq+FwzaSdP8ZjE6o+cgwSdlNJK7hR0WJ87
49hMLwyZwj1Q1JYm8igYY9C6IojghbbUT1t4btopjBrSdNzt/5v6Bg5soPCxOXPEH60MWT6a7wRv
QvKA7LwggeITS2jPe8apzOSAmGfuH6Wz+Ei/Sd9PKqLBILRZIBUxqEjVYikPpzwhuUiVO5n+I+2j
knaL/DMP5kIueb042+mESieo9QI6B2fM/vw9vLPFx6vez7lKh1xAaKag47N68ezQRBjIMWu0SmNs
EbFgIzT3mFLCAygtZ1GOlxNQjZJZRWffY3CDyafqBqnQyxz7SOu14bfcg7T8iYHMLiKM6KNUYvkn
08QGFbfsEia4By+QnQ3OwpN67nhbTrszUzTJcZ2vodMlX92x4/mlRHpoFHdGoBuJMZYFxK3meqJF
mpiN7vXewd2Ib3aTCur2bCZEet5aGhG8S+78ZQ87uV7n7kA7ikI++vS+gTqSehURHPSmA5e/2w4R
cZDpSfeUwNAjJURCz+kbc12gUuNam9qXF8GeLyU8Ux0SW0X2QJ61106WAStgjinDpgWnvxSgcCGc
oeOwUZt2CKF/ZygcqM4Fw/RC3hPw/uoUmGMkxvrxzrviDr/puumEXQ/9MB0ItBG9JASG1C9rtcNZ
K8lvELNu3kJ2bTL8qd5knf+HTlGCZP6reVrrtgMhvTxCTyirq2diaWo5AU4TkTtk3Gzb29CiAT86
pke9P8Ocw3WIEllX4knSRj4hAUZ79MDNeYGeGM+BJnPKvZ+g8GRlSbjn1SKSG/Z63BYcCAZqtFct
vgytv4nEICHHVIN4A26ZGho2iAU7kVR5SyA6tOUn5+GNP3Nn6PNPdovrgFSJsR7BKFN3Yt/OZ9BX
6RW86oy6PAf3m2T8AC4uh3DiwGMKSwTzxsM9b0TPxZZP6ZwWW1hDwppTb/ysyGYrb4v36qW5GkiX
E65M/ic9Dz0RFyzYvCMvgn6BiR6YA0LrK8xzFbO8756VDUVnvjvGd6J49s2ZE1KHgrZueAC0cCGp
naD9l+2GdJkxSh4wErUrbXMJVs4WHneWAn3cxD64ZngPpEHs1pA3ccyy0nP7sXa4tqWre4wqzgKf
/6oBYp+ADO/6aKqdp7bD8gm7wqmDd5v/QFNHO7Tcs7HNC2K1wByrUbey2QEaupwJhAkRY2LpMnyB
4TZ1TJEtAtBhZaJHRTmgPoVasSn3tYK4QI7Wjx82GSwWJPiXMHbMQsrZjzADEhH9t74F7l2GN8Sp
Z47gNSJ31EZL7Pl5g8wrav+i4lXlP4rzbpolx2034+9hwmwsIQbzxTb5Mca5U4xrwjhxKEoiz3W2
AbmJG6bGIo5wmJPAwCTFjl9wSKcMLEh0nps2xRGqjKa3CrDcy34yT0yeW+I4UOCu87bvTh+3IFRW
ZAi/hyqeWTZ2f1wQUAtm8t5VxR84Ehah7IbuRZ0O3gSN1/KoftC2TD5v5o/cUDKf6vYKmfu5pQTl
i3dLBVRI4MrvaQM0nLGNbwsKEL7oYAZ1QwZjgBGZGJrRaizVdeThBjk3iFUQXZfSgW4x4Ke60vSK
kIFJ75wdqVhMv7zztieQ7GN50BtPWpfob7MtigoLrV1la/Mpi8/d+jLyhyIgnUFYiTEyuDAAVokO
//ArL3n664ZbwlXVoG0d22vjmiD4AwfhiajzLnLLumjNTJ3LNpv7LmX5n1tSJHsIdt9Rfjnzd+gr
IczH/vW6VuT5ASFPRiOEm9S3ukgXOnHeOSswgkgQyDjA6QuHp/Akxf7Pe45G05PPrA3xjqWxxmoz
pmMHXRUflB2Ilx3X+ueadg938RjAhi4TA1fLfECx4lrf4tTrOdn/7j2LfKYQoTy7OPLCmbaa/iw0
pIxbWWGi5RWV9aTaDd5eiwHUXzSUVNhnQ5nhE4x/CIF+GT2bFbITEXsytVlzC0wrXP+GqCkuV4p2
+Jm8TZTpy0mMg9PGT7TO+valFPNPy0nT4BshdrT9fmdmOx3pX7bjvIFEvqcZY23BIZCEbSCh5ceV
UH12REX2M0PCCoUV8+wizXOzux9EQGoUrXFqUDMd0TTWSWjxENOR04yfKKiurRhW4V7dXOICGKe3
6cI3/6k7A9/9iBRxeAY84BgSQj4Vli1uTiFQ0W7v6Wij5TMuDrqE47jgvgEzwXWG7rB5zWNZJjyK
0zZvMSxyx86x5V/rnJkeevLuLSitGJ01nKAG6DndXIigGbH9U2vbrNKN1WBcgCJIxZag15QV7owf
9tbi3WcEzf16Av57AHmFLpFMQQNeFnq3l+Kix8gRc+34v1OOf+3h5xMO5lP/fuS2znZEoRbNohDF
gsErJg9BMjI14tT4scPFSRdOFtjia3mxVkqHGxTYrlLUCZNQ9rQd6NlyQQ+qFGyP3PLKu91zTVlD
CeqxaocZgJs1aHo5zyIEUccfp239cXi5gP/hqKEVUVrUe9Lor49NlvTlhemYpTcGOgWatXVEsAFK
mjjBWvcq2lp4bZ/FyB8jPa7IwRQaNThDtP8Ivt4l+fUS7e9PTss9tGYsiZF49kFUlbs/AOAQq24B
ROfiWlL2NJNPRsm1htR5V2XOgmzR2htw6vqNJaM7TPf6oA+HbVx8PccgGZYigXdYSS/fPtCOej9s
8hZCi5LPOc8yMTnV6iy4zbqdoA9m/wkV/0jmZ0eLlRYkfP9qwCjUAq5EaS/b13aMdRIZJsCmBDw4
v6272ROw8Kbqkwjru8UEc71tEQJUnTg8chp0Hmsyjtgp0f2uWQytNhQ2fU3kcvqmE4JqvT0BJT17
d0uVqbyidZU019CfR04quz5wu8JWcduvwt4W0z91UEu4/azmm3ejrUuqbuemudMDTtBfYslljH10
AJ///ulO/7w0Lb3iN6nRzZhUQVU578QVa0yYjO/K0SkMr0ltMulE/0iGwiNr6RAx9f3tiUO8DH8Z
HZXHiZUgWCh1UL0wSPyfA1efyPeZnZ8n+jOGcd/Z4HkdWtukEp5jBYyOa0++kwWjGEPYsXxnt/pQ
JdkLbvGBaSBERnNsVo1br1bXvVk1yr6e3pX/VmommYhEZA15+PaxlddQAVgK5tQsQ5nYWR4syJ+a
orWcgzh/mqlLkmOKPy1125prpEtA8nl9w57i8ZD7UE5BJSCVnfhWhB7bpqP/JVCd5IiaZmgfr9yR
Y1vnPjN0E1FuYKyKA+OMTNKvZPdP6qNil/4FPILCIq4Xg1QpUfugZl6L/wy4tAbggZJEGdidFVlJ
VgraqQ2369uxs90dZRVlvXfkXxI0bly89xvF3/y6ectYjDDVVDS/uuJfcSpuAMyp9tzXn3Bhrh3n
1Yv3zh2kU/mYtHlmFwvm4w9KQEsm2OsXsHB3YPEPmiI0UFxKq9DKyVQpmecipCbxYCAZrIiZ7K2m
oZEM9lRUpWjc6Z/qrBclo9pFMBoKB83OtohsLlBBQ9Jj7SKen8hQwIrNehvLmsAtrPFBrcmPusKD
A/voGIr5V512YMlGyB1AXsajncRCBkhb1AB8IUjYqLEiWGe1wswxbMRMFvJb90VFq4Z4MekeYUu6
4o7VymE7z5Jg+CfS2gwVYGHisYvAb+wOcQsnesANYPaHw7IYpV6kNnFd+4tniSAMQkfg4dKNVKuT
SAh6gygTvweOCXyEf0auB+d0Tvd/+oYwvdkXeg9UrY4Yry3KfpSCuwVGkELVB7qYj5yLccyxWinF
K4xOgfEV6KNyhy+V5aEp6Y0sGrfSmLbJj04YVL24DqOXeQRuwjwp77kF9XChmuaMKMKmG9aWzgy/
VZswQUrsH8FlnHu+zzcPyk7fIupaIox7Fw/3/HYtFKHS/s33bJpR4k8r0zqkvgg3L6e0RPE89bZb
je7UTwxh947VxyFgvJUcL2ox8bled749e7pczk1VRPwG/Fu2NSY6PPTkfUPgjhutS2KHxTf6weI3
tDpJTsXeTWrDJxtQAzqkvzENOebz8OR/X9siJUnRVoOjLtUThx19r1Q2Va88YFIWG68LIqLjMfQq
aBJjjnRH5v/QoRC5T6hx9NNQw1gxYluQqeFj2E0FS2e46u/Lw5R1KMYMyxxkMUIMtLbZ527aN2iB
xId1rMiakbZQPRtPuYdMw4BTkxIO4wKFtxdr/oGWVGkrT3iQhJgiuR5U4iey3R12Ktzyby2neOGy
avx+dYUAEmzWBQfM+wDLQLwjcnt1b2jwyO5gSnR/K3ZYIKwrHzeonKNLcPq5WfXXHPHuKoBAQTBX
aDFHThWz2ZxXkeOF9ncdRH08lzz9Tm4lLOZnD+xKioA7MgcuwZ+Bbpz9wfTIE/dG7MGubZ34biiY
fFLEg4mmzYy1q7/wWj8jAtDBYs9NBMyXj3fWqr85+zo5GiXyhjcJBLJ4GeSh0dALAySAxXu/9OCo
hq+c71yOtcIqs2Q5kc4n7/k2c/eZ6mOIYbkf6ZTG4MOPLUklaL0prY1oLQ7q1lEj+ZmXYSdXjP1+
0c7QqJ6rBZnIwz0LpQCtJwWKJgLchOwJhvKjWA7lCRj0CV8/5CybjDNy7eRAW9rANkXUZRMacaId
cEw+z3VgJ52IvW6TZcjGUzNQ5y8gu3Wvc43wfLzjDtenbvfkL5uDJdBsTK02c72F6B3LmV5TKH+O
amssiiQvH/jMMGKaS2LR/nfbdUJdcIISGUmIX1jo9z+BP949lV37LTEYl+6Uy3KBGgQgvr0cnf4p
tMeI2mgn97pMIV4UPT2Fsqxr2R8KVJUvwn8EgXIEGks3SGccGextmzsw2G64ve3q4uOOR2G1h49O
9AMICCjTHDvCNaPxO0Zkbwr7CfNae92BhzY76eQ5QCVwTwFQopVgqZE8uyv8DOeaeA5EthLOilFf
to9+0QtPr5MAA2M9H/Jjpsej/g8TvNNQWafEj/KqhblqP1Dq1XbGVBiEes4Zlaeh82Y2XxqiHzu+
IbmKHfmH74mmV9qJXKmgziIWUOjXq39co59fB6ckF0bdDcqzb7pi2dLzM5kvgGX6Psbr2vJAmT4j
UNmimskIv7cL+/TLtYU6lXDoern7jvKGg4oFHXHCyN60/VSyBO13YrKVaGEZfc63RHvuASpJ05zY
88eDxrEyDfQ0PasWOFkq7u5Ha7ScVpRcQn+nSSNKPzHywmvBBVQWPlFVpz9zuGmjvcNvlrmtH973
6pVm8WEyZBpzAiDlq4jcbt1yVa5raaP+9OqwIbE3qJfLCcRzenkEYnSQqNFNI4SFUtxLCVQelYeO
Cl7jeg8j/kAH/uwgKxZcf8YBpb4XJxEhMTYbXJWC4fMCUN2HGundym+OeB3Xv7hHScuvIY/hpHgZ
O+zIBP8hKRcadDtJ3MfGXIcQghK/4Xl1TzS08yo+jrr9sIXQu68xOgr05Afn5UyB4gckH2lz4lsg
ot+BSZloSL+tyb5runj+47rUqlS2MTwxdRhsp4NBNMOxO/Qk/kxrNimhNdeapzYRMuS7Y8DJTqi0
47AxXPpFWiDCbISC4phASsv7M40mKKlNOiD+VrvWoZOKNu0OWGkfVahlusqbq3Md8JYWgjO7GGQl
ZzNJVRCUFnLGjDKn4lj/xB3DzmyQcviCToR8DuIJUgPNgdEvr8o2fX8IGw0skVQCQpOC3ctlEhKL
F3rBsEIakKb2DrsqIhBk5IYdcP8VwW14d3sheN2i+ePduwpkflKWfrJs9URXMzMivGtdRy6o+lPm
FZFZCq6N7xk4W/aP8eEiDKQLh879g5HnY//Wa5eNf5ZX1hBjH4E7wHzPhb4WgSssr2hu64boQ5g+
UnuQQSlB/YgERIrCL4KEfKrqZPEYsjKp7QCUBprHpxf8/kefmlCPlikQW1LIAjlF+VR8AR6I8VBN
5BqmMDY6w47de+xmVbtenVeRTwh3E81JieX4rc36nkGTReqap6s/dssVJqH35YTn5aCWZ2itNiQn
E+pTEVU1pdtGjORMhlM/0exqCWESUr41KhTwiNH7kS0l0vM25FXAaJA68BCpKh9A9lwPQBDChmMd
8DNqTgdo5RbDPiR6q5SzSNCfSGHqp2RdS6Pa2yrcHvYp3jdKjG9XmmHofElO3QI2vsdXMqjo0Nw3
CHkfDJBgbYG7x04GmN8+zRoCwGR/ltWYQCPb3nuBhDSEF/BQgd31m8PfAQGTE0+4TLqDrWJY6wg0
T0rAR/ajVI4UBiZ8InZiy6YFXuHMC8jejHvwb1Cv3sUF6U8zxAsM9Z7AiCaGQKQhRzGyumBs0+Ro
9x0Ji/2bMn5Rpf0YMSOPdxCU3fkeYY16MFt6Iw8RsMmggvmJnOP0W9WxV1aYB9G1IlZDxYygNfmW
WQvp36fsR5WF0MXoQ3njrSpmM82MoJqBtKi6D0HWY8D3G+EQjG5q4yNYxypwY8WW1bgGxTiRf+3p
oN+LE9vlU0GuZi35LB4Y73/+ntf0qQ9Ue2IT3kGxTN8SQJRfhhglRvn2hjgSZVql/B6u2gVgt5Pg
dv9nvK/wB67AvDby6mJCEnOpyI7sjSJDhd92B4y9qSr3xmAss2/KTHiS4Xd6iaHsXuc2/1LJ3mHT
8deMWORf+MnakyODpYl5ddgyXuSYSAoSkGYH32ZMNbBnbLJNN9A+5tf/k2lJw+xmfWMraFLn0Z4F
jC4E7heV8ZxxkI77zxv1QDV4JVTmGvgMsXTpHsue0cgyCJRep+C7t+tr+PwqCAuM35aOaSRlQ//G
3FPzlPyMpkEWnVcgn/qTRVYTWP1DnDTXmFEKMC7qIYsWL8/95ZENrFDghgve7ISGpMD6U+2DzNhz
R/l+pojvVKxMNNxWOP8shzAtNGdwAem9gHnM3Hmbe8Uvl6Wrnyn064iu/fVzqtfvg/fet4Ci3V9m
6Ko/D+hUOqOWwH5BV0LTLDoLibSBvGiYM3JHdzHrOH+SW8V6oZmtFXskn0P1F2b+3rOax4geuU2u
IIwy9C4iJiuGjUfFhOYFmwy89bngY75guzH8wPqJ+scN++8J379mUe5ZisbD+1r4dU1A9+F+SMg3
RG91s5lrD7yFfCSZKlqWEyYkku1ZFdXwaoBmGrBWPUQtshL2O6pLqzkVeWjpNLIi1y7LdAFp8gkA
9O+C+4VjgKs3ZpIjR/dWUykRoay39JuX2CC93UzMBJIzo3Ji408RiX+Npm6UQ/NSGm3jFkNTS3X9
Vla6K+z3ErFhye1Hekf470uFqWMkIWpQFP+1GoAVjRbUtdbBdKs64Z/HPg61cx19SyWuogHa810L
1nD9vVxLy84cF5qSER6F6+mW9d+K5wdBvxtW+yOrdraonJN1oZITwCqRl0pPXTRmVodcoq/yb2bu
UxL9CMQ13XGOd6bbT+ry4VtJbiPMlihl0HBHCzvh/lWStFyRgRZzPtZu727LbfH4g15ZntUdcu/Y
haOYIC5WgJ2IX6MjVR4L328rn6LxJ2MpfzgG+Rl92Ts1g8541HhQWna89wFPznpxL5rcRiFXUCCe
OLOtA62FORgJJETfPwAjsCOBHtaEnfkbnGQRoGPoGvJcRiKuh5yNJXJlH3uekKeIac/W6XSxHOe4
Z15xk6WG+UB4oRs4dpLiQseZk9QwypEsAPZKt7OBFoqs8d1ad36zOrFAh77HEjNu2y3mVvK/hf2x
jnzVcaXPubdbZVAcxnLAwh7JN3roGy/r+xUm4dJfIXRU9NN5BJOQ5WmX7QN2Prf3oRYOb1U09PXM
CafCqR+eZiy1euci8repFB1+aKLUU0lV6sJb0txgEu3DxOzn51jcVX4UnlfYRrFtT87xZ+mnUFKW
DkAhTiGKO/pMZS8zubXcopJMpLO7+ZowsMjYy4yFstD/8pSsmERzSvDw9DElY5sxJaI3VkZefKA6
RV3dbx+kEdVrs5TQyFYu3jksJ/R7Aw2ExBQgBuk81YAUNoRf410gzGdQVb8naKS2aIrfuDu8E6mK
aVmKgk1dcRipOwwcrsPjdv7OjrUB7+sc2dzOZgNLDqOey7jV8txYhYZXwcpwL0seaHeDrnUY/EFS
EMJ3Y0OQS3ycTe8yFLfJv0nq9PrbAbElzYye0DTIPWTbR2AW+vUGLiEUmYgmEe1QkMDuK5MWmrzN
iASUuSVZExkT7uYnPdTzpv506AJQvchVlTDBBEdmTtFAGxeI/mPnTqsUh7C//RkWnGVvyxizSply
SYSeH9Bye/Qqge4cAGaeQoseH92prWzRSgXpnEcUbP1PgpLPcFSzeUvjCF/M3X9+OSgciwaMqcM1
tPmFb6xDr6KRfzG54og95I2l2e806HPCi9CENHqLXGTrk1IxMnpd3LUt4fIyjgaNViqRMOAt4R6o
WfcWrcpR7rWnkBpys/KQP619eSLpSF/YZ+LR8YqQ/+GGS1ivLeMslUC1f524enf4WHFG0uTAaLK4
vLBORVNh0Oju9NDhsPipMFawEOsjKtqoAAmsrARuYEhMYKa9RHqKqydkiL2RnRCEqTcDMLzOAqb+
vFkU36dfxgokCEktnXegwhRdDtj3S7Gxd+j1EpgmW7flx66fDwBGQpfCuSwUC0NGpRceb1qvcRCo
+D9dMQvh0lwrzcQ5ZnUx6J8fkg7OvHlFKngiv89caJC/Pq0sgiJjf6U+f0sZGhp3nagmZ4mM1VMv
B8gjgKY5rhzUGk0NHGYt6pg250S1quxOMha/LaRnSmRbp9hV4fWuMNNzh3twAfT05fr7pyPJaB63
sg+G7REhLUsDNtQNaXproz/rm4RBPn148FlLjAztoxbVb91tcCBn9aFVBfiIypmDGvlCuCuaRxAL
1KP1ycnWtGjikBQlaPQTaBTGx30f+B+BGcpfmveiXcMJr3j6cqC49RDip50mbvx9ojU+I5Oe89rg
SPWJ7BOldfvEH9XcmyxLcPcfxrO8EaR5iwkMRaVT6/TN0WvLXLFquE/2gOFm/w//gSW72Z7aIAPP
XSOACambMjW0gFNmsp81Jr7iEgbf8va4Alt6RHgitv/gZKLjbKcNSWloNRA70KYYOEDhYm/Z1W32
GbiPGFVfgj5MBc4mFHTJBAD7GWKzDO1IiWRMtuV7lnlXUvVr3LPCBunNrhsx3KVpwpPfTMXzrNs3
3zcq4U7KWiskzBcBIIbklVqi0JCZxzB9pEkzL37B7iUVfOUSPJ32C3tz2nqyjm4/XIrxMUKXpim+
b21a8rh+rU+hhdVTc7KMyHKhC5ThtdGNcv/S/aKeFqrzNK1ykaA1LStXl5A9IG0hiLyf0IvLrspf
f1tX3eHHEJOZlenBlWyrghkbPAvtVDPRk/hn0KSrCghoVWvRe3lVkwhhbZO224oifyDQ4xrWxu0D
NJ3LuyZHf6LsCbARw4+aK3VTttIilp5BNV0pcbqKKLkx1WXgym4dhYas6j+vCwmI0ubCb42vzL28
ihFa8MRRTn+mMafMz2g2A1biv8WH+jtEdsh8DWEZl87YSKLM0hBzZveLnwkIni5sA8NCjiGakfG8
aILY0SGOi91VNXaQgDNs/gg8cuH+vmVgter3r8mYNlUsHdC2xWwYjyRk2YGh7YrO0uiHLus3LRHV
C5q+aj04Jybc3f+M9gRy+PmUBihCq7Kt4SgsdZ6lYRxmX0sjw2cBhZVWczIPR2MnnDTNuc9DFtp0
lSYQmrd1zA1YPDOzAHyIsrYH1CcO6yUCFv0pWT/V8l73r122Iuwxw+4umn2yU30Zil96IRDyUVh3
nMPXI5VvWE1A3wDBIf8Khc3nSPSRx9NoYzdll88Ruzn3SQE1f89FIpbCrLb8EYNm9HvLbBVYNQCM
1k/lgH6TVRflPj11srayn5cm4sELqEJ5h/Gka4lNdE+6pJEydKq7GGCMcnfqt27A8tILjNNqBmmK
YmNooowibVi2CNjuKD5PCNWjiXQ1cl1+AVmZCJEIIUf3mIG+ci01Z+5MJBCl/phcK+b+nmFz7WrX
khbBQq+9LsBRpkn7EQ35Wq7Xah4ISgJHnfhFdGOYqhzf2ppQc98W5UCQQCd2isFTWp++l7wfR2ro
7VlmgI+nDhnCAp9YC7CgZO0IVHzJNTQK4/CkfPzEYCoRVLwPHtnPJ3at+1YUHu1TvK+bJgKAX2bR
WoI9RjxQGlKE9TC4Xiv8jwhm3Lx3tTtiNFzcS/9s3oxgreaYtEPIEvRpL5353N1hvLiZp3yGxPAv
qb9/RRix2/0KGCo626+NnlkhivjBO1KZObg6TB0W2Jb2uI/Ap4vt/DTz9G+j2QTOtWVUjFdiGF2C
EUAGSlv5h8WCSn3ypfDL8XyYAYcLf98wAZ+w2lkhWvffDZ/ymp8OylcGOuIjgt5RdrmmcOIyYwyV
SJBwIJZa8J4cvcoHwpSidK7XPPzD2Q6OmGG3OsyoHollWljmLi+Igj/IOTxr4GmdKKykG7eYI6ZI
Jj2O2yzXTBO09wMR77GSE2HzwRPmaulALTDgKurSaJKCmXM5d77O2QpouRJeSn5ZloBwNUJn0lAc
cFBzWwK5wy5tU2F3iFEd7Nx6tf4IJL2CtNgM3ExhBznJRVUSOLIwnbeYibLn9GPy2HtqvLX9quwV
9LtLy/wxRYDTdEEIXBPTkDWcM6VHnTRyIpXpnGtSi0advQRNe9/tDBBJCyuQp40X2x05c0Yqeoi9
YFu9g71CRp1115rZOLxIwn8maW6kLDdPEVL5nsqcg5YWYjfRVPY1IZE591ImLFZX+nQvd6K5d2Nl
cbo0j0wcbhhGVuwXbLCMK3JqP4fbThrK6pv1Yw50ugbo/d+wOj9iTvEMmsSVDpEEQ10v615e03FE
FYopxSskHhDgZfCtnyI+7/nd7MdGnVb4vvm9PjlJm4wkL6XDUEBLbgHsSxjDh6a4YuMGlUSDG1yz
H6eBSrFAp5QNCmYhAehcNie2e/0NTO6j1av/hQY499qP3L6qRSdnrfqi3sMobSmvPDYzLybI9Q9h
6qcvNjJTQvz5W5bSeoPI5lapW3qMoLJaGhCbeuKDdM50QKsV25oBDE46TrMqBIwFaQPDjQnSum3v
8PdMWqTA3InbW8DZgX9/dyrhXQDVekyt0wP2KCWCDPgtpSC187VkiFxv3dlvvOWX9fMg09qjZPKC
vLhx/87caKUncoD3BNxWXFhqMCOo7CaU94krxtEspOpZKqSFnZ+TkxCjvTVeX/kZkkFWH5j34JBg
cob9hEnR8w8dcXLM/+s83kCg3GE4zl4IToKKB42FAyhBVFlnGWObq+1wRV8n4b31vBj/ITTiqlrt
TVSCNzOPdHh4GanC2teVH+dTdC0H13iQY+bVh41xDuBZHdtvxgvW48IkHDqyHUt3ufJTUSa0FLPl
mJ2jizs7Xz9EYhsSPcVdQNjIfIgkG7HlYZyKXt6lomq/a5I7OxglHaD/adFgqV+W576oqugemjvq
JoNRVKFNu/TeSeRfUCmbQ4Rw/ecaUYmDsD+DXUsT2I/Zb4pXHi8PnM2KPsZUHNuFeK/DRIxiTE9+
d5FsPni8aXQoxG541NNf6WUktnXfi3P46sTkBDgs1E/zv8xtYESVYHpz21qupoMykABhNjMov4y3
xvUXOtf9fUJQDoHRkd4yDWQ54r0WyaEHgXwS60aRb2G6U7gWkuHy1FfkYhTaXR0H+nMG4g0J/PTL
RFBUlknM9kYvP823clHfGiWhWs6xxYLivw3GHql7M9aXRQ30HfiVwGGHfY1DpBSPMcoojO4UgrD5
sYe+kXMQKytePwTYb+MgQXJcv3qTlB2AM6nHVJ3wizyJuh6Oia0Lib+d3FqKmDdE8giP2gZ/uu7+
j3dedBkEXELTR2jZlqehtNST13VNigs6CkQtUfr+4BWerKIe1cXqH7KoEHetvl3dDpAOVDSVOjDM
vyYtZt4OeW3EX0/DAZ8ntdkAci+ApNkj84PAPATrBQCh6Mjzk1c4bIdiexer5LSm2auIqt6f2zC6
Vpt2sDL5MpemojzZ2PwlR7kSTbjB1GAij5SIwJMZ/i3rbOscu17/uG7Y0o/xp+ZmEProzbzy0CT6
vXtN924vsW+SPzEpuVKimftpU2vpnqq1PB6S7CGbZ8QrGc6+piB1/2+IlQ3t4iYDrZ72TIKdMjjY
jvM3BO4Mu6WseyXHCuyN+w0btVm0WFB7so8B3xCy5EpOPVWCIi6SQOg8h/cm45Cv67/wTi59eDzr
VJAkLXuDghir5CSzCZD068RCNy+mfUblWnOnJZL8fRpVdYZm5dzdUs6o+FLPOUqKcD/LmbPXxSYr
dyKUqgCXYPsxzgPst9p4lVUD0PLN8+0TVTyUCFiqYSi4+m8oa0vRU5QjDjZJLGZc9Mphxoyth57C
PamqQgiYVrqVPdsHohh5tEwNtXvdwe8Y3w1c1Gpmca8ARhgcrEBberWgjbRPJkhYQrbdcJ7p3Y4G
uAo/HA/GUF60Kle3byBfKz3QCRUCpPDRgJZlCrnhK/yPlxhC1sF06qZiq6lNIc+CxbXKRByr4HAN
HO/LcNj13f2lM89lMuycu+cwI2WZ0F0Xq23vKG8VYFrvxJe9Fmw/KE5HLU/M3Hm4WDar9as32Gu3
J+cTguaCPOdq+qspE80QWZMzWoBEi5hCRA097YBN/v4QTz/J533OqyyvNyczunN9Yq3GhCYfrq9G
1XbYRuYNbLk3YhqvvZkeanj5IHMbI2iL6W9vHvbtc3ohDpC6ZP4MfvjFqMVUD6CV22AZ0KPqFeVR
jRHSh7RIfzUaqski68RoZjBbppxw5ggY/TKShrVjDShociCBuChc9U2kjrT2ARaZj7yQ3ogCHsUG
EuVfbXHT8alrZD1U9lYs6zrZGYMTe/aj22FuTSb9brB6HjEZ+9QOu9sm+uyGiED8o7Uf+kASp7AF
QOj9XlMbnMS7z6iCHkrIst06hvxw1Fbc+B9VBKWGTuZg05Q7Id7nw98YSdp9KTUFpeYJY12iPBoQ
2XAgIKHNA3Au6VQkjZ8r49LXU385WZfn3rBAqsQ8sAtXVfdAteKKG7HSn5kUFw9XwLUvkZ3g5iNX
f2EaDVdAVFMNsQaw1T1wgp7AZzpob+gy2xTgd2Ss6gRu1mqcUOnspaGXX1AlBiCDzJr49teTS2zi
Nw+0PI4PrqvJVGpPDT8a9PkgTKVuNwY+fCC7+A8rgE94SPrsfueRMUeUGBICHviosXClwjfPHZbR
TVtGKXm5oBkKxSo4juE/lJaZtAa6rcrzk4vhRaOLyBuYKxUHOJy+oF+jn85nVvF5XYyUUlB4wQ9w
tNX6DQhHAo9aKP0elheXbPhj6hefsNpzZf0QfZQ1AmZCUpSzCBJ2slf6c+hUvcvF5c8tflq5QYC/
mF6SDbUXKGy+CzRTgh/wVQm67lhZUXMxu/QyRCsrxGQNZAmcnatwIkZUBNi7DDtndbs1aK1KSR1p
hyiBO/q5akAgW3tvY6RJNhMQOfupKYDCzGZggwk2RPDhgYOuEsvwuzDY4+4xZYRmrObaM9LIMb3n
xCCToX3UQX7gYwqEaOHaIEs49kvdFavcUb4AambI9y4TDdNnrH+G2sMeGIFWiDBp4PDNgJd8ZZ8i
nT2J3L9oNG7o9i43SnYx1QUhdZlRpTKKMNxQgrg2wk11pI8V+kCd/j1bTpDK2pNxLsW+pohF2VeW
W2aFK+Tu9UarTzHLG2LWF0Hu4ZvRsFq1MH9Go9bc8VsTcmwOSilgLM4pAOjpcYjMpFGsPV/9Ciln
iuOEzWp1yZIh/akWv+oslRRTju4qHoPhaAt7k0wJahxE23cKNhqx1n0LP2NC0B13EzE6CO91ydAw
1SgkdPWe1w73t6sPrjFPF2VYfBku2ykmOcJa0nPdSb3jwHhzOUtjo4Xl9QodcS5L6qHqVmGYCwVV
asBL0LCrSTVgl9CrqJ3qQBFtr0Jp1CTdAjaowufTc4V3QxLCMcC5BeOQSrsutEobJn854y1erAUZ
LM4V0SxLB9hwvwvQRdpnbMLbEwDfvdlyllCuh/vy4OVRMYMxvMFtNBVWr80MQcYhZmf9f0Rd9SpO
hOWZLZ5UiWckWjS5cLxCck+tQIUwsreLj/+l9boAD3Vt2VU27IILaLIoxNI08Ac4xSS8hGNKowtB
TN4CyIF7lIxkH74chhZofj8JgcLhyckISGOP5yFw2I10LoQYRhHM/YK2rredfdk4c4dzz44JMp9P
hjtPauGwMhHVQanqFddG+bvmlgfOfMCX+e6zf/PGyDB8VDD9HIluo3KABJXxfw2NgLYTx/tSm5ty
l1cZl4Lwy4m/i27dvMd60wxWkJWvg8D/DyDUMz/c5BhJfrn4715HaG194KzABsSPjJtsyG0vM8G6
4lTkXipppqNI1nn8+TtvFgtWAnpNcdmnhD//p4dUj0fc0P6bu3NSEZExKo8sAt6/g3GJ1TfnYlXQ
D/XCq967rEyrDFUZcdQmyovZjIkpZd/JxFoqn0ZBRFolE4wHSYooeAn2Zso7Hu/fNU665mGtaFq4
8TMrZj4coK9Bh4FQwXV5OrQ7m/9BwR44panuZqNB4sU0v8VEdkbuimtXBT0IvBK9C35GB12kct1O
KM93dQNty2qPXLr3nzWIPb/K8Tp10JFegehUs4OLcMe278bo4BOcl3tL9oLy5nKhkIHd/yHZ4SGU
FA87BjnoJ4bLWXE2/skYjUHsddUl4uMfDnye7MfVwmnpmnqoR6CQPX5r2eWL0fpNoBZpnb2248ah
/TCb0zx1xuwCke4NkaLmpXo+3fiYSS1m01uA6nJnYVeZckp3LcbY7320Ksj0y07ypPTFII34gfIc
1SKVyWziKwN7Xxu/k3LIQd/JWg3QTvO+jxW3cHRwF7vyo6NzDZng8go0c9DWam20nK15ofgWZHTk
xVaeupxKYPI8/PaLmVQGpLFpFyE7wtFjyfhvO2YY8epJj4pEDRwPGH5pNp4xuma/MzB/Gt7QxpCM
hxls7EGh06jvzAc1g5ebKSReyvxfc6NRfSuxxuK9CNDMNIOaDn57cY91bMyvqZoyNSvez0Xyp9D6
htX8UmXLM5fXuEfj0nqWcb6xZJbf/XnS2+SvaOQ8+6yjUD5Zpwye6lyEqb9cEEI+Wx2QHK3EInyx
uKM0VdfVcgaWdKYqISQ351B8MhkD0COFGpmavj0p6z9oNZmc2dw/VWhPd/tyiNHmy7V2DGF9PLOb
4fO9bxWM1j7xFUrLachVT0O271vgqDnuuIShTIzoQFyoJVwiRbvPUZGI5VxR8PjKgplUKvAo2yW8
RXp3WXxvVcQAc6tXHn7Zb7iAw/zE51W2wNHw1lO/AN7KtUWOTPaYbZXu66aes9trwPzV5ft8QQ6C
ToMrC3jgGSw8T2A1YOPrMKkvDOJa6FG6jYjsSNA9D3UWbm1fJmVWxGmOlHg108rRb2CmfwzDWIfx
mHy/xQNmptptaoEXfSq1BQYzEkvKqhx1XHT5a4GobOM8/ig2UyuBzXatlyd3bMEyLAYsEUccNNAk
OoKOvuVMm+p8vNXFVpLvJKHLqyccg6Qr7o4V0zRyaD87tEjE5qw1pBAo2WE0bLBTFOzsukrCG1XN
sp16j9jE9JnGyEA3ENkARkY2kIqLAy6BGPhMVjFo8VOTnWwvN49ZoTkbeHltlUGGJHoB9Rw/qkwM
0LwpbQAMAVIjuHX8UWyVtNCT006+byznvQI31EqPPZEXA1VQS6amzepNdevM1gxvBIN7PRZlpzjU
oUy9kwxFGKkkXkBsLnEsXVzJcTjBy8tJJj/PL65aLFbJd4OOlhcH/dPJUsrlnQf58lzMzC6VdQ9V
wrdNWPXXeWdVJWm+9QKfvwkTg4N5E7JpFSzv+7bPqwdyerIyMaBHuToYMS471/izFBD7o/GgeTii
IbuDq626JatrCsMP3XSSh0fe6l1huMNvLweE08V5M1vdn4r6sUMzDtC+NFJ5MWt1z/jG5dLUiWtk
Wcu7yN2jX7XOVnZjravW8nP+ONzc0Kefz+Ysri8cmqaDPEw7o/VQpMpsleBTdpcGu/GqQJbRLIR3
DZS1rt4wp5XLMSig6fpMtAcWk5Y9PdCc+NRmYhK70xH1zWS19IvAJyAhWhkjpR6X7cDk/QdvDLCn
c45EXvCzOBD/GBhdGeWOI+HYnVFgSG2wOdEKDdUietMMfxwPTci4LOkUmBOxxqwz/sBne/xnfhEp
4kJ/wdpgJyKy0h1m/in5CWN9uDcDteu6u9j/NCIy3AvkgcUBiWsQ1XrKGxvbgkoRtVZJRY4xqX+r
C8ysn81NEPtQzWBrnGeMfSlZcSNJtIf/cUn7UkRcPkqYENdi9nRd5HWLjuFgCyFNxnSHlCQBNsOR
USNmoGhN3+qwhmNY9zvsv3R7AhcpFYVtnW4YGhDmG1Vzpkq+BtNbKMlm5A5T8WRBOVB0Nu/csGyo
h+F4HlgSUzQ+V7gKlK/xMDCc09adbI8meM5Nl81ZGOqfAv9b0NIxRAqCmC2JNfmPNnr01fBakgHp
+tOjfUQu0PA8mKHm2lkTU30Zda/aPC4udD2UOSIdQ/hTPwg8fMe0BQH/jvkceMcqXa0RCZjqptB2
hBqhaF6cbGlQRRz+6mUAsNZBTZNDzqcXYl14GB43KvYMM07KUmyHEkmBUIxdcrQltu736xcH0rOJ
nrYcwpSX3bnzeSsZNM84ou1iNYjKuMr5pyg2xypuhYml0RxxKLJ/7LapN4K+tOJ/C/uL5xPo3CjD
nJtKfJgJY3R46I3O5BhEzgGlsUc6Pb6HBZp81OWrjb3mBb4qZNA8RA1jCMyu/h2TXGX0YIT85ldD
ITkWBfVVt5p5MhgPOrr554yfAfCkZfZrIq74KUjyGx4gbwCERE8TzeCp7yUsBOO2hMWLnvfk8mJZ
AVKUzKgCUMPg5NDqT5AdvMrehrAPZh1vTTZpU8ix+Z6H+VmQuhJQnvHl8ELwxcAsWpfCgNTXbSJ4
PhLpArYAeFW9ZfJDl+15ThzvEnlqZE1KZM9kOY65XKLOsOIpMKJVnfGiC/dn13i6P5DTq/FwbQGX
6AVWCrUMfLhjXO/JOoVTHrXqT2hLKoIHYx9lID9mXFNL5ocKAgqMAbxG0yVHbOieX956oNfmvCjB
pZMk7QI7b54NYxXmk18ih4T4Bd/awVSHN6Z1ERsO+p4OfjPGoYFNQh3ve3qCSaiQ7w06NaDmPHa3
miPtG4Euy+hqeL2mcGNmL3uXpF+8pXa+z5sla8DNhm9f9kHjdWKr9uN5lGqc7QHnN1ryOGXLYVyK
Qn2qBezM8KvXWN4Z2fREnYYdKCtlPY3R9s6ffvOoRwDYd1ujvvHO6p5Nvk3b1Efqzxc8Ohsv84i1
3URJuWCTosvydgsmFcYL0Ok6hRJybrAuqQvI9q6uI5bjJs50WxgreeYUN1UnJZh+siquQs6FeCWX
xoZlEfYc+gv4nH1KXfKvIsXn/RhpUaKsVlrzP4hX5MWZXe0WZTJ5L+m96PXVxoBgVz+OXjHRLAff
TgEVte7pWgh7Coxf8otKMeeXrCH4IDKQotktq5ZhOsUT6nPGpJwTfn23yzGtB3lUdZYnUpU6czf7
X0VdcHzRmMuooByTuLKAjP/gsR6V83VAcGhEEL27IzeBFhPBCzyARAZmV4XESZVTeZd9GjgxDbLl
MCU+fG8lSFsTSYd2vIz7DpIfVmdj3sRATwmrQPbsLuHmJkK07R/w0akyviukHby7mEhBfeuBFBOn
QHJjB4XtF2zLxa07WqyNV2SSQDN3aLuY/Q/a4SYUPyQXZ7l0YQkRGCX5F8FNkNRlynTq9qQ18uk9
d50Fg8o656T5M07fawNms5MpGplaCLsrXzrlAc+p4b74Mri0VAbszMrT4S3Bx8pAdIgj8nnZIKXj
HhLFs28haOa7ggQ9zwTpvml/LV9DFGVaYwlE1Jb6lS9gm041R7g0WmuClpaHH5GnkN+vhCakSgVZ
x10UAs+zaLTH/hd/sUWrAFjXXGkiL3AYLNq0SNEQA8uGJy6ACB7h3RHZuCbLZCEMKWjiQ0C+ogTL
AuwtztbuscgwRMnHZQ8d8M2y6Jvit9XUVFEzqXeZt0TRyAXhXLbqPHS8kAEIRmc9PRthcg4LxMci
qouXrTJn4IzgOlOEBazTruU0c56DKAp5wewNHM/ADJS/KIbXX0HKviH3o5Zw7kn/pG9+SjLfUanv
l7sMmZeWvWVbjNRG0V740/aZ57fbBM4+5KoTkZwREprCPOacRhHWs4WB5LxabmGa3+C58dyZ+Bp/
U1Fb6e++mU+X78JotfLES6ZN9Ut0dClRaBP34xagCHfAa3E9+P9uhBDeIw0i3nmM4/hY7TncOk18
TLO9rcChxj9tsbztA4SspDv6m6YLBMOpj0JEyO42vHwnN28rI00hb9D+6nC87n4jNEvlpqFixs2b
yZB3Zc3vU4D44TCARcgf/S662F4KKSQtqYiP3rr/CQhOyui7V3dPM4n5Xx7x3JZ6xZE8VS5TvPoq
CarGKgENa2FqWJf6BXqI3FXjk55Dr3mGfxM3Stuv9psA6HQoCivG4Q0pnm+Elip/Hv69mVsoadUI
AKW2TOQFEsMZo9o8KTzzgSpbaqrMDnP9lXPxpb3bdPodaNBRzY4to2eL2zITd+pJ8F+lNwrJtinY
D8Dh48lRZjx8LTDgxd541W6wfaF3fkQ4OXqGReJ3YECkyX7GBQ3YTxRbTkxSz4+xy8RwDLFKww2i
x7p3EtW/sMH8fVjrFoe0UDmSckeigbRmUbEEbIw66/GuDOGcxCcAutBTOqQ0InEaCdZCTyULyuXe
LDwi1idbReFYa630F/uhZvTfoRZIhi6ogvxXAjElZlk2C6TaQnJfl3AZtES7rdpvmiXzKb8mF+Ta
ITnw2My8NeQUXM8dPFwUAY1Q9VXDURXyhIz9vql7FDgeGq7nyWOf+mw2ZfjiTm7DxB0GOGqjoLv/
cITMJ1eEGMSv/jDRcVqoV4vqlDvnV1x4YZmW6X0ZGqkNL1HPPW2qbTRevDbiSCKCmYBM1vf+oH6u
N0Z55Jlndehyklv5EZatWzdncHnUA7p5q+JogJCbpSLQRn0MJIdqSIhmETlu0M9DWdx8djnwTiCx
+siWzzcXFf7WIkHoY0JLBsOMGwrWm/ZIDxMCNnEZP7zyLScAm2ChaaqlNydEnKCSIfJDsqsikezz
nltK3QB+Gl3TTNZPWpkvplMmT8fS2YZB06kY+KE61GUkVcNFBEvEn0effk6qbcMXxTlbnNp7pvfe
ZPF/EziTBh8b17Cgi8f7SaDzrYS9JCZLHkvIoBD5TIvATAU3O1no/qmZqeBPNCBZfB48u/9IzYOa
0gWrP+eWXG26IJmBAPSEAGRwY9QIEJoHi9ya97bXW2yti1MwLI/rV66NXSj9hMjQvIwcvuoCcvrH
xqKvdfMQfnS6jAd+OHdX15D9MHHCx+4uShVLkQGWg379FtPa5xrbmW/kNsOsXT9ul0Bo/aOZqShA
5czoa/RNo7QFjTJGW//ZWO01TpXb7G/g7DDtnOOvla3prETfT/d0nw50hbWG2XJrJumR4lIwTIGX
lqRMFMVyKUOj9BU0vp+fARE1ZVPSg+pJsSIKu7vLX+qUO11ShMSFt/R3LR9bCVZ3Di1Y3Nq/pI9y
dAsSuqi7rwvvUlXP8jaKiR0fL+YLU81oxcJGsvaXfbU2T9M6uc4pI0wKA2Xi1vKx+ku8NozQ9TMi
LGXvA1bPtSvkRkjG+GVXRd2PSDPlMYvoBwF8wZtkdu3oBBCgPHA9fHV09Ua1h335okl4jVz87MmM
vdDGQTd7q3YzCWZ0aiC0cxihui6NwADJXcQWIUjb4g1utvUYjI4nd5v2wJjAmUw/kXK2imj34ShA
elm++Its2lQ9CNagD0Fh6ufailXexZD0jFhRBo3A4Cq1IFLnWu53QIhaEcfSmi1N5zK7lxtNWTzo
OaGknHrFakYWqpDqJbiykIYrCtw26NoPcN/ODvyBr3fwV2lMGRh4XQLLlOUmX9Q6IGMDjJwNVqa+
jGp6Eeyeip35dgjutr/lQw2fW+c3yegJO8fwdQj/gWKGKfbmKJkP9wYkdPlBEvWuxXdUH+V1G1z2
ows4brgI7Sq9NHEwMjWEgG66lHWkJ3KzDgToG5jk2aHFJN5Sv+hFWfAbgV/IqPeX9Mb10x+gsuP/
BT/HyH3cUsebQv0bmc8NaRCnJ6Fh1+0Xpjtmrvcjhm7sVmwUP1F2dtSKxG5Ra9zbfEP3phwm+BPQ
58CH70CbGveNtpz0YQuCR03QpaSeK5gPzV7B9q2NggmYr7xnDMaJioLAuqyjHVERDi1+rSXVGaD3
weSu1Mo2XgIMZBXPJ8dURWZeFI1OHE8ieEsevcmRNKAY9jaJ7Rr1dBUqFU5fa7DYip5/rf4LodpX
FQA9gDeOiKSyKKHkJURgFQxKDRhV7DGPqXJTZ8IsVlT3PQwZWU4nUzPr9ci0nrPo70jYtZCGe9n2
Nnx9G7M4nnRQexDbh6Tb9mNoDwpsLh4VSfQxcbCnA+t3m8C3Zc0TRufc39mT97m7RvMRdjTINLQt
vqfwbk6+obAUeC0Zh+3lSIAA5qf8xmuOLt4bCCnTvwbyeT//6iBzYMa/3AU1VPPFB/9NckdMe44T
1TAWizwQiWfR9oFGyRL/zW/Y3O6r9YsfpwcdaVcWbSh3kOvs5LDAx++bVsl2lvIyKhnDInyB1j/p
TbQSlT9XbN6V0MqgJmPp8RLZokkcSTA4ZCoNWuTq5wTcSn0TGxuGLCG49trxYKnoGAPqKkEAYhpz
9e/69f9oJTdes+FYVk+E9aDEVAOe2wLqz3U9U74g1EkRzRfrPqdj2o5/WzLDIGs4eVeOYoslcbKC
gbhB8uFprR7blPF8v+8aW9u2DXZKSOLH3mY9vzy958GN2Nyq7mGsgqjZ3KoMIo5AGfEZYcNqE44f
e2uFci4KaV94UV4nnT24lWCL4xvlqacBuWcLq0Eo3MUcMppNgpGdjArdZE19awH71yjaX+OZjoME
osPeVZha6IukacdEQTXyS/apLc1nXu5pCFtn+xLJ0y8SinsWrqGwTGUVJ46GCdhj01BVawzM18T/
1ogbZfKX9sPrAXbpHFuyBrLQduRdo8GT/HbApH4oCh3ECRC9OXu2fDabKkSOcFOv+Vqgv4BKN/n/
cwKU6J3Q2CaiocUTPEtuBu4VWk3Et/FPIBTd3uF48WzuX38mbACSq1U6oe8J1CNK3Vaz+gjFJj+n
P2ohm2zbe/M6huTDeLiPRHzpynXLmS+n8ozEiCGp3IFM+I8ecVcbrS1Jp5NgQs1kQgKCMHbcpHYY
/EcugZQ2nTpxWfgAH43yxFzCbfy8BAg8ZUJI2s3Sy1gZvQYTBUqNkHSWhHFeC0tD//8vh1XlQWus
pm0uS4QvP9A5w1A1ReDwT0GGtgX8XqrYNmKt0VL3xbsl9DZgHWo/jDfPbzJZW/ia8CLZ8bpE2T7Z
NgjoiboUqiXC9U/OQUzflnOBtE0RvIkkAX9nHH2kl8S1nVH9YvMiv/wdS1In1F49/5T1vRQW/6x2
eRtm8KJFLS2yzxsFspKd2U1TqzMOIiflMia/oD3em+cJQuEx1KzE/lrSdgmSDZ/UUJNDE11cneD1
jcnNJvVxLz6K3jWfFGxOwRvNUe7gbLePPQ37VwBWS2ladLFgvjM1J/HtKLutSwdXZCLH7uXQvWzV
+O89f354mseDIr4UM2x0QqU3XNsex6BolWg6i/u852Q6+cZwISY21UQQZ/cfLXrcz/AfU1a6cfN0
8SBM1f5AV6jjmCoXUyJ86vH49kphRVdmdNb9Ggh89qr+JS77z8m7+nFRZ2mO57HT/Nx5v1J6ogFi
Vsqdzfo/ZaAZconvYRar6SLXXv8+bZepFRbifiTRrKqLJTYGjlBfefXoYSmjGdtPO4u8ijYIsqn+
XBGATdBIfHaWgM1av7nk6u1/aFd95sWjj09H4AoNgWQVo3FN2Faxn5mpjhvJlHgoQtlMN4on5Noj
tZtF6qPOCCVqdyDgT3JqMnca3fgJ+cK2+JLdlxDNEqY4pAfCX7qwZLODyExFXVAhDP62ddPry5h9
fjyWHhRlXHzz9uiTg7y3Wun9hY3sUv0RYhbN+/70nXsOSMwjNGeVY9vdDtCy0bCn0p8WT+jbijpH
OBC+HQJt2jKHPuanJzQpw/MRR6VslIEs7oLZ06Gctp71trAbZslVtybB9GEjdowv8dzl7O0hZdt/
uDoYMLjhQUxKnu6APRUnL06eSFg8gS94dgJCxXVf1wxLCxhwJptRSepcYI5Ct2wl2Op0B5h5k422
PqFfZHAFD6fK6XuNYr16sU4ftEftR7+HOCJCNYXUh91P8KjoihRGGZwObYhI23H5m/M4TWJbajTm
eTwaRliBi5ZyVjwwVwHWppbqRcqFugxgXIqG5hM09UTvOInZcPrxbdI3v/hEJQqyn04IPQcsK0mX
yz/fs/3LpbxpNH9nAroRIYOorcDZY9ynDDLkmnmjO5hG7EhR1UhHZG2mH1gp3SHmIHB5tLbxNGRC
nGOZ16u5nW0149ArO3Mriyz60t60RswDaWBZByrxBqyjH2TB07wOw3SwI/T4w2ZUPR1FlQ9NHe7R
4H67OkCAWZ+wpHFlDcfWs3Wh9Hm6SkITWUMPu/Z4tMtjqt1pZdOvXpYrqg+XRvk5j/nX3Q2x3D72
Ovu6iZLtS6Phk83kpDPKth/A8WEdBsOiy/AUfsUrbILkJ+E5m1qTIvjHJaZ8dv+358gnIn8Z6BRf
842ckB9pTsbVk623mvsGtaZG0Wz8kc/9p+gLyhA09Mf5byW7veTbqiWcrq94UrrdBPC7D/Wb3+AU
6L70YlEtnui69lPsGEBMPv5Kfq50dVE2xvz9szgl0ZYxGvPd4ai1KYYGCRx8coUguS/M2pZWPBgu
Xmi1nxAv7WFZ86UI5Aj/C+INvmdTIIBQQ99ozs5ili16Azr2XXPGgbYHGDopFEcQ14Zz1LMNiHqN
wrYH8IG7BTXbxzgy0GX6ERe8szyqfG03GuptzRiUKYz7lB2sF6opPsE0qkZNfZjWPC70MXnTHLln
vZ7jNKMbySCmC2akNfSnUpAGrL3bxAzm8TxQXYOLAyTJFD3Zvm4hvA6c7ASEcGX3HIUppHS1bmzO
A/03ZUd6iGV7fIq1UkT5nA7Sugg1PMuk8jAiLc1IRRonZ8p/wORYd+CPLBNx+QM12ApHZFyC5Y9W
YTWKLryc/d3YaZkz4k6o2vM9l0l5F0a1h7j0+JauE2QhQCgzMqRFcDITt7Eyldn6nQs96DLjoKpW
CCPLMOAQocgYrwamm8seVVPLi0QJ3m4E74aCCLZKq0Nr+NM0enJ5GK2T0tW6oxl+LsAZ088z0IKp
PEu7wlypTmCg8s39+L5QE39mkRmUzDtYTGx7XDGq65H8k7J4b5bnot5euAi8zp2aOz+G2Gn4Z8Jc
jwB7lRgxFOqGoRa+h1983BXbMl7oSApVW/xtFtbxIEbzjX27rr+DzePm3PGivHptW0wEGvUjC0qG
S97n0peoXz5KwLNeOdA45EIcWxMxeoDQTo+aLKWQuAGVX7r2ca1jlXsw7veVi1vSjStnlifT1MIA
oeqLq5yEzbb/NfIIYDDGxc2UJTXUHdgmj6sVEdqCgl03zW2TXH/lnR2FETysI8X+WUptBS295kAn
lKecTwu0p4USdK9BydLuaYfHfwz8MT9uXw3HLg1ohDXz8hROwm9fjBxV1leErlji/XOzWjkKXf3N
DqejLmRYV0D/zdRqKjqVyU+dGWyg/Lh2T7D6Idyvqr+k1OxUPRsvTeLBavhXAGaEivPJ3VJCWV0R
P4BP5uOpZfbNcqK6t8rFIIZRm+qI3u7ZmInA4dVidv6j7z5+pmT0xlq9fh0O5An8CQsBWbOwC1Jl
9k4s41oqJopOEhnHySVmoCpiqtTyFzyZ5+DEuXvQRjYUR0eLFQk0rs0snjJJ/nCGARBF9IfXDJ2u
ECs/ULfrA8MzFzEwlZ/4gvAcE5y70IBSSkWR7Gf10VrNgSAq6JxUfKIuyRkxqeAlfQn0QQh6tJL6
REf5Yo/yG1vxqFbn4zHoZvfibk/Pdj6sqEVIxFksheALcQuoDjnGMuoyXdOZGcU3H/hrxCnOZ9vw
FEMM+DH2eXZEvVKFVJQp53jOJ+yiEH7laRZbB0xfPdHTwWFQzwAXpx/jw37uvT14kfmMcHKz6WfA
0cMdaMGaTKjNYbQOjbiSSs0uMnm1W8GmasatEKFp/ZQr+Px0bGFNdJDhyCgaCriGmfrLwbSWzCbS
82DO4COQKmwR2rEqlifxSvhynSagNr8dDjaWGoSzpgjC+4i+fH+AKQ7LB7Vu1hOFR8r+0TzY1DMO
R3IiUChFI9C/g0osNk1WYy6j2DOjFTcwdfSivuDE8VxvUG/sI9/TCP58/7h8SyXCfp5FzLxDofmN
O4bn0WhlNB82MCrbwHQ2WR0c5VUbsevsXWSzRzfUMmx4OSaBR03+s9rdpsmUpvm6t8OMA+D3616d
ccgtpRnke3eMCALEgdJuTeNfp0VMODIwjO2IARdmJ1B9Z1pYMOaTAuGrR8/fQBEa5+4Xtchqajw2
puRwgyW2qUFTqbl+u9S3okgCH/Qk3u45aj0vdGpOZZaJhuwdENEjKPJGUUn2HScTXprFiWaJIRRc
kH85L0L6GvHkZDpSUugj0CWdpXl2MHmTmnmuC3mn3F96xtyjF192td2GABp6wgs3NzzLBrm3Aw3i
oU9dmc4nhhn0sqQj82mOFEBGpNlLuGN7QDVpZ8ResUwmAoATYYKQS+1gED4+ls1HQlH1colzJ4ta
ZhJTTfxIlwVeu/8rDyb5XZVXYJKWIbqQnhI0evDXXBywJQo7HWKiIhJ0sgkeU7DxFZIboQcWZD0k
uTUqxrXK1FvXK416NzeG4s8TjEoIjQ9SMW6v33IfEGm49CmLeV7Rag/qtW6Bw2y+JA1imkpYNySb
k8PPbm33dUXvH354yYLEBMPj7Jgk5propNu1SZQ5C5AMUDiQtPOA0Ku0Qv2CFwScq6T77rld7fUA
Jwoz/adywJ3NFEEYeqpfk502u5fuZxfko0mNPHwJPkYGlM6s6NVqr+jqmPyAuuVoGI2nrq2H4tMJ
NOIPyqhjEDf+uPuHXLxgtrGm7oBkJw/6q3YzXVd+s3NovU9xgVbZEBjkshYHl0gK72MmA2Ye6H8b
19IBeQ1amEHeZM3l+SS3207XpK1MwVflcv6zcdj0loN7zgta4LLdGlJ4iLVwrkOZ7sPL/jDmDqAg
OCgfeO17W4NS73XekJhJ8DUdDeCzU4dp539acAffiO9Mt63KQ9DSpDN1EEHTzSeYr+YdQjv5cyA+
1VH0Zv4xJCSJguY9Mt8nmYfPUogOG3b7OsRWVib5sfI+2sVoog3BcQMHDy2yXoIz7dxXC9Teryzj
pSoazYU94Q77Ft8rkUN35VrylASDlFU4QZXmjS3a+di2S93pS8R3WsC+ImZA1bZ5u/Ro6Lobxdtw
WrEn0vvfCdJk76NLkbOrS4JP1XLd9aHIuV9b3yRCBIUMLIkb5E4vk4cwSoCL2Rgp8Ut9yOtIo5w9
aGjWMyWA9MjzIA3iiVcwRDxcqwjwGeWforSgPk7T8orK4nxNhI9KLSsI9hh5wrbjjsLzkpMJspFq
6BhZmCJXwwvNK4R635pvxqg6UTzPMy7eZVsa6Wu7OSBztb6oIno3pjXXzK6y58Vab/hTyFRrbQPP
3zpF2LVc00kY0h+RgOwGwkJiJIzXr4jzuSX/oMHOaXKbFya3K3A0PWzdj3tMFpvgJete9R9SpsEh
etKvImSuex2ujyjvWb21rcz1BC8rMpwP+iZg/VZNOeqV4ozWezKstm0Yl1rqeDJkFYQdhnnNEf0m
lXCo7XWmbOMthXVZI32qLY0qXrkF8wDj30xZUWiWPv1+m+Tmg4mF0/mZV5yvtPTBOMJ+/Y1DrHqA
TxyfMRJ719JKVW/Z2V+uLExiQ/xG9iA4IvCgTTYEgSaLTLp/BN/sYZx+0Df8nR0TuBgVv+ETR/Zh
cXL01CYpAKhWzle9tMuo2ss7JxZyUQc1nCR5U9p2fu7SDqXqkiit32sCTiBMiu5bras+x9MFerxv
1I89HRjKtMWzZ7y99KVDt1K2VWXcEfPLuvZRngwJx5H5uIdFirb0LE9rWBUnY7uKgJKfinT66+lj
R1+/B3sdembgNxO0OGTDdYPss1WMlGIQodH1Pi497Z3AfrpzeXlklIJ/wIArRTfWsx6cAy4mJfYT
TKX9VHgFWcsjoztKKMXLHmWLgVQhJYv9oyiw8GtSnh55X0Ix+LHXMhyOQVm2vDrLy2vjM0ntzvtL
LTYfAmQ8oqjWqHj9HHCnJX//jv2krwdK66qflptz795QjCK9nRWeDIQLPxrAw6OFmVB+OGCyDC9e
1vhxAFRVQb9AMyr54P/mqAHWq055+3tcc7Gboae18ZQdRYCWm4BE2SO7shWjWHLhJUQadi3TAblB
oPVPNwIsg+PVStJkbRnx6P86Q1grCGaVtuVMa4bxroOpZi1UO5MBWEoowLb4x2+AtHiSg6Hb1brp
qULv5Ldla6W3UXzIcNsdbi1oIAdq60aDy6vNGc/uPoNRRBiJE3b7pOv/cSYFomLWjool2ScnbJxe
SqcX4SsXz8DB0/cNTYiYAFiLtMtcEmlvTbxVlSwGikBxP17TpNiycXUKwwg7/fql+KNF9sDWiJnL
5ie9mcWpH+Og8qZYF1d0dgJTiim5E5i9aDHnR0GknckJ1VIGRnanJLi6KULdcmg1svXv34JhVtHx
6TnPK7L7qcWf0m4BkseIROghTpls9Dg2+af4uITnK61XLMs0VGHxg2PhP2IMaFdW8Cc9F/mbI0RL
lz7jVF+hkbhHLw5NG99Eetbebq0UsrZUfnx4YCnpR4ejB927tb2cBRqju5f3HBzKYghLA04U694b
xe5FXWKYhav/cP293uL7EPHohSObZNz5ePn3LX6saZs2Ral80JZXtyuO3SNwuBA5SQqZu0S0yHL4
caMd5XkMR+BcNzGrlq9C0pUK1albSlhh/I6/pV5pjEaAqI4I3qd3qbiDAjaUb11nYxc9bRIKo5Ey
HgagdaCcsBTTRBi3oLu2narB5wAp6FmqShrmsXNpyg4OOFw1WOBG6cjHOwBvDHXugEHBwNz/b0Q5
QBKZI0+BJiJGm2GXtjXX6okjvpXmTcxb/PnrMwn63E5xwA2QBMLNhN4UVrVIyBzGTkzN4yA9CNYS
yf7PZC226cCT13PjiiCgzo2W7XVtNmC9PrquyIJj0AI+6rP5x9Cbl49Ryh/O/QgXT79OyOkk/wug
THCgZZwq0EBQfA5BrSiN1JTZTB64L1IiVrUo8A3RUAtRPljpju/YYSxlAS1Afl2MjgErKh9HJAcN
t67mIOhIU++6HMPEsFvQ0HSxMebl8Q3VEmyi6oojGwDf7Ng0uzDYzySMCgqOCMDWb6Hu6IiDJiYh
u/oWfL4qVZdUeTNB5sTv5ErUzSmVjxoA2FiEz3e51qlpLQl9h0cwNK6l2hyPc+kPpghuejbc/ONp
zRusTegWTCzBx+gv2lusmNDaEuHT5QvkR4mf57a5OZU/SMyFnNpsqEcAUuVVmkzQn1ddGBgy53Rl
SqeK5wy8zz+roac+qdPECUP5TPCZeWwCdQt3akA+F6/hNLCPMAXyf2wcy+AUmlaf25FQSVd/Pgc/
4BS1+cERe5DuOhr3eWM3hDvTpL8tQPXWstKXCFjwl1yj2vvByz+vZa7/jTiRQ+Hpfjlcc8bFUeCJ
tp186MDiyI3HVAeZyfjLkJkKm5cXoVAF3Ito+MDfHv82+Krlxq/5WaMH50hESfNXOIhHoa9zrZka
PCJE1rEnyWQgtPYB/2zKKiaQwFI8qUk1L1Va3CEDgOjdTf4JrL4nB3Qu2hck5pn0gKurRQy+x+oJ
yh4AOBTBkgqmHd+JJmvml6jJjEkoSXiI8vGL9uTJ+TGjNMIbBtCDwc5Yd5ezUwGqbJmr3Uu0SQ4y
frCoQ3x88CyvnD+uqmePtfyOGYBBnUWDrU/VZwxrFsGaChuDRCbkBK1K7RlmwpAQ52DYb1vBvBUi
HmUoXiLUshITkKpp1t7F9ZUUCMsDMFjaWVId/jxSzt47KiBxGkPOYqFHMPlaOCxNgFbAUaREVtqX
cv4O0I40gJf0MrzjBIzXVNRSV3jsVIWo0kiCk5qSmO39urb1zGbbDGiJnQBLMutt8xEMivlYa4U+
a+rKVMw5XHKiopbu0TdnhxgYrFtUhSmJSVDut9fnC0p/uIc1d8hedpKfXAMtP9euEIGveGlZvZnZ
ctLyH3Oa9LjAtYHFvxaQ26ohWvr72zq3xhIyBlqGVX9Wyn7jLsmyoYbRbva28B0JYBCyf2G3aUeU
VDm0osgIxnn1n/Ce+r9SJBcdAL99w1F02fK7lurPtRnLQ416HNdzr5Ji47QkUi++w5Q7d3rNJm7a
cfccmiG13DnOniUIDphZVKKn3p90XOn8jbJ3ghl2uXRV3ubOQld85gLXVEizG/8d90NzTkkFtUGG
2dKKKwe47Wl7VgqDwDdXix7UGMf9b3fW0u2pgByA9dMsf5+j1WXf88lMv0FJ80n+70ExNGkN/oSE
lMt3p+R6gLy+bJbE0FltLr+L5rNVfq+f/sbt2sOPgQPOq5rQp+tduV+ROJ4vvQWO3ASDIKcZCLqG
FXX6DY5m0I8g8wT8b7uLVyBfk9djWhWuRmnG1Uvigua71j6/HvZXfJCaE+eCwVxIRdzL39RaHgKE
cS3oR9TqTkLtq9BC+5wZujUBQYYn3f1c7VwGACjLlgGaGCtcQe0+xzK7MIT5nNX93CSK7epBJjR9
PLuQEtZHRKpvxSEhLmUTausrHSN9qoDqq7Nyqxcye67a9WhrMy6djhkjvs4HHBAgACYEJQhPvJVC
Y104U4yZj/AhXcQE3Gm68zA2GgmXVzVNCsD8udeC8alp89YaZ93vkklVelxmnzVTsYQGyH4Ztn9M
fQAnWE0r2PEMsQS5icytq1ULbgNI4XXuR/arAFYayDwwePAhXpByuYeIYhcy5hfsXnKl05EpdYV5
RPk3V6lSCkXYCusSlY/UPDrs8wWjGWr720ldlwE7PFk+rtW2r2dtURSxW+cjw+OP1PhH74Uivi3R
MQTGC5RJp3yBtfSi2Q7c+MB9zUqS6JkjOSUdX+Fouhu0wepFN7X8vEO/uAQTzjHuLVqQWPVYnHpQ
ewa6ozzQ3LB2d0Z5o+NL3hKj34s06zjysepJHHIN02Nuef+QLJ79M4JAB8nAzb1edVX++OsMT0xF
dNVtcHePiLlVfUGNWgOJ+XRt+YB6l+1I/1cRu+TOJxf8r61j8fsGq4Xls3KgpJrJY2js587fm9TQ
SQVcRUcK8BSmH7k8tZU6SXEyI6L2y3UMj3GpTFxrbby4iDdaVfQ9ay56tK83NBHck1AG6yNY9Kbf
w7mICeZxtxV376jOr6FhqeDd6BIV2QF5HHYLxidlzF6JNVqqJrR7ryDkRLD3QFJJ40znTWDrn9q/
S6nyea5Z1KdyfZU1tkhb6Z2c0YzC+dSyvu26cmclwygFgFmsPQqBBxZHV2JV48vO5X/l6jD5kR9W
B65m5tUxbONTRAVWGtpnDj8WIxB9rKeumUCYsrfM5J4BHbQrvIpaQorMUOtB89RMWsaOrFBycMth
poA0zEIysyG0l4cOXkduwz6QL64lkQ+yqOafWlM8+z/a50g8WBKRx3kn3zeGkHlqqqelW1bnQ3vE
xnWE8jTiIwfz1hCEPEebI1wJi+RSpT4nnkrx8Q8pCxEhV9mJf7cCipFsZyGVzwOQohXi1e0zqKXl
mmbmHi91hbhl5NSuY8WrExzg0bEWGZjWAVt+8QIofhgAnp3enA1wJWO7+l7RJGAJdkDB1+aKvuKA
3GQJY2nuO7iVJ0wvVCRGbZGyx6Fpc0rrOoW1V5mxjkmuje79CbvZD5j95JW1NB4fpPphaOeLBZbU
x0OZ5QY70Vwh14vy4d6Z7Rcuo9jiINFoYF1mYRo2zWXttAxM6kNmwnHTCko1bUKtKRSXDlBVAtP7
DFQC3Qs0TgcfXnUEEQ9EykfFeo2OYfKDU6+ySBQCUzqjTnlS/Ej26iion24FjNxketNx+baBgffL
pL5WQiZ0LQIk9gtEToi/QKlGeNp835HX6tKD0dkNjrh3+eODSbMdymgLMPt198HDJQmOuFV1llHS
mahbrmaI4nU58053eN5mI2HT+60dMwhhh9rtDEPzZSRteQrZ1ytmH6azbgvrl1iEUva0kTzleKxI
lJ1N+z3YfNShkYPJvCh38ULCy4AZGWToY2jSceSR8B9NUpPcdBCGR9aRyYPycX3lXrVLmWN517Lj
DkDCu0O7dCMNDw7jzvSpOpiHhf5SXS3pq/PvF1TbTBawU5kma5nnyDqDf/RMHkHFO9Zz4KQ2TZ8G
y+SQ7MfkrBx+lTt710hA46RDjwQZ4AfFO8EpwTObeg3wt7aK1Nk1mRe0b325fL4Quyc1VfKGEqwn
68ZV0v2YoN/ujCLk/nG6le3NCfeiot0HQd/bPCrklEBH+7mzVZBcJWbb2Nz7+KwAQflg6/9SZ8Hd
Jg2gJmKc1cBhk6av6ZOHndRarWBEhlciKQcwWkh02OuRZF2Vmzb8bBnSM+MUcDyDdVHtnnSG7L66
sZHh9c4+sDCX7fB1AG8EnqQEQHWug209BKd3EoZMa2wQvSMXrpZFkF7EWt3yi0MaAAgPV1z3bFC+
vSbh+qaPEoQc2JeJODMAhf9qq8o4u7jDsBpyzUo7DAAfxPwwPGtMpR5OhxCNJkXWlkUCBmp80F06
EfA8aOfDo+mls/jtVpIzNzcBjw4dCzTJv2/TaOWuaonF1mA/m56JYmp+wkDUE58rJx5+XNFIcnv+
A2GMxy8iXBIhWQzhOv80GgLIN8L6M7EbYqnRit0DJ5b+AidmcmSjk6Xcb3c1GmyyjmYywHWC1MJV
D9mcCJ0YvTMsSwCD8Hw7A8oryzdNLNVufzG7yyYmu2/kftqMNBHHs/G9B0seKbndgg/AePtn8PuH
BlmJV432MBXE1IOYI2j0Uh6fWNqu1TVD/0h4ODc6tHNeR8BOxu4arvTQxuJas002SjJHKR8O6l9r
2SFHxoFt544ebSv0HoL7qnqHPlqKlNS0RGmghv7q+Alu3Wl8T9MZhe8Gpy0n+u6fB1s5qtP+2cBH
5NQZi5ig07A8LflGnO9FbuFSgj2Xc/FcJ3qUU40iHMgcvlwk3uip5yBYsXGS6LDZ3J/V4DlOz2lf
QFn0qxK01wJxFPlkPYii5BDXREnB3l4xQ4LJyckJKZzdH1xqhbKpkIRFLCYHEhAArIEYHHVpUK/5
cBJSWoDWAd3JT8KRmmOeQ3+qhABc3hwO06bPOBx7MjnaA86U5vK9cq6tJrFfo6n4YYZ+PJP3Cx3v
BOwCJ8uwfJh1uAif5O1KNI/GpHmnIz4b1SRFZhWQ2y74u7f9zRML6qQ/ice13OBnmXh/3wNmumKZ
FJarKLPfID0aweVzi0PfXxQbYJizHDSgYA+JduvpU3rMby45wxpRrXCZHJHrHLE+WwGXOxNfqFcS
q4P7NywIAl6mtCG7z5c6hgYxGthOuk07VCmwRR8yXU4rldlkCBI91cafNtLkmLGfEsVU/AifO7Fz
IYd/seOG3Rl4EShclPgDuQ9442XGI66a99PLmVY3RUozJRRvoiK3PLkE4OodFFMc4KV6xwiJjkdE
53VWNjwn7vlA7CoX9frjFAxuIT4/19e8vdtxZ/kKxa1O3g3jCtXcvyLJIrJR9a7P6BzIKtsuOt5S
3Fm+JtJfEz7kpEMrQ8OOnM3bdit+PjN0AXv/1dYx9Ar7w/YJk4TXCJKCqOdRStifD2YALoTaP/wZ
Uj9SaYZNLHl//8ShgPnR7yHZHdXn58z032i4hHDUoCznbjX3b2oX/vxLi0ADHnAATw7rwdHyTERz
NnDMs7chEQ+vdgABa+rEAkKt+NjM+xyVnHYDhuHgq2YWRDgW11Cxd1rsn4TnX60murzBUyve7F+0
bxRUqCcGC/kDLnWLwvEHWs7RQ7i4AeXFgqUMBz71BKmt2fJmCEyE6fPHykHHfLo7JBm9mo7/f90H
UNDlhrPXG8h8w77gcyxxWzGvHxHrPKaE63fEHpWeOWvj33W8qWoPfVhO7LHvJ+FgnLi3XS6BCWMi
m7WWhHONhehVh12y+WYCG6yfgh8A3nFZuIt6mj0GdZcg4m7bR3N7ZsoaXyFgx4ghV2l0yif96kAR
PpP2HrMB43/MSZUMZT7Tx5Dd/fy7BK0N7IT+m20nQPiXB6ecU97PaSQAU+GOYsNH/zeZ6TFwTES2
bsHvtMbjCbbExG+glDk6Y4OB4bKvZq9fdzD48Olvh9Wxqz9OcZ6zVbloWVszRYm5aU/IXLdJK9bh
lCTyNBrImfhtYJb/HRU1CNv3msZRO3i8hHiJl+iR7tK/6s6GYnqFmUoVJSBaYpVJu86dnu7UT1JQ
JSqeVp3u2yexRZ26jjOxYPzUMG3clXpt1LmNjFyyvGcjW7Ikh4q11KYXBi0YFr/bCadzotQmWoew
ELQmWAHUDTiA2Fn7V8qeG34sr5dQXBFko9duz4TaY8GcYiCinYKc77LfnJGgWMtucvmB5tzNB03o
xofyq4t5NpjJlPLlCH6Les4/P2/pUkSIlw7wCXrgbeXlxx8pVBOjLAELTspeOJNtVuC+avH4DDzP
uHahn/795hzBJRH+Gx7pkJbLZaAT8x6kagkFmmViy/vWb80KkONn74oE3bSv+bTq/n7bAIyFsy+w
RzxJMKtq43dGDzSvyXLDUkB+1dhxQk3xjjlTzExOEs9pkMm19ljLXDvNwru/gETGEpBczZJi2aar
Hwh5sVvFcyydO+gaFNPVYPbbK+ecHezquDGicEnmCKTuZ7g8k8OjeMkSmT4RmJuaMYchNoXi8oqa
GQo/z4OSKpQdEz+BpCaHGt5QPirnTwwE0Rkadhx74dqQ/jdjuu4xcKcwOe+KstA709Lfp+8RBqgV
UeAn6w4DU94tPxwNQ+52Bf7yKdLqIfA1tCQUH33SSaxhi/qhuOhL/3XO5iudIGyoPgW+bO6FBKvl
WG0m0ECSACbGvSM8ZsOaPl+5nV2cl44INvU2bRU8GG+bFwiyXKqk1MCAeMnseejMEVpSuqfkPmhj
8v+XT+D/W3Sif1nX6v66YWxmbkmEn++CZ3qweZ2SqTzzVjBW26IWPztmrTzS49Vk8cqlHpY2jD3T
DC8KN507KT1/WzlC1GOkM3PI/wQFkiTvS4tLlx6PpEgjDhn9EVPaKmEO0kkFLrwIokhv1XtP1Nnx
4GOM7bH4ZmyAu7i97zudRCNZUnIYiSRW7xtcE6YtkVuHLyCl/bUPnxEA2kb7ol8HxmRfMgQirkMb
1lr+B14d3xGpokFTHHTUzFh2FagFLOYuJrjp6SyQge+pIrP3JmsxC3mjOsTq8DuGkztqyNKkyyXR
hvPsO8ObYrbgBBnSnAYxMuoFdAB+LsBgD/oxkpgbBg72Jmx20AUJNQ3v3F/I+JFjgtfQ7DwolAD3
9W53IDGmczTFKg0juUwL1mz6XNrUTErRTCKSNezWQhS2SYNls9b4cE+s6nKggnuCIiSDGoQWQz6h
BM8WNndH8McD7Do359SaJ7WcUWe2K2mIoYEdZEG8gduaaAm7m/R0/RJzWbb3VHIxnEsENKe9XcJH
O6RLGCL0eD+KH9nLFZrpn1VfcoJx7o0zHaNPDkgaOx/kgOGbO/srlORchFYnsRKBCBMofp3zzAuy
QqLmO2+Gev2jT12ZmBOwEuLcTHxPhdw9wG1gkuwn5l3Ayr74dfZEh217aPwtF6Y1XR754gNQ/Qbl
JCyUw7+If1csdOy5j+OV1moum2nXwS3xZXFRjxEgFaaU7A1SumCCY2oyYaaps8LWh0AjntMpMHCJ
IOiBddrCOlbRQ3exEXp4L8hClEe67YZEQ3+XbLQXTbLvf8PlSA3YxjiZDOjHLvQxn8PpdfAl+atl
8jjg/A1CxyreDtjTuN8TqUTAHt/7oUAcqaIJOxFOF/lH2aIahTYeX/DaHQcqcdx0sYMWrzIKirqo
J3yEbhomvjfl81yAQxO+wWEchPp+MfHURNzcvPOEhCZK2Mm+3ZJOswOc+BetdovYtTJ6VLKtU4P9
gpac1YWx7iSwfsm2hghKlcBsCXTekSDQ3uQpoSX9sC4P+Yu1Z11sLnCTKo6Cy1x66sqw5y9oW1He
obLJNqVq4zRioChn6ZB3nYwjLyb9Zycb82cUqpRPbE726wj+kzDYGrWJsuRdh0vvILI+k/AI2Kyl
HOsFXFlrjeI3iRyWzNmq+lvsElLTPX3KU/FnUir0Jy7fqetlInFjLqpz8w6DT0I9qAoBh2bJiuQe
izrQkb6A4Fj5uf0LeYhLFcRGgzBxprcnpd438qjonS/iMRKJb4+E4GgUT4GP5otYLSDCde+7OF6L
m5/SxfGBb3CkkjzDmdBetBakwGfkR0JpUyQ/pFoFycOPpt8I0/GDYLdJL1JG/t1n3NgYXSIIcsZ/
aeQWrX+gD9e83/rECiopHVlZWrapryv6WZ2k8tttlJkeeZ6tIMkxDQ7nsphT5Qf36muUntq1pNtD
pYObLMimE6B4PrHEFsJbr+C0xqC3DZtOyjrVmAZu6AnV5l5uXRB/sIVs68S7Lrw5ssCqyrf3VrvY
G88aOzvoykR0CnhLBegaPXVcZjn+UxCFpP2jDZaYKzC32SNAAv+3ExSlZqAC06q3lY9zE7Mnkze6
7EMEQARiBGGFCx3QA3x4NCtTn1q/ApjOCCYXaxIpW8DCXAu+O9DY5ZLxwCcx8SwezHDg3bx0EfkM
iaWbrKNmZ6eej3RqH91SUhA4s1XYvWSfy7uI9E24EctrKilsheT4Pw8vC1xMg4NGWT3LhwMll88U
YAVzNVo1apvfIY2xpfPQjSpBdmTjBv1sX6/ACHhwOSw9lNyajMLtNbsY/Go+XC0us2TGU0KeSRyw
sU104foOYCqYFlcmHh40CieFUWg68RuH5QylIsL8WynaohF2Q8UbPYnBVnJmuUgT6RJgBr0DSwIF
IFISyL1ubhVicp3N1hPhL+TOkqixW0AYsF5Crn5SgQT2tOQKFG7O0zjONAyoGUp7UL9qLG7P5yRD
fD5CVOW0FEulJAf3s/YFAPerOtAJEVL7qgFLass4j/O2EPBPXcQk0QYQ3tyXmfz4nU2qe7H+9hcB
TPW3UZnZZ8m3Qdya1XaqOxoG1V+4zgU3OhkM9jdAnvvG3QwiiBO3AzvnzUFmqUOmQSRwbqJwnQUj
hX16Z7HNfG3B0FBg5aUfXB20nSEJbDOBZDjKsvucAnfsQvWMtqqVIHXvmgrAtgPJyC/QMqAckpK4
TNfAswpLif13oIVF/8C9zRUyOP0JUOctuqW+v3zqu43hauqD5+bIykeCpaODdV3IFG3ol1z4y7h0
FZ1iSV0w+sU69xEiIpL+CSEaTmNtinVcVyZyB7TVogSq4pEb+ZAe14YAJ92QeKx9KZ6NQjYmfn3u
Ok8xF2eao3ZQDvM45R2umrAx7ujzxIJahMvwTdFg3NxDdesO2WwhFDLvId+7o1xBHCWshyXHXfjT
kqf+E3S6SM/RRRGUhQr7zKYZ7y3/0eIeMIQn/q1ZhzH1PCAxNFuDfAtZxaryOk1VjG60d2rzmZN1
MZJNIISelTfuDCi7Vz0yO05Ebsb2bp3nqcn+n91SiqriGnbyYCKFN9LmxvSc9YfcVJUH6sBjWBTZ
t4UOtKQ3/3kpFYqsrWI7aDDa9rD7fpBxAk6J5OSYog5u7K1k6eJiJpxQd+YsyMRQ4PEv9RheXRuj
MekpsJcoGToWDQCqZDVs1qoaUwT65zhb1W+7LW9nvvCDPK9A9Io1a/2KkyBL6Y+xPiPPatIrfTrb
Lu0pa6Lhx44jY9sW/uRwKvHKyzQEtS1ArKz7qTqnY3g6rXTaTaDF5Gv6xSBkYCh6CeOqC6XmrP3Q
28lW3abkJvjtd8A8BLrxky3Of5tz/dxSvO0N0K0Rm073sj71gV6rZw60mu9jguBi5bYy5N949I2H
0FGUwv2RsVlLTwkBUs04HVihrX9wL14psQr9SIc5BEK5hvY30nw+6Us2lAVGb72E0Gjr1Yyrcsv1
YzvkZJoMOQPwm3KVRRZdQNNiZ0rtaE+Iu7q20Rc1FU/7g3GVisVTdfB3QgF+yCe/pFkfqfzYmCzV
/sxR0Tv8AcVpT2D9cEQedNdhqC8In0iiyTVQQ2lyWCgrz5w+nKDPxFir/C4bTzV1ktS5lkEtTArz
oLEu4yhQIWqqmT5P7Ku5VG7xRjiRWlMLEoGocAUu787kbc66GyevEFNSNbb959hh9eOqMDBY743N
mSRLavxpnNxQ3tp90yEUJqVX6kYTAL89kHwSUlYADX2XqNlwOsKh1NZlJMIeLVVVIG14nt8AS908
GKNdYwu6wmDPhF/ySuTkw2+A3C5yexIF19sIAhMq5HI417JW6HTKI1yy1g+4Vpa0iCHCARnE091E
tlYfjW1Tdxaye1wWxMyzxmpgta7RlI3QyTLx/Q/wsBNK8k4gm/OZtWYyeAw6/t7s3LZ2yoM7XIjz
lJSpWjbBHk1LrTdVs0yHLVyDvAlV84T5OXuLJEx99Zwe2+koDMjffGCog0EztkjZADuafoTRfqBs
ngPwIQJRrLNGkWRe5RkyRud4E/3+Dmg6uP5CMZgijCm0E0isgZSwElpZn6+DqvY8sdL2vJGuAJPj
5/JqvwkgzKG8w/pxQVRiGqndg6cmRfO32F05KjZhYkcv0e/drLmxxmjxCHEag+q5dNXUQ4eR2fUY
M0918YR8ykpr9r2imsdxPcVCSpxoeOSswVfM3ZRuHCSrsMXnnLLNhrkJf4TvBAElQN8Kjt64xL1p
bK0B2n2RCSHkTW2wPzVRDfoHA0+yPz6AEPAxkaj7A/5T5z5lkoeYKHJdk9BcFz+kwTUPGJkYv9K/
vCDHMs4y0CMbb7FVbCXXqTJHjRR9FTIXPdadA5E78uehg7ES3Zo1eRQjNBiuSGytM0uBKP5V57gO
ngz4caa2iMzGDxsqU+GKa7nSRBMSmEyNA/mQGOoyS4hMKXAWjr80WglEpKRV3MkV2j0GN8oRd99g
JGkjuhOZuTZQieVUgwKBlCTgOVmcEkfICFgCdeYwsmaotDtp/OH8cgR/FvuCPb/GnbIQKZwv3eMo
hrnPyQWQyNix+IdosgJcIPQxMXixkeyXlZkZivPhLAJznhUc5zuGmI32dv94PhbwqvGpFB8a3Vk2
36ENpGkvYVlmwuBVYrV643x11G7pi5rpQzfBnPnOzBgiL5PH6vGegMnX7bV7XrZ1Svxt0pczuQvT
AKxDp+gpnNVNeOO3tSMPkbGvdjQTLhH0dfGn9CmPqJpRg+4teZ9iyw2jyYq7IqveCwZEqQe63zmE
8zXADgNjIbJ7GUBBBkPCSq64wMyQiM1b2bR6llk67s+Eaa6wZGJ1OrBpfbhU5WMXpk9Z5TKTBUmZ
J5oYhPFfePVg1Zgob0uGOqN46GV2aFTBimqYhlVcWGs54HBhPk2qR6HYbPULSJ7907uhMKIJccvn
BYEv/CcL+fX9dGJx+vpyiCc/VBpSpiCd+5qKGtjdzs2MCsTfY6VZ9NOTmPurYMkS6WZdy5cFObCM
mC6n7jzihYjT6E6/yPewaWIBzYOWecAUsGlQ9JHmvNkSFZIP9lEKsUtMOM51l8lA2Mgnmp4hkQNj
cv3N6oMPYsU0RoFoynrkFG4p62LF+mMrvQKVL4fPDe3szijHQRJTEG9cAaQwWIkrcGcN88gHFLAn
OUEc+GKFvnxVyQhH8CKX+RIY+0j25htOYaIHnjcK9Mjgk3S4umuErjt8JlExfab3gOs0ON59deNz
YuXWXqjyW75IP1t/Qkgko0Xuy6/0jgUGQTejbhGN3OaErckRcvC6Oo5RvNwWTAU+0d5n5k9A56zq
IJv7EHBB+Vp6VVJg8PHjz0BzwVeSPg4VzcFmBPnL26q6OEo2PLCATZeMnFuXhYSfuhAx999TNsBf
kn3Z47Tggy87ZizJvjfQTttWkWaUsbEwKWF4+6SSeT/yUHcnPt1ZUZZe1Hr716JynZTBunFch+S1
RxiIAWTGZj80FYvr3OZd0s5dzHRAnNvyA0pXGyOIE34917pGMtBWOxbedupU8//rOCv5FGDInLF+
HfP5v2VQJusTrO7ADlSqaQCAIOxj7P/9uKyrvGZKKJiMbLags4kG9CEGUVuGUmgDaoN4FRKz8J42
kQyqjwPf3z/ruorVKq69CShyPV7OIb7mC/8hfeB2ZbYDOsoBkWoUupAO2/d64oFJoEND4btu6rZq
Fjp3uiRK5+aX9hmoSAUP3odOED0lglM2zvIyW0tCveDRcx7wRcNUoYto8oqpRZ+o5F1W3vNfGrpU
7BK3aZOqmT2XqdiQAAh0iYwYgRLQhCM5LWHiBnp7Tmqpyxr2oiA8ubY9ClKze52+I9UCKL6RKhEE
BmjJLg5ZA8GhwQqbtcJMR0+WZ5Jpf5IfwajXe4m/zUZ6/VcCpaxq7mOTbJdZApl6JCa1IvmltTP7
J6KFgtDXI3ixTK+Hm5ctngu4KvXWl0vQT9AeTX3haPylGumMZ0/FjEOQTKVgmQvNjHKNYYQAKuBZ
LnAsEkUSbX5V5NwACBPvBBqhCRcUDUCVSvQnyc28v3LoerQxGLY4Mnolz3iiOJr/0+QsGqntWqoN
MxCTNjVXGygHmOe2O1VgRFo6pFRKyREmJYP2S/IxUgEiOXOV6SdcT7yGanote6bljxXqB98bscWe
PPJe6dFiUd4Gsl+DdgaeV3/nTMowp6OyU3OAyEtbxuNSzKHa2NZl4d7JnGdblQJcWlte91XYDexT
TWrtjYsmNdbiL5/iRhnMr5uOI/tGmghELSaNutCjg/+a3g5k+5bG9t/bnPqQtx24j8fVgPNVQz8t
5zQlWwlajAa/StzgLRfL9AUjkSrNuxehZODQ49nAVD6JZm+/OOhsRWdspXa/MWVTMNuwiqnG03i5
u4bE41zGzPhsv+Fv+jfc4kYKvMCGqTdhhEHy3bBTwlYysJ21fWcFVGhzGxn66mP7tfO009g7YtCr
AcrEFHEQOpmFN6aAT88wDGTJ4DaLYtCq/TYUGjOKyRV/fFamrmBYixYLcDo6bYIhWWuELPCAd0vf
INveLTR4WJV6Ul6OGpItZtP8EgFlGhPLyTEwKFuACKx3fQ+CIlgC5hEuGbkndWP0UQRUcZsY+drU
kX0t33bbNr6JQdoabU696k88NIUSH9EKyhv6hxledX0F86grEnWezg0VRtz8Bj167uyuz5szxTiQ
9L0vTDA90uOom9SrJBqg/yBOlagRxCQQeq3oSziglbGkMAC6iYeVI7/q1j39l6Gw5JUM/9PgCJ0y
uPwC21St0hKko2H0w94NFnjsfkGXWQOuNF+uYARl6DdIrSt+t/WrovHLV7BGtvlyZtBRrZQ4VzTk
qy+DiieWqDEjtSlqrAsV9IjjdThUKpeHfJck2qztjXJth4sjPr4mEcPJCb6Gkt8dwTUB2kxUew2g
pBCg52wQIr+IRoTq4IWtOWKYrDJzYwysgN4IGhYiwz+HWNBdZQ9Ukl9um/M0Ti48xR0gHaLc9x4P
NncTj8D7ZexLJmN9Rqbgaxogux8Mh7EM+9Env+ZYzJBRKOL8lK/G1JGgJqtMVxXmUG4ZWB384w9v
8dF9OWqQ0Xdt/MkqHIHuHCnuzDcocLK+ozuWYVUPjmR9lUy7Y3OVkRxHgUdIxnyR385AR/hghRAj
Spt/5uyWOYjURzM9zMkE7bG85q5nKVfjtrhRYjgSsSR46e4E1fxR7xhsyVjLXIPA9M5dwhFthK73
o7UuLh46fWAQv5/E7UqaQ0Pr0pFACF9TPc/1BO3QPkfo/rKQRc/3AlBSGH1gBQaHIkWgYtoYjyZi
acUvrcug1sQZF6Q1OBrYHhFLRIpSgE/2h90WjavvXFLzhxrVuPDtXj3pOQSe83Mbgb9dYeUkVQpl
MOzAIxPZnuSzksKxoeWuvTcjmWlzsb9wBoBh046BYKMrKXOY1GS2rOqQ3epURWY/BYPeQ2KuYSgX
BGZqOPChTuhc7A3kp5j5VPPyhGbv1oiWOuIzSjNTCOTnF/7UOhXiue2BDYFNIUw4nwnTiO3p4M17
yP5hSSDPMbgdzkM4lkZeaT5lAnzmui0uQSexz0LaqzHAh/RlPKJRQEekwj91h22wp/ylMouHgErV
+Hj63X1vwybfis/Xo0QyllZ5/zTJIhdyAkZmGl8vK8XF4DKdZeN9UiIdz4c7VoHZI2SOvZGjrJTf
RwKHxgP49pW4oMDTU8B9S4Xj1I2OIlnQejAMWVmf3bclpT9Pzs+gUzBu84tcoLuh2ZLEVA3m1NRp
9C2WUuZNjT04x6TNO42m+2og/yz4p4pBH28AKpJwmWDtUrl/ogQaElWW9qnoq9XiLc4pIlDNsRZB
BXK5sKwLWua0y7hHb03OsFfSDVC/k2k9b5vfexMp3fLY9mQZIegFM0K4SPCCIOlqSYdZGY31Mdax
0LX65K0lNrecjvbuK8VUbSE276Y++x1Nd5046vxem0SyCtHjuvsqJx1t3uzzlu01lMlcCy/5zBUU
gu697y1Ujuv4QaPNeeWDcHToRjmmhMsieq8RS5l+rxK2xRUFRzN7Zhs51gPK0Ix03NOiT9tlkLFY
I42HrqZlYhxOVLAxftAwBWSe1D+xzQXGTOApuQuGyBo6ZKn3ayao4vZLq/oVTW5pGCWJGxWVyBhB
uE7OM5MdzqTEtB87Z/7ZzDZGgWDq1fpJLD/dGbaawlUa0qfEJ1LmmemY6FnnguWn5QIi73XF5sp6
mf702iSEgmjV93n2CY2OsNIW5YZk4VGAyCrhLaptgVsFZjW/IKI7aq6vzvpAzn3aUQXrjl5M+gQH
JaGhADSVvJdkYTBK5NIo8OwzmDmmDNpqA8KJ+MS2HVf73SeIzcBHHpffmRmEDvr9ZZoFPvUNH3WJ
q81ZlIowRJuJ/LtMx3yfm7kYPDcKn/gNbgyfi9f0rKTzjrr3ZvZk0R3Hb2tArmvsJTCY+0OBoFDU
ia5xt5147VymwBHOCZhrDhXChAHtYOxkv1Bm9W27g1WIueLX1M0YI0q9IMOdTaPVfC62Joxy+/Fj
JEbQ4FoujR/Q2z+IQ/Vd1xNJSy5dBxWGPE9NIFvIQ7eq62ICBs8LJM1u6DA/2H7KN7Y/TiVsGsAX
nB5+ObCq0Z0gVR7fW8Qca/d0kYpNPK/cBwt8EFoR6csQZFOkRd4yrClGtMXNJtlwB/m/vOtzN2Rr
FLO93F8/SWgV/eiv6JC4yiDQqxrym0kBAtHus2IUfDpVRyLMQ3ipM1b/WCdikQODnmAwtjB/VXzD
mlzhgL9x1s5XI6ZuL+9gO61fCZFN8IaKsocG11PH241MUfDmC2aievX9SWDdqRuncljhnFHrIGsF
I6PwKD2OBOtFOY0WLiMbHHriSPU56CDFCgYOwG/yJ9IWB3XAPmiikljFQzVKB4WN4CJ33Jb7AX3x
bmE6qOkc7/WcsYCIOZXDh46/Ppflx0abgtUVrMjfmDK4/cKCyynmIbrvZ+vVJrGYyzg5/3Kj8lX5
cXsbmqmrVFtYn6XiO0A822030GRDiJWfftGj1CCa8nJdwiu360RViL2r52Or2EXyv0DtySiVMh/k
n7LLlCrRxyxImZDpA1OaOMqCr6ccCgR24o/cD/rUnZyGpkKiF6kE7n6Fz7Tem1AqOIUmdFK57qF1
NLQ/UxhChnLWSTUDS1S/jX9SbwURnsgfU8f1ptLDXqgTb/2jLz3x8VfHrCqNz6h0uVxm7ntF9m8z
fj+q/C0Kfq7rIPiLYkvRcRFcPbdUfKK2APPuc33/Rf7BM1740wIqvcWUofe6a+NrWL6k55/wFXf3
LULvpcJ2psUV0ZYE2KZipGuRtr/jv8BPPuzHV4JdF0B1+ILs1fMV5lKNAv5mxjK3lnvsAtNke2y2
9kH24MdO3keyckZcS3mLLG3ANES2hoEyZF1DQI1A87Y5ra94tUUTsQ4h29zu0CngGAm63K10hCu4
U7JHpXpo5iPHXOpd0fiY/3FQjIY0S2ckcOOJywSpZ9a6oHd5wAN7uu4yra4FSQpVJdO88Ql+CAee
Fm1zOOplRjo68VZGGTK0ZgWjA4E7VeB/J2DC4YzwRcDyquo32Cm/heScZPOZmcKT6MUcK8ori70t
mwVAOwAfBGeeAKBpYvVarbR90jzN5Gq9c53zGv4VQG1aHp1JvAUttUTJc++/Er/+gTax7yyx3bzx
BuoVdJq5WJd5SASx9aHLlksSgpRrBlnL18OK1jFEutBKHdHnZmevNceqCy4c2b0JLzkB+a1ewxz3
Cv1mcinppMr5PKS2z4H/wSoGXQV+73XtY+bynqBD40AZPFVh+45eEHbDX5qmhwsDvK7W47rk7vE4
11HpEXA1beaDmkoHQRDNxsuEsWVUxvh32DP6UWxpbtNL6HQwk/vo1jjucI5VjG8IPHQmMLJp00oa
4F4T62awoA0knRLeBT1xx/qv1I8UJOYZA/bFvSAXOQUQB0B3o62EUXRqO63f1Wu89YlkGt0V+nKW
tGq9oacPsPC0WsBagAouevBvL+iWwuPhaE/tWrHYPWRV0X/UELwg8FkgeUzBvhjMooXTPueLYJRO
xG42acX+UIjOXfLlzPAEcP4I1kRp0/mANJwPXTm/V3mooTmb9s9OGGr7tCaDTyWt/JYlnl2mKBKq
CWfunpLWc8vEBBVZ0zI7Uroo/ZOiHrurtxEyvxEH6+iIa9YWjvu5Wifk0bwW5DUKzJX/KhziGLZd
VD4V25VA2MLyU407aKBx/meIMSBD4aIawx0jrqFJPDQoSy/a11NSG5dVvFqHhkBWx1+InXdcZrTW
p8RC5/D1RA7o4oOhwkceVghEiB6DrsJwIoSVcsTy7nZb4mAS+ZOibIAajMptr+Prb/URWGHTOeFG
aQsaOS0jrwqvLjAzP/UsEPdI4TtqJYlK439HrUVMndbxDB/m7bu17elYYuRUPq2bUzYSgLh7s1KV
5Wm4fiR7Cpd9DnDVbFmHN/Rs9/izETkR2i8rDZrRcXZmANbqABgK7Zp97RwfroIJ1tjuKZqaoiuR
1RyIc8okS55De7ZFNKkF87092WATncOW103cHMbHfyfUdvio9s2jQPl/le46Pj+GCZzFhsh0oEox
727uN1ZaXzqK2H1/LjjXr7cG7ozcoDpowDgAwIu9VMt9ADNz/9xjE7sIg3M3NbFoBE4EKK3+e3Oi
h6cJ5NzghVhc1wDA6MGxuw44iUt19GGF7aULu+Oo5PWDB6JYgSTYCIaxz3Guz+6+/sPcD5yCYAnm
l5ko4MQ/CrODpdN2WTwwWRl4FmhBoKfEA7W2FUaZ1EoIG+ZNeDqVhRH6FcwTqSsH3Ib//s3BQ5l8
ULZ+zIZi4JkCZZ2tVswJzsyT/YcbsXfMgEqEkMWe9nUTlu9dQBeoKuocNGLit4Qg64Y5DkxBsDLm
TyOBrMrGsWTZL6KFVyxWpmw5qYuqPpdlpMsa6LVi9gZXqo+tCKbjPKkWWAv2MkpKYHFPpa1xasCz
yatxLKkTVc1cbz+BvyUXe021dyyqsVuBAAwvzLjO25+SkMP/esvZ0Ybx/MNgrnzhY3X15apMVmYF
I/0pH+jYnr/21rFW6nGpLWKsY8xS9O1HTvPzYu0b02JVkz0QoMDtKwEWYAp3YXrQO9BnrgwCiOHj
8cPkOQ8PZefstgyMEvVTc2K9UQtltsOJLnYH5rKY41XxA8eMTkL7gEe0HHaM9GVMK5fSYWiR+gDU
2Ki7pQhDVE22r75r5RAFXmgP4gS0QVHOxPmrHhBRqKIQiof0J5ZJfIaWxW79P3qSdUv4gnFFfQaL
1ThSm7fF8vh0OO+3vb5CccUl0CrOvw/SjHptLVPAiUHb6+0IRjxNkpjS1r4+5JFFg30wIVx0NM+8
0G7VG5GEIKuRHLsULE7/0l68q5vX2/wX5SMHaFRWKe0jqzabWLZtr9M4aFt9b0cXz//mi9121Oqq
+tk/QXsjud798kzSXMXAwCWv55a1NcdO9A3W+GtAAzEbstNsg/zUgXPdCcsMFIfM7LTYIHKTJW3L
mrCZSOSlSnrsItChBaLMMCHfLsmLJHroSbLPX6Uu+iTR4R1DZDFlp3F0hqnMnINz0b3JQTcMpbGk
wW8BWKfwDQwTH3AerLXd6Wbtgy1In0YjLHsK80OTjlntvUE3qvxyMXiz0r0bhxxwhJbiYuHvZzW6
8FBLt4/OGeEqKg56kUsaQLGPidcpvjlVntdCtqbqvu+BJB8YY6QTNip9N11Co3tU+7UiDLj5tEr7
UskVuB1YgPZIgsFRtBzZb7TJ7RzDIXpk5OuIF14GPaDivyAWeCYqaLrEvMk/90Yg4mUfCox8uz0c
EVnUFxiTNWtEFljDw0BHjPVX4+HlQ36mz8lg866YYogdHNtH4ml1eVJnyjU0Q+xb4JQAf2B3ozsW
b680+/e1t10oJ7rEK6IjIXAbP2NPKAnzb7HcdY/oPHQZTcn1qbM7W/8H2/4+fLH183m2VHGw67QA
7kNAmP7Gm55SmEM0L3x8Lfy3671KEd1It1WWSR6a7oZqziSFsGNZ1MK5w250bdZcnHBYdhXD9id7
gSjDNZAZcehKEZUPBCp4WufrxnWwt7VtGK5EImq7TkSW4+5FyBj69BpY9UBn5dJMxyKy1uPNpliI
x784S924scMhjGCJDExJv3+TKtoh89nWs4W/YFzOd8sZfwFm2uZ+oz4+gRfPD97zpQYassRTFAac
KElUFiEVABKFgtZfox92+2DjEgGPEjRF/877Wk4KIttA5p6uIOkCCoFnIgrbx2pxLIe3Rq/yp3+X
9MjbuAoa73SIWuWrBRp/rWENBIjggn+yr/f2h9Jir2HjrIt4GBdZC54cVoee8oAJVVTfGHw5j8P4
SCaNcJABPuPsxFmMdpeD0REJSHep1mJ08XH+MrF3v51dlyyQblnJmqTHNBkQMlbaMBPW142pjd/H
Kavp1AA7flzVtb4ZetJl4OU96iEam2L4uc15YE+Py5j4Fqw1RYqGsWh5ABrA/naArywG4yAkeHui
w/Bs+Q5TTVtVnuvJYpkVseKQd9lOclpcBcZUpflNF684/DP7YDtAaZQOkVJo1CmQ5kkzdbG14r5e
rn5mogKtJncUtZdIvxLsS2e0wBHZD5kEASc6vneSBtMnL3adFocAHUics6ArWYB6kLs1jdxb7aM4
BqzIN9rOv/zaKfx8CnPfF/3Lq1L0lX12TwAEPp4Ztt3QXgfPRpqw6hOi77VCuMqod1OPHvRid3Fv
OWnQkGj0yCe9BW3PYNh0ZiuJOBkgJFWH8qb4cA/7bRCQXWmo1a5QkGj8znvAjf42lj1JCiteGtTw
deEyavz7XQ924ufz5Mv+1/EkxJWL5iJelXdIu/P1M+rA6XBnBjX4h5bxOjRHU2osttKoJgHhNF+N
K00YmVvViZOuMyMYUgnVeJLVS4C6lDNpj7uUV9iVLMwj2hb2MacRCbn8/t37f34VbFBektdcXdKK
4YZzqGxTCZmb7Le3tQPWFO3Aufa9lCuoyHzPx0+n9LzQxDbMIjK32OVoqxN5UWz7H6URUy/R1e0x
/puX35bKlFJ9biKr4UgQrJAiatyjFvuEFvlr7UAiDvaApJGskQ4bjSaHDvl/YE5cWYBucogmvrdw
zX9BmsojJ36pciScWrWrruD+5MNTaG0R/Wp9AQDWXCcIl7sqphVKNGiQHiWoraIyxKWDSaePLKGc
ZOzoUUoBMjTOvBZ7xeAGnGj9mk6GiN8YvJtRG92ClY/KQKowrJ+G8Ll0WVQe2PIv9XTYot6d69Bp
CPoxrtdaJK/mlKqB7KxBxKvvnOvgVCFqhlWZlL1XHr3JTzBSSYbjAdqnSSm8QilIg96NEAO+xdVQ
TU5gszs2VYbMXYRRDM4uqG6UDDTOLB9q6/JSGthy6jAEeRdqyqFLGX0cO05lunw4VTTxPPIB0VRk
QxwwwicltSJh0UffFDTt17GGox2ZaGcL7GedVy6AZuGBZEgv1aE2eYjYlHEvECfef1Qc2PXTC/Yh
fwjaA2jH3OlXwSGd7+FdA36b55kgvroy9P/kluniqos/C00l4LRMQk1tWxPFkVogrHfz2BGWIQPh
TmpbXD7IPNopIAEU6hN0A+F1ymaC/8FXDW691wOsYnWgV8Oup2Ck/BN26cjlGVp6ufgW2p5EKLqb
7Dm73rvcoqqckoAaC6YSQaTmSPjqwYfKnZskou3/p9Kj6EfxH2CCJq9VYYk5OQ83h8CPXKxuZ/yT
K/GPdDyDgSFgih+5/sckdTg6k7hsLP38GDH62yLrgdAkLQRk5Uk+kemYjmwUklFXpCDHMlEI0aqh
BKJe1F1hERUJEMxUgpWSc080OQww2XWjWDtTR2Wd6daIFl7APaS3XgtqPpnPwCTtwj7jHfkkvfx9
zc8/7Ggl52/BSjcwRFOAIgb47yW9qIxC9aXsOEt81nwwwqHrLnOjps/I4b+weK3i9TFdJRDo3Dqx
Np30j+rQnYUeNTxoUyPjGNLy4y84tRGNiUlNmsZZ61ktjFXkBGSae5bH2Xrd7Ijsv20SD+epUQpD
7tnzTxiAelHrSnstt+hBb0TT+2aKoaMbkv27IqdjjH2jmUHFuinpiCEKGseVAZw8VIepCatFZsTy
XkJYlwRafX6a3lDsMY/B9tsqEQew95l2Z9bWsefKBKmxM+Z5RBrdD/uxvsdWhwcAhdzENpb84PIN
smfMYjNcZlJJEatjwZdtdGxH9ifndgEZlskDpb6GRZ/mTO/WUIRLehuetvHEQz78C6f2vePPFJV2
IwbA5xFIO3cUcJNWJWUgNXgdjsV5APLu238hdUtTtsdpasE4JTlTyZ8IZBfk4f2lhPPf7ejCQXh/
YZ2rSyfYWAu2OnWAgLgkHrHwuf7ADl5nlqJlTIRLiFUlSmyOqM7LNq00EdQ+jIeXOBG6bL33YTJ2
9W0uHjQP9uuCS20H892bxs+OgGxqSWvWRC8Hp72Fm8OPQ/5zscMqMDPdVvKlICr7NX4IclTOS6pP
Qyc7yb/0giw682k9qNVrCanpqBP/hSTsmjuZJ06kcretEs0KtAnGcPFt75QDGxgr/bBUqgl4MXAB
jLo05TW/JcXznneBfr4OKsHSPJurpU0RRPN7pJCp1xvcZMxPyTPIpsJx4fxK565j9jjGeRMcqey/
I24iJzeBssEqZNbC22k5lqwR92Nl4q2mhLJzo4BxreKre6/A/CMbXWEjMqkV6hHL/G1vzTVhbnf4
vb5twdshNZ3dTSVdAjhCSM5fpl4DsliaRwlUXscaMCGdvOfmx7yIadXu4l56O9t+3DXO+FZ7pbwb
knjWNt3WOPk2sXESypk4S4ueNnFHjaqZqmRYXbtDHw9MhnWKHUsn0NGxtYhBSo9bFNxvbC52ugCK
tKsj8SrP2JHX04zfcP1YmDK1b8Wxd82UiyHYbGBSuSxKiU/sigtermaG4BkQlAonKJ8EN+5vOSd/
4eg7PnDFMcMKSo+Eg/tIZH/fNpAC+5thd09aWKYFhRogxgsuzkJK4MuN4TcuaUBg3//Qn1dqW5JS
TAw3dT2ZeKTPOBTL2X7ElFKg7PDs/Bs/tyby5YfcIaEec9/ud/KNVoiuBFYV4uLI2T8x2WH71Ksc
bebLhf7YEX0stWDo8jiy07P3aPh4zs6HqJKdTrNG9Xwh3Cx5iK2U6TXTNvBvGvBy4UToaJ/nNz+N
Fx5Vfntf9Vc3ltyqOY4gA0eIxHknDeXVoLUEOFNRrwdfxecXg/DRDpplKk6iKg5z5azbVuDZHxQ9
zAYI2bIRl9wtdDC/w8ia+8JU842HZ1ProsPC5FuvtvxjsvVAZ+gXo7aYOXS4bDChVnVYBnGcY33H
TZUPCTZMwx/z9kpi1Sn+ABso7zBWWWV68wbwZ//+o0fCJBhHm0w6qLgsHEqhlahZnRgpn6606y28
uFCE6gIWeZ5EkKRfNPy/njTenX14RlzXO4ltJWOMWjk/TGn8GB4FX2vpIccUNlxo9HIRBXo5XExy
OSq+uK1NCXokkzWNMKD3spL9AjJYp+Pn9EbPT42msC2B7vBwK8coLGOYjlgWqzoUg/FZXAys4s5A
C7spo/yHMhwoj8pXNrJamwJ/l8ndarMf+IBMptNiBV8bdol0SwL0oTKDHM6gzHFrxJ68KppOGBBN
CtnBuqiyXfyVLdadsn1B21YQ2vsy5a7isbg74gU0vaR3YomVGrAtLnt1KLxw3pzL4jhixVXlOOVG
lJ89t+sRb1ECIvGzBMehZGHI04ME/O7F0nx/LXQU/8X5gVOD1c/aysCDQOvKrpOLedDjyp46/WMH
7j3KpjihT+ucCwJ/Kozg8EOjPqKsDLe9xczKduu5UStJS9FQbIYmq9Ma3Z2e7lAPbxmY5mBCqGPE
pStOCD3MLQeql/ZcTuzY2hLu9Eb1YAtlo43J2+sSXHTxbrfY7MUWiEp+8Yf6OXqyKImMRMLY9myd
azU0g3byoMCWX0BqVVw5Sk+XCotjlNVsPpKFIUV6GeTy+yduFCr0a4Exxc5Kj+/dANlz70ogkNNO
NE2tvfU0AET/i+7wpOKW6tEAWa9AVoBT+d79TKePjxsAuIalWcvaZigJFlShuY2eq8zpHgMWv27v
tkq6Gw6ygOX5jfzwNz+5qRc/LwaOS5m2+yYqrkKHbu7unMJy/tQxQEqgxKMfWc+xKFgodQS+9nv1
VL+Z4lWqEUVBQvew7abkWFkPKC8m+YK2ids2n5GKjXsAkVXtkpU7gX5pWFGuOg+KlPC7+W7PutEl
4V2VvByfJIX9IFpXXamcoGW/lRoZVl7cZFh86k0q9Aophq99dRjkqYRcP4L0DCnR6BrxCr1ilTS/
hNqZe3bdq3w7rhmm14GIa8cjAlF6fzS2/aD2JvMOhkSufbgWLdaNVoxZinf5W0uMFQRSdY4QMoqu
t2Fd/fZcCXoLfQQiLsvrWDlgKlRcU6fxEsHs0aePctOAWAvaoue7MwBH5ZhvCrhJ3b1QEd4UcWFc
Z9LloLYl1vJ5b+M5fqIzjPZzQyVZqr6mugOtJy6pnTkcI2Bkw7QJf+LpZvRpYMm1GFsYq7GG7r8T
R8KvIQMjE0GViE8yM4q0w0F21KUbE5IQuxImUcmF1Fo0WtrNNzbIu4uXCtI+Z+piK020IwmxPDuW
diqQelX0EhI00cT+WSs2U+oMWxZ4MpD4492T4wI/C31Xj6KHzcHilI4WegfBPR3dtwMUlXEPvwYp
q9n3U4Ei0Z8V1FcI7EtvFAg+vTzBJreXhlFhLQ3X9hbN9XCMwvxXkLhYss3LdL0ntO4nlO+xnlOH
1r87tyAu6MrrcB8Gi3KZJemBRqNgUftVs3Kmr4Ceo9zfbjyJSDTgu9nJ4WBcsKbkYT8onOuPbeIo
qEnvJrNcTcLVxCqDdSYA019q7+ft0GmOw56MOBEmY/2GHznYMn1CXlzm6tL2m2K+IRo6vObcujka
Xv6tNzqwUg01TgbNT2IfVqRToF2Ctq6JY3Bo22wbkf3eMHF234iUpTpCV061o/RFP+SFSPAeErxK
hFHcezdQSjBT+k361tYBYc0TH2f9k6vpBuiYMH084E68/NvNkfT2XVfUuSY7Kc8x92s8O0EIUzLF
k+h8VxHg3X82ELgpBDq9rFjJfAlq5m1kt8XdqZraLX4QX2HptE95obF39/yrMcj18dUDmb2mUi4C
gQ0JB+FbSREcFs5rmeCdYJeguWSc28XCvSmLcQLkC8uYNlbWJhWJ+RNp2nDSqOqpPJm6vJUcC0kK
bJpyXkj/ulb/41z/+fJDfgU19v1gIHhMbbVqeMx/D7DpL/1a7GYl3Ti90k2i1d+jq3NsJ7Lkt3VQ
y9Ds4A6DVKLSYpDaBgJVKwoGFZzZoBeFdVYTR6L/YvMqbXN76rO42QsvLnmxYNoVJT4fXsiOAYdj
+s6unhgY1EHdjKKbMneakYjzl7plubL/pRpZD/LeNadF2zUWyE3dBpYApM4aAAmBF/sJIkzmymwx
zxF7ttu/QzgxcxpoGforCrrXJymw0A9wUAtKvWNa0cIlJdA+zRY5jAaWO7atccpRSAHPQzQIZhlv
UiMMIY30oKCWjtc4ivIdZ8v1qEQdg1VpAjqkfmafiFraHCQB/OgCS9TjhUSMY/GNQe5h6lMpmGjD
8TXNmirEtFDl8ijBsm8pvogyE85t38netMHG4UhY+/mKyVcrKPcPK7HryjCG/h/CY4RbzJTv4Akj
VlJuUeGDF0K/4SKviaYcH+ugRwW2mWH29S6J3iFTrpHNLFwk2RlRGY75N4VklybKPtl9nEAuqWVA
unJM29vLCg7sCtt5qEDxL7Idsd0PSiyYtTHWvSYMTXEcBGyGQ/GlUvOAOxvxI/db2wiEEfJ5tN+n
zyTDTW1KvDHX/cKcKI3EH41z+km2NtLtqKv5tQS1fWpdsFPx5Rx8ayLBzA2yVGyrmGzPovOvyuNj
ziejmPu6Yff4unmPkW+7qThYtnpamV1UqjGPK7hTOCEdUymS3XiK80bjtf8EXGa8gQO48xbAqofl
K/HROpaLh333OBk2tGX+D1VjPkTyh6DAua20CMJgEgSobL49q+NbSqkSwp4CEeaWL3d1InXGGLy4
CYZLxNzjO9N/LiJ2GhzwpduDHbz3YZci27CH2YFuvPBHjOw/MHTdXTOhWQojvqQnd4Kuai0wVFty
iOdth08dYQJaZMXYzK4gAs6IYMtMHXvAeLlpk9mSarVZwsvYoEaPCYzOEPVmR+NDdqMHxhQeM82g
vNlj1Ehta6jav0+5ZiBiJOzb+jm0yBQv6mASAgtR1mxdSoJ9yyRRuhYanzfnw/mRAR9adUsMmot+
kZu9dSmnePO9CGTLvyHou8+22klHi+zqeZqcJprdB2d+H1pvAYva+N51T1VVI65oYK4kRZLZTaua
Zm87eUBZRmjv+Wd3jgD3fXc3Pw0/IzW4+TolEGA0kh4pNlbne2tNiNE+fEsZkvnwKFSTllEbf5HC
vr7xlQa5xqwWWihzaRD98Va2xhYIyWUgKDsza4G6FMDThAEIAqGTjJwJoywP5oKvq/X6tHXcGCPG
7HQmEM8xutCZPFRtIRtWYU9wVFt7SW+Ib0d1SO5vxmkugLgVEypoTb+0Tb7HBD3aNB3T2S8Wt7GJ
3n6rtYNkF4+uAdK4tjKk1jnDZS+LfaFj9XjIpGkkdwqU2vT6cRhD7qA60TAGrxS9m2TbFwBnEa1a
gcamvk6t/jLyybuGyZtxh9/G3852a92sIOqLj+Ww7JUJR7zzWyPBc6+6SqvAeu6rWJDPA8ze5k8z
QhzezSqZaxEIg8nZ6OGibUCB5exaNRV8Dko45oxqXUPFYQCn6a8GRi+1qrYevlsgC4bowMS8P95b
6uvWxaHkYr+yXjuX0jVCv5P83TfGIDs8Xm40b9EIIZEHxBtqRr65yXdj6wPduZT8PeIvOZnVJMYC
2HvaFQG6UPaqTC4/8hqmhulIZcssJspgdAn4O6ae+eBhOAEnugk35doIO1BtaQMNR909JtazpCh+
5nzPtLjGW9LZOew+hrgJtafYWiErTOTE6dcc5al/YFHJiOTOsOWvLHiwRrWQy+EL1p1PLU3Tfu6W
EmZYSMTw0N1ocBctQXCQvtn2/PvQtBcyI0+yEwybNIFzaQ+g7dg+FQLpTId2wPMaPPQQo8Wt5Ohs
rdXMnPoMmdqHVkKMxLzywzi7sKYfjp1q4VNiA2ihCnSvE1FSXC4cS7EH9I24/ZeXvw+0lGY5GFcZ
aicMww/0WZlqXrxrnOSGKuI2SzilpqTFnj3d09AvjZwKjd2JiIA/NIwtT1NXIWB5vL97E0FlntEc
CfF3VP45M/e8H+2wnYbPIbU2Pfy8TQ1LEmtMEqwDiw6yMbYzcDNP1x8IpTu4PfG1Yy1FNRF1eyPG
dA48hjRA0kiBN+i3yb1rQBVUoJWK+pzDY4UCaEu3tSiR1gqRPW603vds1KLqTyVNnmxuSjWcKvNu
rSqAkjaSZ+1f4/J+/yWxM9Despzxcfxt1jHO5JuvXDqVnkpGw96mT6gClzxovedvINCswcXWqFJh
lEaxOS2152ntqlCJSENlEsow3B5r37W2j+Zj5/R/SZDdMomX2n0OOeqTqDW77ndHOByQqH0bzlXX
9ak0V1oMb6w55Xi8yAE8D2ovVj/PQ9nC6B8HRoX2+yAInr3hXn+zdRA4+dm92bmNQpkSQ3v+RvvR
XYziPPZzEcJv811wfW0lYZKAJjA8vhuGwwadf6yKTcAseWIw7Swi8jIeYrv4JoDED2Up4EWfwpWS
z362CinRrdBj+OLD6CeCS9e9GUhp0q+qtUmSumFgvJGbPW72WHBKPYj++EvUDkDLg1D3rOBSOzRA
vvJTJQL7dxqLhAVGkfxnYWv4WFwcnt5pHl8jYopt0fSaLHXZn6/1tdoLgeRdL/ZAqpXpRrplc9YK
CbY9R2/265INCZVNOfZWx0FZmDI/zw84n775NzECDta/M7XKM3HFZWcKFa7LfqEW6c2ihoemY5rw
Li0N36brn8w0l//MyERIFPNyBIaTpLkFWUHluD7HF2tdlFj2nlkmyFJlfYdyZW7qA8FrXm2Iz6BB
UJXaGukDDqpUwdo+buVGLBATvns17gjAz86tGSEItMxs8u/8MmJgiVp0SceEq7Ito7a35KvBeAi+
6Voovvfcx8FqB69KeBi06GGlrdhvgJKblvHXLxiCu2iCmaw0w0KD1RavZUpQAdHp2eDoGVQF5CHs
/XkAPju7p+TaqAg8+g1B4Qz29U19+CYhmNW12PPxNn6rkMVv7yq0WuD0e4kTbpuPFlNf5W+EDovo
sxQVhL8EflCUxCsEswDtWVPL/ioCkaSNbsSzzEG15Y/MaXJtcYgNE10lPQbaXlj7mskxwfIeMK/y
Pe3C8f1bDVLNQxJxYydWdivDNpKzYKFlVP7sV03GLH7Khg9ItCJoEuYtiR1IZLyM02hosiC/B7vg
+94vKUr6f/xUf5RnEGkxMQ7Asw46pOVmxbbAz5L0vZum208JTzyeTxjxPF0ztfgY9NtnC7fFfPGs
P6oxiUOFtw+8vOV6FAxj9Kp8rqo/+8EHS2oPTbMU2Q9Qj82bV/4VFeim0rL6oz5wofrUkAGEuc1d
PxR3fEz1+mG0+9vQ4TlkYKp9gGVhKJ9gp07TI1Hd9tAasH35nBW5+KHtS45Yg/78dunWDKtqapfS
fW3IXL1mzneloqStqZTr74PXv6z8BGFU+JYdtD3fdbJKSSn16NgMnx/iPiEpl+801r/G0vjWaXXj
zCPp4wdKXMK23Qf1Hy/OB8u7N+U+Cedpa41WpCNjbvuvWzn9nCtPH5ahGIgZ+oBFU1ZeUXPOOoLT
GrAAFEeEKW7vY6NZdTHhe6vYVnzLG6qbnx1LRCmbxspaY+AjOfZE+wBtckYw0e0j3ibeN2Jzd300
UN558v+99HiXHc4OJX1bDKXS+jTI7hvHBKLifXdkZM5D8IxP7Uq6zmepQfn1qWsVn/2cQcbIOycE
e7Q0PAxgoP5LMd9vK2KLmQdRmLHoA0TbSXy+rRvG9SqHCGVJ/fT5He8qUk6cnTl5UHbWVqcaN8/c
YF57g+Jvbsdi5eYHyeoGhET7EQiSHjiTVEdRUs+xZOThxIlr03vxCaEUOCuTkxQq7kxSij2RJuRh
rTd8RWp490rvufeMGwZn7FhzdQJn5P7F3/TNhlVg8qgH8NMmcQBVdIm7kMqgPeZoZ5O/4iLum3sh
lgpMyHLkqVtEeNFYjEf01KOjLElBTFUjOSD9ISZdrWaqQjVIs7ScGUvC3ExUZ1+1fRmhQSIVnNEZ
zQJA+BTODuOF9dmA0plTXaJyEqunLI9uwzqRTTxzA0ibpo6R0gIa7L40BG5OuyJNrp3sdc68tCGw
xbEsW1XLEmLpaf9FYsYhU+I5FCEwMCq51BU9Irue+FNmWzGBhLEcxfd5MgiPpqMFUhb4MQN3HY0p
NysD/F64VuPrVvdpLJrb4eCUhPJIvRrLNAOMUjPTuqVO+3EDAiQ2RzHlgtTA2hH2n49dvTeJHeBb
VUvXFQWcSUp1WKRUbY2/Z0K1FOWtkoOLZyktHH7KIpHc9KNyN9+vHPZDAjurPHP5ZiLeXU5GP1Vn
LY2mRe+4y2axCgxcQNYifYx7EzDYWA3uSBiNbl3j7blJ0IjQN+0gZ9aQyN7a2pwtfuR2fax0d1eb
F8zouKLQ8DnbwO86MeYzr/2roS3eHtuk0EQIvN/rPYKAokISOyNylWQIF20aIOg2dJXhRpeTSKwk
vlMujTNy6ykL9molekdGsU1c3+ZCsNPyB8SWFkee4zrogohsKMUMjk/Q0Vb5GWR9irk/FIkT3vy5
+bjO3MhKoQFuV+PR35wf+9wOZLddH/VNp+wT4uAhSy8phP5c2Sgib5PvTOcWtEuBcWtHyMtEZVjJ
neuuBjPAvp21r00miVxnlbM3hfrV15DW6mfOjQbBSKPJdAxkDEdgGnkGebkLG1kT3tb28vTuuOXu
moH+Ugmraw+4EnfN6D4rv0V193ULe0mhdjjj+Oh4+m9wNLq+2bs3DfzT5eB2JmBosDgbCgTNm62a
uSG2275w5NT2/GS1U183IxBMK0BhWhjbLE2FKiKhgqIRDaNGaWdoODLO63R7Sa9VBYQCkKQYeFib
2SdvOwjumSiy5hOK8RXqp4V8i+gF6DRWZz6woKjk/nDPXfdF/rMdnnVqkYDflVZ5iJ0HGyikrn6M
j+k3RQdJdO9BIp8fGQrFwTbBPo0XKfn/HBAfP7P4ynJupSj1it/U5gJWVdeFGSjVGceGkY6nu/VJ
scqsHHLNpWCyqmxO2bpEnYV+frOg63UbUKcBx0OHWSwP69qSoV/GVJSMbc3cj0gqtYHf0RA7sOwC
9aX7MaAkmcLc6BnNVVYwYl7VQUhn6ue3KKp3MwcLACMsQSe1gLgsfsnn6kGuEzThseAWkX+O+qm+
YNTXj1QOWDo4rfJOrP+SSmxsz0bPshE2+9+qTh/Rjxg9+seWgNnxjREKLUNhVSzKdpiQhaZFrXPg
wQ9HHzm0GdiOGqYmtZ6sO4l0pTuQ/LTK5GfwA0/1Gq6sajlHZIo+yj538sWYTWsAm+MNWhetB7+B
DlUcEVFh/YRSQCVz7e+mnKqXuSEP2Y0kqt4KssTtgoE4t16ftTjLSK8TAndkvf/Ot6Nmty4qa3lp
mlRfz5J17l5fkhfiVjG69AfroNQmZ01ZaNPSK1d/GG36hDE1O8uSsaAml6mr1gv8UT0c2dnI4R64
OLs1gSjCFMq7vCVkXsdfApAZ9PhPI4MgV4zktpy6ozJAo6Xy+G0Q6OBwaYqnTNuCd1QRF+tEzOrx
fV/6+chtL6uXuX9teK7KLqQccNa6U5XeiKnVHNw0an2FcCJi4LU8W1tknCzNTwFNKw2h6o8F5hOf
tl3vg/DNvQHmldc6qnARQ5t6XEQzxCdJnw7r7tQGHXmK8745bUyVpE9vJfGoFSMDaD/3XmzehcQd
vlhxiGneWxWT3dqyOnfrDmBAWevxaxhcZb1/mIaEXwc4j544cmi+ek6GT/blaDE9oYVsOAD3fLL5
CDjV3od6TB+6NSQMYxv0n0xSsf2F5SROzieMFHB/xvDuz3rHGMxNUvk0bQr1a2IRsLZCD/n5H9iV
nusM66z2fu5pava3nl9z1AZqz0CJCzKn1tXySSGv/uEvyXioEwtp6CMvDhqxzzu5znNpTVNwhhQ5
VabYj+Qrh3WlAPEckRv0OUVObvQSJWQL4XOP6AG9Q6BpTe83rbLYM1ZNr7lMEE5VdyCoouGu6YvO
F0rI+tCfzs+VazZu0hq5PgOr6hPSQPtMbUwBMrKBw7GYdyuURIqp5L1taqJTF0qJ6C+Bb6ACYuTT
J4/HFuv9swmvcG26vqrF4Q+PBeAGt9Rc2k531J98pQkshRtWXLSUdsAHJDAn1gBN5jQKKfOfQF/N
gUtP2UFKMNGnqqbuovSPhUrm6E6jYZaK5kbWCARjrXxadwV0GQvJfWunYPZMuRIExzZo8nLYw0On
rrIX0QhHYtitV0267pUE4rKnE7a+wiT1Gf5DYWkjYcbnXnodCMjdz+YrW/69+QS9KzMA3sZYHMyH
Z6RAm/VuAbVTkAyrzoYB/WnvUDN4W78nOQm7wuLv5l/tkMtO4uZ+nTu11X/AvFMnpMQcTjL209vZ
4cO8pK/puY76OuNCQxuFyuMh7dTjvUsZzAogEKpsLNXIrgQs9On9Im8tuECpyRWnj6vxXYghDkBH
IFQiMaNS6xzCWaru1vY0CrDqFA6PT/Z9mai6U1afJt7MgSHfXp1HI4aCIFlEItWQ/twUl9fP+H40
qMLPT9IWpec+WlHq0NUKcKsDHM1jqdJ0O5u/tPiCY8L69WLF1favX823HgDxyKh9g16mnXbiEsv1
ecmS1GjRpX8WDsZ6CHsVAJK7dEqioKLZocY8ZPve1IjpVyJy68OPbbRVoI2AWKUPv/HNaoORRoPP
bJQ987mQAlZ05n+Iq7rJcc1QuXL7vnSDc+SN3Vp84vlpPxgxUUiZ4FuFZnWnpPWEyZ5rTVLKbZiQ
0tMLIuRN7XIL5IBLSDXao3Z+/TXaE5GWKq+PwhVKgJMs3zhk2xlQDC/DZiejY9mHtefEooj6FFuI
k96VHgYnDzNA+CcbDwPM57MwJO0pgMV3vVukZadsS+VM9Aec2gzf7pAWuzNAm/0M/x1nchDUxGXb
gz/DEmyirAPQMD1MJP2k+KQDVYj2ogqUhRE5p1+zNuh2/KJ9uBa73/QuiVS0JavttJ7UCSIWnvji
HsA1NZOioyj7U/jMYPMmhdBFmoxAZM7vBQIdLsifVhj8Rj2xMD45tbHyzIB6de75FXyxjTZMIXN9
T/wvb577aKEL6NhtpG1kR4SJj2XGgMQ09fayle0O6xwTdkH2oYFElUu38N3iwXbQ2nd1hKoMvzhb
oDy6YAFvkCwmISIzxGnqDgkHgBH/hgC4i/oVDNMsWUuuIQKBhztAtSphtOSJkj/VuJYOU/MYWYfx
KE+HWnxJgAT1jvMV51YUzhXlg2kkxH5Ifc016Q8XEQuxkwKAZtI+7LPbFDW2gDY2FRCZoZXB/bhx
jJBlOCufVXK9VRp7TJB3AJdKfCju0MjOLcTKBK8sfsWnyCx68fezhTC7s0/nNxbRx52puv10P9ZM
5AAU8cGPaeDuzic42MlzKrSlJ+NSluFwYBBZOerXLSOShNPRHTatrBkAfrPhfWiS2XICV8PFNUbd
/Ii/k2KUnHkY/usO7dIG6uSbiNKLK+jbo0gYboAzXtIpcUOrZGrdqrSDjX4YBavg+TdFb5rorAAP
hht3ql6na6oarDsCMEyPIDz+cfpEldldLj5jPzboP+XqzApAosINOJLq9ursVGRooDeAGAmrxUbD
e3pBLDTp50zOUBGnMld5XQrSTtG4K/LRyjw5rLHl3/tOBkmMTY/zgxubQs36559FtZXqMUqhsO7L
L/Nw4QMK+BOTW4aobcSJok5TpM6TH82KMVJ77O+IQXgmRvrRwZ+hA/xGxJBHySFuqj7RsiYw8O7G
YkzymffPRjpx2SVLGjQ4EIcbpGwwvTMSGpd6UzOl8nerxBCguTQl3V9YU3CQcmSFPyX1tni9KWpE
BKuN4rBHG5ZdKd1qBBVsZ6q/wDGS+kuJqaaaSbB9YmXV/hur/Oy/HAXcaORXv7mNlcYe/Rwq4vVR
2l3Oo5qgfPVYqsAYPp3JeaorLYjbtb1etuqKQdDbeI1ICpgLfun6qjhxRQu3tCEG61khHpyNZd3j
7lN/gmGNENfmSwP3pGYpm+LbDOCXoNrElqohi59Oy210QVPipsaH9JlN73POaYwG/fSgBHqGYAxS
6lm/2LfIMO2IB7DYwzZS7EGyG/0SzSD9ilEVy2GKfmMeCFbT97otLhM9xSg0L3B7SZPAt7n0PsWF
n0XTUb87zYgJSo4ge5B+L/VY2ei8xUzWlfjUSyTuGqG/YXqpOFvZJRzjImbev4zyd4U/AChw0kPe
cqHOZPIu9pQ5pjzzHZvM/YDlb70+9vTTnU2RcyRultl3wwOBygMB+rTzRfVQ2TT9dtSMROS2vgiK
GdTl9KviOYiFwTettXB+Ka8RT4wRuXkI0gxOE4eAiPk17fuUux/uBdNtvSbVgaqJF1N5+0oey5PP
hQEXSlUZ30tjqP9RRxF30tYwCYwEcD4BmUg0jefETMdcYs8CN+8IPQweDUWufkWsXDgdro5iEeCB
RAUI3O7B0FlbPpnwASPpiBTWFO00jYW2MPx/OAy5F5Mokm6xPt7AlrC+LTcmTwHmteCMWNF1vZow
dF6I7gTvrfYs1D3iYHKjY/0WHtucENynDNrhvZkdtE0zjkWcWj0dw+Najh6j6FUA5eYFVol8N4qy
gTK7NtzfahHXEyv6fM5i8vH2oJ47HYRJynHEid4ANLZotsT08//8fow6nJqb49hdxpWgzgQuI2rC
j/CElTdwWLNjiTRoddkBVRoaJRghAwXo6AaqU2TiVWNsuBfiEO9naxIPOUNFUw8FQT00HrgAX43g
QAsTn2ppp8jXziLYTOIHhnSZ6UIVOlTvUzfyMYEiwNfdXPO373PcnI5+3HmN67+GIfUQH/up9O8W
ANbjg/ipQ1v5BnIwaKisN6QhFABCAEkfDmMclqZ2b9XGLxN/nDTqBZtdpBwLe0nUIpoQ86M/XPcb
RTyAzVQoCXB4Tio9KDi7i9ApDHjNV7m2VQ1Z8j9+HF/hNfLWuT1mTGfQ9PqSv6q+XJaZ8f3YpFhT
vjMjU8kVZ6YAaWvdOByV1NPL4Y96PLkw/JsxoaoMu5hA9pEMYQ/YSqDZ0eAjfW06KgTjlc7K2dN1
U4uKKN85Nl61tkRtkpa+y+htwQP2GoBfmoChpChSQZqUkW9v6X8BZwqORGkGoz4sXUowkgfOaEie
ooo/XE4tnyGjfrXIgufNu5BwXxFxVXpQN4LXjhkr+qD6Nx93XfesmQK7XV98oV0QCL/tTM31F+AI
MrQsL8eHaZkXK+7UrnzlYadzMjQTlkYO8VDWO7AaYacm2ajwGSRxpHUWVvv6tPRJ5Od7r9Jb3hY9
OynKFM/pgZDgBehfp/TvLuLJ7H3EjC3EmVK95+LawkIH1bioqbbDRP246MNI23juJapKPhKuzN9A
i8kFaeDRm8dHhKw79sAFLHQiNqf/bo4tGkUT6lWw532/U2KGfwqM+7YbP+1eNerubn4WNKvNRfs8
eqWkpI0e3yiLasbkY3Vq3gk4eMLGBVowcgQaHJjBJ6ZplyrvLRerh88H2bhkQehLNW4wwTrv1c3G
whQDwynpTi6CX9T/GfQ73lJyfHKgXtxlByOdJmdChWGUnxJTqn4Y99Up0pwnP2WCy6L4F3OuFZTQ
HeyNXTBR4P4ySVnkXw2rNDqwjV8zMWz27A6TuJv9KXl5KrGWpEFOgpuExUZhRHmfaU2Or4H5Wm4R
bX8NZQo8c7/y6aiYiXXxCWNcEMtfYeHoAoF5dIWcxMO+2pruW8IoLW0H/1mqnxkw7HmUyfkBmbkD
Yijznd0sW0uWVsBOeBbGEQ84Kyj9+EohL49oeXMrzjI+INNmeg0SV1MKboMxuqSWrYN0c7ZPXyBX
/UQtf9LvURwRbUR/J1e7lsJzOjU41nhZw0ha1bYkEnNoo5KChOz36SyspOtC1L4Fc9Sjs7R2Icgu
138dYiPSVHwij0h/AabZcMjZVr9dddStjShetP2HZ/7Ft7NaSQqzApFyKSNgUnn0cFLGAGujzMXc
IiLs+rq1+bLDerXsRCI+xLVh2UJsdefsjFyo+2PoaTsXbINbnXgJfmeoLM3DN/E71nlm4Ya7ZJC7
axmdfCXUFBw6ABIcgvplGeIOt3M8/YbzJJjJIhwHfSC9ZnwAvnZW/jbcHlKwNoap5Q2hiMgLorwi
Zb/DEapLTTL57LkNiIKwhtrv6Q4oomvJ9yU4A+Ysehpf+4PBbYX+RQY+wUHqsGhzPGVoWD162cOU
arNU8GLdcYCfDpJLEgtkvqU1CrvcPKyMDjOgPTAC3/VwjOvH+1/dm6femARSIS33ZSguemg9Y1Ou
LG5KFkJC0wTfM7BXEahPqbGProUUsXMKnCAgO9H1ECYA3fHwnLOZe7D5Pm9MhUlv6io4MUGNTO1w
Ia/epilVFDvyEKADQIhckwNUPdRUq8Q8v6qfjNyv4XgzF3H34cn+CDjqkLnbIfs5FW9k7mTxR6Lx
pHVXU5dI+Jwq6gz7F0xLITOpjLliyZbK8nhcMrmMvrTnm3OODSPMIijMWlQX2CpGHjvnUS/VRWda
qY+4Szd89Uq2DGmNTpoSnawz6YFmphVyON07HZoBjQF3H5mrAl3kjB7zn3Z70FotBSIBkSJbUjJ8
xXz/qZUhWjMSHFWh70V5NiGsMrNGp2F0e1/mwlv8a0h9yvNIEsIkt+BmN0s43Y/HyiDBdcF01aU1
i6M4gbKm6DvTjbg8RXNtuyj5OQCWiPNd1dEVP4QYOZbxD9dxH6t0lJmkQVeOqS6J+RvGvjQwW1DC
jUDsvftq6VvWmlpo/r1I9SUND+VJCIYt8O/2i/RMkLJ3WAZtNJoUzTE5cIFZfzFgSAAchAv7djlH
UUoAKUG81llryOF9ok6YtR8pl/ATSnnJ9ppUhXWm+9TQYkrUUoU+o+gy3UE5BnS4KMO1OCUcvVjg
iF8LnTgHVjb6C6xrCFcxO/F1U3xNpXex6mT9udIHjMKZaYOkkhLPOMW+rJ2jmMRGXkoMBjR6DcV4
8/eI83pz7IxP6w3b1g6hLeSV/n5ssGDH4eo2ik6e60Q3zETzcFukLUoPpoaFPHMCOjnFffTd21cH
quPuD4S9zaBp+Gkqt6Jr8EfdCmzbIzhIPps3n0A4IRPoWxH+Ql5k81zN2uDtDxxIHu1x7elp7+Vh
z2ppmkpXBK4QPwoqonye3SDA14J5hkkOcPIGvjO26H3CGEvJPNY0nzPtiFziUAEF5hnKOtaHPjlG
KweVRp5gBDWhhXEAOXQNcNI5SrG0WOxiNC6XzRWovbM1ke+g4fkyOaJWvNo0b8b5QY/BxdCooNlp
hK1ziYWcsSfh5cFYJ97nGal1DLF1L69OhylPMsrx/6dEAUBW7mJFDjK/t3haZosWFecPEyR4zwWN
UQT3gbaLEwOcnD522Pgp4wRCKPkWX2mFpmlcWg7afN4ga4OUZOsKcMQyO8hNtz+/MdbuK2mtRyis
VIESJqILFZfhT7dzecbefmADd0O1YdRVg+Q0zH3+eYijOKgMSYVEnEL4C1Y8DL5Xp38OivfULrvK
heDn5qBOOerWEVKGY8fbzvQC3dm977muFWSVw6zz35vJvNd3zqZA0MhH0EklE3av/lGNJz13nNPX
XrDw4eiBfJ0r/D08/WbuQyWoDpbDqZzHloOkGoJCXdFapWxzbRFMR4NLd2/Tc9dEiSTsQBiIxwwb
VndZcWYyov4e20paJOgjX3msNSOZ7nZwIxMPCekQEWKUY1i22nBkTdFUN8zIcrwU6gYq/62Ot8+C
lfDHhfOytKqs0g6gYpgC6JUjXVNTSZx16JvVW1+Fn7E69xTWF+Mr6RWkUFjE8DpjU/5bn538plbE
qyP4dQU6VFsNkSXzy9vUb6qhtT7OXlzrQ/UCxeQO4mmGVOJk2A57yUpwNw9MpFG25xjh8p1vPBfZ
oZAx4Nl8Iuk3H3rnEf6mD1yFv3EzdO2ubz/fZMmfh9QUiMEClHboyct62bZflSAXEWnsBLCycoMH
EQnrFs6LAaVBrS7jryPv4sbaH1K3en+sgVNL6+ftWJgHf9tgpIr7pmDI6nOyDY+P/6mIJSH31QqN
bHbulFx+XArWMxfOJmYMcKR0vVkgnPcBobEUCQRR1bJzABdvp7Uf4kKFGyWWzIeXZque7EjpaFCO
2GXD+TxbDcXM8hr/L2cX81vExkI44qlbUFkdflPJIrH+MTCLZouOgPns9s9ZWmQ6YgJhYNutlsS9
vT+frUFzUMZcXH7i/6zlBdGbHfCMbO3OGB8oUc8F5PxFrwR5IUY3hD2ST7D1T8YmAjOMJw/2EF1X
PxWNp/iqWMgiTHq1S0bAHHtQcGEosDiW1p0tkp+MfUttm1dpw4eLpLDlSQ1kRgVgq++gfaVtUveI
SHgYBjq+RpuYD0QvQ/MLgX3U5iKHoyY42d9kJPt5WJdvgxREGMoABVaxnCBwQgL2qFoDTZ7Sp6wX
CvurJCeGw2N18bEWWatMyeLOVXIHroxq4sK5uQslRFwba2C79Lr3FFEX5F/1HlunUSI+Rd8q6MCM
uJa8fOO8I4MuaUwdZI1G8IEnYb/hs4NfjkOoMrSFcDSJ/usfOzr/1DIiDyo8IRLQbuDgrtMAcg78
Fc+ld3V+augAxLKp/UEwLAreGrd5mQa5shw5NYhLTaEEzs1rdmHKesZJ2qbe3MPxeZjLal98aiM2
6R3SQ4smM1KkNkk0fssW+gQ9+uxUECoabT2VJ4laaRooWPhqpMfeljohQE3ZE/PZonPqNfvxwz4v
jTibLJcLK+n0bD+2OoWhpxNq8pLR/Il/jVJ8nxdKTiIba2oY4hS+S7z8gRJuAMWpKlymRhRXApJk
EhxjFC1rjYmLoNdwcSdCIWvlVsdAN3yDWSyUraxBBGw/EIvQnYluDuWbckekAvRd6JztdrxhDTSK
MGc+0wsZlzmvWv819BP3iz1JfkbRvM/nyzZWVtD5H0YWgbAyEmZ8VvBMevze6qv71SdFWXVbAEcg
kHUMp2Tr/gQ6xJy5QVwQlMu+GNIion/Id+XL4CbDd3qawUanYNrhjPS11larTrK5I0ZSEenReQeP
tumDSDg+97NDjVSPn1NCi921/fyi0L0X3E+HS0XqphOXHLhbJ2R/2pa62GTh+e97VkYfJ6nzFSMF
Eo7O6Bq2Twzx0WWr72D7C5e/s7GIMslgWw3u7y+wNOf1XVl4UO5bOAgnrKSdKnCMqsnp+9txPZEj
ZJ2NzuGdSHkk/GcxpAKi+7JDZkcQgiz/W06e8Bm5q5ssRiXnePzFuC+bQBG856sasXUby01sJThO
sjAsKIrA7e2WnFFOVlEfYBbHReF41Z1vZPCh0T3BOFKbnP/fOl0R7IuQPDSP7QQfLkC9beYNCvnK
aPL2U2gDGZa15569RieynaAT5ACywPBVM+hg5vNpnWc0XbI1KtC2tKX1hVaPfFTO0SgpnZaIaozc
De1ilMVxVjUIt2ZvuoPqz4w30yr1iQrgaQE4btuYYz7hhg4nExFyeljBi+aDXJRBYo/FsUZZcT1B
ZsljLxbWmuaKmuAUEyu/sta1wEyv7p9S+NeCzor2GfHvi9lYhAAJeJUKqqVunu6lIfs9m/u4yDZl
llg8CVC86cp2B07t9YcUJ2fCyDzaY8DuAKtg83GkLT6KCwEsJ212UsAMFip5hFF6V9kqaLzLAOm2
kdNFT8XzbU4LMD+EJVSEYYZkzgtthj1NZ0eUBLsCeGssyEfx9bT9XWcJgZydcvaETnAPgKrnrtmk
Ms9MNWmxzPL4ZPlmK0XckTXbo3QEzB5pBpH20YsjTXd8ZnGd+Eb/dPjWPDFs8fsY09T6SOzb7Ui4
5tSt5DHdo3c/9jnwIk5rL3jPaS9uiP4n+o4lXQ83p3Dd4OaK+TWWIOa5EYqdz7MSImUG4h2TOCWh
uH8BZMQg8rGZEHEHaioEaXepvjQYWQatO8jZYGPZjIz7ar9U9bAHrjiAYY2Fn2eEYx9fczufqhAh
q76ywluKARdJ1vZftZhX2u81nSXQ+uPVycdTwmP7nI13hXtvxffx4Q3YBat3EYx0ybk+APDHsnhy
QS+ciC/CW9tTx4VDL77t4T6zDW0/URGXdJX1MddyZJr8bIlvouQ0N2aNYdJy+4XAQw+DlpvdZQxE
O8Szto8dnX8Hd8s594UEBH3oKU/G9IhS4xe5OlW7KrZ8gbHR0VSs0o6pvW1b27Gvus0mrAvUMZbf
OvZimEjDrpTK7X46fovuhGNoQXceeWElkCAmwkVJcDXF4TjDAONQxjQoCCPmqqbA3c0aTPT2uq33
aPcPgk+K1/DCwit83tqKlZEGKCqJ3pDRAbxlmnDkOdxbPehJEX40C4HrJ1qcIGVpPHrV5snsiOb3
ULKAzu9pSZVllF+gArn7wE7psZnF44cJHMgLvDCciTPgjrklYnPXenbwKnzVIOOwzz3VWy8RPf03
Np+YdZLHl/7Ej7NO51/TcA3YTGbLxchoy7o1mEkZIzxXmr8JC784/58XCQIw/gEvYj65cZWkvcfz
D6HXwgvgJE1XlsuersDcME+cCKqMv+DEKRq6vZKz6Wu8lX5mJLOXnEnD+VkLEltTJ5mSuHAyErY2
wYuUu4MQHtmVF3e0nscr0IbfVgTk7i0ds5Dou1vkgeP6O5f4Jqn0QLoWVBeEuxIlI9DBBIFyV21i
mJgTcFi8Db/NgRG1lzV7298jzl+I1qrzfxiOmGBpTQSob5SC7QWBBk8fQZlcxLnfUhK9V3muRX/6
Ji3xT75ldNCA+yYuRbjFr8AS32xTwavC9mI8rUsVEWIbNPITixTAINKk8toxvPpPxB/VLBSDd4yc
CKlXEDMZZa/b7v/zltf3RPOZ3Q/B88yaSFTJnLdc8wP8DdEqo6xXUkJHBtqGfHRVGZ/u2fSpGgO2
GYyrZwo6E9CMqN+mp4xcd5GP6Fv8mOeAqwv2Wi+seYu6IdxmwLqGyrMu+eZ07Vlllpe2ardx4D0H
ASIKlIZhzO+uFD6FECeaHmuROX+apI1HCC9Ci7f//kcLCJoRDAc5ENnydoZMMDybtZEHa0L/KH7W
YTCmVmNpQJQR5OylYyfYggQIp95UvTQomOnrQAMRWwbHUzPKi2s3pKqLy9eTJqoQAgbjEKWl677t
cJ6ex/JJaRqOz4ke9Pgq8gxtGrg7V9c2WN+sUlY09ilsmoZH/tBXU9dOo6VtPeNRFsNmBgQu5Gsd
rL6lIQVlSMZcAB9U1e8RgHPnA2bBQ0C09hehdpAnjI2PTYUKYWuELqGQueMVIgCBRAbKeYUAyjT8
Qu7R+/oNKdREiI9iDwODACM2bJITQoDEadfsrMr1CF1NA+YdqX4J0BXHsjvB3MpRAQ/VSUEUlt2o
WjhDSsp8JIPZoeHwpmdoPNWaN2VubalLmxr0eaW6LROCBa9yW6POCugU0otzgC0LF9/liaZXVv4U
NYzTbxebv6g1x3RoVl2Ly4K8Xpm5yLrqtoPwlx+ruxOXBvlvj20rQ/MPuQBhFGxoNzsx8PasVEBp
cfatA2nDskY6RteckAsSstvQelB2yVQte07+/2TiwfoxH3dbGyTLCtfiYrpgUjyOrrg/EAw1IbTy
A96StT4scUuOmbRuI6R3Vq4J4IdLQ77tgNZGaWu80tDEl3S/uCYHeWi8SvdmK3sdZ2XekRvq1sNk
8vr/+P48I6tn31eUgGgjikW5O52hsS5XbnaOQ+Wfr7AohDxSIhRMGXZMxYWoxjvILpdAgNKpQSyk
RlcPccAfeMqav3KYoYxMbbUHmQtmo1pDJtdQ464jK+5vQjZMqSb+VbjCCUz5nbKAltleiuxzuG4u
IodDfOjJmKlq2p1Bsl+HL9G+6zPPV7I9Vsjo2WUQz1wTjV35AOz2Gm+6wRXy45LniSgGiRRYbyVW
5t5mGoCaiay+2VlON4fhlb32/XQlQvHyBPSpf1WyvpWUhx8oW8rk66eWlEOmrRGHNndbZ2oWbW53
5p/wW56CGpojIBC4mFNBNBUzFKWUGzfoddN7kenHpJ+pg0drG2JYLVmqgMiiLmfHf4mNbfCaDHOF
VDYIoW84/vPpIcT/WV8ZRRobFjVZUTQbWykOTY6YiDhYrIPRPaPTpllzIN5jxivYlpxNNFABNn+9
kRUVsjBS815XNxZLWe6Co5HM0cxg0IbNtbmYDaEDtYx0nhrhVHVuIDObwRc4B+N0LTpqFEWeHxgW
Xn5KcRPJSbqrHm0vGqOe9Gc3VxWIsrRgZQSIyM/n9yQzNCIqCcebaBsqVcYcZiXw/dZKXATaEP/f
yP/RxohH4zKjchSOCSDqAbOF/QY6ho6FIkX9p86QZw8RtumgnOx4I9m+aGk39a7oQQjkMSMXThWR
MwlxonEYbZ+u3xNLNloF+wX6Knovopdf+0I0DRe/B3K9NwWMpiVTJfekvkt5swp5Z5Dru2OQlFAP
CSd1djDHqJSyeSYtIfmPL/kAHp3hr13ISMk0Z09VixcLAHdemx2oedexHyL2FwuGa0yaQDapRbcG
RQ77cTbnyNc3H/2iekDO0tyeL87QrMBvySYkJdn6mfLZ96Eh6UVjBwy5uA4jVDfyjzjO8TDkGqR7
BjUwOn9rEK7HkKqozjA7K/URA4Q46c9eE3v1PgcfJugD9UxwyE8Iaims3cKo3nqdGmXTar7SoM+Y
Mgq7vKqaIqUan69m4nbRgiEIajccN7+F80RPexZnBzPjITBNVRubzN/ZwbQHVIGNJDAc/Tv7VlzH
M14S7DnEEgdeVHT26GRBsjNWFaRCCSuEUsMPZyWq9/Gmj0tZZvxOzR1wgmT4MayK6i+G5i04LhCp
61mIlC/VXAUVbfIR1MqXgcAz2VKtun2XoZVeszvyeFTpFXq9JGFeTGwNb2X/ovoBc07s2SN5UYeI
aOuyH1BPV399Vw+aAZmO/NKyQnCCOg8BbHEajrMvEIywP0Yhuu84Wq5yi//t2mrEM3Viq39Erl+A
PFC+/EORWN+qj758zINbp6aC5WhqhapFTdDIitPoCJk+1mLxgsO569VsfSBVkIWrOtOfClE48F9s
yLhlkG1zEHN1B6njRearEhOmrDN+GqPG4WBvDObwd27vivJOhSHn1R4x5dNeEa2caDk8tSZrkCDQ
Am3lbV1wjE9FqItW2IluYTcwwQx3fL4f9b8MsKoQuDnFEI8kce0CFkZzU6iS0tWVIWOLYD3r7A6A
rFmwklzypmY+wk/CvydP5wE4VaX8QjeeDBU8Ala2C8omzyf902dsL2ueM0IExUnztOkB7bEYBq3I
mzSKVqGY5TFoqtshJLYztooVD3QAizncLKRL50dWEF9a3utBxzHWYj9kY6SEBx6yYRuLaqXsNkFM
GDz50IUAptftj2xNIG68vORPxTc1QhfTQ+/0vOSrcWWtpS5vj/3qe7+qud9aWQjOyX0HbvUquqLM
N0ZDpXs94YJjcc2pdOJrCPLz+kz7nmvdAuOSozMoSNoJEEajFyS3q7fxZjJKaMzQwXfFmZfCZcQm
V+IIPHvdHvLdwz2DCQgd9S/qs3CcHMaNAd5t+xUS3b42Qbcz5jnkoznotgdVki5W37rGH1iopbSi
FNsxBIxSB8n1UPeVZ7v/0zSxD7a3Hx3/RBj1k2XOV7J3xYy2RU24MyiLbpnpaepb0Wa05Z2/eys9
hJCg1271uS3xLX5kAWXmhzja/be0XewTah1UsUfG67cqFd36vik7Lc84KEK9s1jGdbRMhJBrf64y
9MkBTGRPD3zJ55GBO6NzexjauK5g9fbVbIfVUXTqIViUvDwzUryPFeo8e7yK4xl9D4Vy0UF+vfWi
JjgikpWBZCwcJtDqpiH0pcv4s+M6osf4anbzZBlFZne+6nuBJMvAfUszg38qbG1C2O1gGlGW3QbB
GKbWtqopeFM+DMmSOjBh0chzpm9XpJUncOSbwnZ+QtYc4BQZE2xRL2yB7XKnswNap+vVm9SSejIx
PhVFEpytp+VTPpgVD6MkWtCjbbhGhnjg2Pir9jl7qjwIWfgwX2DPBDg7mJZ6bofjYE5woSWS3q3a
ZKEXPako+AcoVzA7uA/1tLD/WxeHPUtB7YJ5YkyLXYMB84oCFazYWSOzVXmc5sXm8qN95f+KEI1V
HzQSTdXiAXxjMO8tc4oPDS9jk1k+O/rg0KQQfmTaJbOWugy11ewCWxIjwcp6+KiICwh0RbkOi5cM
28Oy45UZvU5dqNnY2ot7L7hg7AyhYEJXRmbDTWtIG1Acb4f5DYd/eUpoVXaG759NHSA9mT/L5w01
W8UkcQUTjQQ9lKaTWA7epfEtqbsACrWqGbZlfvvKjT0uRlMX2sl1mzX4/oOwaWNUMxJvIRvNF7I5
NrIDtaEmmJrH6GGe7yBHzfSZ9ZgK3f2GKzzMI7t1RX3LRacjMrdxgraigi3f7uAe4b+0TnRqo85u
ZmB1YyQs/eTGu8KeOaqitBE30XxCh/YsHUVlqhW/lsdRdazprlH6xv9wCkjUGKNv3dLT6BTUFq1X
pW3QOyduBN7rceLlh9tnotPT0pL2I5Bt6fhZ5kQQMgTobUYhJmrV0m510AnWFYL+eGY6a2odyGEK
yY6BvY5HniFqQTN7mtCS7bAQY3olwrHzSp0N8J5jhcCeMoYYZkY6miv6k0eW6fAZ9l3mvWy2pMKC
ed7jedUg0bNBMnLZ9hRrHVXlTKtWcHxKLzV4SV0TlYjdm0Y2e8UqH0AFvvs21Iz7TmZSo1wSN/1h
WWrUbG3gRjMSBY8NtXbZrycn23WYncHF6cX+uNa3NXUUauBrmBmEmjz8wksdbpITGN+7jZkoPUKP
56V1KIg4YjQQbj5Kvoiq8uCqTXYn3tmYL8NDnJJV2HjLvouWudSsyuIJlBoRRUlH/jOSNoJi9qgl
V0Amxg3ZmW6XSr7z/KHOzdpBr9O3IPF0+M/EDrj3oi67vBBbJT2DV9KpHRKCg24YJDGbfvMHV3mp
Q5AY2cWGdgyKPF1BsITK1Z7xHiimASetcTnDd84MKe1rGPNTYjfqf/c15BagiIbKGoJDyJG39wAH
i+wYOQIE51qCEpzDPjbj9PBCAje2O6xRQMMgLqqUnHCkQFXsrDxrAaD3V28qh4iJg9wiqV+5/J6q
yoV6bzjKtmTNUH628PxkVdSoLjTN6ku4DopyN/emmBDHse9DriMTqk35JfPeeGPebwfnN/HD1NMG
dEuSyZmxCkEgrZ3X9N4KvZMKv5omaxA0hQNyo7WLnGwisZfVhv6VFdIJA15MMyOU0LafECT5ofhf
AqcCEQWPoyu8I1FuxK0/50VX63a5+z3msg5SluT/gG743aOQfN3fyxSjdLzIAMpaQDo6o08bHzKQ
xHD8MUIYzPjd3rGgX/PB3cAgCM+TinQJi+e9mUdtqetXoKCPH9Lhu3YdDw1UWE8ryup7MJo7ueAm
IJxVXXxojGTnUrioh44jxPpoLzfPqzyQl14x/OzEQh8oGnoAviRaCs1fgae7oSttKerNhS+KU9Or
d7Tf5wno1fSnqx47k59vU0EOUBTFUcM779tsurv8ugxADIWHyAZ9wusPwQj9q6nxTkvbkkEcrwqX
NiuUjNACT8DaUHD4aJlmz6lHsn54dZrwc5Ee6H874FfLfPfgAnqRiDUeiJ3g41rY+ebkMwS/BtrV
SbeqtTuajX86wCnKr8mcsvtMolz37npIB2M3aFfv41Pts5Kax1XiPZmva0hdj+OgCZjjeYXK3z4C
xKeHeJslR9rI72TmgXNhPlg9C+IeXLX3xmtP5b7gj11KkTNUblS6sHMdtKS8NHxLGrI8FendqAFP
nT61+5xx3lGajxJCNbZaEYQm4Y49eSpSsM5PhwUnjdjj71E6MW52WiXsti01OS/Vl+OZEkLZ1ST5
uZpqkBqexUFufcsYJXSzE8zuWBj0qI0bB0PstRUM9RbvsAAM6gdIrwmFJQUF/I8d/RkLOzlh8LWd
gb8la9PZIt+u4gFIWYj++V5Kv2mGSeEti1t+fLiNGZpGOvXr7LA5YOFrdAOQLtY1JdiObPXIVwKq
IJdzEn33MaWJ3oVFwJJSTGCe+RKaSQWPwj67oKklt9Lz4nNsEwU7xt1fksDzu5dw+zXd6fgYCu+/
RxIOCnvkzbrF/JQpRnpVRWMGjBupoYmSNVwRteCAP4Bj/nN0NT6sgKWYidAYdXFhoPZUdZ1fCJBw
S3IOpAYJnS98ec+m5V3ZlW6KrTbJdCi2L4UUAWryuUXMQ+H6bhK24h6zYpnGRmDtUNhulk53muj3
nRR/UNWHvrcqowK6u5fyNkTEvlH0q5GI7o/NCoxYmjGuOoHSeFrLv+dw6VxRX14KN4fzM+Ztebe0
yB+CK3ggMdZ4UQeUDpey+bthxGoK7WGLDJfVgnMWCi42fH5ACFDCkl5HvbuS7ZXpSlApFd7jMT/b
9Ez1Yy7KlGQ39WMDVosqyQTELK1iNxpfr//XTGSLE/tuyk6AfM6d/tot5OpQ8vdedGkWgaryMdwL
3My3bvZztT2xxbE7XH1TGB4gGSBwWy18ixJM5nccAB5lkDWhI0Em/NHWQW2QNKM/KGd8ttPP2QrI
ATH7bSXJE10UbwzIHNYusYAZ/Q08MhbydqahsJb8o3bIihiRP7mpvAip2SPva5vsWZu2yhPDGhT1
SbP4NmSLEf5XutLpnureZGeZW94s+7iTi9h6+NlLu8brTzZy8FMqUEWjzQkPerGR/tS4Jg6y0PSh
3+X76c+BkaJrDgCGPIhWNxPDy+NuoOcOK0vTOi+dc8WeuexyAlN0ViL6NKg/fJmOgHmnBS5ducM0
afk9eszwIKjBiO85RNEnAnQW3U4dTPHXBuNjZtF+47hnpym2qAHUFYnjMP5Qmut84IFwUESpA4xt
jWS4h6vXMSxbI5OPwt2r95fXLgLclVomGuBC7BVxTyqHTvaCK2ZyrF7nNWi/CYUeO/Rt0zkOIgEh
cGOFkD29pDoNB/5JS4u0Zh8uN2DPo8Ep15IFRkJglj39WdxSXwF9k6WT10EhM7pDBZoKKMN+/lf8
V54xZdn3eNlHFpE4afr6PXUJKk8NG0IBAiSRcBEO6cCDTw9bz7yj+rnGyhQ0/Y9PmGS/gcvEb1HG
ewHnZPACub+MOWWwzTopzBGxRwgajCa0OGt1E2NvQUmFg0nrUq9B411P9WX7QUdNb4M6dusDCyWa
HzvwdKhTBR8jS7R5HVnoKwlOoT6WrCXmQwGYEYPb8ByviBh3Zn/TZpEed1N34waRWDEPGrY1w4v4
TD2UFd0mq6OP1RrzbmfyRfSSs30s2Nl1W65pM4Wf9k5A39OQPS1hwXaYz+JMA8DF5d74JGFA01bd
9Pg1L14Mw1dMS6vn+qO6biMDJHvHbheREPs0KMxjoOTzkZxkHH5z30lz82IFlCQeI+h3pGRW2rj2
AwmV1BuVFNe7qUmMrOh5GFj20ZQlE1A7QjIWBq+ERJ9sOQiDK7Cg8cc2qzKyrETbGiBo/Tg8w7fc
1ml3SROtg23sq1XdrA6oVgRHMqKRXYpVMATFZl/KTXtshdzv1pYAndbUOHPo4KN+/8ZQZAPF97re
Ixr6Nmz19sqhBiaCAr3m6cDbPJncIF5Lh9LC+pqGsq6zxohLmruo+fqp5HvhuPdvvgSpq/HFS0oL
ZkTVimyUMO7/L3l0ACRxqZA7lu8G7gPabuK/CXb7WFe5HcbYk0AmnDT3pffYvfeVQi+bu9J/uHb1
BwRFcI9M8wPDqtvar3dfvO/ZyBVtdgRiy9eDCQqhI2Cp31iwi92oh9MsaSUeIje7cj/Y9IB8twvy
fnAaJxf4k6unWBwjrSv7MXqV3pUGMEKwCXxD9nNpvvrkjuU7Deq2p46/0pE2eGXHKHaHT6ANak8X
yzJS+S+jQQ+fH9162UPNpZhQ5rpJpe7zFns7Kp5k48uqfCPOQYHEe9nlm6euE9xZg2R86yLWZCBa
QE9lZ0HyPvsmgsl0k5EUMpDLZ4oDHNPlHs07Eyu54rYqAsFhDpaHVNWZlcEY5/9fxqdZ0zWUoIpM
rpKId4RdY49xT4KyhOr4zIxqtptfQjdmG0AtTShquNdTZmg99qbNvYOSgffth6xzIYZhmWk9lN89
kVlc6EM7ZAg2AmuZuRIq/zXJedcvYsBcmae1iuHVUzEUFgx3rzYlm0KSRoc/d2zIeXDidHk45qan
sLfEkThDurcY+x1Uhss5VEPH94U0/eWmhTz/hhBaVGPFji30YtogE8Yx1djuPvrqaugJFZo7+FxD
/RlrDneAgBD8YvjSv4GTIllH5SXrrLj8FCNG2QNPyMMh3q3O2JPuQmtF+jKKdIvXBAbi7pH4wcC0
Fbgqv+vFBA+Y/QlOX1w2UKwxThO9sSvWAPgab4slO9cCjoEtfwP0CEJXnCMQy5Lb1f5VzHixjUMO
XhvSzor3GkPRBljv0v2HOX+LK/MhrePs5rHJ8N7e6twOBuwJggsUjpTEoSpFsbMOQeIfw7hSMwHo
IeNIBpub+nkL0HgqM0u0srtYj2ZAzlZ2KevSrqVO6xzCYiUJUk1ioip3Ngw7ghIPREy71qiTcGVN
V2tBdArJQ1u4VkBfQgWJgGPCVDRkU/kM3Q6V0AYuwGb6l32ErCcVSgDBFPxUIFf5r1tyFK2Lboo8
1NO4+QZ3hDI16ALAlWERgGjx6s0uKouTGn2szj8uRkvNrqlgkLjSBZ8B94MTAKX+6ZxBcY1cgR+b
ncwVqoXOxs8gBZRr8EY2g/++jfapJyGGGoazXm7EtlJscyM1+MjgDQ0AMJcWx6gH4UZAuptpknXf
OQFkfrK0veDmGz3nIhy8cOonaYzrhF+XNwEpFJxxkYRf5Cg6YoSSSPQUFM7xNHhjWbxxMXZuqPQC
Q+uKJcKkQJQncM2HiVkP+FATe27UuhkXlQxoDB7OgTvinLem8cQDD0/7ez1iAXE47DWclqZvwt8y
utZQdwrf24+/5Y1BODWoEjwOm5EI6A2By7ieo3utNGQI18Pvz92Uy45pq02YKPCHjczU/s/GYdoI
yk8ig423cDj9/mH8Zmg7Qc7eyIW9dDzzivc/cVNiDg65kFE6zrbJVPwe9w1s/HzprjHQnLCQwxOT
Um561ZFsD5gYnLNNKfM/xWYuExMgewvve/m4TLcuLBbRUFvhJByBvUQ/ccAQ/ddFFIfgwaSY3jW4
eh8SUN3pDJ/i81vCQk4/d1XsTB3BTq39jxSrwfK4yjW93ElU14kSIkhSxvH3oDCBozBg5/AVsUAO
rOlxxlkOHVDbGDIPB+sorCGbWKIoiu2dOfOZkoCH8scLshSvUGyceP+yD53fEOP5P4O0AKuehkFt
FVe2OIa25RW9Qejm1XopzjGkwylWzkRqV1fbIlOO+T1aXQNWpvTSYP7q+Krgm5WQGpG0TOG/ruxf
Y//kkX9jew+duSHyWXDzjDHe08c2fOm7AvQdlmxDgN2gd7vxPbmdvlW7MAMO1Gcacg+4UJGoSZ1T
0rScY+zKLjnNjWeJR2T0MwyKIqOSbc0bZNbgoJGWo07CEnRV1a/YkS2q9KyqDXVRVpgd9NEl0hCj
TtS/6dLPVlDhGxzaIIz5loCjnA27LRxrS8NYioFSZFdnN2IeGOHSGr9cy3EitlkeSNFChNOQpT92
9KENV8X0G4zUsGvW7tSM0ur3i5tA6PdFvrJw+TwTsabeqBgPoqlQK8/a84EwqmoJEGM6fQ/WA0gz
cAdf2TITM36VNsP6o5SvsYymdx6ZVdkJhBAHzRI2WaN2yNaBqZ9Rqfog1NvxDQEyqNCzw4bFyQJ0
qdDgiYwoT4Mzl/KLDIBLm4q1rIGIS6bJqivH0z8n/v/H3SpbPk/OOy+rihntZMqLD9M8zlTGFv55
blpJvMz/OZvO7DuqhLNGtXFRO27ioUf41z2QDZoUhgwT6+cxvKCzNWVhhq8eIUr1oSofeDMQVCa2
CAN9QGB79PmyLZZt0s2rAdQQZadFInca5vYYCaV5V9Ka/FpdriAm4wbgoSqPXg7zmAAKnT86BDFZ
6cEN91DdvlwGVpC/rpC/5vB8KPGXS6dChaODjcibZzhAl5tb76WFjJuBi/K+uLYVVbyU7bOU04fo
hnUIdu1kImji9uMxlOl/If2Jb5AKjQMrfUN4s7ez9Wd2t15fdeCAXX+6lDppdc5WCtifJnO8hGYL
3SjVWE2DihQvKekIvi3+PT9VJisZMdg+t4UNbShQ3zC5ISXD55XxnKKvp2zQeXi5vtovldB+2ciw
uu+t5zhfh3c+sgwYXehMjXYFXuYGYrH0cOURkUsqKGHgSo3/1cF8j0TOvL1+Dk6eAiLbmEqacyhm
qdIXXtMdRc2PdiCKceeDD42xiTyihyRU2s+JoCeNwEQ+0eSRyRJJXOHyE5xsDwSPVdzDstV57RNM
kaSrFBVxG4oAC1vLi4CDi2KO4/UYWjC3H7ZtZEPLDheIsOTzY/X2JHuWOD6lhEYl/losV21uj26P
P4XkkLrAEuaj8IpxlqwLGeA7c7wqxNhr+3mKtRrCj2C+FwPSciwFHhYkrw4JCC9o9oZbpjwJ3aMX
ID6TV4QEuw6lbpb4EW+dLsiSyCk1QYicSVLTqYUfCLdsifsYGL2AgVr/+etfMo+3jh+vyLYfB2cZ
He4LTBY32qr+5gh76oIee86xZRiqPqkbSiP3lN0thNb2wXx+KBUiOrJfCQ30clKV9myRVQseNRa2
x0szJFR2QA2mtbZJRYhngHxUwl80G0vYObVCRrEN5laDuayLB0ZN4Uz43sFfeMERS1zbip4b9C+5
frQAUiPyiQlCoBS8PdW71zTRvgUSphr2QbPsNfOPcS4Tgo+nCweBqGsul9te1dAfq8jaz6vtVRDt
JkAy8VsWvYm4IS+F11vd+q0ixPSCz4rqBHvIpqSW80HJtj2OPs9AVwZgO3a5m6BkowgsYaS4/ii+
l0M2AeNl9ruUXfef+pdqyNdcxxGzUG8EKe7n5VGlA+y6lWu6E6wlzjsTauUsDRfWKC35iZou3eWV
teUmBb1YaKLmdl5qpZEnOWT8OvdeiJvFPbic0vL80RzpvmUXLlBtoiC1Z0HnIoYe5zP+hZdTyzKQ
VYKe3SuAYKAhDFDPQtonzjACPftq/6vrzUGGYkatz+Q1kZE7RLP9NT9lGbkqATcBxKRCCsKNu8zr
Ctsa5evbpUTiCBwCjlmO33GFoDMk3tYOa/eOS5ET/nfIn663giDJIPNn41uXi6znqC1hbiCoPi7t
mEjDQwtSpgHMyqNJXAPEADoZ0MeQ9ZUWOf9qMC36NcQfZczhdkLSTAdBfii4IH8VF9PJswe4ls/W
oqoJNopmBjyYPvRJALkJNUDLMG4bCWIqpt3xaxUoGCykNSruQB+Orb7Rothlbj/DmgvrVvlj+/54
rFGFWqG9Bf1u4zABehF+cyv9TU+aSbQoFl5X+eo6e0zubTB+jaTpmDGT4aFiGImCJG4dnoBUL8/y
aJcM+B2crGj3dR3M/xrEfomuGyfqM1j1xTdhTNKwL0ffpVL0jgekp/cd0vFh0zvCoFPuZ0KsoFcD
3dNeQcO9X1uPN6FHaO2suQZODx1IMIKiZUt0Z0640kx1V6fTwYHJGSK+3kiDp7RdUlDhzNKUjy2d
4GqVdOsB85VkP0bfuyj+Dwg1io9ffjbeQ0na90p1BZPSMXleI2uYctl6/2X59MszUqEzLl13v+T0
/+XV7IXa8JLU9crxXNkVIfouTOyBd8e3U9666m41xHAiK9fpaAxSZ0WvD1onGtdhvVUeGFDvuXBB
MGlvHnCfGGddd4o8rwERlammgqltjidVbHTJmK/3iuMHu6xzP9X2rmIWbbBausAMTKbCrB7Ued8+
rdBgrFKkHaE55uVwrpEUNKtLNGniIjeQTrrhwep4f7Izx1Hpc/0kvIEC8zZUBaEVpda2ZtZ7xuug
zAPgylMUFY/YooJGaqrFHOpI4sIPzAC3XccJ/Wr7DFM9NCcGLztsL/EAbllP/p/FjUav7w+KJsEv
VGM91BQkhYO0qYTFy+NkDuunKsU5QunAbfyQyZk2NfX30ysWsafLOYnsQd6JLML4HtS+5owYExdW
rIz5rBZ1HaiXqLE+7yQ+PrBUMeji7N8n1bq2v2388S3eaZgyk703sarGoKLyrdkti6uom7/6RORB
1y8xvu8XfjEAQVFHTsRPZwXEEaL42ZUxlULHhq4DLpvQnGnXmWaQ1UwBRVTRpxxKqX+QJdmGyLMK
Z6m1Gx49IyUq6DXuC95f6d/XlM30eq0YDJUuhhfFoC+f1kvJKzu1d+/hohQrECScr+aNfjz35GcI
j1eCSBv+IWqcX2ZgTqjW+96YGieVAJ/mRZ0N32RrLIMw6duTgd6OUpSXpRQ0qeYnOIlJ48iV/K5I
tpDttUsezrNezRaXNjfJAPVUhASbGo7C1mw4tDMueXoRP7ynHqPpB2kOUtQdxF0XiTNiH2gOLqaP
qc0ontQRE+68Uef78ONXjXVPiX6TIIjt7XAzF+FSGw+k/U5g63a67xffvlrhCQw++UorAUIvCujT
XxO0v4YhlKXJohvhBDVcjVzTw+cJIxjFOB2XCUbfC4CZak4lubYGrjnl8bXlhttJTIHMifK2eE7c
N5KENAc8mvhuzKXGSrswJPJHIeM4rTOkaFMS2RhoPvPZ4EIGB+DC9/TfPHuKPm3bBVCXHSzuWtx2
ZMctB7I28LeMvudApQtML9MV6GT2iZOFOSPP6TBhhziD3kBwML9LyU99S7XtA8P+aA5AvFVswl2W
dmv/V2vmbDP+a1DYAJF6COIcdpMXggbcCBD+9TMsamIY6fUGcpt+1eEJZDsp98U5fbh6UGGukO6f
ZjNKtx2wFwYVM+dwaVlUqrAx3y+vBciLDanr+gm5qNLRmuu8Dm37j7U3oJhBOLl3+QrqMwDKZBGD
QWPnWLmEyNfxJKCcwqn0J8RrULbNNsT+3tlRRhVpGbYOhuDJFmGaY4Mz/JFt4zDJ9q4M7dSl8sW6
nfLOT5LWGMI/3SbVLVOmy5fFOoHgSwj02bEgUuqQ0D2u4elUG0Ee53otxBBmKvKIFgklLnMkrtDu
Fz4KHOdvWnmMHd/pFjh3quZrrkI6w7+VYc0Uzlkgzm7P8zm+5AYoWLi0+KH8JKe/JLP2ZWmozdHa
VEasfwaBpfEG95emElW21fHCs0bJD11DShovlrnYmoZjFVA0gjJDNG8isdMHJNmKDNsQZejMyyKB
n/IdLwQkb2RVp32vZ/9ZsVXfCgvnWQ7qm9X+R+RViwbQmelRXgXfSlDGKYQXtVSe40XhnZG/i0hl
dHnIZwlaA7xnN6p5a1LqGKcZuJU3dqF8+W8ghhTzyLcVlr3NFpA2i3zdHdbFUruGKCRAkKC7CzlD
EKasWbsW3DJ99Wt1Omqq8InfJs3SIg0s9oudHG/h9BbLTuzCK11CVs0LJeWYJPW9iuhPYJGjEHAh
TU9CXNZjar9ODpGDUFd2m69F1Fq5VRiY6TO8qqG0zj7/p4iOlzQxI5zeV2wayGNHFQ+naMi+K7Wh
pKcJ4CMTYJsI6qZX4sGk2SklkjcyT09WD3dTOw24yyunTx/yoLv3TKGbqJYBsFF80Ip+jW3T7TKN
zmlEJIp5GzJJCkI4/rjECWI+X38sSTzBPWpUd3plfYv+ovYUh2RzcM7s76yDKVkhBcYA6TUT0q0K
lYmLmQYRxncsQgwiziZaexlnjBNj99ustB6Vq90lPrJ0DfjdPYW9mn9LqZd2Kb5Lp3QYipodXbmN
O5jtCXyi05lPdAeqyleJARsOvUHkzsy7Pi0rtQ0LcVLQvcIAtw/RDtfzgni0TVxxRxaPDCVSs0d0
x9FyUqLqlxCy/Ch7eODDkXaAd48yflTX9VrEBEcGTkG8PJ9VJHKQZiCPAu7h0d5Aqc5NJVFkEtMC
KYm2wbKridGD48un4rWlWz9akRHjTCvyPaA27rUyngfy5/gNbsbEkZvkVTxCkwKNUj3xgWyKeicC
pCXHxVtkTBiTaQ873UyMh7qwpZUPi+5+SSYUQIoSJ5qxEs5dZP3azIQZkRWDuABswp3wiiiyjT2n
ta6wT59i4KGXrxdCG/qMI3rDCQSPGlcNkYoCuhsHaTiEe9eh44IgAEaeHbMKH6lnp5Ku8J2XCK3E
do/SjozUkrYnITaBuBpvgeCS9GeZw2nNmjciIZGCIpqzKn7BxC/qA6aKWJgErzrbSTJukYA/O4Vv
ABUYPC1UzGW1wyZDyisIDMa8Q9H3QgVdwFQp7ED5BbsE0GV5hqxGrVHpQu/tcXA/opwRflkSwZ+K
bwrrxD62noDVPk6xjXu8GBzX5/zyQ7Vt7vSq6PzSdw5yJl+nce+IZ0AJfK8oUlLJKTzsL/k8DQKZ
SOqoMF53ezhfu6fJVj/9dBxjajAYOKu38IMiykeoHA8q0x9FS9wcatCAJsBjlDNSdEVIj875tRLT
NOlsze10ytAtW7SSeFk0UyI+Cb2JVrIq6VsPB3RuOtMt6BylrX0Jua0Dm/nUSAaOwWbQaHypOp+j
ORPMc+h6QZ2k3WsGaX0ZOrRCSTznFb/5BTrZ9ZREhqWdlZS6Hu8C7asI38+H45d0HLCuE/hhwzV2
sEfGCAkJsNZDs8Gxdhvzx9n2DaKRS8FyQ+WtlGx432vpA1q7prd+dWnrvElv8hAhNZFvICsx2p8e
lp7F8by5W0aFnU4I4FfP8o1zI1/c3ueTU+TNaNYReEzuo4dUt28tTn2e+EOCNVjxGizrYMrIgB9S
3km9Cb1em6Rn6dIRRlMdWz5GfGMICDuXPB+1PqW7ODYopOqMeCUnlvSJTJjTLxCdl3NqZc3pZOlT
gSBBx3ilHY7yUUReyZbyuy5DmX5O9Bc7eslwatuyLu+LTXiJi9YiF5MmbaHI9eqEodccxjTc4eGv
SPP+aMg68PPTynRYXMH6MRP6LszRxqxj6BmptwJma7ETiWv6aSO+KzELsXSxvXOdkXkOvM1D2zFF
nCFkwMAeh2EQX92d3nV2hiY9tooy7/1eB5DvNob9I3EfT7+GKZ6eCoopEzQSnm/McXqW5lQj3G13
FvZWEaoMcURIA4+85us3X1Z3AtL2PEOfE09thpo5T8ObKwgK+YIJzGkBnkRYezkyvkdnFBVEUNiO
COeY+dvtuRmbYsPQG3eSTR+WJ2s4cC8lpK7p+inUZpQ7Fis6fQsUpfn3htY5ewuw6Z5qI8WIOoP1
EDgyZQEZ2Lu1TpdIDDf4SOez4lRaOyFqr1b8eCzjdWa2fbZT409qvnRNrvBsRQz25a87neyhHq48
jXvPRi2c+iWb131qRWMKDJWsp8hP/BhOtU6ZrgLilP8affDQVV9PiAr+CUqJhHCzOb9RzYwaRYER
aXNiPawjebI55y8n2QSe8Ys17EosPnknCoRekyU9rkf6+CcRfKTt2tTFH0+QzDtQK8WJZx7lICVt
L5JtJIL0Na4KYycOk0qRM9MYQE6byS590VOpDnWO1jMWeaEAgD7q5k1CSj4Vnc0Y6fOYbGwsTcws
ZjXgubTrPFoxmAahteqnpSAlGgWnKgiRkUrEGjbJjSsIgEVyV/FCecpwWPFii5lCFS9CbJoquDpb
JR/dwGzuR4Xke1DicoyWlvisK4trCGzGgJ5U1CS6bAqf5GyDdpitbvEjzcs5fV7KayF8vwoWvD/0
xAA4Ik4AcjZlF85TCzrZU5UsUqgw4f6WfmaxKV1QeOPbN7v9yy/C6XYw/htdiezwClFvyhJWT8ry
ZbCTg+kyBEf5VWxSgapKjqS8qDxjb+0CisQYVxego2lmMYdbUYqekVY8tM5wGxQ47rFU0ApK9Cku
dqJFaETf4YTg6cSdwulq64lounl1JGYfDbIYlYK+8krHG16armGYBC5RNpOw9B+YaHvLgQE7xnEC
yM0QanVspsYtmGsUQ95kT+Ksn+UwNkrMXaaipEjOcHm0OjUIYiQEkpAAL/ZqMAuyZG4wKj7C+cE3
Xmk0jsL/Rx26SC7Po5M2wAYZRyTXALU3TH4fIs18eCYU6Wh+fpzKe2/KRwoM7+dKNM7DQD5BuzVe
zpODvcMDUTB0aAY05QzW8ggVTIRQjYjOWZmKMjx1T7Vdcdqj3Um/oMLM5CLIj51ay8EATr1TD76I
y+KH5c3HnYnqIjSuj0ACKzxRvdod52AivKnoKl0YtovazoTSh0bTf8XevHVzkn6+ATGP3sdo6auP
UbGpfMVchSqu/TWIm8bbjB4QPkAFPkP7QLU3LrlYLTkVpZ5EyhJjpk0ZC3Ilj4K8yD3ULKNFwpFf
/90+1oppBj1pYBruRe/Q4+OAIRRPEGPQryujrgO+KjHndjBVKONuwWAZcz9JrhKh1KFC88mkSi0L
ul9fkbkTCOj2p6r9nMDvxJlktgO6nmmlFj94X0wgKJqVHiV0MjCNnKxLqKX5A48fXTtwnbt5bIjU
mNjcXmgx+EjDpPxN1p8x2SnpMincNLtvXC460btdIbfnQd4KgyX2yz71RMNoEIqpmpOnZKZCftx5
2KiZ148Gw+Y1ADd0DzcrqnAmk/gJfSLvd4Nn9B4WSARiUeKJhjeTX4cB1rUqvfkc2exNXxpT01vL
XXJLjj6bMn0tI1i52PCTw06sboCDt8ScA8+vVYzB2Lug4SkjmkLCPfChPJ5oTHiYTVK6nEiHyUkR
duUR5mqqq6pWfwx3AV2OyDyzHzxKTmAGTECp7jk2AAlr01D3cwGT229Txrh127zqocHWwFs5MBlY
tKu1EBwJ6pmzK6dt475MuXSB2zwYKGKsqQb8yGkYNrFWcm7YujDBY72Y/FIvSh1FUcyhRencKL/r
wDWHSycio1SHqycpx1UdIlNFqpNUbJDHQnT+642xJJ8dA6lWKHgG3BaePCaneWC0J+9yXNFIxJ1K
+YqU/GrGPZdMZ9cTd8f8T16ZPzf5l89F74MzIYbxma+OiDk5cHUCRAYmxRqoXgJucB2mAP5fOJ9H
YSFB4Ad0SaELsajsyH1AsaKNoQ1JIygOFDjJYvoPytJ3emV4kO6DfyX9Plo2h+i7ekVqtt9SzjNw
+4eCDH1QJBfWTCyNGgG4Qlydo6eHUb6dy2sqnFPz7OOy6Up8dK/IbtLgCCZ6enYSYGJ/BO0KbRDH
rgGu+8wMUVYWbLSvVt9Hc3kIw7NN3fqQx6ltGbSmZU99K22ujabT1cDQfYTolrpeJW7XfraeKwzU
SQ86HUEFcQsY4MHyRqKU0831g01pJGbKlq9qQSjc9mH91DprcI7MkzKAq1w++7eCbhLtmU4tqA9H
0+UlmWNJOVdzQ7v1Y40lM6Zb/thjE91E4rN7/AWOObb9AWpJ2dKSQVsww75WkQGw4uks3oaM2IbK
4FN0G9rAFJ0yEAEjIRGzYEe7wBzgNJ8UomjnjxPGFW2C8ccv7p09rXPNNB6rcXP3zoOOf0EP9lJQ
uARjmgG7UAL5Wd4kHr48/tbNtUb7nCYudAqYVzpk6lziF+ZoQxNV1OOI44fpuTR4XkYkSkWZA92k
Ld6HTKHswV8l6fedRc3OvINrqSgC5+lpsuiO6/bWnLX7h1X3FuMoyFXr47UEenvRjuNVHc5rScv5
EHHR9kz2/BcUSK5a6eTa9CRiFppe5Qp8reA9TkaSh4XIDpDdY36Ld1gw5wdd+PuAnwRQ1e4EJgjz
o80aO58fC1H4NaCf6eoN3fIsGODslelmAejQDs1t5MBitr3Rnz9U18O5xvBkXiGIuvl6xB285+c1
AV0TtMyF/XKBjmjYDo8Kl9BBLtqjNvyCHWRHDiFI+m+WiTZViBDYtqpEflSBkb6XMKQnqZkdWg/G
0NSLU33wfCQxnUCwVnWz7W/RNrMMBgoQsCHJ57iGUYztP+A4GZw8//VtPbEI8TGVWjQYxKKPBqnf
INo7WjSEZAoxd+nvIEKGbZIbq6IqQcphraJGA2PqHc2mxGYG+Le3NDHBfGjy8u8SV41Y5Yk1H6R1
+W0aE+NRaUMZJ7BZWkkFWG9G3D/Bok8owCI2GEacVdffKZTifkCma+rfxLhEykF9/o03AeFnbI+R
XGLBst8nwt9rKYainq6LoPhhSBnCIMT1hYe1jyjjYK8odXaPEDAC6DlswG1a4plCjPvhMAemM+c8
DzOtX7r/h1D9mF2fP5JsOKOXAUvLmrToALFEo71pE1ynEL0mff554f3eN8wwXifa6F5lCV1t5DSf
z6N6e4TSmjPbsxYlDDPzjdrSAKLCwIhxh3XQmGTbTODCa8/vJZelBisV2kI9gCP9+Md9ZvCUrssk
q679rRDZs5caeyoY9SgygvcrjX8OXfQXIpTkqNcImAjn8+fB2271/G8oBy2PUc7yoIyttrzTHJXa
1P6SLBsfZCed54cNFpEY8XHFBzambmzuh4tyeQzTVKppjyKJFYZnpDyUfCNNIjyKdH9TItCrJ5km
uabyW0buk1shBxLzHTnxlaGHkHC6MyC2XCj+kn1RU7e6mWY1H9+zWeJ9OlNKhw1Ku1ddFwfR4mLH
JAUw5bL6viFm4lmmGGH5kQU985+SIdtYrS642O9eVL66DK7DHwCX6aEZZdzecvuk4S+B0GzV/YyA
Un8l9N7hLru8wJwheH3ClgJadGoIkWBRDFu9bGWZiy8oegZJo4Oq+YlhfUFSVlGmpv2opgmLv5eL
NyQQ/V9KpGTZRQYgbU9Sqc1iJ74VizM/2NdeGJrEfn2jjfZ/YyGsVehJKvrwj8XokfG7hKfN8IpL
MrI+sw67VwPEBDdT9w5ta4hs4LMns0LG3BKVtlx0BeQUkRquUQoL7VSZTyi9w5brMk+BpAxj5XLF
9l9nV9A0dAbwG1pAS+1f7H2ZYhFk5hWLBfzIg/MdFKEhfygnZdpSk6XfPDKCQV3yp27QRxdaXeny
AIwWnuWR3Vg7+8m0UUke96LP8Oz5KT4jFV9ljltzt1mhpiSXYcSpyDRnIGzop51bTy+MdOjuitW8
0bXpnYjxCiumaOfdkx4b9IaHB1kyI8Jrqg/2yFjd0BkTtz1L6u197nl6U+igI1TvA57V/1/Mf9+9
ZQB2W+/T0psOfei84aqsbA0aXFIZUy7OamOUmH/bmcZO5STY3E9bTVsLexIAm1OYyLkqiXmCzUcQ
WHle+AjUWn4B1pgQ04grjtNHavLIZCfvNL0Qr46Emgk5srbWvgajkCfihlfFB0trTmSKxKj5SiDU
sj3nNBsWD6I8ahMqRwy2GEijxU2XJ2ay1FtmgS7mELEZbzWManBbUPLtlcFh3LURDZc+fuJjlYjW
T7+yBrQw4v5jKsM7faLcDkCES3pV/HTFAJBc2oEdf3sGkTdu3wHMHmLR8DGgc/OjeD9rcFY+LInt
9CeiqYtmhj0rusOln8sZd/9ZTCXGJvJNUTu0jCElvBHnhj6WruSFTzJEZq42maLoLIXGe184jCU8
ypGhfyoecYIEG9C7q4ryFa/bC2cVLIEaYWlwnWehkw3IVM7L1GThWK8S1Va3yzByGonYM1snq4/1
KBlJLuQ/N/5xM/EqArTBBjapirBbyzFVpALIRIlQFxbZGH7JPgbFIOCElgh81EmlArYpHgJGvBe0
rDijqFrb/kSkYaS1CEhrpMSwsSNCLKkI+W5QPSOW9l4/KGKlbg1jmRN3di9pkzsAYh8LFBJYUh7I
hGBtIuYloOoL9Dz5KsWSIQsMgudH3j2JFSHM0kTbZObC8gLDnmOLOR2LnrUN7lr5158NcSJgIQ5J
4jmenevJl+sF+fac22BBFuFT2l2OlXh4LwIdzTPGfAKnclng/VA0Cnal5zX0qqeRBC7mXtLgdLmx
KcxPIf7EJ/Z1pUG38bgQPGZAO7BKfrZb6hhvRB2rG/DarADGcXaiZG2aH77wcqMLkMhOrq0JqnTB
oJgz8r9oJGC+nrjH0OwWZM/wl4w2zab0Vs2bs+CrjVTOP83k0+lKskAfHmXTmmwF3pzatAxv1v7l
ijV4DO53T7Yb+K1vsS7u/iDq7GkLNwInwQLHi1MENIrUZVD8Ykhnl+MjC1WOTckGSlezntTKxpZ/
1QF8uhcNxQuAoJdcSQcBUpu95gvBlsp+VmTGsVDxWtIakxMleI0WcW3veeVn1APOWBweopuSJv21
3QZTsPR6n+nyG7biqXxhYUzysvv4pD/ywtalIHN2RTXNt7bIxs617aZKt59rpFzGsDqfti7k7b82
sMKDoHPIhFtXnOkzvCY+J+FIy6/k+4PTo2QRXwcA+sjeEYj2TiYKUxNpW4EVsfwooqtXFCQ6QrD8
2oB9NE0I+bGTY+SnvlttkyCzJp98ESxvwnfVIs7vyluwQrZ7vTlquC8zHE9j8uDOVz4TizV51VEs
Zic925YI8JxjdPunH4BXlN0rLAruWNc8Mop+gGHlbzia5pzhzgKoSOay99/e9q0ij2kE+NEFhK4A
PEQCBCZ1uA1pySEd4+ah0t6uxpST4jVymVsr6oJBWozb0Q1HB2APxY2KPUhLVERlTRXiIASeuW1B
nwFqQzlq9bQfRzB9PdOskCi8+tWdIGXJem2xLRSO1ZGono6jAleJFmh0E2ub885hHKoTOqeVqvfC
bdLDlkJzQ4afZlnTn06MbtOGg1rO47NrvLBpIxOYjSKh8BbHVJh4mnFI8F/nDt+FMBMlNpPCcTDI
xGIujgbk9TBG7HhxjQuUmdhzbvVI3AxVLQnc0gahOduhKv0bzNJOrQnefxMG4N02J01+0TA8Cyrs
eVnuL/1wsb7eJJ8IbnyJY2b34YsDpkDH3DicAuvNg5KPDzSeFVBKV6aIRF4NuaxKadQRrn7G/tJX
/VPCYTru0MnZV+E2t8Peu1loB3VMs2JF2ggZk3IzQjv/hwLDBtcCGEvzuCSe+/LTqgF0OROhaAnB
rqLepnZGe/0ygfuruNOrLSvQs0uKvq4PmFt9OXwS7gsY24AGaLUtvonCChH11ftRhlYVAsHvugCC
FPXcn/s2s+kqj6vlcz7ufescZL8I20o1DQ5lVB1Bx53OasHR4Q7iNxTuhgW4LhBaI8n8U4RkivKQ
C0fW0jwQPsvh5OvCU08E2fAFLhpYCnzahy2TyQB2/2Lc+8MxyEnXyUvBEWGwx9yQ6PNWbhQSt5Ch
mdfe64wmTaKPPqctu9n+xOeNIP7y1neMftKDZHeT5d5fisLvCKxmqo+PJPs8efEF7Xcd16qfqEQQ
mbWogdNXtr0vqeAFpm1jlCZsY+lm9G/meem1hPQZfiFHJAls7P5RSZYXsFU9DXjxD2ujk6SudYAf
8KONyHwdEJtSRwuB7SHgOZopsW+PD/Hg1iUm4p7/5HpSQHyaXT4fxg2v4BJN/aAx47N9wrckdWJU
GOrQRu+E/ur5izEqR52GZeD6QcdL0EdaWNsNQSNAO2hAe4xFOzfJbGj0n/SFXZbrfldM5vfq53Td
+on4BK58CTjDZBlYXhdqXjiL4ON4II+ya0dqv8ep6nPORn8ldSgJVDZRe/uOCbTpyGpcakhgww6u
bk8qbyfXpM+hZ1R+bR+LzP0O8RFf/yjB0mBeUixiEEb5oUVt/HrAGtjLQpQBwbWZXL/pvyRYbi2d
ecwhyKr8qv9PYBSp1dFBS9e9EmujP4MCTz7mwQG1YgXdovKqQr+0/nE5Tpp0/Pxmb6ZpJS5ykks6
/B+x9xrLMNrCD3OR+4PJf4buCfvqJTRaGdT+GwGun3Of1FRJMC4kMTpikxpn/tS6TmBqTaHvO2NB
JNtc+B0GAqSHUyVbIZ8RmYqgvmx3BS4Y7NcW/NS9GoMuCs5NLzNUygqKE6bYdSgCL5uPgYxGxaSd
LuBDjutJBHMr+QDAmbZyK5Xi3gFJhxEmALtTV1Frc0Z7ZMNMJ3FK+GgruB24H9VXbE+Wshp139vl
J4MSAeGc5Ml4VDoydVVeU0kj2vlQ/ihVRaH9KwcMEHaV3xKIO0pMtQgx3LB/KYCfQYGyEqEv5BU1
rPDzacA6F8QLRokhv4CvuBAaO3iSAsc+HjcoIK0xvvADFfn7ipkGDGka4QiTRjGPoa9kyLOA+eAk
K84wOQtkMMrtP8HR6aDiLtxawLEuxcMDeB58pn30vv/vxQmwgecJXUaBgBdJ+KpqKmyKSCma5Ucc
x8vo4bziIeuKVuvtzbPeAj/9V4hmJ+Zul6ixug8DNIzwUlUUjoJ3/EuB76xF5vzh+MKOiNDGLaZx
RjCOahgwh8T6M8ckq2rR+bO/p3amvdRC9YJh6u5lrZ4u2fc/fUiChYH3j1aJwmy8N/DhS+LZA1GR
jkn7cD9mdo4F/pHzayCG4jVAOW9dadzPbVRM9cgb02An3FANUY5kOXpVU8z0B1kdg1pUDI7QIt/S
SGb8OjKNceSPRfcCl8Z6kllsUDwvnF1Y+6xghAiS/ERVrRiCOUcNYBTaJH0H98Pqsw65TFQLROKS
uEP0O0v4X7iM6JpkTEpsbqOXkPn4hCStEuyfXr9prNoFy0tKGfGlT62fCJ1Ks0ptCVQJQ/XOBZbz
reBm1D2Qy0BFh/ck7rtBtU9Y8cRhe55WhuvDOTAQZsaeixFl2iZWZRuzsWeOcIFzjKcAzdV876yd
M8n3Swr+dt7xz2bOvP1P7BI4GIbbzqpSdgH/NFRFh7wyJqNs3vw1hDLiYnf1QBDpNVTyXre6GgtY
gygSVgDAx3H6QsYpNl5Z4zvO/F9eE793Em22R6m2YpD7/wZ9EGIc6R5r8TwomrrUmGWvJbp35zNM
9AQgEPjMV8YL1BoCXmK56K3Xo5t/w0w07QyMpnx23V5U3iN0vN6hCWHBX46LCBD0p0OwLenPODTd
zx5nH6EDhqhuAlD7vN9QRzgJY+MZFiRtPCDJ+EdcXRZqRFYtJJ9Uz7FUhCapP35PTpJOjc8fwAnk
XufQxxnNzp+l0/e5GdH0Op48paMzgnG/2+TGm9TaT6aLWcxnOPipEFl2oHPPqelmQKxbBPBDBRjZ
dILQKSePVkYhOlEjguEyA8qcTn/nlaiY9zwWPJYvs9ny8beUny5o7DlkNtmDKM0n0PGrWoAeeZ8w
vFs1+fw+KS4vKHLUrnuZDSNCARxGIHyyZmQA8IB8QDQ3qoiShQHvEq3yxuHUPuR97ObjkN5h+9fJ
S5d5CQKiu0cJFK36VQeo8nwPF8psjmKDQqvaDHDriBha6SIWq80b+NNP32euMvsybjF+q2v1/XTw
VmjM0okr+2aq6o9y1PyH+pzWiozoBm12/BRdLyiGFS9jPraFZxnvNubshpcoZwp44Q2OlvmFA+BY
epnejqyo9qzChidWnHi0aT/vsFGpoRgthkf5pAqXMIaA8VUACURJf0ytN3pMP9Eu+lu9aD9zKux9
ik//Z5Sw68NyeomMICcBd3ab/31J8JCybwOptXZtbv6CSRDh6ZQuBbU3IOUiolhFFaajDcb+OQac
62mGNCO4pCqcEpbKLljX3V9tPl9FrXPZ3UpDjBfF1fRP1UvekiO/PZ1U+YIb+i06o/wdP1VB3EX7
3PL+X4lvKq1Mpru0iqLTsJLs4Xuam0lmJELvcW8/sKD0mxbvroj38vznJXLG/U5gs3cwv3DykmUw
5qo84DCzq0AGT8n1uCsoPI2ES9qcUUKUkKl8921Mc+sdhMvNgAr2UaLPl0Jy0DSAdvvjNQK2XoS+
3LeRDSxDhQQbwUIwvP/igqpn4uc6NUTXhFIkW6RUM9meA8n1skxs7SSMONQwwHXaKQVRsteB6PIZ
gyUyj0bO2tbx8GCWqN+6vOWmsMf8o2AS4MyBnnpTbkpxJYZp8Q4/dMPMT5b7U0QyCS0nem3FrTZr
u5wnz0dNsm6aGVbp4icHtbezACEu+DhIGowh0oSD6y+jDphHtmG5vQ/aLCH3VFkNOBXUV3vaQtRP
5u1io6rtiJ64qxzugFkbEEfXakJSrvDwo9rdPrbO3hMeBRuCQeSaFiyECit4mRvdLCbv3y5/cehF
PCNUnlebMtVMoBLYxOVO2vLNXINW/uKNFGT8UwqBFUPxS/JCAwWGksWC5sKv7bUNJluMWC9XDdvN
Fwj7h8cwWu5IK/HHA4jzOI/HvXVASQPy8SZKPxa95LBYGw09M10l6wvkoP0QCuXBx/EoUculuesO
Q+7obdpuK21KjvNXMlm6WeLWwQWjBXo6fBW1/9waynKXmDvaU2rRAOiefBmImu8usa8CimuZ9KeW
gAVar+8ztHn71dOvszqwqK3Sz26zEHT3cGBocTbgoiona9xBJlDQuEiM8DluZMwFnlyPMFneUZZ+
BhOfvUDs+21spDkB3zsxZ8j8yb1HkL9YKVM3iCQ9XPXKlM3xMPyftwmeCvCX0thcAYzRUZBHZ68w
WBlN6tsCgIxgSaUNoSFqM0KawuLcWdxXfB9ihtYhKTHf/7J3MQnH/CE64+/p5sUzBmw2M4kyXyVN
1qCP5cbJ6yMhH27tRD1ny3cmFc3qJSu4Kp6RKBzfnoxNog/z9fOYf7yIM2RzEdNWOI0q9OzlvkIA
sE4HPFiRLlDvCuoSf+bvmjAotxIG2pFyaYOt0p2AbWS6ce+zrZIWHrqMVXr09kZZ06/sjJjpIqHe
DJQGHESN5u6pxmxeSvpqycckP/oX4HX4zO4btTe8rnZtzsJmaJ3Coh/jQ6UO5N/q0Wy5qomxoGQd
4wT5QDdeRSkZMXKsbwJ4/uSVg/4qdIhENDAZtF4G8kVfqhUas0JPkPTsHvxP1oeLHQ+4quw4RK4L
P/cJR791q3VFaxTjD5KiC4xE/0nTvTPgLvZEZtfbFbtIUwWNsIqAlSmKqHYqXtsHlbE7Jhx67RAm
Ott2D5uxcox4Xpfw/zqnblAr75m7yKh9XAQApHJuBgyHi8rBjgTFwMAZBe41oqMY0+Jtqwj3g+iw
MJ97YBLq8RpMMTIuEDwzUtghcYsT/QfMh4ZuYJ1z0ChIumBGwqOKhIY3nKGp5PD4wpfSUZx1EY5N
IKhDLZvktm6Or3+ONC8Gs4wZMoQpAZuif/7l9d3eIX59OHFAUR3YPMrO9yaVqcVESylMJXLYl9Qa
LwT0r6K8befD4cw/j1XDdaQfFU2g/wrAW4CY2rAWjUcTSrfRqV/1w4GgzvTWs6xIK2RqJRjMM+5U
IivUIqGjxZEZxvZcFM3HQg+kkmbpL+W2G9DX0+LkimKqRENxcVY/iPk3uBMPL2yAn8ggiE+jsNgJ
97E0fsHxBTD4a5XJAlmDyynYj36othWj+1cuu6zCd+M3wm++w6yz2KzN28Y6wLhGDfi1sDhGNyiM
vQ+ZP8QYIKihKGLebO2ukRQQcHVOvv5IIPtvfK0jhssaPQ8yj2nSFU6SHPAgg+VQIa83ypeypu62
CwyUIwME3GWR9Jsu6QFH04EJ7kwPeet0ws8EAfd1FagMX8iIXC4b55N49BMxXTZKfd5MAZFQ7d0B
yOy5Zf0iyvAaXYVxu6i/aDh8d67wIBeMRSRzbkjpsE0B0cJChxqXgJD2KqkNwq7xRR42rM0bnN9z
qxC7g9IEjtMIkpgIims6Hv0bIfTSPw3GkDVbx1v0ylfSpEferMVRPrq+7EZ6sKA419xG8e/IQD6I
V+fZ8V+geEiEbK+hwiqEtDRCEVq0S7iCuypdJi3n/TnaHqmTO9z4/xHZyf1Ywd22T6xhV7KVbHhx
b6Tm6jfwumnLeGFwkes02zJmtmj5heOnE8ELD8hakPfY2Ll+mjHMElXgLr+zvPgKK0oE1gpVa6K0
DB1HAI0QoP0xtZQCTwPS+i3x+b01clqqFJGytYTgbnigOI0qwz64d37zZXdkY2dbLyqLP5YE4S76
T1TsvrOVJNNzBWIZkei8I4XxNt0UCWJ177M5P11Q70XSKPUR4mL8g6m/+GSLctodJljE2fbhCpuc
95E/pzKRCr0VGaEOecp2s05Syiq76g8zBxBgrRy06ge/0mo9n0gCCW7/hU6Mx9NlKhKZwlfIOq8v
md7iGyPbZPjZwoVLfzr/cUo+Ae/XiREAqRWJAc8bHP3KsqYF1WPMkEr9KzhBQ/JV/B2eyS51sbpA
94wqlJfCO/JXoyuKptEVQFhkQJFa+9/afZRXVv/Z4xedAgxbBlAP2T8MJokp4YlpfJNqtZzBZhoe
MbijlLTtR5wobmrbO3sIB/qRAQtegU+MghMC1DFcp9p1HHJu2HpCSfL/bORRldYsQCN5/rBLbG9i
5IxJHiLkBxMEdrjJfJHeoz8GurI+VR393Uv1sQJ7j8O4yBM5iLDgIh55MeeCBhn8K6DMtDneBDv/
yP8B5mnbW6rvRwWJLzo1TTGSg+ekGlPsFfiTtTcO6hWZ0Jhg4ctnWFwRLlkaA7DeFs036gLDVPET
07M0DNYzsw1L1BMHuXBYYlLahabXqf7L9qZFHE1y9oMw64rH0b2SigzJhMu0uHzkDL750ZufekFT
lwaGN7qSmyP7Lw0C2v2WC3xhjcOWzIyt7Z6+Xib4JpFKambRjSYC2qtXmA03Xk4SnnVSRpOtIg7p
l/UHwYQrXpQqYt6qzPG9AtvbaZRd1tOKIBtFuLnOeLa6gumE6637lhHEhBypozogdB9s28ACx/eF
z5dwbJRyK2FkvsYNHN9Ys1DG19UYR0LuX6zjoqz13h8sns343CuCA8oA4QyvRqrsU43h7QD1Kq9S
qkAFN5yvtzoeg+M6vwy2+Q52m2NoLl8VJ3Z93q/TGGrf23H0eZW/qEzHH+9+WMZFG/HGBbGNFm36
6/PvYlPn/QwtBobtQf0xYUoUw0BJW4Qy84ZF8bXlE9UP30FI6TWHOB2pST216XRg4gZSA2zIu85c
aPz4H2n9lvkaSRQzHP0p+IKbc2XaHlqZKbwMLZWSEUgql9JU1s7xJci3J6A999x5nyeOvXoiwxZw
zr+MiCFU4QroQoQIaBy09HGvoT18X7YTyViRz4KXF6zkpoCaptro/aSyuqn+eMHSw9yiasR4Ajiy
MYer4+8CDGWgyxJa33DbmTOT3Aos8c1s1sd98g4vbyGRlHJwSgFwR/M7bSVyd89L7mRoDlRDDMR2
/Zf8LNrSURgiCueYj9d3zrpBnES7XICJYFxQS/TKPAB19YR6BaJYh0AGcXTpd+Sme/MZK/ls5Yik
JdzmyyCQZOCnHCMDMStwws7v0X3Rt3h6pYsJjxRw0pm5+8jOlmYQ4PNyDqbndpX3EQXfh/GlmyQP
SDQktRj+f5+DqrC89Qmh/feCcUANHTPN/FN7urPHQAgzT8dd2/+pOpv6h4D2IDxe4GBct0NueiF1
zt80RfBpHsOG+Mz+kLJebKMgr2mkWTxRkDnTafLtEIicb6cTHgGOTkGW6ulD6hkslamhzxJ7s5rV
EcnpdeH9FuDN86oShVtYK7vnX8CQSbj6pCCKAiAKo1qTGAeEYudenwClNuIVm1vDekddF2Ytmm4f
OhDGJE8f3Hmj4NuBqPGxDOwpZXToHp5QJBafiNfNpGXdMZIn2pGyQGrhieIk8PfzuCB+LlhXq8Mk
PNtlOVBhELd+BTHOvaZcgScNfObH9apaem0o0VaxAU8tjGCjgWoVk3i37BE8yeiCtrUQBNQOPDgF
ydApltHCYAmD6PftRmIo0Fh+p8s9E88QyI47XLpyJIgN0etG/gNAjbddZNlpWOHv7Ee4b/kTyQHt
q/pA2iK7YmAqTokdxGqIBpuwu1mkFjWoI9lTH0PfkJfunestNtcqrfBb1mhYnVtdUHUEsRV0/5AC
GkAvasxa8IU4uLeVkWR/qtmGIxlMvo476Vlcd8lXbE4bTKN160d8ACsd5ipoZvWXmo1SF+8Zj2sW
7az96Jr9A2+ArPHjsE4bLQag9XYfeFAi2Xe4O//F0OModV+W1b/+8KLDRi+Sn92lXlyYRrrkdYjt
QkL2RO3tUzHRtoKkY9YM94JlfRJndz2qAWrH6NN+ReA6LtaOAxwFuwNaUfZ7D4fcLSiXvtv5gDBV
6P1H+rI8EMEf/s+OLK3AKUmiD5Jo3Qv14mQS/1Pc+gFGAjP/knzJvV70MWAKNPVIjI+IHwqqcmFW
93CxPqSLuU8XS/tPpNXoRlmuuMc3tC7ojFxSAAV4tpwyAndQRbBPCpfDMtZwF+qsUSJmYLqY8me2
mx89MzsRWtN2gQnBda4rdiSLi2a1IR+mQk1080EllcUxXnboeSvU1acHlJclR6cRwJVFrPqU+YAU
8TXnxWlGCymcdB82dMin51jJY0IF2kbuMe9ZgpdUFcnBAQnx/DLrMudBfCRyrdMOGpStaNo955wP
6h7WtOyfvJujdelYVlDTa7ooKzfNitm+Y1UXTrQIR5PSoqJHFPxuptCpPryLWAlBVTUdkFKE83N9
vj5xRHC6BqcQMXpH8i8KSNQW6N7zlZuKb56oZpIuIHUnIIbLR67+gtCVJYOW+WLM7I+3U+BhstF7
BK9JPfRB4ZkHLJk+0oD6V7H70X/fmwDsMOJiRS418Lw0aNJpn9FNXMXQffUGmzaBOejC1TxpBGRw
BtRUEQSZR5vbJtyVeFN9fpsuWyh0xOXwVBR5sz748hNSi4/5hpa9pC9m0e8WG/KC+sGpnRUYF7ip
pZu0RBQ0AzAEq/g/TD8PkaxovKI5YMnegBblxroURRdUk3i2vxruG6TAPr24qzrCbdkIep9ieZZ6
InV/iMsZqGu0LB+DHhg6R46VRBYK6iLixDs9XmXWTkV29QR6WRTQoufMk7AxQceZsbofZE6xwYUL
PGhs8r78JLR9zw4f5u0tfxGpC6OiJ8/QJYumSD67QVwsEwJx6nvk3F7GEEI/YXh4bRqNmkVlnUjI
AwndPMxBSelS3j6eKe7mDyMNsa5tz5uAmXWIpcbxCsljiKuhQUPncjsrPA7uD9rimzmggJOM5CXb
5eeKltMi21pRcds1mmDEq5kZG06B8GSNrU2Svil7v659WFiqH5YsRU1QN6pVKAyrLJCI+SYCdx7y
HfxrDCgnL7SjMoXHsIcXJ8rKD9YiP1w3wKdZafGzS+7aS2N4UZIwPmW3L9upPyPSHIS1LOXGw48T
5WgrXbTyOoQHnzPJrkZKRVCBkzFTULEEsQPu0clxaMppHu6FcKxPOVN61kw4INUTJs9y2N0R4f9B
KmIzIc0zC5ZYxkb7HSRKASNpOVdwd1TI73zo9mM1lcUJ+CuQR9zRJgh7L5p0fWdXWb+e6kWc8r3s
vwzuW9eLZZ/evgjO8UAgVqVulV67ESBzJ4LJexdutulmMAmdHP/E9ymcDNV8PcLqsScu3uFi0u2A
24r46LXE5AJHZ2wCAbqiakUnQHl3XV2Wv/Pqx9vZbZyrBpcHfWaUeEg7D6VHnjKX8UkLR5B6zjdU
E4PV6y+8T0eKjkJCtWadGmxGVAfgxX2s7TJ1wY4d0dTmCMMpEzlp6KlXeeyu5kTBVVsOG343vpxa
r/OolzpSto8gxA4I+tnbAw9Ojj2NH6VQpIKxygaIhN+50nHri6SUYPfiU+H8Pgl+qhs8M92pwdsk
EsJ39PNb0vOZC6tLWwfxfyza48snyW5+8+X+MplEof3JrcYcVt/kNlMkMgN0l8gpY2aRUMfs0jtM
U0e6UjV29iWX8s38In4BGA4SdDwK1D8RyWqfgd5i292IGPOL5Q956fRxlqkvU5abYayY7vhASgEj
NQx6LvJvsjTzgxWUCkdVHAuUTJSK3vw34AWhR0EwgHkH0tV9eP2ZNSEfnh4OzaEL3f/lT2qbv36P
Zlk03babKMi6MeHoIuPz175lV0Ml0Z8qe3pJvN5FNA+5WVBgDeitsKVM48t5yDP6CHcGQN9CQyD2
OIottbu5Cdd4tdv7E6HUh6nGDiJcSbW6rbHTLaGvsOmxTzd6GgOwlz2XJh8k07g2OcKVkTVY/8WP
qU/1ellHhMa6od6qMp+5gjz4Ov+D2QLY9RHnG1Z89PMdwu8fsmvwOxya2btSNIqsvtKJ1Wg4NPQ+
PbaC9/BFMtGu980y9nSPWJ4B3iyoPUgGfQ/W6QeSMjK9GBp5HCA/3Es0lMMqVsu8g81WZQztAE0C
8bFh06YTx60CaOf/1WLPfDV7gQ9Xg6HGYd+rgF805bL3nWZLuoJjyQLvDEmn3PYnw3NwxCejoevd
zqa8VN9Jmpsnsh0N17RqDIpKW3E/i7Y1T0aiACtxq51NK6ypS7e2DMSwfZHAMAbrh6oR9dH8LpG8
t6M6hgM8rt5we0NeUUEnjAFcMfE7LURDBbRwGBDqQKk1z6moz3Gxtugw/6Mjif8Iv4h6/XOV4rqQ
XhaPI9pC5lteEw4Hrll4xBCaAA29065j/te5eZFOy9P6oW18qlfFdgwehlDbU9Zk9V3V1reVhkUC
xEJRijtBCR/awHs7gOUOHLZLkqunA1vPd6DuvZBCra9myVef36cU1CzUJMUjcTAW04pRz5ZaUT8N
v2MF7rxLL/wDzLoHaA4t5hveU+OFuM7idHAH2gcBLCkxv95/EUPiro4nmpZ8S2PtdM2NbgHXZdab
1gW7DQIvwz+PpbvrV2Id0jfy68JeRNLKQwUcsEUag+ueEULNMvSOatB7sikQ0xq+N59gCsTGnyLF
AWJ4kWy3kRzSxgUdV3Bu+uBTyVDofkILTZT1wGlvaVRvm0wWfj9VZ7klKv8AHZgOof9nuw/iV4q0
n7+CqRnYl4On+z0eMC5j/qSqf8v32yEyfX0WmaQttjPSQGCsLGTggzMzqvUvrHPyIIPsubeJnNHK
gppjn3YOqLARHXRWW9MN/KO6PFaArA6DQ99RY3Yi0ZnI2Ygqd76yPfxDYlusgqS//bb644NBafAn
OgAdrWLY+C8pJspUpNLXbrMsO+MLuLu4nDwtEvo1hjSO7Ol0+CKqV/7H9ukRZVN/omFJ6en57Cu/
JgaOPxK6UdTea5Fk3CibQdmMksVlhvIYRgiFFgvpKrURG7UbXZ8lL859Kp2u8JUMKbGRz+vb9ihq
rsj1z4ycZT5AGHews8j3d0faRuHtGTyy/Pu4WSHWByzqnfFHjg65WUDWDyLfNuUpa0XMZHbjaiVQ
JGSO+4zn4XyWBB+16T//napznkiPkfRHEKT41scDexqoYctgqVHRGBaYpQIWdi9RNIRzg7pMfeIt
UVt/mGUEvCOjLE7Mb3ayyKuN5O+cprROH5cZaQDlNnDtOayKfQp0YA0qLLdATQl8QdZAplsXjHwM
+JIFYlrthHy3C22aKmtF5MNO2d7QkGh9XS7fDKQE4HOplPN1aYnMUDDWnCgdewb6r+csDdVPNtc3
Tb8cQXLB2Jq+UrwWbnWE85HdHgEGBkTYPO7oWrVJ3MJPrD0Kldg58VfMJO/s4GScAKqLg1X2rk2q
MKeWgyF8fsJPEHGSy/rN0B77M6UKPKK+wSpSm1kKYc8xsX+5couPcVoHjtUraRjFfXcge5b17vzo
qekaACots6JvpzBBFfMfMOTStmkkLD+VECGf1wFf5NveieUMu5LDyRh9y2TAwgyMGsje8PQN3xwM
ThV9uBe3cpfUxeDR3Lag3QFtEsCuKzwchmCtcpPvGSr78FeKf3xNmuRRqBuCrQBAaAnx8zI7hmod
eWR3kmjMXtCKJOhLg1NtZgie4Lm/BBbe9aPQgVjE22TAmLP/CGeuLTm4Hkjz38ZbvUt/BrIClxLq
+M0qYMCc7qmqHiZwe/jcSUKUnG/7Rmya9U7EPiRSRGaQmllJnRdr5D4hKUqdqlq8a0APpfeQn06n
oXbz3MBTKaGmWaBRVDZYPGCjDhmH2PuNejlnecmut0zl/M+zKwBJC7IEDg1tTw8Zi3CdvxMTohXk
mif/0FgdYDKGS96BcxmeFLP/2B2IWOCGR7QtEFnWowrai3TC3/26YCjdbhIKcPQ84jynf5Adm8hs
xs7rFUUK0cME4pbWNH56o4RktDkstlUY4J4RvD40Vl4cOzGR9CU3cwxfxI0UyiVgUG+O/qm/KQJP
5Mr5NwD6LpvAndP11EBL8fVBwxCOYFmlfSLjHMLajsr0nhMUCibiht7xoLvsrvQvELkOpkxubKcE
QDRpgdD4tN6CxNQFPKU78r3IHs7f2IYYT0BuBC9jq3W81ohXcI9RqA+hV+ydMVF793GkodR1vEfn
iqONCl+Go3YKcpzOb6losgyoKFs/MuGI1lPLTIHjBiFnLzWW4k5qYEqmc0eYI+vAGZlNVme1EBKM
ggPdidISvmPvxJ/8fzTsuC/qH1jiPn3KsoDzr82yn5r5cshhEKAmOorB1xzXKpBKugp1+yo5y9p2
5nj+DeB1Rh95micvwZJwRw8Q/AqEvxcnqIaqnHgoZiT4/Y8hu1KYi9fXbjUdLpG1LumEsvBcv2ct
1mtvsiYBqvZiU7EuW09JmmURC8SQjJ9uWw4pm1MVTOUnzmh+35+T1cSBBnCROI++p+j3CsRTyJOM
+QBwWCG62bw0yqWndKUSt3wyXldAbo9MWNZ0MZbPYx0DOVZvgn4ZY+4S65Dw2tTSmZX/BgTPZ9eB
7w9UvOaMuohDVvUVqT50M1pLm30N0Vum3JUEXPaDnq+e9ORF0/zvslGE11afBtcLhI83EtDlNYvw
bVc2TkQ7a4dGw1oDigrfO1NXRIDrTxNcPbgH9CoPWkcNItp64rlVEXobecIpTt6aMyJE3xhOJ732
FEwQdeza3Zur81IbtnpmHE9Svmzb39Yk5tx7fFPdZN6gvgb4SWue3C+W2R71AUoa/N8PEHaIy6Aw
0NPC5JGlhgJbpqDERrgZeqDUW4aLBRRVrybQzAXPwtyG+ZF+5HE4GGOQkOAO9NHSc4jxyWyQC0OD
FYDITGS5lm+hBNsB9YhKCe8FxRG17Ta+7yyMULloQIyu4j1ik1peQR68rpC2hsSI2aBMh5Wz2d70
CEj9GfhT9Lj+GEOJ+BfIuZFwN9cH2v7wioLW4oaaUUefcBtjJPSE6+n0TySDDbWDaLCBXqZDKfAC
LExKZCfTDWnKjQIM+ulJGvwTJkHFLaZ8tnf78T392V18fv8rfX4oz6hd76+F9ai8w4fQ43WCWMn6
o5Qg32Jdw1bc05RL9thdjJDSr8CCV4Vj/PR/vsX76EXZ7REvWjIPGm4iVrW+dTZL3QYXleCtaiMW
V0BiA7EtbREF4MFHmzqomdM89QNBcJ524BGX642SdTtFgJgsRUE4fRpOGMnUH/vUsE1lOh45d4jH
DG9/GZx6XpyxQgWdJn8XpVi5EO5v0ebHYSZqsCHy/cuu2xKi+MssmR3rGWh+klUim/GdtJtcDrjE
VlU0m/BCTN+2pX/bRkhqiRODhzNZVXtob5haKJ7azQGsr+arllgzpJFLx3Mw3FM++yrs5fL9DP4b
tHGRRzPm6+bLt7NxBo+xdf8b4vTwOUZEcvF7EAWG/mCiqQJMsIUxm0aH0BsODv+rHLULT9MKD5Yw
4QvkKhybhIYZCWV2d6gqy1lMV42pMXj0lc5+/6wycYDwwiQ68nJNYoB2sR+tJzvnF86HT9NukTcK
i0gWTp9qaKtolaHd9/SqJ2ek5vY92IP+fpf8TPj20nNl7WhEMxo8F6RJ50A71PjcgRuihrMAAT6E
MbjDlUOXhKveM6e4/xsrh//gqDMuYozjw2NC8TMDrpMSzm+LzXTITOcxUZiFYOYsDrKhVzA/QR+k
SCPMZh8aHOvWlxjx6R9A1c1xnJrc0mrqAOjOceHsq31xHobe2d/4S7UMjDCk/kRUm9gYWHtvqz+w
9qN5Tvx8Ca32mP4Hf1yWVQ5+XOC6KTIdAsCG+zm1tUkw0HDaCz8DDWebui32Js09F95bikHUlFEt
pM5E2Ezj6NBwwNpk1LjRhRfqFIjoJYYEkreotdXAO0ar5VWoRWV3I1oXwqNxulWecwb7Qh6ySNEW
Rs/v9MCDXfyEoT+qJSJUzLBDWB0IfcTFI90V2oZ5d3+EXaAVFf3Xoe3M1flw2QJyZKOWbt4LAp8I
zdwc80qT6SCda8kEG6NLa0l63okG9Ubfa7md8ORzogeM4lCQDDagY3liwuyPa2JmmzJsbIY87Z9O
+YgGcZDcIaS5+9vureqhU4QtXIfcBgRqwCOUcz5lId9s7Wohsh725sJLA9pkV/6yGnuA72JlQHa2
TPTQr3rQvROPhOsdfEHBt4bKtf5N7zGrBi7sIcf15ekKhXHGMNK7yqG1npLuoUUFnPWbjl+hCM7Y
aLVLYTnArx4yGwBh3f4KoBewGZWbcD7Wob/ax+kxoUd+3YoBvDYs7qv0dzP3Gr1vxnWSTeQv7jP7
hf4ZuT/ogbCQca/PAIgwOr9lV3KwfbADQ2fVBZgVTedOBBwrECr6YvrGDvEiPSG2YeBg2G2XgYXh
Bm0KSxZuYa3Hu3BebZae851gIXF5IPnnIxAW1iiiL9/QXR0erj1M24pizgKL1OFD2U7TXwKcv5/t
srOBkHA6iem6h7RjDtJfGH2Pn6pi8a3jg2gqwRTxUeHM5mRXfb83yUinsxZrkWQSCq+wTG/1q6W3
jqM8RCLYWo2xyZhO4DKI1MSRr6GNwpG+lDSoet3n9QpNEHAyrTPQs0NbHwVi0SngvyCvRjlvkGyI
B/CE6WWHZsq0NxDn8Vd+H31Gg8Gd/f7kY6IL+G3wW1K3s6OJj8Wt5AaLUIayJdZ738eWsxpyjH1X
Wqa7rXtP3mB3qS+QBE8QSM0ZAP8qaJs1nHycNQMScUBC9OdiXrAWhqMq1ztpOFiTL48Hstp4jCWY
TLdkq261wSGjbRExwNaxY2L5gJ3V73SyRyQcpqjuR3OpVbU7NsvuXE7/VXaK5WAEfqMf2+R6zyNF
U4ipupgmwwyEcL5nSnCVBMVxdtGAC3ter9Xc6TeL9lU9VUBLBiaQojE+glOSGpDKHwi68v6C6rBq
6MQcXHVQkYBUjZBiRfzy+DgmrrcBktB8XUqX6AWwfKHBNFVuFYWK7NJjHE4b/woK2oyJCUx/40/K
IqvbLL4+zu8s5g++vCni6KTHcvPhTmubFjtlzhFiG6NCRwXtgbjU77fq5eMcvLuG2lt9/fQn5vWQ
3SfuLzPwTdHVdCUHT7urIyh+HMkfADIytPcq0yI20ZRwpj0H5opFf+3+aXR/LaHn/FFxVMh9ngCc
drnU+KXlElF7cN5fPbcvcCmKfVZt1X0dclfZMDeX3QxJ4dmO/5uvwpQez2q1UAJ0gbKjJg+4k6F9
4AQcH4facRgwHs3v+2eF9DQ7aTWgxAsbD2ZJfd71FdIm9mYEZ5zv/97Qtk2Q8xCOb9hPWS5hkb76
eFbraDwNDOUiUysSlNRldbB4ZbcoNSWX1gtamovEFFP74tSca+hNyTURxi9mt+S/68nc2FjWfFAO
5OXNTytbQlFSiG2PjlHBCXQc5GuVsE0Ek3iA8xFy6khaKKEqt1xlofgehhOMzFWnbGukqPC0S5DS
oK0yOTkeFT3xI0hxieTg3o/krVcF/kmJBlmKuNByKEB0w+qTCg5C7swHkRAsC+o9btUlmcpZg/XK
5X3nmu+wmBt+Jdxw5M+EoZC5Sg5/h3FOD1GwlWj4MYOx0bMem3LgmH1cGSglvqhHIRYoawDWUqGU
5zxzCORnQJHYfo5SOAOTLe8y3q2xF9waJij6gRAHEVzP6MhKO5eV+KpXtIl55fouIm9PlhvXYyVU
3Rva3lajqpmtYQndPCq53iooobtZ6Ui7kCt38F4lae3Qz04gS35Hhi6er84Oqi9/apdly5gvtuna
kyukRlILCQ2nCjt5dczqj+BKjMUkXAD5V0JrmdpAaoCsVAVYvinFNXRDiEoTRW6LloNxUSJgq4lS
ndyEIfdSlKl0OgLN5kZqzfmd7J5Y71lyJF5LA1j/nmrK18sX9/vNpu1QOaE6qy1DUTIJJHZ5LgQ3
3+L2yVmmmAaUspPZ6dBLVPfJOs/QsdWEt6hxX1deb3UQ5kvrQWT/Sahz9uruhDi6j3/AfYS2qN93
GfREpEkJXhaTUe8/7N3A9xf7F4rNyjM6UdU4AFpJrWvVEWTcSzYme3EwREDPsxctbb5u3iAkdnTt
X1NWvq5x67Nx+4YTAKinBdFj05DofcPFW01OuwuVRB7HYYa2NFxfa8W7DJC6GayfFlrYy4/Wfw8Z
zKU6yBhDdxQ99q+TZWtfp/bsa889GfuZ0VOVC/BLzBp7IuODyzH643CGaI/iQc3vs9uql+gh+w1r
xH05uB3LEfcRJEpp3+T5OpmWbfvc9rM04yVon6jFNLeosejuwovJmKqzOSnhsG9F1bFqyFEnSBKM
4KlOI2jvLxgYycYkLtnD5475hDp6tDRA4TX7faJ1lNFHg5lLUInOsDoIachXTuGU+yp3s+KIEjsz
dIHVTm6Ln5zvuVU/L4OwAeHTdN8vLaAPSoaLtGkHyD/1DY3rDw3vMSZrR/khZiyNlQXm+g8HB827
SvaEtsF929eGmvgWw9WPvKCO5Y68EeGrLfBTojoKQ/EmCIR9Fv/aHjjWkZpYjotWjKrjThxTtakY
AzVB0UpoDl6d251/gIbUU2MHQgItnucbaepODLTd7PA0Fw3EViL+rHNZ0TaOXUbgGOGY0Was3HTN
Wlv3GRr5NhFlOIdmwU9go6yfLxGlXE/HXfIhwnJdbtwwvK771tWl94OQz8r9V1lXfl/NjHEjxbEk
lPA6fmhqu9XHn3CzUDxHSCw166Fr/LWtlLqNuGcEHFrVSyy4M+FAshqBh4rlodcCEpnUg8PvH3Be
BOQGDUHxO24fe4hiOf+hW8R9+0IN1D7p4vD9Hq+vIx6gL05gTnDHDU7afuMWAUrpg+H5Gu4awKpD
2jNPni735qoNDAwOQCUJ/Mvg3P3T8NcIH+/1Am1vzdpu/NsWG+KHe+XS6zoRyb/R+P8YZvPyh/kf
0wvFMjFbaMsCM6hufLsJwcGZUdQtpRURBN+JsC29XR/BiWeYuu0PszQD93g1STxKKiHNHpF7EHdf
fhOTYeiKZwdoPM2r9nWs+bq3y4Z/6BIGpxcNPNyaNataaQDK33tNqNVx9QeXvGJOVrqMyMjh+XNN
oGc405nKR9W+UNh7+df9ouV87a0qfG3ecWh7G16I+1DflvGHvGws9hcHXUJYOVcKZW8AiB6Kl3L5
8COOrlVXflCWak4Mn2g6kbyElbDxZ7/Bb0AJBUvTv09B41GHg3DPZhdUAdKnXvl3dWMgrl/0j/yS
tQmXdToJturxS5uO+KsgIJph+ApNOrru+eJX4EcwbFXd5DASRrDp0K3GokL1SG9uy7Ej7nxkn7HY
XYnF0o68qix1niV7VxhzJNFXItMSddB3VctlTnjw+rpU9+iy2Jd6rasuNrm/UpRvARnuuh3N9qbU
CgaRh+46XuORCOHGWJmPaTrdP+QBAm50m/Ve4GXlHHWlbpAVmaRh7UGpdahryLeMoyMJTwyt4s3J
iEmxbIOjPhXUPgV5DTxEc4XdrEyG+qmlEXKB2g4mnn3zj1PzO5n7AoA410m45U46OkaS5KGpLFv/
/AJ66KWM9p5nM6tLCAGGsqFI4GIl9CfUEWK48u9nz8md4n4+0fIPjcTaH8wci0vEZKs00F4CxMnk
gG0oDEt6aMQEnFQxZuPTZlHipnBqKpncKG8T9oOgvXGNx7i/8sPzoJAh++uSiMwhHaUfeCWOi8qo
128vHLe2hHMabdIj6uWmu3CbN+qUFUZpABxiUzyeIplwgqK4cLeOM9SOjTzy7xejoaHehD5DPvpK
sbotftvp4TQufOiJdIG8XmuE0NLvNe0PysYsH+S0CT6g3Jaqs68+VQePXprAGThxpqoU17NpbhFV
ORvsZUoDuezaGZabSt4EWyr3c/v04fHkQvyFYN+HGXN14VHDmMbn3MGTQGWpkxHaR58kNEpoUcnf
O7303uStvyiol+5qDDEtJzd5COSSnm1CELWD8DtRyBHh2dlmkPHxPPvo76V2bhXLxX1J7cPGP+h+
ZRHDkUJ+9dqSCAb0WsN8h4UnFflEG5b8QEc5uNveZHSTLw6o9SJ334oIO2oBjplpnyKZCnUg2yeC
4WUeAaFu6IREUeI/5q5ue6Ki3ePkJ46nfmzcjKlmElx4GJHQsMsclqNAgXE+uXPRUj+Fw2LTowm2
G+z63Oo0OKXPw6BGp6jnnt0lT+x3Rxw7eBtk7oVzMxlRepGoJRl+iKqrjNg+Ty97F5mPeWnkIOVf
26QUoJoLhqMeHZJWCkasUucHHAHBmi31GDufN7PsOLuoSOyuZuYCoAKnIgwhoxDcM0eJZwGgsNd7
lNAYAwa+Ia+prrOG49QMTR846cxHKY7Bz4us4+/x88u3IjQjWS1oobLkwL8NN4iuFV4dWhsHF7zP
/od/Z85vzxFS/j2fnkFrGaTh7ALKkVh2sQzjlT13fJWlBzebZG5YtkkjAlOMOxJqXJOfWnz0Jc6E
PMSA241wT37/e9DcV3IwhJtIPF4sl92KoECYNpzMjgV2pa634ajbt7QhT7z7RNPZrbcSZdqvT5V2
2iCqjPO9hmoQIAholHASjyAYUObVr5tLXu2rMqGLmNvbqcj53UfKCQVzdAwEmkI8XRq2L7rDmHci
QRGdB9GX5TY2gXSU/jwyPwUytBmrwqZ4nzXHHuvlCnesK+VoStw5vtEex0SowvkSeWfDNw2qvO1x
4SUvZ4rm/2crEFbgFAbgE6/gSvQYt4i615e2Op8B8CGHyDSNtglNxvMNv88wr/+ssN6IjgxokUyR
hGNvaqvad5hMjiwwzRLOUexHEschM6zYKcT43P81FXCIYaKR286VPZDCFfq4FGP++k0VRrAG0FcR
PZCOs+fBCvY+nte4pXtwSemyidApf8MEgUru4Rg6yawNnw5q25XGo6/aAKhxzQErTPwFwD2biwpB
iitFBen1qZuxjlI0v+uCokN0eg6diulOj+8f381bx6PTMyY9SQQ8zbsUYEz8WRaDc43Gu0E1YCLX
Vcl5HhXsGEigfZVRehb4IPHamkpJ1AF0+Zi2flCtq0LF1N0wF5KRr0stvFzm1bNEy0LSIpFpkxfx
kby/H1kFxnu54Rzq2uSFo0w4at9mMdMTzIYldUjGxeSmHZO40Mh3WbxrbAViyVBelz0yyk0nF4N0
fv8shAFaOSD6bKOTePRg53lLUndGCeI+imY4Smoh/+w9c4ognK75/SRFrHFP0ZsBcLMzO2HyHCtr
mcijC7EEGSdtbNypQmk/e60wfxJKFGCCJrh9YG88vE0HBA7x7l1Rjd8USeLm+IfqQCFbn5MO8zau
yBqq/lRE+ECso2Q9G+iJBYXKT66y8es8Y1hRFrj7PAlEvN/oBxUF+h02V19LbKvAEYPXzAptl3v2
fcnMIeS3bzXWXKsYY1VOpvQOmOWlW671+x0lT+VECs7rDOnsrhnwomPfc7Hs6C6ysWClMz3AC/EW
wlXyEUHsLYzQyGNwnFfWfVIxgR/2gS+CgpiJz7/49YmJ9TIhewmbGjw+X6A7zm0VwZPSHoqs/VrW
ZtdMQMsxd4sNqJ3zjFIuKT5rYaSghbVp72ksKmL+bhAdNHYQkebemkmKZtWItJ0RC8ZVNBGZWwzj
+7uLMImW0N9kAUVf0O1oLJY6zyLZkL87O8RlzmUJIgDUeyv+3C0UTfK1DYDo+exNzszGFOWVWQDj
t9KfBYmo3R2JHX9RT1X+kkpsAv3sfKdiDgJA/WqjpNCrb3S67HFqrwpJxWjymaNigHZmdCvwwPT8
DIOBsiOrB7jS6hGHOYeHU7rW9tlTFTrFvLHMgog+iNx1jbbZF3R7m6H5lNlBLdZ1F9PKJsmO+G5J
YdybJieOnBQr+ohg1AQPlbDBqHOocZCX2xymu8XIOsF17n92CVMlX0FpahhKirE6Fpk6UihC6N4H
DunOLMRNWBDANfTJhO3bb506wQ2aNhqLkM6o5lXfFVkBJb6ayQ2yhqr7oxL5uR49R5IJ1e7Gln3v
Dd/XyCoeWN7sudhzDqz4uzRzgg3ARYxYt0O3VQVbUC0HL7V0MmU2RlNUS8ZqYF7ZD/oAkZyczw7N
eIzIGexAwGE1xZf4jVyOQc1+mx3/3eA/IdQE1ql4jO3EwLgwuAnBL5Ohj1EAbyH8EpgELGQKb4N4
I6OvSC/qg+ksjzJGMilh8Q+rxzve/r7asVmNdQbnNjMHprDJGve124dMlie4tA8yBTo2WodFsQyT
cU/rq+j92KhpA/lUhiyOR3JiR6bWzaQOqiWIAyE7jPe9crmDOd6qdj8j2POjG3AhN7HwQk97try2
dq33wrC+Zjfj1cmF/7WwoIrZVOnkcAcCHRsuAwsW9sBuhxWOFbeRUWLnv1G3Z81Ie2mmP8DUsHXj
6sm++X5cIjXdgwgIFsoeJYA7/PM3AkInCxCyplornlVYu9woGfMeOqPn3eawq4eVi6YYUqvatp+C
99HvpRY2r3LeLQ8sQDieQINAd2qPLprLIsNOrmM8LcgC4H7rlajoUQ4SdyoOOdb0GFt2ZVhZCCL6
zX7G2GIs/8tPvP4E8T+qiFPdnpRnDMeuwgG4D0nU6A2KtEM5sqicUaUEzS+56Q1drooC2Qak0nTw
fraUAPpOktCsG5lUDkANPfPJcHmCwl+PhNVLHI0TQx79hr2okyGVpLMH8ql+y309FFmzq8rq2Op/
tW7Z7QOwPeJtqK4QO8QbhTocczKVMwdTFSb4I6FpS52vmHfWjdWlzuHtMo/4UjTA/a0CxBHL8ytM
T6NCm5YFu7TtcaDTaBkWcWmM9g8l108iPZNdJfu8RGKAFet4skphqikYtTFJeqr+S2KQXtMauHmT
ma/I4NZlhnFRp2ViiAKGldFHY1gmkGrdnfV7jUm7xMFL8DWauUCkuDN/KyDK4CK4hxj4GYiPX/B/
OQssY4h+J2SpuqfLpGzGnBOC+aERRPSC3p1w1UNzZggtTcwt5rAzehJ0fF2fWWViTUFnHFQ7QBBt
OFEYg1Y/v59PETo8XIWMn4a2INkFaYX3xzOeoc6+IPXyE9TssMgZfLtBU8HV5p5Dp88obRyp1ZA6
cpaxB48NsXw2il8APsLgg2FjV7KzlsvOsrOJFKVa77m6sFTFjzO3eOdwu6ejw4iCuaAxlkARZXCf
yCKi5MESnHrjmPtD3wTu9Dy7rHhEDFecFuCaBbRGkFi3Us/COzsaT1dXgVSVmACwcX+VmxlTUV1Z
XBqruaEbPOIiT49wIi/l5Yf5hxQBk3bCrk93ro2I2gLqhyiVtUS8EweOHQDg0/4zCezYdTiqV3GI
yMtC92LGC+c7AfmHoQPBZ/AiIqBOzppWBrZ5mamHjjhpE1k3fsbCxck+++NISiq5dK1rQMWNJqzI
+6C31goP+IoJncMCTrzRx0WQRlAiGykTlypfTUoEw7ePknAFQBpimMiFWFGltGVTEKx0Q+ZhEyZm
UdxbbgqsssVrQBZaF2TnFl/ZPPjv0ogVjxZvKN/n8nwFWVeYiOcEs7yC766odMX5LAEaSAcA8bvW
xxYGit0nOkqjMEZ+qsDPik3Jm+cyXcUXJGt5IzhPGJ3GmhlVR0QNRs2wCU+MXHjZHqsxN1t9yUV1
7WUfeDZjiQkA/XxLeEANL1g0lE8SyLBo/sa/GmO43BRhBeXyJukjQT7n4oGUGH2IkXd++rl8JH7u
X0zeEPZM8c/SPw7fO7/axKMv3D5BVvMwU09Z7UtwIeHeZ6PCrawBp5WEWp/IDRm1Em2L75UHqoxV
LzoNVoQ34hgD5acMxgIxfZlligVIqJQIYSfKF6xjbY53pedSr1TWe60J+bO6FpzEWh8Uwlf5ZcVu
ZPqyNlFbmNmjoJevoS0PBuPqhAREEsoaoE7o9u75KrVYMsE6ZUP09X+rDY0liBNVYh0/fckl8imY
sL6YL4qAgtEG15PVsowcxu1QZidDB3xe2FS5kXt7tWFdpGFRZh8ZXqWrkWXSomiVDq36nftdxdCE
Tq/hUXH39Xe4JEjxmrHSDjYT8Yje8sc6nijg2OD4Iw8DpQKDv6Z+SwR2n1dePXhaxZfz8hOkaOjU
3DVTSzpRpTm2sQWW9Kks+SvF4Oal4SXNtUXIEc2V/cYz08WwjUF30dzZgDQSroxYG9Qx+vHW1xIT
6wEpsH0OORfkqrXSBYa7pTkUHOL4HlDkY9l4m5AXTBPxY4HbGzwzetZscbc7vVnsMrbYAdMA1K06
MwtFb7ZT3gXpy5TvVGXATYXQC3z/SYxbOWnD014kBfzopWmWel9zZJzbIhpM+3oIYY6Ex3I+a2zJ
QEBLeC6bKWv24nKSDzIdRw8KxLl3cEdf30DC0RBZrO/Ed01bLp/J8zB4/iTGfkrEJmp0kAC5KzsW
+DWBHem4T2kz4Ix1h8HKAP/5rolVKCzIUJOozc1Ny9NSl6sMZRnrKoKY5uwHnGs95XMJZqfxs+si
r8wYgqkUENoyS6ifxBl0f5mjNtTDa52jleabM8iBeN2kwTTQkEIxRV9QPptsSLmGOPIyIYRK7/SJ
RXLhG9N4HionlWbW3ll7iwRBPEd2XctXBJpYe95D+ThKwIfUqw80iKzNcsF+ECyACIRcldDH7Dys
Rkyrqz6gcmvjQPP49dlWa5A0EZdMb8UR4meKbn+002ldTkrcaYVbJfoAgvxYGyBcnqqknH+EUshS
X/0y4SfPiYD9QbULy2f83EVzu3tdKsmfXeQazRnyLyuWjNuFf3rvrPXzQ9FrFNy3PUs498b4JRkw
Yd0FNuJW7rnvdWJJbmheuJC6uaBJA9VukbsB0LaNVjn3v9ClKRVRH1e0ZBJzvoBAU3a+vxQbwVPL
fNnhKMhiJakLDyy1hY5CM7y0HdHE07Y8ezW2Re3LzUk2yymytRBA8HnkizpDq4em+fjRfiMV9zk6
LguSdm4uKwfVQjvX5Mm93FwlymiPs6HPbFcJiA46zz3ONop+F4gpjvngG1QfW3Uey+PZXIWy5C4V
gWmYGOdMMQ4Zm2ap/1dJRKrgp73Ud6I+SsU3vTCx4eQ1QBlLxMFyZbme8z2aw440aKNOkIzy8qaI
XdFfKPyBmEYcM8CNbQHVB/AkAbFTMO4BwVNVPRvHC2OVpZshWtoJjveKKjTIBiePxA7TVU4lqxgT
9sufl6bHYxJW+DW3yeXhl218XDVV2F4T1/HpvV8rS68nVmv+IzYpKdb2m2L4pNGhetY3x2sOR8ow
sC42l2OIwEFhiA1maaR2f70Jao+I8tFXXsEHzS57z1v55bOIWeeJLlCHeb2cnnfLnAceZPQjI9of
RYm8h0XdqdZlceLJA8VBogdYhBfJRNg2rJyfqFa5MNS//os4GM46cFFz/VNgrdkVO2HTkQVYX1Ev
kRWeJu+Z4WDBNiS2KaT72ZhVCmL9htoy0audgg24c2UZYnlBmu04/OHOVsYeOk9qx6ibYQy1Re4Q
vJx4A5sfbD8mbDQQ6jxbZNg0be64xtSLcdmpvnLUn9yRcc2Nnjur5H4KLCVynyVwtFFLKGoTYXNY
HWALosPrJRH6CyxDzIPRNhYDJ9qD639MwTHUDn2TjjQlXHb+katTJrpYbnQignJ1i+UOxtd/GtRH
Yq5tAAo0s6DDXsdNcj8xmbBG/LhK9CxAJ+FRqtG+JZjqskbPmGDIkBIPc2rLhirFfVQX/Vr7Jnl1
+YA1BQjoGkGOklmf+if6NhjpL8aJsYvaj1GqViFRO7F+wGCE5Lw0jrPp7NZwin29LnZvh3p/yKO3
WMAZrdVn+ys0u3Lql2ec3mtXgNR5E61zKM0bEwPnNyDS4kFwYnJo2V2n2RX1js3Y/pDQbfFUGLf3
PHosCxn7ZFYnW9zBlPQKKgKHyLgTqSCqTfIZESE5sMwEveYMIEb/4SKBJ7mKPoYiIRLdChMMXR6u
7eIqtZH0+G4Dvr3dqHgBuVGXTd8wsYwrNXnhcASPNcuTEm+A6i0rVK9Asx1ZMdYMZFAeW9m5ywCs
vfqAKwmnDZ1iMP1i3c8QUkq8J393SqHovdU3jfZwDXAMwRuaFJiTh9IizcNkxN4IQfba/vgm4LDw
4KNFissbaPN6gYujoeqD9dEl607ac68ZZVQmUkppo7ZGffPv2qOk9vurFjFz/Gct8iifJoq962i/
huEsqIcrxrzeH8YtvH/VMyUlGvLtNLGOOvo52BT0UY3GXVu0BgO36JMWHZAwtfqIEGb/cltU1raf
pGxxvK3MI1NXJQ2OIM0uZLZ0KL/bLxPH/wWnqgGd6vTPc5QUMaXofn+2hKGjgRfIuV+wzbd0qCZ8
BFI2uAMIr7KCi1Om1vCfcYmub2vk3Wu64tz2oYTW4aEeSFQbrIfWam5koMOMkC7UE+fQdOiM5FVT
H9iWBBGDFMRiWl5dxAAuPAcM7IKIwlrhUHtsD8FkvH2WUULTUb5s4kiqfqN0k2H0DTYoyfiaTU5E
v5MW6usj/Yi9ov6WFxuSJs7z2PmJxqGLgeDdlIrruPFAK8HxQgDmyaFOzIrdp37Z8KSoJqaWEt/d
yz+LPC2d+GAjQVdc7rY5KmjbUxFYkFKLOUnzL9RnTAHkLo2ZLZZF+36EKsUqdIBzKrgBxVLl7cxx
NJRkPn5IaS0ySWBRuX3D35rYhwnMb6osQ2HR4pqKl09KKcoh/yWqT5/z4JMgf9Rrwn3gtcPg953i
72WrkgfvtVcyOmYe+Ayy/SGRJoUVQe+U/bhj+U1dij57DcwBHTGK6T+5WsZf7G4EbWERQdPSIqMa
s5VUoGSa616YCYEu8tZHoLavYBTviyghCKUG3pigOmN+2oLz6VDtB+EFZDcLZlqG1TDQkkjtuAxw
5VaoX9vzK0w5c3yOKOZcfswTKa7Aql8gyiWmfgDA/7wBfLnk4O2C1A3l2Vpr0QnmfyEkd+f5TV8e
0MQBh95jwSP9y+5biINwG0n19qy1VOWqRKa6nzJr6gtsKKsyk6SKxjW5OJNLsICPsPL83TtpYQV4
Pm1lEpK3Odhb+BaFVCmEgVHquW8VJeVtF2a7gE9z7t3ThehkQ4G54/zVve4RHrjvlPbOnoXf4wpx
g3i45hCZeqP+jiNjdK1b5PHHRMPNjLzyu7Ua0MhhKDeWiuwQwDUk4YjkVJEwoG4Ee+PSzQvQrPqo
fgU/ClMJt9MZZyKZZRk9rjkXgq7ytNPu3Mr6EgifL3XDzfaH6lSUxsdlyZvvCnOvFQ7TBiE+orcG
aoHXBJ6Sx5OhksMQHxAOQaWqIvI8KFJjIOiozjVa1G1TR28ebfs9ej5vhpF7Wx/qK2MKwpRcyf14
iXi98MpboN/WXFUhP8e0OXkOd3Jc2DGCC5S/Yf7MA1Qh38sTi6gqp5MC3FgfenenoTCo52NGcXlY
58n/PrrhFwvAM9RKGcCTiJb5MxL4gsK1yH3/lQ5ZSrcxD55dPtKnHda+O31+G45NkF2uMppxl+bT
wiRtA5NIVYZpbURHVC2Sgb9fdIfWxO1L96KJ8WxtYPC+EbCKZeZioPZqHJv573106miX17xKHX0A
xHdFoZSZMIIezAZrGnad1QQiKpSkwog+VJWNz6K0tZa8uDUAhjSwVoUOnyUM2NHhFBSYnniEcv1E
PN42HVbkdanMV6pkupKsHbTYszFaSXYbQZBapx/efvBO7vBRDplhezWqGqOzUDGQB74lylDOzlzg
OifKs49XHhQGiVZUpg7dq5Ej9Lep+GoAuaMKfnCGvCQwUYSIvhhMqizOdPRu6alPgGj42DbKxTJS
u/hbrWVjPSeYh7kPAO35ZXirJoYKYt2g6UptdZ45lGmKm9ccPk2LIw6pilxLBcKVOkeHUXVqe3Tg
/SFHq2y/6EKYH3uIt6W3NnEhlrvmQ8p2oWFRZfrD7CyiDeME3kQvIwOe+BLlc3F4NWYmbVe1809R
6ZsZVnliqcKOBZXTkWmhLq61RQQ/2ZKViyjptPZFVVv3V+uOa9jwtYITmni2OxPUj4x9iWJ5XaHE
SVXFxkBQnfLv/Ys7HvgkBbSJYQ7jQuhZK7sb5EshFbHqlBq9L2RIziP2uehxiU+s9E1dqqTg66Vp
RWORjiOmUWuEVGoYsxklGBuhPCVU/8W3afypJbZdpUfM3rZHVcPB+GRLZ3Yg0H2PjV/zI9a2/QPY
QVYjv9p/teat+cg8R2U99sIEvhV7h980DhH5xoxltm1Obra1ZFaIc3H/EvL6xn2LUUVIuNjnFjTW
eLBSGb/XcKO2VVpWyZiN/Z1ZYaF/lTHvTVg1qXNh/Y4RmhfxQhdrOAvzf+NNP9XxsgiyTPXn8VDp
IaAE6pMo/ZQDLPf8VE1iKnBrxaLkNcITfbd0q/rw/3mSfiUx7zd07qocOu7nB1TreytMmXMAppoG
R0GE1rYTwFijXAsQcsiMV+Ta3J8xcANSGrIHl+32dtMzGcVv64Gm0RYW3VvQjSaobgpVGC+UPBcn
p+xEFRxyl3CxQO6Z0PkkvATvO4vZ+cdwphqlWCFAkrJ53R8VKW2LJjp2yg/iYKnFE2ZXiQLpq7Rx
p2+KfbcSDkCEF5Tto3GBqkxre3F1xXmnFSv6GA0rBjy0R5RrqKwka2cuBhm114Wn0go+3oBjdzfV
6RZKC0Dao9SShn9SHudheuFhUcf70zD6br3LRs6XKwOqF2DxOGASUaWhKq5e5cNjr2HOTRO2gb+a
xtRDyZ4AhczwOz9eorUda/ucK9CqlMeYWeYasIapTOaoOV2aHwAY7XkSLIudbaowVGYPuTpVk0wU
eDoyQidDUCRSpKvDDL3irXwpJcU10swJFxb3HHcM11VW9csLs1dm7sMOwtiVPH7EhfklVs5CD1AD
YMFAEODvCJkN3HpQpH0Afj9VTw21prhJeF5GYdDInMgU+CvdyxaKNEYQB4YTL5VCz4gm5vTQZ3La
ih8GjbKiIV0UA9c1hdlB43fcWJaEFQTl5+CgalxVxa99NKfRBMRKi7fvS7dPSl7tbpkkarMVKsRm
Y+zOSRVp/7sUuk6lRYcyCN0iGSGdUvGGRimPewkZzshWRBrNK/fdzWUiB8nS+1m8Ul4xQ6quTw9s
97IOgQ9rS5WEpyCLXk56yzhHRMaQXld3N1N/8xczuTxk2dhP60idzg3E/aAft99OgtYHo+poMJ2M
i6mutjdYWnR6kmi40mftG89dDR4g2V5dqJ/2h1nDI+jwGRYYz+rzsqEXsejxe+zaQawInbAip1tH
3MGyr7qfWTjzM352kuNAd7ncS3Va+VsINKIF1Coa/yZHDRguKE+3bdBWNlfzZvPaklGRr2nmm3H+
nMhPiVPn4mk8wusSiLq0PnAv1fLeNdxHzsJtWADC8Qjouday1juA2oXKzuDz4gKR8qh7XvXkpT+d
cS24mBn0yQNnJrrcfblSTXnLyao3yRr6mkTDqww6nioQGky+miwtElpqvocwxGzzC2oSujG3Tfav
w0ZrsXCtqEaeHEK0R9KlpbqWXJLflGHLfA/y1mtYf4InrHw2B2QS/0kEzKdMXLMEX9CMEvI71Awj
4l2I4uTgNds7CH182wPirWVjZ16vor1OkVx6IdQgr4AEhOBwlmsd+EUH4M+dXIu6Kw+4O8Fi7rNl
2Aj2+7sezeZ0n4BlJwaftBxTmy2bYviv2eb+NjNImmTVbX5fcqZKvOssfHy/jN2Yrn4j606GKOki
1RoZPERK3bY/3ap5ypfehLYo7SXQM3nzMw2LCR1DECq8LX0aspcRD+VZV98G/r906MielEWyVnw6
iMvq8rxqq62A8utjdx9vAJrpLMPDuGSFXPmAPBnoz5lVj0wYVrwU1b/pe6OR/6iZxrblfjBjBbgw
mJB/dcCklzTsY8d2+pbmgqr3J9AfuaPe0HaPjh+K/vPLrLk4Z/4ba3JFnHvlC2t0twi3vGKXXtZ6
GoM8ROZRVvhZavdwDnFtRZfRK8MRr37BCyEGRy5F3EdaAqXbkbvM33K+u2obSCrVV092OaVBVmax
qxBTTLlAUj2Uw/Fi7g5/tlpK64kkzf5i89zONDW1Lo5ZagE1pzj54n5o0g3EDPraUWhaMp2dokmx
ZbhDXlh56bDgb5Z5nsd78/4lk5OArcg6vFsE12kYiGDhERIU9bUd0heP5OvtSBF+OpWe7JQ6jk5e
QPBWTT/I8dS2J8ZySt6Y3lZxFWGpAa/oVFQGfC9TPvXPRFn42jGtZ1A5woVRyF/0wItcnY7Ye6Sq
jsuCupbOncX4oDv1JZBs9wFgOId6zdoNdBSMzbPBiXg7Ev+S3s/YHxUrIQGMUVo96bjEUW1rnpra
/TBmWHSmTLTakJ4YKTBSq1mwwBc0TMJ79ebbue59iFLHiOPJc7EhIT3seYpr5tcvDqVgnUoofEy6
YhIzc7eBquy/Gq97DebIA3bYYBoiOs+uQDqfUALZ8AMlKBoQJNT6j4Pmwy+/uV6rRFQTgYaWWZd5
PewhDDE7cxrrWZBvQyLdFE5yTEmvRrK/0VHlfSMnnAqwZiCtmpOq2hFAjDv9MaHuRLdPaEZF5KvP
hT/a+wpt0zihLRjvHPPUTdoyfA43HaTdF/YFEUdsNeTN9fRMiqj70kVTqwb3GLz6F2/5Aax7kczz
axAof+QXfQ1XVkjTEtT+LMWiwOQyTYBX6QBgiPnv8X6wpMUQhZGM1HSvelV7yJs/Gop0AIyD9DwG
1Ao+xoaxuY2oXHR/UrKqPAIsZseaxqD5cab+fuYy2xJ7SogkncMILjxGy/5xBpi6D6of5bVQ1f8v
9gIojaX/sVWAtIVJYzuMCHWpKKRG8eGpH/Dcak334cIIWtfPaVVxouXVPuD6oG1Bvze+5fPmx5Bm
QItrNKoJXMSGBm7FqkgW7Ljtk5Hn22P+W1BZhwkSPdgHE+8CV2tkxqHcgoTrdR2ow4uHjJOsLLO3
IGgI906DTnmKkjwEh0rcau+PzYUBVWS4h5up9QMFp2YbI8xpuHNMIg2B6VZKeReaq4BHtK8pvv5Q
4JCTlWk9G8+r5od3a0Tq1u6TH66BsYEE7uygAItUgINoI22RPfo0u550OsvBCbS6rQG4j8Fw3mvX
Ag/hILHB0fZgKTsnr0fqWgMNZ/Mk1XZ8Jsa6OhCAkCl5du9MxVglubzMKszKhj6aAYTasFO/zbcs
YOSvIORPUCLEx5A3/9Il7mflmJLb4nAirm8zcftrPjTNOhXqNeDb8BSLqzjZHg5+/5D4TMzWYL2w
baNOX2lyFI5SaJkF8ksEFxC2nnyWVxssABqgSAFrwAb80u83yj+6FV6CLeXCCXaOehfsJfh8P4qt
J/ZPNagzoAd+tY+ho+OcjG+Cqa+t8O5FQs+FjW8sOzentcjhuEeLJWeoMhSYDwdisUdNkef+KfyD
ssPNlMwt79YdD2HFax2tOhodu8g3+NbxYtBIqTf+U+sT61QNI3/MTONw5GSrJ3elzjxnsbUEwpNQ
FUwYCPzTakrGEMawLPhWnfVB9xBGWlyTpJLZmuMyx+u9tikmgzeTFyb+qtDDPcvuEtSSJIS1jTGl
zJmRAT8qJZ17sI20agfnRKkYViwtG7k2Ez434BAHCLaM+4MD2MS2J/pe5foYmLL5xb5fXxBGndqZ
/LJQNXTzbllr14cV4oWv4Vo9w04ugbYgw2B5qqwsEsGiFVO98qKIzGfecu5HOL9XaznSPM4NyteA
MVEQIAV5OwalOUbHQYDQ0mXARxCnOKfXivcs7RaIE/dLS2FzEDmlesvnLhlqw0Wr5igKsXbbAbaN
Ss/HRLwr+qMxObrANwekrKr8vVx3xCLg6p7krR0N1lnM3OYgOE28HCD7F1W1Pky+AyprTnfsCD8A
gqB1neVXE7DmNhKH0m8rD9+z9f/BXhNtq9zTAXtjtAISXdQHWzZ8wQsjW3l8/YB2BF9qnP0s48Hq
OvUipKgDR8J38CmsWwhzqksmVzid10psKD2jNWersPJSNmiUpUVjFUoIo/xGqSHd45uztsuwFEKX
Ejwko9d7mXNeV2Gvs32dj9i6bIx3nmUEs1fjucVBW4jtLsqfZ7Ag6m8VSzLdoOIAX+y7kHOWXy/e
VW4Sr0P/y4wQbX1/pWSc82eQMlVi/V/yquc0gSAe8evHti5CWd7ysgpEuXFI2QT+ubOQ5CWJbyy0
2ApD/RmwPYsvOHNds3s/UXRXLAlBbNtyfZ2yyvayeUci20rVCcLRiJx1fHMZejenWprGiuzJv35j
ca/zCu6qdlMtBzDUYyUx8YW7dcH42hqwoloTMtuweXSkIrirGzapcbg65TPZsIMZF6j6yyEHvWiJ
mvGyiOSUZ6/cHMaktLy4N5lSZCgdomSOtmSiHDzmddHh7ANEoSt5rde2C1yc0/q7z5VgZj1UuJni
HhOI0Hb6B/C9hreF/Xao/dHbpkMTGyIMKoTWjzYEOXxWHWGSsIG4aJHj22VF96CxpCm+dbioPMLv
7kr+594xWrVToDA8q0Y+hpHZ6suv4NJjZv3GSorHGFWProoRJMv9sFdk4F3EPOiuMEwvE2zdJPJ0
ooUmSZTEzfCL0FMIF0KBVbMatlXqwM6zJpF5jkwRNudXAJ5byi8ZsIhDMiy3/iVlry2AJYJOJ4S9
SuTTnoH092ljW/f+9celhCHlHcW3Sz8fLHx4Uud8zbU1JNUOXHpz8IDoeLnpuYrnICCpNK417xn3
3XdnNXkPjuoA+/FddBcdyOErffVNaz81M4n+i2h0wuO0JwbY5cKszyiFTl2nkQ0KM53diO3g+jty
bhteetZXPxAKIY3aCeB8fPOVXPofgiIQmoaM8/vFiltFk01cdGhuRk2+GitXKr5LAMQ/fhVcLduz
UAHtpFQwFMCStSMTZOWgbHSokg3z0iOjwoEI0OTWMpwoEelBOUQBlrFpsBhhkC3JL16dWBiGJfba
2cxapCkg8sFbYnDvb6RNJyUCq/EffNga9udNWBDPSZOHnIG4xHJJ7kWSk6N+HV7DADIwsFIapv+Y
AXGjjVtyE6JVIQ4sWgNAlEdOZHBDaJgBm+bjbr/ZF9ZFYu49qK1i74NFiEDdQtNb5N1Nei7sCieQ
Pn9FgxTzr4rTLWtJZn997AFgHFRKeibFWkQqgbTUSavgsTnOQuXytDX/VVGRuspjYX4LBeVecEGn
CBJnE2p8FwHAmGomCVyIUAbe+xd0aMgzr1/kCNAKtGMoHP9Aa3sqo0So2kiqXPJrcEOG/Wm706Rm
ju8zGh99cbQMKSjVfZuahTjwwhCXGUlxafUh4vPlZxdpA74/YxcAuGVGNJ76AxUf9fkZbNQgzDBp
NpVj+6TQ4NPpJO/JhpCOveiMAveBzFXAKsovrWCUELjIE/0K553sPiXxQah+mQ3RCQdVau4qpZKW
v83jQSnDHrZazIHIs5GivUIflVZLOdxwUuxkp4GKrj+RjnPtb0EyvWBxEa1dF5+i/oVPPIsvmNPN
v/NSv0N+oqgyudALkxkNu1jBV2Q2NLNChFdlAns7lvDjxaJg0P7xWoISUgaiMl/dmL+ATvXfw3uF
u5YKBWRtSOl/e3amS4RtCbFziXdGE+jQf393Y18hAruTHrFLk0c3UInpk0pOsnXOHz5a2G8xxy+R
IyeqPcvETBsSEne8P2Ok1DiZJRULCYr4sUBlPV017dxvi4ArKaMtIQTQ7w5qAV1nqNfOnqUzpW/6
ZeziE3C0uftfKw9M5THoVs9PwNWDc3j1wYuhORCckPR7t/8dPMCqwqx8FPtzRY1JqupOz6DY4bCv
f5wq4ZHDaduNvv6U+bovCbmVMBeDg20ifRBpMpNmXX8W4FbdzGxNVfaYP5YCaUPpOYIRbcmdwLr5
xFWAfT/s1H9ExuaS3eFFFlwa2vb7zcdBfu4B0zMrtLOuDrj6F7s0Am58Sp79D/m0C6hL+Sq980Tf
y/Vw+LB+YIktKkud/RtcfD3jCfDShAvGTIBSJRI+krYSyX63aKspuNZi6NF0l5YYzz/hZFChDvMc
B4zXahVtNbP1IpcW8+XHKBpOqm7584/CqnlGVxv/pO/SFfr26t6sCJ1lKM4eM+C+cN849REd/5rH
UUbxHvUpxVsTU15U+QprW4GAupgDJzXszsSbdv5Q0xfG/aFoL7tNtX+yX0DIvEsUeJB2WZc8VEAJ
ecCu1t6UwSKY5SvbAxl9XIl+PAwZdFOdkiZsUB5kJ79JTa/EMPT0ZdGw+mW1cuDEPO+iyjE/DpQw
va7vflt2mMA/P2g/FDrW8EopxTHpmsFD8lmgvyBp60+X5Sf8UfH42VbGQrc7aTb/klogxqtiCTFD
dWr1Y34YwA+LnhM0pefmDOYO2ADB8UCuh6QnloneueLen4P8ABRboOVnp1q5MtZthR7vlaOcUwpY
i5DUhtuR4Gbc2dIXS8AO7uskUjmF57XOLto2grVUui0DS5h/sVM5kspzJQhCzMeUv33lA3Ux1f+n
fmv6w+LrWtp+SymjQgRzHcS09WnM6wY6UT9S3znjFuy6wvP2Sfn7cNFKV1OIlITl2HiO/URoMmBs
FDJQ0/2qhDQBSAixXCm8D4t3ihFF5UUna/MyRZNhrcIBfKPuL4ZerK3gYBiwa5NnST5YczdZ3cDi
Fcz3PNR+d4l0R9cK54ruOrsfKqEuP97FRLZ/6Jsrpz8hGrZ3+CAFo1FE0OVK3Uo7m6v3c6f43+A1
QUBq2GqpEa+cxH3+l+FRD/E4fUNI5vgAWMQpE7zrsseJNmWdc4K+dt3UDI5BgntJmOpA06VPWp0m
D0yHb+hmdUymaAYRiKyggEdeRJlaZvzQu4XA2ab/J/FYaw7IPRJzwrt0GI3+IuELB2cQdyrAGk4W
YK/NPU3pxFYGtwIFZLPkH7GaE33z9P13BIc6CbGiNxnr+An7yy3IP9VJPCFSlWPGbVz6Pkm9baC9
N7lVaEyiNaDT+pIDj5E0V+k7zgIAympdXHQrj8KDqBXxnvHCSNRRW7JY+1kuqe5FxJWjcnku1Qth
64dO82FbRa8YHU0jkf7ZhCVtxu4m1WJjMWSWXbf67+c/firiAqrs6+YZUL1o7ZL4tZTRkJKr5jRl
/32b8sQLc1ofqoRONwXyhHhB4/un8c09SIEKf2YGKxe6q4teZswGHdxLiVcBtBVc3zkBFL6xGjqs
XijaYTXcrY/hgbpd+kxOHDrJh80m6n2lltwh4HPnZxEvWfv/NgloNhVuaggtobalEbV63sG5LXaI
mLhUTXCGji65KW5FLxKMC+tI/EmnmUvLb8AXMnQejk+0wkACePTQ/p/MYv8aWb5D6hGEDKkFeIO9
tapGYV865ma7MxL4hRgdjsRWBk66Oz9fizjIltG6AbwvdDZo85uq8P9U+ITTxxRywDAKciYPPr1a
LH0Vx7O1liixVqnv0b31bwedKGdMJdXHsbrXzg6lVhgAkYKeEkDBxSbmCLX/K6zqrYjUedMP4vbr
YTumYmubERs+UvQbbwfU4K2VDRwBz9aUjrz7z4rQcEoKU2ZsKTT2+NFAA68jkCYzfMA3gWDN+aYM
JNbLC97KmYFUt5JkjU+4pdTKRdBHGxK8XrWuxaF3qWfvBVSWbwEftF9ZQBnNDfeZ66BWRDnRn+GC
GPLQ1GIcHalT8Y4fyaUQwgdSPSBSMxtw/3CobTLEh1AF0v0wFRP1ZSL8+vtbPonJUv9wxNYQGvcq
sVVvsaRiZcfEdHXS/BI6UHba7Yob8xduo5McAGvYpLmnTIhpdTfqgWQAv3UGGtM7hYazVE2M8juZ
sYwroSU83rRULMB086ZfvAP7lagqamluEh1jPOeUJbiLXWhLLn6jH8b4rqw3tii0jBIU77pZF3v9
a7G146kGZRNOJvUbh5qMDMx/ya0dBERRswZZC0tXPjZE1xXUohRdkaoqbBMtVqfrj4eDqqy2ZynI
3JbUPcUHBuhduQj6C5SWQE0wQFbyp2e12SuFGdAVX+cGzeUcV7sYtGjgsVw6F1C7VaPGM8k9NKfK
17tLTOGtYiisKnzxnr64G7/Wp3kOyCQ29egN7YxG1370mEHn0a9RRMv3Rfhn0bj6vt2YJ9PkilAk
aXV0eOzbSlx9b1iIWlL9UMilehNqr7+puSlnBPXMju3atX3t60LU9ztveQHXPusePaWO7yn+WBeh
i+f88gKE6A4css5PHiS3p+cGrwu5oS797FAaCewrG1CCxFG/xKaTiMVDnT1o1YNpy85y2wzNjEmQ
eU227p67yG9O7Iy/Gw3hy36kAZyzcNqvjtqdaRbILRKcPGYSOBlr73Xwmj9ObJerIJHFWBvRHmim
D6+T7irODJjxPVqz0LW4Yut5hLz1XIt/l6VEFm2SMPVq7VY41tiz2Da+FPRE33JVXJgLxCd8SecL
mf+y/hg1Ik86c+apgMxTKAWFILKxTZU16mvlPO3Ozw3tmYyyhgA0NUloX19+4PYQbf+fdoc/Yjbn
PorNkQlsoCsP8pVmI7SGmNlgaS3nunoQMfUGoRP4CJb3gMSUbgZHn/sbY2UiUegkK0PU9iZJLT4s
zdG28TRClVa8Llixb9GiTOaI/gyZqw2azlC3l2fEJb8UdVR8UFZfvJsM4d+ReZUR5PND3Sg7CgGQ
ZHPPybaOkq8bZLi4Kwl9wk7GYmxWqzeMDiSyhDwtwXFWFS0kbdhXLX3+iJait04dimT0RYOJa1PD
TGs/zN4QNiUZ6ernHrqQ8MwqUgNn5WeCD6lRJfXWxKqKp5orstbPcGuCtg6Rc6m5mmfhanS/u5IL
bCpC8TrayHwWd/oSbOAXyv+9ospItKeH1M+PUbonj5+gqTYaAnA89VgldDVhNnLZiW9XNY2I3kfM
kOXlieO6rVAPKIrRt8yQcjNz18RErhh7u3cOPPWOPtXo+8dqUa4VDWNZYoB34d79b4inO9BPeo5c
av7FbB+da8Cmih6ziGNLZ+nJNn1pJRMeOLCtV5+HNbJ310rmLk+TvgMIuM24mcv0fAdA+UAXefTw
z9fZGGkm6GQ8Bvf2uQfTq7FVvDwgQ+BOSvui6+u376YDEdHrp1aljHFB6OczaKYZ3fAf/Ypvjb9u
UDr8+1LkIg/oiYfCH7NP6+1FNVWVAEnxK+TECnK2oaFdkYH90szXj0URuAFDxKfaHd0nXqw4Wgfl
dyIdEX2uXSseokcG49sQEUEIKFxrolSCfsb+rJzImlBMrO7Ud0q7BXd2qcjfBnHd5v/xC+Jzp2Pj
/iK7Kdgj9dMwTbowPHEubcCzvC8PAzPfA687t56fLFdteY0Kn87UOAdc/CZADQtJXfYqS1v9V4Z4
JDkFl0edfBbgN11w15zCEDKfpUKPBWBx4UE7rZ/B0bs2FdwQ1381ANF9yrUZ+bASjzaY8ZptOuT4
Bf4wOFN97X0XeS6UFygRrLgYRcuuLK3Qv2mMX8SIygYhgkESY6DDTltULIaHCAeRZKbXdpYsamiZ
jEwoPEeEOsX/ZuTiTkL0VfqwiQo6aQAw9sGsVjDd1CgFQJUA3vraCpN7UjFloh6h5dgax5qK2Lwf
B7HhHlWjRQ1p2uq4yrUqfC2P2/IwvsabwEHZba9hcypzf99eQ3I7tQMo9gx49SwVvexG1/zR5DPM
swY4oBoYJwV+h9ogtjpCi8ouDiCXapZtg9FTjlYmSGVsXSnMwhQJ5sBJti7TKcOe/TMujbOC+Lmb
6WRlFULS1FxEaENjGKyPO7XYtMaWB4op7EJsIKFgISOLLFv9gy8b5zMEm1sXA8v1CP5CvZKX4AI4
LWaNUawc3AZ3knLyPLlrusYwR7qvgC2QBCKNKdmy3K2Nc+ImAyIOwwe2Jf6lBEhmVGM82y4Y0KDU
y1HDRXTqBJd0MmLklqaa7aHkq0qWDWfDV8SpEDL7wfdu426aiNMFoLXhQkjc/qGWrGgNbkhaHt63
NkK6fXyTbU50SpqDy7AJCyFjAHYl3gHGRpDH10I+zYhgKXcR0gPG1e3vQt6YTTdAGWVIOom2n/tx
4tKHg/QfZ3qE7zAAWMuGLlSZjJvQ3FXRR8MRYafx8wTSkYExMxpC52RHwir7UWANm5hskpoV//vd
d3RGopeBCSsVlqkPj+kNU0fqMqCnX/ZC8l73LVndr29Xa3d59NvDDshhnjY5qSigeB8BphT4ZvAA
uh5jSfdk9LTO8LsU4smJOl9ba/4hf0V3w3STtb5g4Lh/P+eZ848ws00X+UnWyVpdt+JaT/nECWPa
r1mTRt8ijnFScj4iB/l84eJ+UsO73p/DZQlaGfxO8XQEWm+5AodiFu676DjUS0OY432k2+od+Dai
ba9ItbH+Q4EnpfAN/79SKqOqUyln3jli6M8g4zNq0NSm8l22xTfQQv+KIIIKnlYed960HznNMlfD
mmAbJoULnqoWjVRFxr29R8tUC1XU0xztiWZQ2/Gvx9tgAhG4NLczV/UrecUbvck2XW74eIl/33et
ILjVhuyEMqwa7k/DvvAkXwnAUZBlSlu6zzXddTxF6HfDxhzuMVf92R+JwLoZQd4fyI3UkLA7+IMg
TBapTkfqn4aIqXAKH1+7eLeLZnA9BzE6oe3dwJpa8EtCCWHX8Gvfjy32zRAEqczIgwn+5+OM99BY
c7uW0FvpMCnNEhwFq/X0HIuUsYSUq+r9reiEc2j4ej9L14NR+Xe9lLvdIJZzCOmFVmWjX2KaUDZb
/9EUBmFGCUjIXh5ueja/dA7m8cKZZLvjWawjtVTX/tTxWgeemDhg6vspPIoJkNXP8+LmT9FAcFft
H2vmutjNFVMGtST/3FyiDfwmw/CZ2pk5JcqsoZPmEsKrV+W7U1vCB3cdTx4CCsPabb+MoiM5Q9MF
yK921bj39RqW76BrgQKO1LY1Av5DFmYFETwWV5gQfOIssLjREru3URKCM3DD1pxuWLzR/5USV5ro
NKJCh0UGDT8lvjjClhh/MMwFXi7EWvJv38+MwWqr5NEz69YaNvlg9AFVAzKeipt58avmvalv3iZj
V/jz1hr8jVLNwhBL1MghDwmHLrB2PjwS0rLtnJgiK1wCwVdCCkNoCpO7+M4BPagQvJVLKruOe+S3
PNohKAXHO5WvxKxjjYHn3njB0JEsLfsZGPARIKhGGuyLQzGiCgBoy9Vfp+WVH0k6Feokuwv8Fq0Y
0Ph/njRgCFE/xXMVUMwnNblikvmk9ytQ1VWG93xjwM1LPrM/IHsIofd/b2CGF5zjumtoV2G7S2pZ
/vVnUXX7oaghJfVSJnyu8Lbehse70orUeVDVkbURseChhSyZ3fW9Q5ltzmhS6dzf9lqtc3X/ru2/
PanlZwQzcc0b3xdAukaxMEdtOiIZ1Cru4k/+gXlzOC/H4zY7JdWj37fDlnS1H2dBMnmMAp3rqxBc
E8zUYZPBFrR6GkI4rvq2ONseDGmXXwuKUwH2RIS+ZgHaoI5Vg76b9nF24YeTZMd6fLztV7ARenyD
TMuis0+0WZ48bigv1VmKvuzwvYqyyneFguZIimtsgTcL/R6zWnHWovYLN0mwahH70Az4pYQ21pvO
h/SEQvKLdOgOv+W7yZNOZ7tBGZvCVw1NUVEGKn8mVaZzOhYLmvztK/tjKJBpS/+op6JJ232lHYmo
UiFOaLeWMwj23N8JFpxpyxEyQVD0i2tuTz/MhKXPTocZvfJg80IFjVegx8K2c+aSBpBU7+1xxw1r
Tq+yl5lPVdadHAi7SZJfo2+16nERtDT/ZaERTCO+6Yb9CXH54o9VM6IxFv43l0pU+iF4rMa25xoT
3iwavvZnuI/p84k9VXO8ZY3O1l78TymvtXJIJKdRAvJFOukz9afZbpXh6fdgHKViHj2MW6UAB7u2
z3U3axSqZvoDkoMBuSA9mFp+NVEjTik6U1njXo69VaA48u/Ky8K5uWD5QWOw0KRqtK2xNguOzmqu
7P0HVzGNZnQzE4fHGVIUKA8GXfTD4J1yfV37XStsD1T1DJ0OBdCxwarIc11Xdf9A1ZhKLDJeha0H
9HLBKjfp6yIX7PXMvce7mH0A5IayhuBNUIHJy18mpYfyESSTB3SXp4AGgAieiE3jwtd1QVS/gGIE
XTqcVz+wuPjkUuY1f+vB6MHUcxmwon6V/cIOvPZQQtEIStLAHtArYWreqpa4lcdZ0uJfp5BwU81N
6IZjX3KlaxKPriAfbn6Po12+q2Z4Xda48epiWnj6H14TnCUNKDEcP4zyxwp3l7i6RffRGFdKnyGG
Xa/NhkuN1geDZWA2ayhI0Q0RQZKeBtWaIe9u7nEFu9RvDp4b73Oz5A5CWodxgXZXR14yvz6gJ8GE
cnjY+4GnvH1AIr7DK7sMYZ4uPmxTyDygfT5z37tOQldlrRcQXbv/bGdGBfgEfC5lMftSH/Gk157B
MSkpfiwEskb0TP7eDd5r2ZWpWiTXiHnUcJKOcKD5TcpLdc3AtX3xBO695ydG7hhkL/p6kGZAQKfV
4O/9VwSYXtMDOui36ow9nSiKMeXpyKPcfdTpxsl1mdekvnqwQ2GUnmds9alpSDx/bs+LiG9f2eAz
pf4gpMBkM2ZO7v7Z4oKhj/sKMo5JUuiw23X6Ip5Tck6msLxj/2/0juIhHZ6gz+YcKCoyNV1NU6eg
XGLasQKdSbU6tWTdU8KEZaejoH+rN/KX0c6bc1AqYbu2T0al+L6BggKaygNRko4dQVlDriS9W4EI
h+fxO9VSrF/Q5BuC4PP/ok4cWggnQ5bgjSUb2Jm5fSOE7Q8xkyU2REE07QiQ7i6V8iOD1gUPrxTS
rUc6ArR7dQ1UQWsQuLlcZzshrEb8Od8TGEQJ0WRvBD/wuYCJz4VwW7awfzyrqkBEox6EAHsaCYyU
gQFVBJSzYQnuwZ76o3LwVhzswci+eekNa6VnDVLfVdUtwJ8iK+ruR5U0VZG2iPY2TLDOUmcMLY3r
HpMH6HzAlBP39cGApxAHYr57e3zZCsWsZlci/INnM6ACuFsP4sJ+jqGpxpK3f7HQH4nAaoh4ENoP
C9zl11D4UoMfBZHrjoSsS/XUA0O38dKSB4J64vhvbplIIc6cMnFj8b0nih5rTF4uk+uAXP018w0f
XA30C47W2luEFJxgNbtzbGv3KqZnwBb9jJHk+LGo+q0OVbTllZ79RHP59u/DT4UoFYXBNNjFBncf
whyF/lGIBTHB8JJeEuGLUFGZ2x2dL9Bm/a6+0qibWp7I+viCHkp1D/4O6sRNmwmu74f0CbcObFQv
x/W1dyRNLJUvzTG6Kh69P2nkYCxo+RdzrktnOLtOQAFUppT6dTaHAQccPsv5UCGYPMuJc7x/+Rhh
v9grvgVyBUCl200qBheh+9xl62LmB/JS9FAvwyjtFtACVYkw9LPQV18yS9h/beeUiZnMvNRjL5An
QUhfYrLpFZE+12y0yB7s9/3LryVmzKwBLGISC0R+5Wz8u2TADxoVEj5+OHSk3w3XZuGqrd+Cf3Rw
OJJVnmTlzh0KB/2CCVFxFBXbpNp2DyXRiZamKQS0hebhwSlRs4YwN+363c4wBu7AIwrgKSFOjKyQ
8NYCE+9BtpwAmo2tIUSF20XuVavjYNl2ZPTNcwNVPWmL90UzqKuTNB6STgn8RMHfeJTSXZnpql6l
l8rTNss3S4LPP5/x4U+NL2FdrLiWPxaGicpuP38kOIjuAvPzRHoA7ILnhKaN5fXsmy5nxrwp3DzX
G3nJt0DbbylIjwXOIjZqBUhlEInAhdI+yalDRsH9cesjkpQawiMSKPLRbY70ww/WvzL1KbSvzSUc
WE02csiv+9r6jF1hPcut4X1Moome6duXzLnybbUl5IDp7hplq6aE3dAJli169GwzbGSj3wzN1Cl3
zViws5JlncMQor9L6RqL7441+ry0j9hkP02lSl4Bk15UxT/n6RKp91v2y2LrL9K2+JlooG2WZ/8o
55R/sc1E71HJ8QWdIOoCInPIQ/RONnOzgXr+uvUxwhHv6kbNmJ0B+ryS2/S6tLQ8l6s0LAnNKqJR
d7N1QGipuWF3l++S+IWBsEBsZHnfPr1QiJ5QjfAN6AuMERiGLtS2a16wL568/BVpLbAxnam5CoYw
WrDpND2gQYBvSbbzO6opfqKlTN1CbLpFQUvf6vIEVTzH4oH+/i6RmzLJogBJYodlHQN/7Q5ULHcs
o4NCvnu56ak0Ae27BdRVwF6KzFHavzQ/W/W/FjhPWxT5Od26AKgWacS2N/V76jHyyDI1ITqdE75w
t/nZ8YbdwbU0OYgaSfA51s6b/0pFhK+OH3gNbKVOUqaodbNsy/zTRhgJ1ceaeXrN1FtbObdx1nD9
pXoZXGpp3UpCT9fE7o57mPsjPt3xK6p2P9D2kC6pPtDHywqVumpB2U498reyftLvcekLHnAi3jk6
K1dMgtcPGPutY9MkWzHAc6wPL/V7Q4nhOCJG6oJJU/GOW9brivE7erWDqugeRIdE8PVlvQN70E+F
Qz5jWy18Dt7zse0leUbLiaJFa8b3TSvUkTGSURHpm5f94eJjflWZSLg27/lRKvZaJjw18v5ykip1
0W7Ynku8jbLk9iCFPcypupaGQiV9rIEZq/CXmwUsFaQJvmwzLq/CJJz/LgwZ/xl6ziqQ+O3h8z22
49OJkFIQ4D/qu/ni3bNPUIP8NGIZ0L/JnEH7L6tSudTSaf8ajpbYj6AH2JrMHI7GYiRYFHtyZGH6
BuTYpsJs2A2t9qGPY5wBoKMJatuoM4hvzwekkVJjQvHt1ISk2swZ+ftRQoaymQYDLd+d0IkzW8Rh
0sO+iVMl8NNkovxpFgm7/FVcqts1pNAsLLRBph6djp00w2dLioyI3WGPgMo0hN4S1GxS0HV27Ybi
9ZXNXDIh80YhyM+IPUfMEaFQZmVE61d64GdGOMkt/if433wvGHnTFKtVW4vMQwLh6nMWpPOBs6zT
zZTKZvpK1EyuCy6/pUHAqV0UaXeh837QampKVnfMhQ6b2zNTEpAyM3H77Xzy2/2RUwOv5aaXelAE
Q9OcbY2hUxUswE6MRQWv0YIK4lkcEN3z88ZZNSQYrflDDmunUqetme5nku05eOMM6Y2J8BOBs5Xs
wBzEnZvRg5WraJ6ZlIDUvmwdWv5cEojEIn2CD6isfftsm7ywD0U5FGLES6xlzMOGkVxey7T5VuSr
QeLoOs+NvUNSiuMA3MDslAMVpudkRgJuh8y+fJA4Qp017PMtj/1q1tVvOItsttj5lcHRGi2kiWTX
ZBbizWBTi83+btLVvBGLef3+SOVNOQFO7gk9vonv407JZLm0uMpEqiMhfaMWsU7IHr063aIUfIru
uJVABFlMFtviPNixKCugeXyiRPEvZZ5QH4D4UTAFjtVXsNJIqaA9Ih3LZTd6hru9Xqg6wDvnQ1Xj
GBIs4Oj5H+jx+QhAyE9GsQ0GLFt8QQtr9VpUatJeZ1kJfEJ/HtlVKeO1O71jD+w8uy0MIBDC/gE1
NlOmF2Jd70PfoMRuRrp9wVgORaZCEC418VPgXmi+oRitr0sucipRLZeIQDdy8N0FCCuQRQXZ7mRd
J5CMeIlKUqH8bTpbVR5yVIUH+D4gSrNLzfFOVAB6wj9mdp5Mdl3WMx6HV1pogWPPjbE96L83i9+C
0bp/dfW2nt+XRpjPEtj9ToYIAugG1AONQWuBY61/VWyhXjq75+FX0Q/tFR6mze+KiQMXZyHHsKEB
+2v1QBTL+YeQDCatl6kL2F3g81NkbMyhZvNPSEGSSnVvX8O8fQhIKz7ul3z3ISXFO80KeUA838V6
lsnbM5HjHXWsUovLmRa7B1lhfuxunr8Z773BR2pWWAca3LTnglzY1vgD1HdhQGvcdHDBQIQmkI8+
g+u9gd4pAnRQVXUFdGDzXB0d1jIAl0mjx6HapHqSE3lFtJwIa9W0BWUmtxTjxI4GWksg5HaAwsBa
OBWnv89a7ProOPh81Bq5NIlwENsd362cD0/DmWyjI61wmnM7MMG2vS5/zX9dbmKf6ORnM/C7wzom
4jsb+7Je/VZ6ADq1x1qHWYe4/YcJq88YwNadLBlAsrCwCmQ4OHlPnr+vy28wviFpdKFJ4DqGxp6f
4EbBi8b8TCv4pYzf48DvILN93aRKhBIwoQ+dIwXp++XwtzBJYHAMjK88hHKXvdScwAwp9tFQ1nXs
vDlAFWqoFc8fqRarKrebKMNU7ztU3YlqtHYu2Eug6KRRLIgzkg/R9vPgyu2K2x+GI3XmovYSOqz8
ULN1l9Dd8kbVLBfDGmKo8toBYd5xOnC6sf615drmxupl1+gdQrJJ9vSP8aINLciTOib0UzMzUSoL
689D/vK3Ea5PiaS5j3Sht8AN5IsacT06ZuZkNJv8GC3ChNSs0ru7KQhMJMrQfedUG6T+3yJLjXYF
mqXZKh937JPr1+g6CUhwi2+14ZjUB9Cf+TmMV6/o73879tf3TsLe+kXuZE8uPZ9ygINmysVg9VyJ
a/bVuH7dB3UREWGlYH77Pv8D5PkW5xZ0PwO3aWkt6/Dy+7cfOvebfmS3jXQ7N6jhSGIJfklTyydu
skXeNlMyrOX5D5e7LYbMDbldoZKLdePp8YeDar27S4aIgo11qgDh2limFBsMw4InKkqsiD7sbtTb
XD/DL3PrgnrZnh2oR9crFsnqHADwIB6Mx1gKTTrUkWzOfXkgMgw5XdJjVPQ1CSPxfMYofM7E89kC
HyqiB1ckcdgXbfC46pKxzJCeb9FG6JXHelycq32kdHdL7zgPOZpLIIUixgJRjMpzuku7Wulee1kx
6wk7fi8DobcXcZGvf/N9cASDyUyMGwLGrzTLKkfyng6Y1IKz7KLJ5OgSWj//r8B9TEkiy/dL4soQ
3iXVcZaCaS1+EDpcxEEGhChMPKkwEVCtVIqnsyGu0eROFTYqJckY4lrJx9IJdoR35PPk/unNJUw8
tBNvlCAQcAnhutZVPyl1e7Qs/3WSM+gG+oJqzGBteSQ1LcS95+fSQZsPu80t41ylyJFN7C7p4xRX
UUUs5gTARt9jgXIEylMSYeM0Kv3wYvxlzNZ9kaRXcK+zzyCw+gM5Z3w4iRRgGMRIHsKusKgHGzz3
caAmY3yp7jKMr5q/HLq3y2m2JI1LiOVNypSP1oYWpwpWQnqHtf2eXkky7vfohA+b7FZwS0qKrJRq
vbuOdcqJDWEqmsAtBfyyP/5kz+HnK9VbQjWsN34qqQvR3h0yZXAchGeJ3mxXESNPQB66xqMCzk/y
FINU/wxUtqXPXVxGOKDu5WVC3uTcxTsujPGrsC4rNbDDuWh0xgy0CptvMf1Y+gkRS5Ac16aHfx6w
6B4GaY802j/8b8sY070K3Om8DJ/yL7IexOM5TntzhgPFKyySCDB28DWom3aQmeH14Q3jNLn0FdbN
Zj5WAWal20HYTrCHrTLesadw2B6Qrday0XZIc6t6MJfCLCif5EYzhRtprKCJt124P/LA3gF1V16n
V0++rZng6Uuj1URqg+s/cOn8MglEfwXySSnGmpmNl3XwYVs9+YqFCffAy965wLk3rpT/wwAURaO8
+b5HALxdMrL4ODnbW7KMFxw9V97lEEPZW8LUiT8Mffs2a/lupBn1eKTJRHZHgS0BFcE4FDbEKFBK
zKGVMCJIKlzBLpn8twFJqUjrAxEABk1E0871MvM9hKUdVarWsLyV07cLMSqit+bPCtl6y72t9bls
EftNr3pfN0krCXt/My0AMY/fJv+zqfr6DAm1y/ZVUfZV6OA4tz7OglXOhvqnGCKgOTH/XfqO8wh1
l5XGEVfldhpZIWU3NEuHMwhlfdJNYPjtfR6FWsP2MXFc46v2f8ZiZ4P8LYY8ibz19aCAxgIxUs8Z
uu4PePJbJKPbUHQXSxsnVtFnrar5MTzz6K/UVe07LFMGeB8izbIaeHNFJ87mn0CT5fmM7TcsbV1K
jpfIyMCtb2gXJqGe0keGL150CtYftjL4CiElWFdgxSEErRA7TeuDPa/F4ODbu3ng4MK2Utw04Qut
XG1yaGrvcX+lUsmbs9CQNUuEWf4rO8yyhk36KUelViu9FKs94oXx85N2r7KC5cyJl5Qfsk2siDKp
rElGfYy3Nsmmq+afoX1pvv7UkmcvG2On2utIc5Oa7qZccWYZdGuXdXIn5LWm3d6ADWOCGUuIMH9C
9xNxX5JkRUkicmgvw95dWmOUdgAsot8G9MAkzaMtH6r91KnAowxT1VQFjU32ciDDVYYySgxwnUL5
YWtBsMUE6VM5dAlPT37HtLg7z8wO5a/KBsL35HXPEfk1lFIMe0iXu7FDYzCLWhOYKU0ItExHW4/C
6ymB2sfNv2NnTGDsIeod/keQt3mGThJvwmsj176+MnDjhrAAfG/J6USB3EoOu9cxZtqqC7jpQdrx
9WnDawsqE5I5LNlIJAUxim+njY9BEZbzvFz1VuJOPQFVbEMSPGknCaCP5gFV+MazkT8VtuWUTpkJ
LbnH0kyeA9Mt1/BhrOZSQ28mMCp1G98Gj9uHMgbcXPZlYNiKU55pqrDOQDrXCyYDloylUbkGj9ku
g3ZXvlkaz9hNMAQY8bOjEELUsPfsGLa20qbex1N+34Fl88BjqdiGA6b2pr+wcm/IUWYDMNUw1Z8Z
0rc3y/+TRiXOCZJV0Bc9oqaoRGIbNcmcWFVomlJyYLemaI3NuX6fBVFjvDpvSjbsPK104Oqje5y4
YX7Vw/mC2FOfgRKl4OHoqD+aaUAAw1FsuilkCyuTPUacu2UKrJfwTs/xNnJrAKGtUPXRpV9S7NCI
hIK1a9YES0giV4WdyENcOWQF4f4SbPEul1Pggi9jyzqQOnAPgS4oMeVzDaCedvDh1qnhV+8X6S1Y
1szXbevShnA6Rwu9XNVUtcCERHajxhv4l1jw4TVJk/a1+M6i2GEASHaTcsUzostZB2W7+xzoLgzN
1VG7Lvy52JUMCW472n4uDxsHiakovrFXkVkjdkzjWKFCmeXsiDXNxugbbXcz67WePqEszxKYcxf6
UT8XyDwdmb8wOqTZMFWdIRLTDnli1+n5CwWRwlMxxXGksAQTbuQR2rkscdezOBbPXLX1x/5uvgvk
iq0g7czaOgQJVH7bH33OKP8YMavj2Kpc/9zo3kcQC3ksFVGnmvCkjBaqC+B/OhO1znseSp/ilYB5
0FKbr0Z3N2zy9sRZ9mUER+CsPbrGEXwUCEL/QeGzuFnwVn3Mqq6EUwSXKZjyt2hZObS5RQtt26oa
ChXa/wkVk+/4Rz+sAauVqRJMnJ3q2rKI+gk55VnkrQQayx6E0qiz3vmfv2EYdLhqjlKZS6ckEbyE
XTKrFFegsp50J0QI2mCkJ0jswL7TQBIoTyBX7cL66EV55aO2xZEXRnfZ87YmFFG+xfbRsCc5ejmk
Ei935bB1BXL3bzXDXz6scrKYD5DdgILdj/rZmgWAIsof3R8K/JQxMpSZZOWhxUanuIirnP2itefy
DShL5EQ9+5GqhqGzyJQMjnFxDiE1GMnl3OQuBaRDskIRFaztmiQHVQWcqLTPYtMqw9GASr1xTGPQ
6MJBYS5jrYChOmBqgUeAlctciYQIgkvFt13jEoa64lir8KBcKMXyJ27719luRzPXH6yOnbcbO+2u
ceRyieQJKPPyv8F3Tc0kPttBkEaLzM5RsofIlbjvJgOZmr1pwBMFM6q3dbIt/eVGY6gNGs7SFN4N
KqUuZhSBNu4xz7st3XbkI0syeIqKngIWSWrKjrOz+X0UGqOAGBPaaYDOso9uCiyhSPxMBIwl1eqA
TEm0DBQZItNVnqKPVLMF7hl072hI3O6nfJvFrYEp/j6vz4z8rTHFy7M5z47OmbuO3LiPH3vunYoI
MJTz5ZvrivKEVownzJ7n+1LryLY1I65QQ8CgOFwEdUKNGaWlO3BguZkis5jWyCpf5S+z3L6+mnR2
1L6JMfNnfGH1PUlkffUGQo6O2SC6xQ0VVffVxLQBH7tBkehKvZ5HWkuc/HySOgOVfQzD2ZMYp0PD
Cq+X+VqTI2Cqk+It+VJNEr2si3k2uAjx2utKugGkwGygJd5qBn8kYjx5pyAdmMvVEpaFY1pSs8fe
KeL6L+wI61/li8YuBmVuAz/cszHFtjUcNVEuw2Ia/wNaMb+RgNxDvw7QzB4JqcLz3eXePyV/q2/s
oVaYZI0xCzuK6e4FItl9LACKsMp+fwAhnWlyZd0UgJCrTd68piSqlIwtZOd/kshYMAyzpePb5S4U
CTwv0h9ZQXIXI7OxIv6sddOK0txfW/Kl0wumYzQURetQytmIYcmePdmQNK+y5HJ6fSADlNn2w8mC
Ic7/225K8pFWADjqjJS5RM9kf7J6UOqCUgftYzqCGc+WB3NjdU6uRCiwUzVBk856U8q8bTKUIclv
cpftO2tKVxmXn5PFiDVmsJ8Rj0EP4B8Cw5OPvRubKpi9iPceFk2GTlLVIiGQ90Myj6kBPHfM/Urq
YWG1p/xepH5vmyakxdeqSLP+0EbqOTtS0yphBJtxEOb29vMHF5KZKh1qbIDQujqkJ79g7NSlnEtc
iPiuHfZPkdRG+Xzaah0MF1jP0hXg5Wwl6Zqtconl+XCkeEub4miJflmeyP8MdMIWS6GXizlAdSVJ
YA3OrxPQCamSmPEAHPzvaciDlBhbgvvvWVza77mdOi36eCBqN8TIaK93Jt/mFBV0F7Xk3ptt9diG
M5MJiRy/s81WGNSDquW5mDzRLgo4C85+QVBl27807s/Nf5QumXjUMOQS7KMjFK6vzbw9Cu8sQeLw
xHBsLkcr1oedA3T8qPtNkWL3GeAnY9Ps8dSlxKJEMM84uLWqjUPql/yjKAq8PtR0bFzC0SMOtMcq
/mFMiTKJm50VbvS3Ga/2PrDWbqvyKMjr+bvcjqJuOcTQn5cu0+dsWkx2YQO20FKe3DbCxr0Kp4zh
c25/eoUyC6sYm40py7r0KG1oqVfKA++DAgFqY2EYncuKqJ4LY/zDsLy4yxAl+tLEtrnhyz9KZbtr
raxsi4zYyQ/ByaK+2YfVQq0iHG7e3KKgCVQIgCkO5PyXMz7lg/xJ/dsp3QKWFfX8Bbb/Y5g0qvu4
DHBy2iMiWbmjBtOs1AUqd51HjTu8RHL11DvrBwQlY4KdtuGb/fnGKAfNLCyE6Td8lMGMUZ15YnIE
aefSZ6kTlOqf8mjyV8Mrt4EHiUuZYHfP5CYD5d06V1l84JVzL69DD3D42f2SFvup1lnXmKouuXpw
fD1kKXd3EJy2CbAw3z1j0w+7JdlZP+i7OY6NkLGBmkb8bhn3uCoj9dHrk2NuEi5jiKxhEQmwnrqo
rC6HuAf4bCbv+4riG9XwtlYrSDtv4G0q/68aG9wgLKZox2QyeF/eElZfJZUSvTFsgI6LUiJg19qb
J3X3QLRvD0mjtP4NkvZXZKC+92CPjfGqWBC1UF1CVpKcQsvFRQKMEqO2oWc/RdzpRFfaJCbO92Az
JADidw+73aInkhMVV/0vPBi0KibmM9wQHtJGFXLIf3PNp/H7FSEatErtDrGBWAts9ilJRMC3/ksk
EHA53pVczKD3XQXjN/8BB7TnkEe0nh/zOTzmVotmjDri8wIqsxUWfXIyxT11VXySyUrnPllx4TPW
zq3NlrBTjcsoEfmhEdsvG7qnrXnpiReZsAzcj5p6AQ2EFqbtp8rU/5QxmSYP+wDR6LRoWUsYCkno
j/CvGiTAZeVhxPntJVLlrt9eFZ4GJLPfPIhGEjAiEzhEg5gmlmb7iWIo1yw8cJ6h1kVupTepAxw3
6/H8eQDsFuHjjbzYUrEEy/L5VZgQ4H2lrukWFsIYrsHA5vyB9PjHbO6K7yKjIALbEZCaCitMZc9p
99IiNVB4v2gQJ05X+MoQ8pZcc96ePhJZ79r1znQg4ZQFLJ9ySgg1pa3IFu8Sqvu7C38idzVSSeuh
2ygUJAKule3aey3ZecG2tPeaSknPlNe9jWiFUh8Cv+J05IgolQo0QTv8Nn8x8uQJ4MOyfaRdMkXq
Hzy3/4sphayMPJOi5FkACrCKoqRxAql2IfzMK3l0PjsqQIox6iqj0lFa3SVT2+tXdoiVjb3HlrV0
6PApqw89HShhPHUY8Mmo6Ymew0Jvap8BYnWargipyIlYobMPqc2R7oLAnD24Kn5afpsmaGialUjR
sdIkXVIsLjCaeIY+zrHiWvaGIvht7DkLbebXghOkXp36mFTcmxH2DGMtbRW7nzS6tCEzo0iX0iC9
zaE8Cv70ZNS2uuXtdyU/dJB98li/2YHMvFVIbgXkjFTkjxiAndZTwX+GX72yB+tfcGoI9YMp25iO
ZwupJ2+MBJ1NJQnQr8JWXk8hpSqce3eVRnpIdJsK55/irveQKTzqa7Rr5IGxUGahjaAlaUSWFLOT
zVbxQ19UNO9j8nlf9K+tAUanvkfBf7R+ybT4BTYk5HCHr6aJw97gU6IBnja9mvXK3QfauVVCKRR6
dzig3GsbZj0Ym8mGzEtos0M0CV1pRdR5LT/LHiPlqw7AXkKqkjaXbuULJYv7Njm3rXnOwQccEC/D
uZzNY50CWAunWIGKS6we++njSb7mBEMFDIaM3AFL7BEEk13YuqbOWgoDFTFa0xmvzxp5zFXNs2mx
UabR76VpWAJqeLmRf9lhgnew58qpCjdsMByAjyhRjlNi2hxRQlCqA82X6zLLgKYWZktVnjIAO6W0
m3EOV3qW9BCyDUB9Oygn5ICSrscozaQwvDaAHRuLI9mYqhp0f3vX4c1I3/t8qr2bk3iKt8FxuKa/
FPsotjaLven+xIIzATO5BNhbu8DDCbJsoL0EEyq8CeJ5XOPDN3wsUFOgXf31umhCNRXch83kWOot
sh55Am691BjQ41nW2aPdfJ/mi81bheVteK+jkgYBSf+ah1hda9+0+2I8WV/wXPCU7r+zeSQeybC+
znAMB2c7eKSh+HpiKhB2yc18PZM2fg2Bu/TcCMOfCCGT3Y5KnNUFl+l2K/1fMxWRveUYmIKZ/dxS
Xpb5uJexE0irYJLbQWL+6KxSDoTrQljqOQTv/zLnuYfp6baqn4xMnZC0k9s/bQWcYeSeovMH9J9o
cArBESb2P23QjIVQddCXWE5HOtVTLHYKQSwP/yKrynRCWQiFUap1I1Ku8NqbECZGFK2eXfQhraRw
Zv2qJYsCGxmppq03z3szuiEDkj+HrN/Z8s+EzQot3XL8hfgUKrSVQ8wOqz6kBXui/J3vLTGmz598
10uPdtHn1ZepOvJynH1uyt1ANEx7WghrEThDBT8WqWowKGiFTnMkNh5OI7SU+J+AmQgJ625cukpt
5++WNd6umBqZRaBaZ1OSNSNvb4f0ik9MCSiwMC3K8AIq1zuLIOAf98DL0QrydY9VEbLQI7TIo+BE
LJg8wQdX+Sjun9r+NrmjLGIkcJMte0AowxLFtu6lTKX6iD08pxjOZ1cJlTiDt2E7zYn1XjW9GH2s
tqDNrz/X/7Ouu3qcY9g+FNPtYOx5BK+8vZ8bGPAvzz3J6Ze1mabUNQ6AIjc/6WiYfRdG2hkL2KPv
5wq1m8MYB/m555YJ/bUlqf2sBdNCTI/AzCG1aplR4R3760Rz0o2496zEzpIoXDkHFGboxdZGIzeS
R/+FwkCRZyKLQfv56RMtJorbDoopkfWdX+EyWa5kZi+rkmM72GZXAyrX2qYZjv4QjVTDeVVqFn7+
NdlAAIVBMmPP9XQJnqedwBHBB+IgAv9t7uVAcazOrbVyQ5vD5Erw+JWzqRkejhGboNiBdhvOyceQ
EXiZ9vwrNmQNc/J71Cgf9BPdoLMXDY7guY3/xX6R9wIrltPGIATYsP0dLqw9bGBNdLsWAYnRypWr
KAnIcal7zkJu1ayPx7T7NdaKJJgHaVZtIHJc9vUEuzGXL/rUnBoWa1ECzhskBV+3wU2GwzNuqBIa
Vlhit3ON4tKLw1UEA1feRakqx2bLGqRVxZhnAruLxUK/sgjk0BBex9RbUAvoijX7kUjyKJQemxbC
sNukbL3oqxUOK5cc0tkgU5yrJ0lI0yQKNDIz7XNGgCIzfpDh9YdrZeoKLnXghpZgjdO+aUGVGfK8
Zl6Zy2OwhXkiwFG6IDCb49d9OlIFNFn1J8tsaIEOxaEQ14RME75ZKkEzpwEtnR0aX92tYFh4zTYS
7wKevbSJLSAY6ZnDX8isHW80QnEoNlJua99GIw3zXB53XRFm/0rert7C3hCIvAbB4IWJfbMwgQ1N
PmrE/zh+GNTy6fiim3O0rnuQ27hQt4SgWY7TydQgEyyxoW6agGH83ozIwHpJKiY32MgpO8ESRC/B
bCG/HMbLHY8fs0b9JaurBEbSfDmms9DvjIwlf2afLe9bllA0BsjQh0e7qxMoFkn3zRly+FD5sEwu
lolsAdIanvB8XzlqRXMNP3ZZzuhOxUVTuoGUtfutAxU0RSoDFgSAIRNwaWkp9mYohfgEzABkyUwP
AnXx/Mco71bi4Oy2pz12Bit+mJJal40ygmqxvUEAK0HfpB2gCaAh3POqpgLCWFmYMQu8SbUDSV4X
4t0DprrM+1HWzglJh+LhsmjvpnSbHx/OVNhW+clfxHPWDcgMZrxaPuFhP4asgFq6vpsUB0Vpdi5R
OTKM6hpJl58RVroy4F/5EIaAo9UsDNfGD3mEJrb0albBIK6lX0Gd4YYIH+WzunoZ1ZMjPnWyR5yU
LnTekIYjfB9Vb0z9xxaj/0tAjk+gz89dakptTjJawQcRW5FOGifT0XLA6iSMxbHxg9oIRa8PXXR5
7zcYAsYc/O+rPNbmfNqdtMTS1RCdFH/TanJgKxlUBavPKHFd8Cxu2jqFrunfnyKK8VE+wCFW8f8Y
Bkl7LaK5Hhf5Sy2LHRtuowlR+2tU8rKMcfwO7tb3u8AgVgch31iPqJtKtUDIrIj7rtE8W8oOVzLM
6tj+q/VRRoIYfGh7iBVSyDI1MOLXyLvfa/YcYMrIf47cKnqNCaUBj6DrZslMERKQyzHPaEt7fEVO
XuSv6bnafnBvT2AFv+0sPt/EkqdeQI4RIotTIVCFmRj7kOYnJGs4yC7jaFVCT67DpihJzMhD3vCL
JSoectpPOCsJkU3V9pZPoFAzniAapL1f9bDrZbd7RHFxTv479hXHKlb6/3hdpxn2d8QbMsa6nAqm
MPNeDLWxgyZcAKg6Dwgg8pYpHrQQT/K0JISXT1xiUHN6gppJp6cdnMgA+tfnUyJJeluUw0joXk54
e87yL19mU0SVoY4MEWVSsQ6hbF+lRDD9fv8Gi2GWg+0psoKMhAbEO9qza1JqgMzU6qGJyCnZaT7c
PD70xAkZ9C2KJ6mVEMk4CyQypeL/K/UhFgbuP0KKTfvp4dnIafF0lC6ajIM1XtUCN33k93eSSZLy
Lq6jFI8uHzJ4IcqlJ4R2DnqtZa9EJCOoCCMlKFKEDOWdPsFAJ6KDARzYZFtdkuHGknIzZ+cAAwhV
gF0nt7PS3O0cQWdZ1+1J4+P0LlNvGyGDYlgSav94mBLDnGXbj5o7FlfW7HQBm7j9TZgp36mRuBkp
3/rUb5ZkDzmKC+ujMZph4vsAXXjhfF6ooKpyE/xXs7nTHaRIdRWdIp4nYE3V25YDTGSN0bGeLIYy
8hRUWoEEpQvwpIRxv4EZVsY9aV/UajbiYtt8urbuU42UKHj5nA7m5dZVk9QXYoYRzwU6l/KmJ/xJ
9YfpxQSul3BKikPHBxBCrJKupBZ0mQin14uFg0Nva78LUhK4X0v9IhyRVWLNYuBDyUscxul9PM2p
3IQVm5YvWRb1bkoRqwP9swu2OHuRXhLtGPQXVknXiC324Y1YlnuhfcaFQSMaxtdYfBSZV1JLPJga
Hzv4nV8T7S0AMiyZSbRRZaRJk4Pc3a9NMRjOTYdQWTSmsZ5uuxnSUdTARlXyu21jf7bP1uJPFNmD
7cyGae8zQamqlQ3Jl70qCmtE0Ovs6Vttvqhl89eyfRrm9bMukZs14jHCWl/S3MuBH7IU6dufC0Cu
794WCfkXYhG7fNbYfMhpexIIq+5uJ3Hhk4elwmKQWSXT9WxWnN+0eMxjwOV7USRb7Bcww2HNiwO9
tiJG1t+9lPOGoRkxzVyJfSxefSAL0VeajraebN8yTB8J0DnaRKaOL7awf4EvvnjlcGL3fsQCr/bV
MTVa0byrZq+yyFf9DMsBMXm/zbJ9XV+SI4kcO/fgsZJmpuqp5WHU8JqJUj18yW2XgrNgmfajrZmW
AF0mTSFs4owXQ/nsO/Ob5r+sL0u4DypGgmvyb6WCBo3DJo743Tnu4Aqa5fvTiqSXeLn8mr3MfYYi
iHoCGHdptlpBKIkN39pqRXnIC/bUe+dKJWZAWJpjj7Ha5Uo4Zts1OqSLvQ34iUw/QRUljkhshJQu
W8ob1Qc+Ec0lDehSlErEF3s/MofYzoyZCRz6fnjvPFDRZViNOfSof4/gdM3jDkMkdRUu5GDK4yZT
NDNazn7oXB6tmp6xask/e2/v/Rlm2XA0d4gPrwlHHfu+TU2pwVE6TpfOZXuZ6ck7CbKANwouF/5q
p93HKTjDldYnjWZj+9gQeqE4aa4LLSIillqAf49Uvp9ygd1E1bXWmptW/AzVYmssnXkHztoVEP+J
F3mzvrAVxDPiPGiiPn6WAX9Dw8SAKx1dhohOdYpp5PjfP4XBDnAwYU1m30sR7KCmoaF7Uzt9ox1Q
1LcfO3oqvFWUAhz7/gNrGkcXXOWp053ExA6bTBysWyfVTjJc0Nyc3tl6tMbTKi6+gEi43kWv6jwx
NYbEIJkz09e49Y/5FAfX9Jx3SGOXW7VZf1cGiI8dzMBvOxHqCyhGbDyS4kJfpWWeo4P63cJW4A/t
01oMPu8gwSz2FYc6yNG+6OPkzhp45vRJH0YGe3K7I7bMRpe//GG6IJ0ovtBIvnN4IBot/KMtLOgX
/3tZkxGXm8pQqFkRWq7gmiIIVqesMN+Qyr0Mi9h+27ShV2Tfvju/hjoxNKERIgqAFEqyD+OIuaY/
6518/8LRFJ06cPf/dEwBwnixwi7PFSxkV9Y8UvfaEDNuu+WbCpZR7+yrFNQb2zp/W0wcIqKcTKr6
L+OQiWdxoCbZDKUKzW+ZSpE+Ihv2lQRQ0twvXy1iyLVJG2TX8cLlHfZLVXrHRym2vha2Yw0RuMeu
9ahFoTX8bx2jRFghRTy41ub0x04vzw9YWkvheyZFUcoHLYRznB6F89t4z9aFhQXuI4abtNvdg1Tu
m6Emw4MhaRedoX+P9Jos34vPaiTuxK+CdS6qAmrMFGriGjGdV88QCgPDT5bvuB4zuBLyJzM8L3FY
ZVApzmplQ0kirAgp0u6z/uJSHj54fFC9Kxc/W9rZEQ+yHOqvG6J9DNLbIR3/ljaeCbN4BqRQwjQN
v56SE4SZJzq1825iyLMTnPCsr8OiUhh+mYdi8ZSf9JuMxH+lfQz2jKhv/fmpkBEIjtwaL7cKQEyi
EEIv1sO4BaHgTG8IkAceio6tIF+TKMp3vipEww+32jF0Mt/5vH9tdTst+35EQ/Vrbr8vAS+v0zut
BOmrqqrEPhfEuY5gzMmSCGPQMxL562i3w8tvxhAOU56DcpPxmUidNBDKR+N96X6Mt2kZceTsQaWe
jPpRzLzbXAY3g6qD43RjskBOzqf0mGc//VRhguTXA/kYKS34lfNBUz3RPPNMPG++uiBlqi1mEWfc
BqObW2pdxCw/cYS/AzzzHgNjeA5u3I5RwLIJKedcX9tK++cyrtrhQMqG078Vv0NTOJGOpxpcWAgu
WhgpsojWIbL9sooh1Hwe+AdvFKQoWku93dZxb6Mkqngp6qyML3lE19s+WixZJ2oMJppmmHyBH9vs
DWXOa8CE5olTVxcqFCTC0AJdkqCLiV9wDiVMkJkdTdZCZ+A/NT7kZO8qAABZ+M0Uvlzu9iECJu7k
CX4eRaO0yjB4Vy1A9119j/CpyB33Um0UyKgkKwEWhe9Qcq7baUTgxcnMNZi0yD0WUXxbDmImSXTn
qXKS6l0M2VqG7bTcTBqCy3CXZJB4s8MVo4bmADBirxPrN1QBa3oH3Ig3IGzQWIFEM84geXQafQJ1
53XJEIOQvL+iZhazgnVCCCV15wC9Cw/nO9+Sb2zVDBSSe998YmFYvyFSmrxbaCbN5uNtZ9MHdnFD
ZY0zeBRuLPSI20hd1+oGIB5qeBAweQo5s3lmudRGg3tw8Sqj4bXziCrzL2xPJJF75PFDxZaTc4Oj
XoXWrn99bfI75AOPvV9iDyFAa1mrD7E4CbjFZxiomVRTgcJ90ZXeKXdJ7vbyvz4rN/pe6b1xw8X0
MVh6yu0c+shtC3cmf/IqPoNRe8mNs6OnTc3x7ZMGfYAnBt/MtT9nNtxP7sEtvA9W4Pq+iRbpugxV
cTkOCYpitGqoAP+kLeY+DEWmfXFYuNB+lZidGdcIdBOwqCjdpgx5zzqIpBHI19xONum2bkbi9gt/
OpjldykN+WSZyhuOcGR4JoxJ8O/bmfFW2p4w5B2j/GgFHqv312dY2PKWSw3nvEYx397wFZJ6/RXI
GAADVVP14bymowa/cavR8+A795hAJ51m4ZVwpPhrVBfKltwwNtCjG1hDWFWP+A5ierwX8n26O854
7p1CMVUhkBqHVkL0u/8iNSkBEz0Z1IPRw+zUjxUo7AoqwY898fzZafW2MMyg0jE+wKmFtdCzTaHc
6JubGxF5bVlkrUYIh55yrJJMguMcv8p5udw/GW2woJ6fvHjDimarFEGyMCpB5xiqXpqkxVNAFCHE
/E/R7qw4vXDJhcv6vIUl3Z7YZzaGLOPWAdmzsxbfe2JgY0LlHn7Ez4JvlkcEgRZ8VLpOJKJFMhuP
0kpvxrAJt35PrftDfRhbc/0KCujQ9AlrMPiYe727FGKHU3YTd24jypRi5L3OS8a3ANZjwadfm3RQ
V6xj2ZykI77iu4NwwYjnpmxI4Jjibn/cwDzlrfPV9AZEbklVP2aOFbBNqozVS87OH4IXZyeNTnkf
x2pQNPcPeJz1gXtrELm24w+woVKyiWqSDY5+RaD6GaCk9Oi9ZLYBEd7fqqnqaOUQT5gcNWr8IX6I
ftFlU8wbcJEnCMUX30E8KfhNYRV5Eo3dTUomweMxD8g4ce6SCo4qyerz5nluYxiBgACM8bKUjQui
RMxlnZXrvx4C/AUZONmz103vC1QW/WPFNjny6sAtFE+UxFA3E392dWA2CuenEdV71fUEy7Fyfb0u
C9oVIzgeHWJc9EGdJklKbUDdh5GBc1IEr4EGS7lSh5QcNjBvP573p/pGR0f5U7vAalZHRRgPpr1N
TwNOH2ijQX8pwTuyAoNVb0z4H3LxziQVZJfmDhTn42jz5int5v2qWN5g3FmQxnvINdi0CfgcsFfn
NyLvzjDi7SoT7ScdkMc7mYzpx6l+LGZURSW1AaUQ6CB+iuJUxg6yPsqV6Oq2bbev13BvCyr24P06
It5Y/4wihmPJs3+lHHASyphsPkJUBWt6gn+fiM9JgpQ2+6HQ7S4IlVrhKyHkxBQsk3p53TOjkGeN
YN8IpWZoKAi0o2eJd3lmFUU9znjlj90j47x28r6Ipk68N2k7G7LphZuFfQfcQh81zv2kqDPIJL1Z
b1TRrOYUXs8g4VpMdef58ms7wcY+96/vB9PjXidX+aAEBWeuZ9hMDEk/P9yrnbe9oDDQs5hOEOdQ
LTDvwTQVGmGc+o0H3SisaCkNXF8tGLztVZ4nBoqCUK8q68JHwQWNDt4LmZdHYLvNru9Cy+Rxwbc8
YYjzldy9SCUEThV1hAM72TZLaZX0QyTb+CBSaZyn8zmrMfx7sfczLgn8KwKgZ0Je1u04r718GtI1
0oiRroocpWXZ1BF8CpkCoRP8EJGy66zhslAFwEuVJLJpnoroAaKnerjPMG5jn9SSu8Ag7Nd9noCG
M39VAADJ4J7KzcNMOmqZICqWcHzkD/B0OAygFAaT/ND2PjC71upZTvD3cdiuS7seLzhBQVVxxw2u
zpAcjgSiAASeCmy/on83UwtBu4J+fON/dyy9d9uEA9wZ2vQRtxYyHwWf/wo3B3YvJHryrAkhk1QO
mRqaRHTmmMGe8CrNVM62p5NAVKPILVHQooYmlJJLAgSHkIVHfBgsURniGmLv6A4nBW9vgSNrnuTN
siXYG6A2epyTjKYvxoyWyPc7djMPDhmSn94QGj80i20ulZug9bT32ioFGDka2WYGV5r86viT1evD
esbfkdIeroIdsxpcXL0Xu1oGuNJGut3y35hX0qW9ttUyLoa8i7pHzmqJmt6QjJkpfsVYwDuebbVj
qN5zYBfF/wzEcedCLJ05Vfv2DCGcSbGCTY+NDcGWM/oc48oOuPOcYvD1N0kfS2TpFhDTZd9OUPlV
Oke80GQMRK8rWju32RFY+UG7BHPmt87kv00vPY2DMPMzxzWhlJKoQF9xln0vfZR5GDsl+CHyOpuq
YocYnRfKqhtmlPkszz/6Jl9DPdIlDRG/lzWNya5XIjDZUFGz3xsNed3qjCDasRp7sI9CFVPnnN2u
f12yMiSrSXZ26uDOG1dQ2npeKLtek55WoOtyq35+SXBek2/KRHYv5PgpQi9fH5ZbW+abQS+8Wei0
H9kuf4JSzlD/DEPIRUXFQsoZAU8kmPX6qQHghm979AvHMG7/uPd/f4NoGWWSy2pXb8GFmy4eQNbV
UqdexU1Nev5xnJ0BrBUoaEElqyvz5crR3O+xvsNf+vP1lyBwp0zABqTgMbmkHQZW8g0+4z9lQt5p
T6cLQ3/caauQ0//MbcWBWGWJ3eccrX2EL8tH5ozqsvcZanMPAK8B71ndbggtE9Mtb3Y23tLMzbf+
qmKi/dyHFCNZGjqetNdaESC5sdyb2e5Yy/B3urk1jvf006l9wdRPksD4yhyJRtIY1j6ew9sFbta3
597QvcojQCqdRJ5tBvBwsgBsy23/y3xGcYuFtbb0xUpw2ugwXw6IOXeYlZL9PxxWuzgy8OsF3uxM
GgJL2Qv6zhpMMZLimMjZXkocxsqxGrtlap/9w10RQLbLY2PRt8W7n49eP91krNW63UKxo7iveETk
RvKQnlLBqELvTTiGlo5a1nYmiasTwkyDnX7nAp8ONfBsqvB7DiCMArEb6e0aKtlGQhF8oKmbQpdw
7rCtx1edJm6odViQD6olYrmYpQKb3bq/8yvrFmsLmKFLeEWXYEDgf0+0xZteBScpjDKa0huY+gEq
jZrQcaB4nBBR2VSaCcCal5PP9GEg7lt02MH1yHLB28ixOJ2YnCTH3mUOkDuzdFAUE9DpyQD7QpTT
MIPmC/7HX/ogD75Xr/RNw2d2aRJzDT27O/blgoTAPvNtqjM/uG2pbsIrwytfCAl6kSdXFymjYtqo
oB+kidrvj+92ATmEJarhzA+K0c7m43z8rkC3bsIKGZdXFVJE0inBeFCrIGgahYg6KrZzH+0P7Kuq
WjdPV2fsvPyNcKnX+K1pMMDWdss0dkQVr2LHUWyvxFroqzB1Niy+qvdHUo8SBo/eA/2Gku5BwY16
qtXDdfmwnqBQ5mjPi771bN79TK3GWbBGvWlSpxAMjL00EXMkRondT5miw+oBTftBHbMc12zzxlJU
7SDr7xz9e6YjsFqTMqafoXJlqx/KYPu6H8OTp6AnnPyswyD2YTiW3R070u0OIwW2lBVFLcN7joc/
gkwnmhlNFo1M1RwWcDxok5jqZYAx9KkxLG/dMaKjzL4kSSPeB/zMpzRg+PJcXM8VpkR2jQagm+bp
8eTH0YpXcwHwTajxDCXhHN+d2WnkhE6Bv3bXOA1eqbD2fTttxphX4XhxwaQKAwcVi2FYN2U0zU2i
UZdsUMFolRXjhWUgY0ETBBcI3fMyL/LEOxa6Pm2+oUMhywP50i6oHhBGH9/UVXUyYvxU5r11J9lq
WPhYCEq5NUz+mPrh/9TywyDpPAm3JD49iEQ1dYwDYiBjyqx6nIPr+MZ0EbZkytG2XQrodKBHkZ2b
lOoVAjGrCwN4HCpdKui2q1cUeioSV/eEDDZa1juFvo3u1Gopqm+4s1/rWDoIekYranMmU2BPKEbe
ctcVz3GEyGl4bKY32YSxOLd29dfA0ToVURYXiZFitMbshGuxp8FY7FBtr9ywYRvlmh9txErRzYnD
Iy+I5Vlv/5TJvT8CzC3gTEwir9qZvudPfKfkgw+F/euKJYgWSEKCV+fPL+XIf/zP90EPoSevwCRH
pqYs+GqkaVkYiIIz2gI5aCcQAsWk0CnaydPpgTTIZDWwB/Mm0fUTwjE1D2Z9fESrQz3RI61sEscv
YrZOdhiHHquuyYYuhEOW/CygeDA+iOu6HOms23qc7c/vZkXIERsODeJZKpye+NDzXC7pc84crg8f
uy31yuiaWneEbqgevcOBRuclChiQ6o9yjbca5ZNqeEmmxaHLeVFJfWpoN5k1UMxXEz7oc7fVLOl9
HCkdgDeok8c/2MShyzfcV7nIDO8339f0HUqLGGvwKkmWcIU5TFFRWbMlBf/ti0Lu0xhO1gc5fGnN
JNwif9Ui9YI2NrCC3UH+SLD1ao54Amu054Z/eEvM+cfkakbozmC+/93Mz+2AyxKNsU5rCN4vNPxs
350yB2gNS6Sl7b/DQuUVi8LdxUwjIJQSg7v+JRLNm/XBrjpGpfbhFzMzdKpQMV8jVcqt3MpKe1Ax
Vq90tvIFFxXtdu7jIZP1pMC3ohcbO4aIHeMDaRjS11+pThZKq9rf4YZk+1trq9s2Mqi42NNXgoB1
AeCs0Qmgtpu7r1uIX2bPqi6+t0C6I8/2m7gEQCHFZV941riUaOXGQkcRX3unZ3CqFqguVE3QlGEg
Mv8MFbrcgOZ4Lndr4b0tHKMrv8eboQ3nPrF6/EjLTTL6tQrwDKhuP+ltKF5liFxsUtG2DNFUYvW/
P7D7Y6WLymFtCyaCwoF1W0nJwAfVICrIOQQBYEOoYsozFKl3SqgVRFJ50wQm52eKxWVcVgZm9Iu9
PQettLYcn8AWwEyJDi0OUo0cfffAbsLQaw4aGFWeMICzXWuKeuZp8OLuldzLGpTu11EoecKTLpCV
l+1U7zG74d5xsj/0UuUOSBccA+BY/TjS1PgrMFiGYNtkOvgPGVw5/TarTho+tVMCbecAcPjqJM9q
QGpWipqiGLg+tB8JBQmLnVL+HfwliO/uvdrBBwtxlzXNcxr6BEmjAxLHOxrMgPDxXMiiPQwspPFl
6Dy7BDZqT3p/lgqhehS7rlj00412+AYq/tOXpWHQTcxHzApzVx8BDocWTUBgdPhdwh6HaDalOYiY
QYxOBsqgI0BsbE7NoeW1xNDMAOozZouAUz99Rs7YF4WpMSC4T7ZUjFBCqNOGt4Mo8wEBCz+BsRVW
0h/KZdNHR2WwvA1bF8PnzExIiRPYAp2LD7mmbLa+flGXDnIzOKyVA7Uon1U5gvNVQve6sKsrgR6c
sNQLWaooNx6LmnBlAmU2RfUwRAv1S6ZvSlrimDAevckUCEutqxBAV8S3cmKYpHGEcvI7gicLFaWT
8yy8FG3hzitxOT7PKkbAERFEPjIdQLB+IUGQupA2c6lz1B6OpnM+Q3IMV/z2boAcGt7IPT7par79
csmOmRKixpU2Mbb0uE0QD/BbHQ/2DX7Idp8YU1aLXXl0y65lhuI+Oui6budZJx0MsNgSNcOM+bgA
tyVuqpq4Lv75E6+i3h8Rf6IXdDL3M+O0Tmgy0WhBp86U3ybQFvCm7Fcz2khrHvNBSYEM/zMZ+DyQ
o84rsEIwc2wOmsRT8Mc2xeo7u0DavcuxR5+hwyh1XhQG77dHCyee+TzftgHxRZQVGESMpRaSbVx/
orSV3YXYxQQM4zOO7OLOqKU2pmn/PYudZcWAAK5rnGdhhEgcPmvOsAS6SjTGxRIsLmdX5mvP9gmu
IDrU7IEDK0BQITwMeTANW+fpF0mBZoR4envlJ5QFKFFRwuCDeYzKOZCqF5qTA/qJPYq1AlRnlkNM
8PaS2h+sVmuKWYHSUU9P9xsCqF/1kteApfYrvvYzXZNr0TwLN+rfI9vpKiHP9LoYfmQbGMKeEp/C
RO49xGPWk3AWP1D1Snt07aqqDkutG0aJo2JDu8FolxdGl13yZ4BiK3KukeDWJGiT6a78sqV9kM6c
MTQu4rOivrTRwuxXRyguMsTTY7USYIn0TAXhJSI/U1FxBrFF6ymnKzXUIyyoquWG2nvPVGxc7kfk
X91TxlupEHQXCadmCXZOSoZ5WJ0l/bmvVMboP8Kxr0KsYOn0ejAO6xHqfjQnZm2ZRGJZbM6yPr1u
FsLQg+cvljpzeaCokg4mSieWj+aDLolQQetFbEWmrdHoV8keIa4SlUd1wMWYrpfl3pPzhXCmw2dC
AAvU7bGRj0zvsuqj6pvlaMLObeP2yQ0q1OmaVsirneGHbt6UfeWTYaEHeaarn9yVDmp0Ss/JGeK+
+RG9xbbvptlTyWE96B9V6juW4IwgRjSUEvvbSA8x9EFwR7dmKaC+nN1YB9Rnb5Tfv2jFyAXrnmwl
8mrVLrY6H+DByi5s98/O7F0W0S33atw6kHAiMtnwcCBEEe4eqSKxlDNdigLNRbpYSCHOjP5dojv+
83zJs0rSoZWIT6HtSUeTJR4nCeCxW6GjfdRNKiyflaQOL+3bTzOLr7Te7E7p5pqTsQE9pLtF6gbK
Vp0rhXxF+3QXwJXdW/2jikWG+ojA/IMGzwcsF2TFvZnpu+GwFZboxigzmSuJcOLKtwTAUjX4a2V+
Tvcs0P7+sdl1wrr075mk0KiDmsxAEobduErSodb/OBAYC7CtdppjqxLcStX1CwHPJ8bhFQh1umJB
kqgpMEdUDHSRx0MBATZDvkkXjL2HgtZqkpcqPjK/+a33ZB/CYZdy1fBuG/SuTY/cz69okiBCdjdM
8+x27i3spKXO9rxiiX3hG5ptBgBm/i2sjysxxBRIgBa0v0K9Xc+dPm758YQqxIuwWU6oyssQNxz5
3dOntUgSjfsjUGcFDPfm/WXXZQND4VLIHkTfEewWfB3brPQUi0n0wzQERnyMVMB3mbW+cJCTH43C
JgGGAnUmizx3LLQZiBrTlXMvQLpqUEzDqTnxhvX4E0pQ5uFC3YH1Jh2psLQJE3C9HoEub3iJqHYW
bbds9mpxseFcOdJrKtx5UMne2AS+An0MJqLf2BGPCUvdVoggXKygnpYg2/c0WCdP0VwnnQ5vYzOT
U3565kUs5dBgI3qNmowx1JfZtGIOhgeEtg1qmW8/unkK/XIXb3ltGL3CxEOacNrBvdcP5XVXsAYG
t20lPWccJocmjPEPImviQs2pSW74Nfu7Wcklz789TmFfO5Pq+UfmPrC+8PhlzOxvlsLq+ursZKxS
rUmYFl7LwXBWqzKOtMbrLtSURU9ZmRkGl2a2xa/8OpPQbVXll++H/Y21qhh8HyRPZ+lELnJbXIuJ
3ywjjMXMEEf60fNOxQSm6+U8tDmUI+tS2wEKLpaH0vYW4hKIPvsBM9LS5GYqL20XKRg3OGbLjS7x
z5TIpb3zEundr+R0viewj/Zm+Z9CbNowZWNn/phYEDKTxvZs1u/DO14AbMnAtw4Y1dqDIzb9cO07
klfKYFi2fx3jsV3nNsddJORskdvUBy6sIGrke3HRb+q8ujlOtnnke94JFAtUz/zTPrUY09uqEgsv
sAmi7XwUw8D/9W30grJThN5dHMtMQD3iohaytuxszssOMOpdX4dX2hB8N8MOtFO/5S2FP92+WYeQ
NcSvp96L3LQl7pQcHdOsMUdfNblf3dRNfoepJltZW9DFgznrJGTuGkbxrwDHesd95Io3lkCupHCr
7LIQ16sClxMTI00TwuxZTh+E42iGAiVkx0jN9vOJWHvzA5Vg4vBT3RqVG+EE4p1q9NwFncawrULA
1H0VSCQU69/TH9R05ZR+DYjDuOmSbSmFmVQ25cG0EhIf9YmB/bHxRq235MnmJE0JTkuolu3Wot2f
Vbmkw2nwyN4XgXkdlcz68cmYJp4d4S70PELl0z/UzgXZdiAv1m2GM/i9B2ACTLm/+uj+FGe1alY8
GuFeMvWBUxxDMSJV7RLWqOogCI6vtzHN4rfGlElZ67aIGxM3vRhTPqELOPU68P2mWMOPskJpbd4o
DNQx9VL4ioRKXwryrQ+DV+J32zW1FxYJt9wWXwfUHgW2XAgkFp4JmZsWDVbsyNfFMxXd38OasxS5
ol7SEUOrvKITKkXLoobdY5VgKNJzTh17KUnRyzC4/YaPvLuHgWOqQ3dWhxR/Ub3HhTVHPIdKmlvb
edpKFXt/vwQ9XRpH9otbrXlfI3JCjFcfbSGy5MFTk1XwbUhCymWjOLk3lkZ+NgRYBpsRLdk9Vl6m
uLfThHs+V3IUwppdYtde2uHjHmUxJxKtxtHeL78Aqugw6BYvYDb7GY20CC1mpp7oJ7P414lZRKxZ
R/YMZpLQixxharMFhaPCHxf1qxPH0dcG9XhyvBAVvwfC41ytf5TCMBGIima4fWXLePWAAOecIZrT
N+gUx8bL7VwDmwm+rq//KkDuE9z9KeH55VTvcH5v+nPu/qYZs6AfSxDg1lp8ytCnk0AT9ZtCbToJ
f36oA1Jn3FN0lPr8znKAyqmRUSq9yfSj1hHsObDYI4qYz9UNhGz5uNVENWQwNYbV6RfpgOFrpER8
XdUdIBVIL7/HTdFpMY+gze8f5whmgNMZSVgLGKMShk1U9whovb/q3KTW/nHMpbOufFuNzq3vVJNT
jITIfxHeghmTzHlmYkYMk46blZ7x1NEQFvOwSCcQEzIv/reIhik0r1fj8+1R7xsQX7BfOeEmLZZG
biM9ROVf72MX+tbrIM4cTeGILTjvq5UlcLYAgPgq7OV4CaIHCld0DKPSMwjWJYjWTSoCtr/vC/Rq
DeK5A5ip4z/KrTeZhFrcp3YAIGsahD9h9dEul47z36eQTJ1Wwr+R5NZJ4ykgGBs1/1uX2YlhMnmh
eTX2k4VA1FicGuZcpVP7lNqoI4KS2KdencIgvjwoLOa6KfRgIY05R0I2QOE//4BMismEduvnfako
T9xEeqUxu6InY5iMLKx9Be4a5qGY9zTfAMpDfATVj089daRJ2EjSMRSW8iywrMa6qFc/VPuLdWm2
qCgNMCq1J0gEb+qAMSSCbuhaDAWeBDyMzUaOzGhFaorSsh72AZaCwgZjbQ+sZxKr9VawkGeV3fVv
x8KJ5SsBYbfv0mO9WrQ/cZrhNNOzpOcsXSnEhQ7WptE20NJ1O7Lnp9GZL53nKthGch/Su+8ccT/2
lNvWHXSIYkHGyYHmkMHIz7huABRtdD+1346AFgSdNQBmQGGCnTdIIrbGuiN0wkN8XjpU/zG3+E6h
HmG642Kh8hBpBiMiezmA9RcDim2IcLtwR8paYbdXKRqX/E/XY4AVzOGCbKgSJ9VnM1wSEee2f1nu
Rt4faayAMeX1vnQNYXitVANnSusTZu0YQMlumrhlQo30uEhH72zmGp5oN6e/8mf4lVf/FhAxM5gn
nnAHIcSjiS5GL43gfo8qPAmpteWWQuOkhX8gpeiUghx6SKQgqeO8UWLRkh3sHDGL2Y6Z3csCUiKz
YqABpy0NyW34XiPwBswsmPmmRoBDLP2IFSa/VPiwLf4eKW46jdnsFpyDSTZa6Xo8ROtbdA+MNDeu
a7LtqOmeZ5IWY9Wi3lLQv29f/HlNl7375cDUb6QDXP3UQvkQJRoUmfN0+X5sbpaUMA0SKwMk9/F0
DxNqpd6SAqrbIlxfJHL4+mhHRYCZRi8chqhDmRTJws644AkUXzeNrl/1MJYEuA+EIaBlHT5LBUii
myJYnAK4XAFwO4oOtxjC4nlQasbPRwYRqrBzKwXI4IU+aSRZ4UYfINAAqa9NUBzVHJ6luZthrAc+
Nw7a345kBxCpMrbiv11iM9DxweltIFK7aCcdmDSWXb+ppdtQSojjZdq/ORrRuTk0/BSOqd4t8iBK
P0W/BZpOd0wWM3sI8lxC/O8SVIRzQxM+aTm5WRsTjV140egjDOwQ4mGyUEhaTlF2CINE2aDnazyv
c4j/SN+q36XQopoNBZ6lUj8jxzhBEIQbCcgrXpm2Fx8tyj4KgW6NmTHQle4j3Xd3aLG9DZulRo6o
kPyT8ql/Cll+6moHyy3gQxZ3c/jSVVURMxgtE633TaawwXt247w0yPrw+Ay70RiNzt6G1U/9eYVV
zQ7ppezcZFIbMCKpEaLcq6//tVsKa/WOXtUBoJQMJ9V2dWLeN6xTLvuWgO8LwfbMTaOeMNB7N3b1
7EeHESNLey1pJP7LI7ee3i4DZAsqq6+uszOMgU4O9ENDAwOVSvuvMByXjDIG8+87XKvg2D4J5ZYL
9LJv1u7dQduCDFWwIM0ouOwkA65VQlmV6hxH1NojgCaD8FzZWZbtZ9JWBeA5Y94Qnq4vo6BBkHZo
C4FVkZKu6jKDEDrZWcyt3gt0qKewW2UcoEsq1feDAZCIiG3E7ITxXn22oGlaVZgO8BrQ/IZEG586
38FLcydCTrUG65ZmsJ0kDbgLNz9tEj1tU6ZlK5F5em1FQO3NBR4snfXlfSOc8HAssHvlq0PEh8hf
54oO0OqGsPnAOjhGbgJREIWwFqpcqaCrWjT49/Oj5a/TKv5s45a0T/MtqvHhP9d/U/2S6z3GQbn4
pCZPYWB+bnYCiEZFA24CEZILqRPqxDegQYXaBPVFgI21S6oJMr5+IkSU8jq9UygTpgmOgbyzOx0K
NZUhKys/DBf64MR6yVGcg4zlIowLTgEBtvL0+vDZH3zeVL67hhMuYckSeXQRnphXmMgXlFDc6E7H
PMOVmhggI5Md8iOwDw2ySJbCJ4wlz6Rir3OF+Wm8MguGPevjvB5e+hRTF17j5aWAN9Y/Iqpofwu/
pekCVCpWfTZRwxK3LaRW/KuqS34pk0Nh1QopB7FtNq2GqmDNo4T/d5H4OrcHVo3AmYce9+I+Mj7B
KWwMCXgyt7VGqTnikA9nSh+XWFTD7At6lgJQIrG/2Y10vBEBp2XSs8kHbaoFkj4s485meEMbwMx+
aF7ewBYQGFyC/kMipTEj7U1VI765pavVeRwuQDJI72aM6Ci9IP4G2h75sorCTsc5rtSH0tlblD2s
cHyY/rSKyH87QVpj+ea0qxDl5G4mCdq2Ts5eZ6bOPqgTnnqeH/sLAC4FxCejGjWhrQHmd/PAWCqq
HPEG/gxLqPkVWVc5x7fUcYg4KSwnyVEEY7S9I6uwnp0waDGp0Jy284LMRbWBG3N5DTrKIRMksJ7T
saC8/LM0AReO/rWqdEc1K/WPX/E7izipy0q83BbOk/E4ZgWOWuNQ+GJWamxwBJZQYhty1uiBhFey
dDNUs9XHHIPlUp3ByLkiS240xUN7w0NtnXAcmElJTno69FWf5P7QR4PURLwcbR+fxlKZbJl0Q9M0
QllvIKgOitz7EL8JN+hUl8tLVeu98W+OUnu/bn2HnZyQxemgnOEwIAEAPOFFYWLDyqfWC/p8xD4e
/+q/fAvcqoAQmfO7axKKJTYLbnx0yV0kCwItDltJKJhG7krS23l/0cMN4mFQPykBb9yhDb4YQdFb
HoT4H4PeGEnQVxoEka8I/OnimADVJRlQ3Xsqyxk7k8Ke7cLkWcGro3jV/3cfAlR5sSWglmdLV/QK
THfdbggYV3IFRX2i48MhJ5hVpa/lu3ROsQOW8lnZsCTnaXcPsKX/Y9GLVEH8yHBCFHHoUosGuTVV
98Nib9vS356N+09g6N3Aik6IVZexArWZQQm+r02dhmRvHYP0wA0bPH3QaF24+o/FG9Sm9FNaZtwc
iVCDchQrcMvaVoUcbcjxTSPxGApTzn8cnPMDSb17vkGbtGS4Kn84vGJFoOfs90BINm+n7XbcZHT1
jo/iKIZByqQH0dW+jgKP7jA9Za27JIgIGlztiyIN5TnQfORsMv2qXh2NaLJIv5xd7NRDe5ra9V2H
PEm/b7eD+Otv/3IOEKtMo6e8kIRoSuNeqXO+9W+LW7EV5KSpTpXwL7XZCUc294ffTyJBWSFnjqAT
7Uq2RFVYrDyD6/A13GE9uOaBjJi1VzT4suhQ9rSXwhPSxqdWM7Q5b5gXL9auPduFlmVj2INAXdlF
ZyREK4vTi//GrGJeLBMeaiaj+I5NhVFQXD55wl53pi13GpW5AWNlsyAKPpPE5bZ5+zYscO2QR2K5
TIS8KjJLn03XeR72sl+Ak03ZefMUqLTtEy/V9P1fXR6yjixOqkPhs0zBNW/lrDAQDZtves2NyQ6A
FATBLix9gFaxniENwKIcR3b4q0DXxpM+H0smreaIwK7ym4VVavKa2td1NwVW7fjvJdCwUhXQYscb
ILrKAPec60UOxnSVMebGgZqh6tA31kwD7NJwFJ/ikXqu3WgS5N0962FrITA1kJ3rz429pYVbDN0q
CAkSh8fN79lHTfA1yPk1dH273CXOHnU+r3hhNIxNu58nVclX7PQ+E666HghCjwyi7IDRAfG5fL37
wsR0k5GWqLMVfxrnOlfOzQzAhUQaiOxGHnpp5rE0DBdmKucDO214Q6SyjF0flf2bdZJvqUBQ5vq2
TVYIDaGaSHYzFSVjIezb9tqj1A7RAYOzHwYxtr8eMZlyi7pnGRJdoALBRv7TCWaHc9E6yvSzeeqQ
6VPrbMbtjLN9TeGEhDAK3wZuePQWPRbwiEMerSg43fr2sw2flSTWwdXImXOgx8usrnEuPs9RoVwO
X8r6kFyX7sa5SDSuefXBX8GLQ/AXrutpnxeMlXamUiwrqA4p/xZnlGNElTRWxH+UR67i4u0PSw7+
F+9psYxroEtHCVUWkJUBqZgFa+TQV3yC4Y7p+feVRakUHnYRQJFNc8fYEbs1iYAKZpMvojEAz89Y
vXHGAn0XrnQ2T6maoB/U4ymeM+iYIKoDQUJ31sSS4tq2w82O6hEuZsdR45EHgf7MF+lKX1ZBM5N2
mOhLOQ3rDkpiqXI8kRrR1NnXvn5TSsgbNsEFZ+cnIuX5A0Du8PNibG89rldvGVqNaamBhjjZRBgE
J/9veNuw1JuX2z92NXJB9WZW6ysti9lgo3hXDu4EFFVugEO/SWYAOehe3hQAmc3L+IZH1kZ4K7X7
y0yq8GhK6AkI0loIDmaoXL3KeJ4ZADixGCccDtcOQcqudNzu8hmvRQa84gCEAAIhU2BVWWaw5QKR
V1/m4r+yM+HDisJEHfw8H/ZjGEPTzMmIjvS4CZtpztTeXmIYXDSDY46XdrVrgXF/uMVp3B5xVBmY
sf93ilxpv5YPr0H7n0F9HUTWxYBYxmLd4lYPWTW0q1JdLKnPwhxv9oA0pRO5tXoHbCjlQmhileu7
n3syjplvx8v/E8j4/ByqG465kTV8Kuj4nJqRrJ0ZIUo+UVbdvpO9Byd7B+4xHn6XFmQWgzRMZCfV
PrCH/5AKk+CH8L57PDRkeI1HxwAWYLVrQsQNIxWY29XA/kBtjr3ByjH6D8XC4ZunFJ5VC0VlGPCR
7U6UpvIO2+97fp40KKQ1htDB6lGZHpB0syG3w3Ghu7uUBEBQwI/vDL06lVkGtDYvRPPfIvb7A36z
lOrvYBS7mhK82mVrdfEizlJClNyLZxXpAIPy9/UEXeaYJ3/X8XV8AbXoIjlUVLDUMXm+ZVS7HzoC
llMXr6AqD9ZlJhEpa4xxPapaeHIRRj8yH++HpM9MLfDywjBU5S00J5nM1RCqA/X7e3YDWOYRycv8
DxYacnTWtqD0VjbyNJBOs2ilMP5TD+ASb0iFCrC/iBzIK1BbI7l/gNEGdn+r7q/dHtdDpR2qs1Xh
FdIHULXGbK66kg8xxrucFdPJ0YvvQvfYWvsvQDPpMxh9eRk1DoQPu7bLQTsqvN7ztpe4ovOYqOMY
o8GY8wl64ky9gr1PxDYPtvgBCvgbc6aFuPMdP30zkTNs0USqOY40/6z8f7QjvrnhQD7uF6WafDlV
9YgFZAO1taQvrkvacN+EPOW0vR5HuM7tnXlWW+Mi6fc+Z6yKSaAaKAmOuKY9JDrrLslcbd/OpWqY
UDhz+RytNjup3N8f5tOQFOdVEYVx7n6iNj7LyCsk3bo9fnhbEcMFW+bRSHwFeo8MD4F0XT5nWmYf
QDo3YR/tKo1mrpm8XRYp/9W2v6Ww9A4qJISU30gTjPSAQ7fibGKFc0fE5EqW1TJb0Io+N3ITYGG/
uDcbQTcpPFtg6w0XjPY0LLhobvsF3DyI4N3hnidVlfFJ+gGmRbmW/khzPRcGLBZxDIF4UcV6VuHA
taZVxZRTxLJRQvDtRQeiYPQG4+SgAzswfjekkcDCRYR3uxJCN54VR7v1aw4tO/X0ef3FKNu6RkZW
0u2N+W9LKm01MOgJjLojF9C//d0j4AN3BqBqf8HY0sXTLY0Y2+2C7rSsXv1hKSeG0Ocagl27SxtA
8z2XkBvi8/ETCM5PAazs4waKKXQfoS17+9bzHDiPbQFS8oio4BkGYQC3cB5v8mCxzyi81BNeY8Kp
qxill03RGfAZILmrBiiGbQ4tUq3ECUZxfUADPDFac7HmWn9RLxCmJNWaeF3bExq5wzSOSNzuvoNH
JCkDfsaYCkP++pHRPBJNoCYpGl2xo4wMHaEjPLlWQUgeQlFTZZFTTcSHYg8wP9rEH/L4K8R9rtmf
DUONNC9zedhlwUp8ixk61/dUzvjPADNx5JlEhKT9Q5hKz3e6MBUp9Sq8b2KTl6w5vRAPJQKg6w9g
P2KkQ+J/0EvyUUmLalWy70TuEjLkQ0YxX3FBYo8PrCd3Jw6WHBWIs2Gn69WX40xrgxF8l2qTIxeR
MZNXp09Hdu0jKiVdXQl+SrAohAjh7NHMfSGj/ybX60/wAwIvqSIp93IL1+SBkv1q21xSW6o3bN2h
mAs5MFJkP/kru/SSbHEiA/hPzBkjlPme4GmjqN2FUdTrBPa4fOu7FrXWqPfQ2T18f0ccG61qAia1
SzTpV1xLmLLVBGssqA+HUcZ9JEloe9wnbtnNyaLrKafd1Zp3k/j/Mwvx4ELfhakg+ehJTDVTDS3q
Z7/HN1r6Wpm7iaOQg/BVLc+vEXrWoMgDSMhxoLDm5ky/fXNbEABE4b4HMALmWSXfMZZz0GLaOsAU
R6bQ0psZ4ykq7K/cWsSUhip2O2jGyTH+hkD7G3wvv6y28MzC+t7WnhC4iR4HvhdimMLWkk4gguWB
Ob8hjD5UfA5YXp2Ud+9htzm+W5GwkV6QVjbEM7E+Pk6pQ50FxuzhkAC1XRXb6ffdd91Foi86ondZ
qWrqk1owKPpe9EPNTkrpz/rjejCFSJkwx90CwGuZRAx3UH0TaYcpgrBGp1nMz+7GKFLLdaiHIOpm
qbvEEESxKtxTJkmYhd5VPz5boK9T+NLKk7bvzjGa/iOataA9uGRNUi6XK9BgLpkh2COHAMx7CXFJ
juhpXq8CgC6JAC46PDnokjFw+j7NMcO5PsscnExtOM6TNBuZal9FS9BZwvONcGJ/VlyEAD8jZPQi
FMQzwLKrqCIls0zSGWa7Ehw43UuzrMy+vueics8GnwZ6PVCZ6ArjJ/V66k2nG8xxsLmn1G7jgiRr
3hb92QxcQY1jIfTrFbLKEo+HBxOxyDtAeQHEUfMMKFOgCkrNQ8y5MOPF47w4Xzzek8WjPJaN2KMm
fkYZaVwevBE9arBkHA7Y6Hq2raRl3K2ol5xOpVZAZb0QxhRnDVcVEssjtHHpMtixS9T5x4ySoVbG
QjlsIZdLQEicUKxYcZ0J5XktvR63eWYpJLTFxILjGImVOYOI080B82uZGmywQvYEvAhyksWjZEth
nlc0Jgau/S6LEHRU+6lUGd4MWJyqesTuQyWgFqgmnLrFd6Jk1ry/z7cgErMap0gLzveSJTPhFYHC
emtNoR1/EwssyhuQXYeezg8OVr1SPJx9a2d5BaS7SYDPVakwzMcc7cfmHSg5d/9ax4KwMQhL1zJg
fPCLHgrkI+xlGhWqw4/OukFDaA0imbznYQRBogBYiBTuokDM1UzYu0MJQ0+xtvQzg3C+pRRd+Ln5
Ev4jsMOIraq/2TshE92MqDDTxDsouuLKuQRGGuT6XEvdCFx5K5RfGOiBEy6IoNAQJIvIHo4V9QXP
dvOI0qaMAOtOBO7ZyIscEkcb9VIUKLrX87MjZT3gC/DbHwW+DwlckQD3MImhtI7BXMfv3P5kknOO
7ue0755jqI32OGbOTrcGy2nyEke6DoA4Q0M8P8MK7gseB4P3AwyTRU0F5fU/EBTdS7FzxHTUsrgO
E5HJFNevpNh5UL6lbH40v+Kr0IgczOeyQswM1O7JXNXs87vzv2vOzq6S0ZNnm3pIbGmUBaOGa7zt
tf+KDccdn8hZNXezDwAGcAdihyN1rlhDG+wJIMFrisWFXCbMGW+805FqH7MAMUDBUk1DUBE0ZhQj
f0FCGgE3ds9iK7nEZIpJ8qsmriTM5bTga1FCvCmlB04hkg8ARmhJtLVa8cngjDO3LpTShudkm+b6
uzuKdDpUgQmaopg7Ipx/eOUhqy5H2gUL6Wf1Z1DvxGku3aBy3MGoBTFmLgycxPjWrPWLEW5EdSHd
njPX8G/6M4Z3jcGAIby/oFYRZvDOAaHHBenrTDgI8O4iMthTRg+inCyyQ6RWWr7TEKlDeWYKblpC
50qWIc4DRVAgEPF9TGg2GSleatKaTWAop7hHqh8zV4lOHOL9XEBW6Iv4AbMW2fK5ARPhBlPH+xQ5
rcx7OW5dTu1G45HMARweHHPoQvFrjAfpXwMuS+TulcDFJ/oH9wSSFUqXePtm7w81q/aQKQTqUF1/
YzuzeWVavVQaeDI/lraIvps9mEDx+yLlbVUa3Vv8TJ0i7mgmWlgQf4nbQqN4EC5WmkQkWmT5vqAy
9m9l8fbq2sWhQuTX5xRGYKVccDGAsUzPZf9T23jtcbBfJuMYS6WT49ImJnA5ZxzrR1vcgk2wmgc8
00x+9RPLaV3OHPl7kfyYaaLjFhfZ8hCsnXTrmLkbFcH0Hk7CrW0Aq1BKCUA1+hRfEZN9QDIuhU6C
FN6n+uYtje8lkLGKJqql8j+hmDJ7udcMb4kzuofgmrLEsGSruF/hm8kjEE6Lbx+JDVFLXQJ/wimY
5q1JECk4yBGsORYy75jPje75f3Yh1HXW3tO8jnJ+pTqOBDRP4+N2EhldWNss08R0DYCFzI+BvUtK
HQA97pOePPLnYw2uIHz+85VqlPGLmh6JN+kqqxGCpb1XEmciGiXblrxOGWg2rXIpfM6TAmOAVU6d
kCIOMjm5wcQtwOHuMylrwVTJxv+i+iwK79qHfs9VaShTJp3lE+qoS3yBzhbQeq25GnaiVBifRfbv
fNEj30+kCLwEjTBuqHPah9xtzyxdXskHMSsQdhJPDoKmJayxYJb6yrArPzkNjXQvnx9sssoIIqIU
V4my13yFCxjrfv/9py52mdROpDTU3s729xPrtMBFB6p64rc484iD7L09Vx2kpCsg1yopyHaUw/Fi
w98bqfl7dok00xGR8AcivzeC/YcxOfzEo5NlJBYBxtNOCIgl4yH4cu266PkdR0yhNQF0tNDhoh8Z
nSBGaKOOQGkW0fg5NDjpsZDIQbrxVFziKsR9DmJlMRk5SNkHRYGotjOwAjPdBd5r+m/4SgWuIpZz
nWMXtVUhOpZt7GV7gkY5tB10btRk7g5yfF3yEz3AzFYNLKodERETBx3Aad8fvEB0LPiezv1PNY7R
DcAOm3lLs5GNOKCafa7NGcnUldAPEXJDifgQOnE9TGFrFLBtSRjLaBH3Jkbx/em9SYbyMWiQZOoW
xsVc/QhKZYXK+rvPpbuNJBG3eQRYoRAOoNaX9xlcua6tOMMef5AVdITHOBEkbEooDKvyq0pfwNjM
AZLRn6FQz1z5aNuI4ggiNXIJn4ODdBrDSOiw43TsKoMEbDgUd19W/HOHKBoDiavwML3FWCT00bxu
DJSXrhe1H6m0HwTgyYfzZQ39KAzfovyv/ImfMlxgyt6Hnqcd+3RYBxX8C9UNVm/Imxu42KXbuCpg
dQiECFaJWnmirC9Q8d2VJP35PH+bK6fPOrKlMiHTZ71DzXe6UX4OhuIVMnbHkmXVeAe+2WFgwYaA
aLsvOKLd5ezDrQ+HJhkw+SxVCblNu+hFgg1Yx+EGXMOZdjX+1rUq/2+iqkKtpylVD8Vlfh6arUE4
24mp+z17YSiUlqajHDHL0qcu3XfZNpwtQzXzYdWAUtZQ3IDCVO38t1hlZ8ta9OJleLTDZWQHLh2R
MxOplGdsA8FnD4oKZy8rv2BDfD4DYS6Fq3VVk5D8fbhG82emWCXaTyjg9aXokxJ/lT7yjQmT9Xr1
2AP95RvMNdUN04dSTiOpJJseSiv5M0ZfeYceBC006cCdFWFLbQlhjHFV19CgIex198kURs3e2+EH
sb//L6Tu2e75pq50UmUYZ773mhnpM29koXezWy9CGMaXQECD/TosZV7s67XfmJ+f/QZzc55a33PO
Z30s3GAHmgbpWPM0EJuOPl0rbk7ADSVxhDl/+Siem1Ew3hsQCEOI5B+NTQ6PHv3jMJRQAZR5JVoV
IpXSbZpoivOMbDKZKiVnAkhpA49k36os4J6IY7rOuFVx1fXOvtc6lCX+6TNXeyd0sUxVLctYsJ1l
yDwJt36dE/UPP9C58qHulIpRJOUenBjLeb48F9cDdmhU/CoxbZ1rMUpHLOZCKlqhAumuooGeLF48
MisNXbL17toQ4R0eSyFKg/rZfur4Dan6DAepxTK8vEfd4lNjYuaLDrKBMiVrGQiZqNUwZspAOJjd
1TY3DibF00eyG7nW8RgrmUDbHLraKvlr9zureJ3WRfL03LQ+0fntWLkLX3uN49lUPfn6gVg/mtMO
cbVhAHSdnb5/e8J8fLJlEpCBzntPeIeB/LFc8/R7Eip9d03yib+8mzAnRV9snF27SSXxN/vteCMf
qWMJobssUMYpy+v8TbjbW/zM3T0VbB2RaQJ8ZBN++xjtPUodDAmOfJnZbM2c8wi+l3rAQtGP7W+a
/3bP13J7E6gEfu02l0W9YJS6jrk7/uuPwsEpc+DYLmVoxEQBs2ZRE0jm8FkbVOQhuf6hHHvgn15b
69lp/6vXuHywOTGcu+5Xnz3MOkuurqHfT3fl0lfMNDS17t3aCHGb5uANdeuAPubIpaZWmlR4IqXz
Bwhma50XcJWthxX7S9BQxAw164d9CK61X7PtwXqdXGfYy2c0PL8O/2jDFiTzbXCf3couWW97V5qB
PEkW+FyX25Ib7LRkG18LF29piBuP1BJwTTm5zIEetd5I0raZtbw52mxanElwrMHAi349C4YSF42i
DkcMOOjfjjEJvIh/TZXG2ULxcCO26GYE++KwCM5vpYRd/J2J+Ca7YiD7L2hHj+TVZRvH6RCNmYo/
nNFH3Ve4tkX8N52cX0/t88YcdHSSPVFv6HgMr1nwbTGGpMePIdEGi6XbvBUpwF2vZPx3Mco7lHYo
4jfPaTai3kBOcdhawWo9/vsF04/oziUWZtlUw0vCF+0H0xOOOBbDjejYHu/MPw6eLEc2kecTKELQ
wPn3z9Ti5WTXoh8SE0t8CpmQFZtZb/TGD1mIJFoblZatsJHCBsC6aoamLecTNfZVkff4Xxs7f2IV
nSpRobLWrFa0OKN6DHMtYm5PsxlnVfLbN08ctSOZdKKWYg5f1bHnGrqlsRLOr5HiWxi6E9QxFYvj
xaM1lDTAUVI1wYbNld8zaWoe7OMdUV0f5xxRumCflD7bvHAIa7RDPjUOfZI5o62eit4pFAQ3xoFo
NyejvjvNN5nNBJ10gLJM1/2q8IVH69cEXt7EECqEW4tCEDnr9/FTRTjip5XxIs5ss8179flXwpSd
qBBe0shYLV5fiJXAmkDfjr67rURlJmBrO+eGQb6gcJbIXUGEbo7XPNIffv2XzS2xoT/nIQkxeto7
Yps6l0jJTu//83fH/n51SSmDMjs8Ur0fGzgdqAeCmlMMCJZcx7JzRTgGeKJJMWUvNwgQKu63c9nW
X2ia39yjqcAGCBPTiXI7zTmL0cPxRoNzOT6gwPwyKuVhpVivMKXfSM/VgkxNEcNUdZuFaheEXVuB
lRN5A9aEt2T/kryyzij6ieklq/STrVoS/hXCqNW2Gdk8acY6S8U7nyj/OcjC2G5hS/VdnV/I5H5m
dgJOW0EfgdYdhsXOSWz8n57rBjp9ZhwhJTzzKXe9nyYFIYGx4cGAEd/HH7muKk2U64SWTGGAZw/k
DTIFA7pAE3j00x8Igp532OGcQGIltR0tJycftz5y2+C10DsNAJNyOaZUbnO1tzOse9+9thUZ2m03
3dL1nzZI8pWA0dqyRDGq3Vct6G5mZ38LTKCSSyrwswISLBtUOg4PnD6iZqObkpijZd1E+4sVOzca
Ka6HeQzvdaZqjWp/IaYouWO5uAPuN50UCrZSRaao0Btc9vhEzW0aZXfzMs8z4pr8ARgBSjdGYelN
H/kpE5UTaIKiTuvu7N51tt32BpSF+flarUmCpXrduewVJLJtlRg2Kx8en1xzqzBYNb56eYCqQp/B
9JhCjwzbSCZqGxKO6ry3MOnNKUfsEif818VuxUhSNi4x9bs17H0zRE/MZxXPBqfd4jtxgkeFA4qg
n8R46faXOClCtsvuXA7ej5Xgvyt6r9FT/G7N2JIM/2DIy83Bc1UCXOx6ch4c0YoWtbAClrJdS/ss
xIrWw/6SuWrwTAw+KFLO60t8oEEpV0qSgOOcJ/lmDxFRuLTEeyOE52RVFI6DTuw84hsxHCNvBstv
2OzHSTtP73LgWCyGYZYutwYksEXvPI6r/wtcu3/9XqSPBBvZeiJjrrhQgqqMgkGDancCGlNE4pDW
BPV6c/oKRzd/9V3YHqe4NSHn5DTw5WHGf7hMiNaxNyyqysF183AsV+VO1h6wOBBLXGF4B22NiOoe
YizZ1XU2H5WcuES7p7UmWc4txvjVahI8VC82ZkpM1FZOcNyv08Nb85TlSowAzwM5aOJiTNmJZvLU
rRPPzFup2wBc22kI6xdUK+CECPcLaIZyrCUNqpmyizdW5qJJZ81HHdn6WTUH80Lbn34RaXJTVlLh
ic5/yOPwQj2pp7vTQfe7VobVOjw1KLeUxepuyy+w78thrGzXmrAzsSIHQkEQEQLhwyKPbkjQGWhs
JAyZ/Pjnon8CgqM4v6/3vaiO//a1TUf+AwPSjnpwntixPxD38vx0kYi8pp5GywJ1Kj9ErCypxItE
XUwogN33pClnWSJuCnhvEoGzQgiejeOHeCehg060MxFpl4XHqWOEFrGZtJttyVjHFzLYAjifWSWA
S8DEUGMNNCfNwGRoaFXvzRrhoM/gpM8e2UC6rVyLoiZQFrfQzHVayaJG9iVC5nrlnNlC0vjVLs35
yF8wsde0HpEahAk847JhRdWI+h5vS/Y4gy3y4ImJc3JAYd0LHMCZgIX5J6BxaI4pabv1TSi08mVq
Id5+uzumoL9GftPGJTmkwTPsss4svcVXISEW7XaPysGXXFDfSlIYPRukGVrSSL05yQ0pefo4hTyd
cHu7OW5Y3ehTHBzDXpCMLaYfJfChCES4zZHGvPHxpw7op31PuQmT+1NQ7Uc/Z7n8+H0kzBmSxAlK
NVoriSwxqlunjkw16Wk3d2jbpj/pUuWT3Ljvlg+4a2Vv7dqRWJtWbpSpGm1pjQC/wGJwxbutA4A/
onxJq7NqQ3OCt02Z3hP7qQr7W36YJJXr35m7oZFikn6vh860rK0CHD8tI+w9iSlFT+yqzszCSbdL
zqpsvAWAhpBDg/LWNNg619iqa05BFhsOG0jI2Jwn5zXpaEf26qqV5ad3ndId8NFXfDca8GmmvEBP
rnQsX5fQDHunnpH145hYXZBqYM1OSZ+d2lhZ4XIlC/+4IJQ0LkvasRUOQFajJ4oTCpIUmT0OED7P
ro6pD7fhDgrxnrf2vs1EIyy9/dIvHtdTYojpygeq/Twe5WjcsgDDsCRT2bO1g6DulAz5LOMeh4ko
vDpkusxN4DipWVFNY2/XsmA7hjtZgH2K0ephwlO0aoHmnlAV39w7mSsQnngOMA9qeMZnrwUu3VZI
24o9nU50o8CI/o+wuK6DJsb4WD7oOjwYUVlwY4jEQl2C8gOQZx+XI833jV6+s2VS45RA2sHgoId7
Mo8woyqnyspSQaoV3Nmjn6R4qWQsOc4DDgOLA5ReqzNYPsp+xg53mgRZcSbUXS4BU1SFUoRbk1us
bbKjwiVBcuhmDGiNI+9n19fbJYIHJjIpVRvXGa/D3b720n9EnsVtv/XGQcx1qIwhuRqHPay4d1j4
sfwGPH52TnATKgS4vSDY3VblK0o4dwDVYcDrsT91eClFEQqagU5dsv/qypGf1w3qhBdDqGINqJt+
+UIeRajekvrA5H7gB05Ez14RstuC4NvOf63Jd13/OjzHew+HnG0DmaHBEcx/+NHztJ5UrFIxb93b
cI2v7jXiOxBzCap9txePTuyhlkpuHXBjRkG3JAkE3uK+RFOtxbKuehPtkCkXiLt/6W667Lmf7z2x
qNvfRyzu/DCWIVabVEFwOQ4DT2ipFuR+YnyqWB6F/IphOIcvWX91iowjzZyKVX2v9YcjJWWql+39
O/jVMt/KBWRPO0W9BY9xGW9OJbQ4e6VTdIt6APpHQpCrBORUbc5jblhxRQRlg9z/JcUVjoagV7ZS
n+tzpOzYFk6D581u4/0/RSnn2v4ZMN2Tohww8mxXaMNOUnSxeIR2Of5rJa0lO++1vdJRUUBiTIvW
SPqNWq84M9FeKs5XcDaCXJZDCqNowscFunJ1XGx2yjotOPA2rqy+2uURR61slLtSxUHm4HZWKtVV
bM7HWVJvu8zvsGRKTt8v3hYk5MKvtlVbD95ktfsOYfT5tKXhxW8W/gAj71jiHo5d5Q6DMb188IEl
X5VSkgmdiSxEks0ymbX2rTOet5llxWWwiwJ7QI8vjGroajGtwCV8j3JhzO9kTvKJS8nkNQ2+qIjs
WLU9eNjqwKwTGN1hvN8y5qcjEsdRPMMLQRiplKmTlH86J7q4ViqUKjAu2derzJse8SmqdV2gi7I1
Vws9pd9W8P9Wffe6C6DV2qUQluWWEkxOQ4gjaf6I7b29ufZBwx4AhrsWpHzcIppET7MPCldI1ReK
aKuNtQXx9BXvg5w5Rg0WGtiQ8k25abRBZ5A0gS0BErjGU/izry7YWaBX28aKO0nt6GfrtzWJCxsX
DzHiIj9NYufEJyFHE/S7LDYi65cHuYjWAKjlvM14f8QjPbE73pLVqHLMDckZ+2pTj+9X1JcZ/Z/L
FfxawNTFWCYQ7dTIBY77tiQtQL5BtrJ5MFpOSAjUxsb4NKyiN2SLMyXmdm7X4RHhBZqprtw55aYx
TPl/+b5X6SZrZ0k7bre5hvIwikYplrkIc7weK/CVOKTbiBWfmGIv91eVIVLRWbQFxiwD85N3vH36
BzOBsipxyhJPaSwevv7LnkZZxoA9gfUfufKbQZlgxlK7h+0HG7aAldoNpRB1P5ailOvhWJLzU1Z0
N9f5WiPDL/OmelW6AQOWKfvVn8wlCDKYZOdudSLf1uoH5u+WP4vDFREwUpHbGMAlExbEiODvxbB7
Fd8Wllxvwwr6h26OvNjYcrVHDq8fcqj2oJBquePZcrBKYiu+EfvEUWyn6WDmK72xuIk/WSSv6jLt
CO3lutlS+4X9AEW9vFFTHwFJC1Q5Sql2Lo7Wf1LK2Xoktquyxvz0kR2kdbd95ALpp0wONJWXFuN/
qxpQEVdBmaq/Su4c/HHg4cjw8l5tF8OmInfNmMjC1BBoUtTR3sE8CmCnD36pN2BGbr1W+RTN48dl
5pbwswzYso/aLlZQu54gTOJMLeZF5tN3VJCRKI+ZXE0Z07xrRJrQF+xYS5eq4uNAxoKS4RooEuYb
esr/mBlG/eZ8gW2gjrlNxsLHEEFH/kFIMPPIl5IraIPvsBuY9UHiJcNaIQyKp1lbjrfFY4gOqJjz
RnfjvSyckWF12gpx2ns7aUs9D7qhjpIoV/5ATbvEkEuV/obuGcVhwuPLBmrKXRmF2dkAxLxnhXrj
iraDGQBim0mW/ehQiUG57gI8mQe4fLuPoLUR4SDVmAcCRUwSJo8CHCE4QqqDwKw2nBPySgYmjWAV
JXreeYNmIAcXNcb07Gn01i5TpE43vMw9qx3HW31ysmz9M3DzkqBJBeKUWmDmmy1cXqPmlTr/ZC4r
FNAGbrFD7jy5SaZvQMvmsZ2Ji6GYIHHmFRWs/yovfYGjCA/qyXoIJHt4A7nc/hVCL//XjBaIMek/
AIsK6a9wQZFxtk9tYB7/Uhg/X+3qArRDcM5UOufIjxpgZA4y/veJma1a/g+Lp/pT+DTgYu/dlpCG
DvZTwIz8Fr5+6JN2HzV0uTND5Ek5Lu/8owfteelHxlLXA7YRCTQZ5Eqi63B+z8vuljrABQIf6yx9
LZfuZOY8NXnOqMujac91XO1v2ywpMUTHo56dBWmSxkYftSVKcPa4rMkdw3BhiEjA1oC2AtIc6YC9
6RvJPtqImOFbnQAZiB83zatsKlNueU6SqxvlYPBhV6prRxk3N6i5MVI+06Xr6a202ocB4wB6/7pk
ynrkwBbwVCWFy1QVL5C+lnfWaPravar0KU/QImjsIbGV7IjYdAzqrBtG7OcFueOZPY0RpOA7jhQe
GxMyhg16/nChoHBrwOPFbGAhY+31SSubywG5aimF9qy/nJ+14OW+UFMmluQ5WXkOxCg7AxmDFeif
uxMS+qaL6tED4qUQS1nls5viGWDtxTSWARgSELkPn3rr1v+hBWkkei4bHs/dodc9cMg16YnAOtWd
DuZLmh0PTbmnjMzyii/lIGCQ9Ue2kCG/hbQH2JkG8c4sX+cdwahGv0slOWlu/4hBT+Nr/rykaW0S
CQqeehIl7Z6aXcMvSE+Y9Ysk7f52zx+qSEQO2PEpgIH2tuxQNEvGEquqSmhXBdfqCY8cayKyhgL3
3F0EiOuyEAuVSR4IJ0aXdW4ZCkiQRUHj1bpU1KTj3SPWtOkhM0BNNhtBsC3pnwnN+jEtUvElhQK+
xJuATU8+8yLMh5Gpbi4uBt/oOTRN3EUSebmWS77eV/h/gtLchMfDv+Itpyp4v80RUatFLiJxlj41
lU62w6Bjhwlx+jIPP/KE+y0vDd4pYvA3r38TdKB+ZAP9Uh3sYnJSNlsTP0Qz69Gv8L5bcjO+PJsY
/63HepG6eitQBhH4eZl3bK9gi7+UJlh5xAEQWQMVpjBki9kMqhScvKeCgW17hzXFs8T73/07xfw0
i58o/fMAmdJgMTP06DmJ+XzLDipY+NCZ3Xss28PPHWUKxz5qLtrL+WTwLKS49455fzWnfrIr9vEX
1Xyou8ZYGC+3iZccEOgz7mieZzGaDwDq4IjRD2LH0HIcWdbhe7IKFIxuzcy1EvlX1ELdQodG6D3e
abGbhjfLirmrLs4Xlt34kuB82RFQ6FdDrYZPr5QtLpR+7WwW5krnrKwHMzoJyXnwFUDci9cpsR9q
93f5rp/U+cWqDqs59mA2FFT8oBwwo/fTBbGaiQutuUh/h4qy2P3ctzPnCNBut6JGdnG7UKaRn5OE
qWTnUbTUTAqfd7pOJj/efB2Ac+ymYDbAgfuaBVk458wG/Cg+EGrTWKQNBcTLBcDd4GDaYn6MdMSe
aIzgbwTGoRc59vtYoFZRY63yhwueeVlw6qrhUFgNMNACkGO/72x+bvkg6pss6nwGWvDcgRdQotb0
V+OY1KPf1VzzahwgZbOi9y9cM8CEmeBIF1/ewLA3wrqa3NcbYKA4TK0l9HY5bg4+X/Hv5teH6+wT
asXgdb9SCJlfhy1W6UwQD6g1wrtvvOITRYWKEdOzeipJB/PmmheHho0cKvKoR6y4vxJnbFgK5nnU
yAy5+ZFRUqR6MFn4zEVzQPflcxppmVOSDFQDaCfo9j+6T5CCX4ccNxoxWyCVDRsi3WZK+jRi3rCY
1ypZLcAlQXFoYkvg6SH66IXoIXpmRbK8uGphK7nSEjjk/Tyg0WwYuSth7D+fF4It8uJ2BM23iKbB
grqDBiAW4g1p5i4Vs68O4tFlE4PB9Jz3A/euCDImw5YFOhtjl6aTEruCz5xkBMu29sQPfUdSLz6F
3QBiQVolsjQ85zx+glzcHaVbMC8CFGaqG2VW+uvPxU/pb7ulk0AuTSDb5d391GF37BSCYLl6J4u4
NSyxfdKN7ij+DHGfmOabcRJKgg54IzmYPSzR8oNDuRAsKV52wE+hruE+SIevYZ2ok2bSQjcPy51i
UTd6kEj4kJSDX6yxd1L2d7z24IUtvHIBIJ9KKhynME9nMH6DHPg0nS+VeyUgXndDHypoSk94eM+j
6nek0dXzXf0ntiNj37uPgSNw5PNz4fpvz25UYN7+daHGGdbiiHbTiDpC4WBoUg1L+oj++32osdZX
rNLu0TcphhyD3DlWz81sLtaf3yvRL2qBG7u7rmuwAza8ORvhswiUEcKPKe3k7AZQKnnr1fhDgXTh
UlxMfDG1PZ432TBgvxDz6xcGgKGblssobcsoPDHG3o6repkhNOJTKM2cEQvMrSoufDwUeKIn08pS
+B/sNBzMPYUIwIHyeuUnSmWHAG9j+sNNTuEXGeeuHj9qO55Snc9zXsTuUFyutS5395vn+zBPDyfD
15gAQt41YmLnOmn6HBuV7pb3cVfZtRNezrlPrX5pqa/8CWQLY+8OQvbClMeRD/ilw+vu79HxqLuV
EhnLltcyN9AXqf2NZs8TGf7ISeczZi0kQCVUDGeSjbFkYesmjYX0osb+A96m9SNokVV5lrTdU1yD
bJozzj2ooIAB0lbY/4WQERQK3FyCAJthlihIZ1FnaMfxAotPdVuderDl0dKf7HWbINtPOwK+JhjU
LB92PysKMezSKE76xg4zTeAlPZDoiQxj3POyEQ/16x/jl+Qrg3wNarpHSgZMnoQYuzLeslMF16Dl
3r06ntKHO+Co/i9CWiQDk/fCwvRD1iRMhNOyvGIlh6gtGl4eOOsYKCLRvWhsq4MLnVj6kPc8SZNr
DWoXXaI0229CaMLOs4OfqQWMtTyIsSKjEquUtHfNbTVe2N+E195ZQmMzUz/QLlAhxpzUwlhITfDf
Sh3EAte/ViZHmXqbB1Id1ZwD7I0jLHVdrATYtxnvPb8WPlD6DKwG3i3lY4NkvouhnjEJDeO/33sb
fuOsIfa1xP//xecweFhw0Px1TA5f73qTOLh74H3JsgtVzHsFBve298y+6qZAPRNbqYORxAPC/7pN
lVhIRzohZR+e1/7pFCHjArJESkBSNlTpNjJ9Pf7uT2d6uFItN9jStBT/w2jE+54DJ8NOwDe4o/RC
AbCVn5senU7jy4sEu9T6V0rSvhHbVjDSAz5RkRN/JUTVIPYwN5FK8/OOnpj+MRv2L9fZH2w5z111
6qaMoHPGE8CxrSViJFz3XZvvLvuQOB9SWoqA/aelbbknpYGMvRDCLLOY3xtLhXtv4ekzTVS6jkkn
1Qgw4ZoPFQ+CM2l5WJuWhZONDRK4eVNVhOa3ej/1kkO9J3PnjnykKb4LzILgIolFTFGcKTUlSfOD
lyUFpcv9NcFOzsMbTig5NLrGzzR4x3vjMVsSE/ki2F9Dhb9ROQg/0rpB4JNQxroRldeYO7LDze/o
B1qAa6E3iXg/CFPQPwtjF0fgqaQ2EPsv0/vT/Zu+04sJtJE0Wwz74/LIFtLPITGZ3RtHxB6WrS9i
e0bhh8Z6Cvg59Ruda33kkh6ksgORq6FtaUTofo94j6k/5a4RGgl0axlx6Qxp6ivF7tShpM+sUv8J
YyRgQzWWyODV8QkSQVEkqIqZjh2JPQV18USZew1fFFCtAp2Dfu3J8NxyMMjTjd78i2eSqtCXsppR
xf5x95VB8BzUR1suz+bxR8S1qC6AmZ0DERpwoBBBI2/JI1t+PI9lzhgLBKtUq6zYOcIENeeSS0aU
LDIJdESqHckfiCI1AiKLaveMYohJSW7yYBZi7d1FTdc0ydxt16vPld9QOiJ3G1/I65t2L/EtWZft
Xs1ekLJku95qrmIHjOpnU6D0oJeLwbdfwPBW75KLEKGxzoUBi0+jfrCjsdXbgU5xBQERr4ESoUyn
N5w4uRAy4qI0CZ6aK2/jJPrrXTDtmygyXSMcs8Oa9DGLPwqxPobuPJYuAi8d6ncvAvJgRJr5oYgW
M2x31++zKNoF/B/VUcvj50rei7dZH9re7J82ORx/kOoxauN7Ta6no279mCiCMvfBnlXHd694VK31
z3NXk7cgrefZ2uoHQQO24LiNdMsJvCmMzZ0l1qDAWmJj9WSos3patglsHmcpVSpLzOkZ43NGLOyG
ZE2rKf/CEqqz8iM8hf1MCLi1W0FiDBv/YrWn650RomEELtFHvNXrnHO1mbKY01IKOHZc74R6dO/z
qIWX6TBYrg6FV9bwHk0xhzVjo492WhUF6FQWDab+AN0525Q+gE8tu1sEATOz6rktFelaA2Kd3ORV
Gcu1GAnjH7zc+Ai/h/3+MhKk3m6o0QB9DUdd/ahEXd3/PBW3ZmaPt1IWzO2mdr1Xgku7lw81mTCT
3pQE7GjyFU/kimiFZXL28zfEjT2FGlk3cWJXrKC7SdW9GWdsrAajJ83xusjZxc+m+jXjDy2wyqv4
xceBxDnBItbKm+/YrAdophd0EJJ6GLPWHZjjaRw0gIWNuqqmC8odFgp8sIhpsH2AmccUCVkRyaAd
D0B6TBhkxhno9ZGduO5XMJCJdV9F9QwC9RU5Son1lYJtNH85d1liGM3eDVPuEMuZBsIXAqW3XsK9
KJhhTB9Xc5lFgu8QzKbPJkRazRaCHvP1phC0YM260dVAA47StEVYEch03D5ksOEDhBg5WaPIjQsT
+aZ6yrhI7tfXSNYeaLjmDDrxxre63ILfqmWu0tKXgFiC8eEFCZrkMBfMTL3JpZeYSUyJAou1eM6+
yK7vlM9GHopP6h9SY5sRfXkMs6nO0NL2k/2+sKx86SxkG7EmgsDNRrpLs8T3JiNW1KAD5FGDgyPN
7sBBblfyDtLmaTka/pa/nem10dUryeERoQdx2MDPzF0vqoukR7al0BFEMpLX21nAVlDkygH6fvLM
9SfjBxGVMUq4yEEQBkP3PQedsipBEx1XFDq/h8Tww66llXF4qFMZUErVBa3bqWEzqNjQBcjQJ7dq
lSf+AbRpR4rOZolZdkIclUZLkMMSPdE2m3O/yCrSePIXJ+psVaE8Kj7X0YZPz5sgN/XAkiqyU5po
9aWSnlKuQerFbB6SfXuvtt/0DIJzCrZI4tS7lOHQ7n/BhoLKr8lr7867RI5DBz7hyWWaiU+5AOy3
ZHVfBnrP4GBrK7i8BUESXpXzEojxPweyTTzBh0IG2id3DgtxF6EFxt9cRO72/ejg0tYQNwZvL/C4
r8A+ZDropi0FZRv1sKxSGK8UXPtXslpuI5VOstb5ZJ4Ei7Q3yDjg+a/edWP7XoRkUxn2Eat5cFNE
ANySVzRb9EqncjIdgGhUVKIUu2QYP/uAnaf6AouH5kFLrBnEW87vFWmjwNVg8Y4T+3dv/LnXs8Dm
aJlgSSGd6TTLJtT9K/D2LJmSlPC8qRemzIQE1A9r0Lnb2XKaCWgH3kKW13Kf3ptss41jGz0fDyHS
Sp92YT04WUEQWQ/P92wQV0xElzRl+cIj6b5kS12iql0EPs6t6fzZQ4yn0kIaQviRoCE3GvdU41gL
xJ/GgiFxHoZXxSHmeBQioKz1FivVrmRHZE5KCC5Y2Zvyiy2rukYGYNNPL7X8IzCYksqcRG+yGVQT
aMVCo5u9UQ1Z7DFG4i2/FrafrSgcku33yaKr8FxM6vawBjOIrXWNcBBk2e3Nu3FghEE/0qeprYYm
ebmmjPXXEv/FEmg6bbZKeXF2g/z53aMKNo/HDLtSFGapS9xk6O3ixv0YyRrkIYhumoFDRGqGsai/
e9U6PnSjeP36rHFKcCpYMRONrjgsXHviyhiBK3YEwupkHxOFPoaBdHjqkKv79nJZ5YujW0CcGu2M
56QJKCJLlvS3KSA0O/OqPQUTQMlZegKJ5xmDzVoaWnp1vDAUXJLhVZSeKZNz50tIWpU+NKIYzx4Z
8TVM+m8TxJzjm57o3b7cf8UCXkokncxQQbRf2DJQU2v6VMQN3xAgspJMK+URmRF3s0QyzMNHP0/s
cwPrQQNH4UyGECVbMhUsUwdVNDvnsALDx+ygDy7qXZa1S0I1D76zWFW5qnCbkQIMAXUVqx8t9try
z7HlWaXHSGQ4KAp2/9Zm59FaAK9kwzyp3CJ1JcGsF7zW6yOzQRBCp+SNymapg+K5v/zhLsLVEcHy
whUBpj0RYxxIb8QiFtMYXTjrInpNnD2nED+2AfJ27/pDYlgfGxX+WsoouQtL5byT2J9FH6CP+VOT
2uQNAVY8IVNsoVH5DU15A43JQAK57ZsEpUM8BKvL/2Xof7aGjKTPYir0vwM9Rh8AJMf0FH2mgc64
aE6HZf5OidOm10OBVTbmUGv757kJa+bs8gQCzvMTGu+6CGVxj7aewl5R0B4Eqi8nZp2kU9WelIBc
S0/J3YWFjIK2waIhpJtz9y/SWqx9/9Ni9Q1ZRXN9d/J4VgYLI7y6o1Vebxu/UaI3Z3RzbWX4dT4s
Wpru50Q2EhfdR+Tp+8YvJd+WkQV/DmbmgdAfGFNGwz/oqldKWdM2J4gWBSu3voUpdjYPEYxEAXOQ
NzYcRuxpHhMX7TsucAZtWBr4iYgeOicTjscWwzyptxrP+9N0gWj748CDgSJi+ZuP46JDQlVPhiim
C8jIqa6fqA208VZ+VWFGkhv3zR+qjcBWWKoPtT4+3++ReLVpjfCADoQjbdHP2hu1uHvg5YtrEh61
Xoh5LRdgnBqOgFcd+1r+6zZO1t9cRQ+urUynrc1zh11M9bWvK4DEzVA0E4AcG4ZLuaFO8vlUBk+l
nHad6VXnsg6JE4FnMIy9qFEgYMRS1MucYpnufXw8D+r5v0YTtOlpaPEHCmamMiGJTW1s6LMUnreZ
EE8vv3MbhzDDlxT96zuw9j/tgxXYNZDl8liOilKmSeKtWgv0hllhAPCWdm3pKtgU341COSgUp+u4
WB7udYRmeoOf1I2T+URHy7BNDfytpetxqmaPx8A0qE/EK+il/JpaNhOkhKCKaU2O688SWE8awSQD
MD7x5VaQGshnzsA/Kt8iMKte/q648uocUAFfR0wrHnm3pZ/mL7nH2PWRk1F1Z0M00/9bm4KwdpMz
J5N2XgHVSlyCQYWZfnep8LMJtu3qE7McSPXBmVt/tW8BkJmNvP82eLzOZvkum2kPyy75EGKwJf8x
FGk0TlfPMoy5RCNYtlAX3VSsZqo4/sx2bTwGQFfskm48yvmkrOJoUpyed8WtGzZplCstrFfCZCRi
bVsh5EqSysh1QOp7aR3w0Spn7nL+qfblFfNxXpKOkJtV0PfcS8WauxFzdtZZWYl9fMUtDqGdufad
Y1VRRyHmqbTNt78ppcNA1AuKB0lfvtdds2gqKJ7k4laBGNrBmzEt0BZ8DcwXBUrfnp1RAUxSlG/K
5qZyYJN63uL182dm/zLH8GnS6CkTGi8p43G6rtJHzOy5DPMxSPrmmD3sawPcRBIyvrxA8YYqPJrg
DrK0QiLbUTxhudI6aH6Ox5z5FG+EnTq6URcYCr98NUOJEKKYASMcLVbYF1qnMRbXWyYUmRGU/udC
MzBZpdA88V/BGY1pNQENgduUL7p40HOGtq2gqdS/ACR+9ChkrtL26lonuw9T38IN5cDM3eJV4Zyo
ZkRxaoAswDG1PMJlLbSEQRE1I0I7YisqwrWp8NzHQBz8lXXPlRILssj/+a9+RWMuPIiUHQ7B0mHZ
4zx8/ETU/RhC6tWgMW8+o34cAgGf67r6RSxfYGHqosW8pELX8A/CjzbHPFfuFWFxu0d7S5pip4Xs
GN7w8ULKqm8zIavhVQZT8yTBkc+Yet9nUoJ4pzZ7HUv/tUrHpEVgacPTN9MS1BR/kThKyODRUTgz
e7P6QmOQdvtf2NI1KgSEdqwu6OI9iJn2NQkTtFWnfTgJ7/Y2y05AkET/lzHwPa9Z9Xf4+Y/pqVmU
75AHeSvN6+EtEbfM8WqAfSQVhLTzPoRH7HHfSu0fs5+amyTwc+KOwaTbbXdY+Lk9b7RRS7bfaThQ
yBHysn5CvwH2kjxLP7PM5Lo1AJha3x4kIWumrTD3hxtwAmuxsw4z9RDJNzZnzWigYYWjgraNgC84
GAqSQfAWz8EMMacQ+xUTidfloto/DMEEnqyzBWFIiVpmWyQAD4/FJ1i5LAzBFDKfD4REMJ94q8Ur
py0TyVdScMPYXCbgUMgnDmq34ODwy6JVGF2kywqchXlGI5cu5bQad+qs9n+QLWwg3ZCyoYeKWQDK
mv2go9usnuFprOVXs5+OUeW0mFEMrQ+AgZa3/IHNCqsMpEYyf3RK33RkTyptqU4VMxBBo2vDzzju
6jxKDOSDgCTP4DIGRHQX5bvyxwVDGj6m7MULM/YafYOWUnFJ416yOjj0EkeK1kCl1WWkAhHHLtbB
HQN3qS8wUYHp0V/RT/dYSBbRYykdPxGah5vgV/59kJaDIrCBq9w9GCR4MfSBzjA2jlBinyK8kwBq
JFu55TzkBSh8u+XI+2rc5Rbfu9QGIoHAhPIxCjTkheBxy/CmdCEJjZg8CQo3RToekNenjDITDgLn
OGpHOBXfyz5bnF2JkZGqm9irVkyqijg0uk+ORAnzPAeIdFexi9XzeEVGEIUtQgsW+Y0i2ioD9gxi
shIgfesqBb3LahqDIhDwo30OrES9eTP4vhz/G1nyArrNvZLmLK1V1w4YrNAjy2kPnYJNtG2v4ESh
wioRM2c4a3gntf0Tj9K1VkhyzBFND8s/LNFYorui/4YRXzLGmWw/990/GXW58hqu2mYZPfijMspz
GBtDOqGWK1EG/OcmYds63hZzmUW0iU+3Y9AFibQnXsjAo44wkLW5q4U3u5CbSzg+HTCrcrrwJote
R+XE5y5h4wnmirUtAvBeCEldLbS7jW3+nSXy+ebRcMFX6tlE6TQgiM0/fgTXCnbBqM605O3QNHru
5csaLNma8WvujdBD2+B9Dyr+D/xNq593Zk/9nWhBDwMc3NLWHu6zfg1RwzWB04l8wHfKfPycoikJ
yzCniMVB2ZpDuXd7FbaDBNIMLUuSjSXH+8DMB3CBR2HNuJa/pstTldCUtMzkWsETrcZVeVI+Z+OX
dZuQVeCNpGo1phIhJUXC7YObnZ8V+ux/leBjQS/EHQKm49gk/ESyfpXsQsTcGOmRWrLxim4PV1yr
EVoVhLYSsnFhYmXsrcwZjShIfTawlN9+fJ6jZFY5S26FOOoYq2qxEMZhIlsjcu3sPAe161orNGgJ
utpCtrebkQ8uJQDcLvK1XyRmdyEloO8a1RZWFlUAHnU5Z6zqC+xM2gbXJ7DYuwIOKYISeG91eLEZ
4XQuB4rmMDPG+AH5B/cy+O4mKz/13Pq2on9+ttzgJPv0Wh65ufkl9du/exK+xdJ5f7mDe2xdba36
XIFKw19tT5pvMRxiQ7V660VwQ3B9Pv44zFAZqDiEKadDTT750ZT2oFE+6mkrZspJS56q3qlFgxoX
7hh+NzkpCt6HlRa5/Lz1P8mgkD8B2xvvK3+x0WHO4yAb3vPeYeCW6BFoQFUDtcgOhTWQNvJQ5frk
yh5GHuKnnuBI1aHaxJDS+pQRtmTkb4vCiGKrTAg4IQM7xFSbzA28iOd9FAyEwDBXwVi1KSleMHUq
vZpIJM7lRAxQ2enDR6aEsw3Z2cbw/JmvHv8BPb2i5acrfP4O/CIS8W/lPxA5xwGAZ4/wzkdbj1LO
9pPs2wu0RZbp+qE7vvwCIliPr7fzxd2hsfd6S2ynwVHUq5pgIFZXlBTZgNisyQ+3b2uGFpF+OjCo
cqeH82ifKCEGadlQsD0vME1XQb9ua9pph43LIjnOwbUFkgM/pf3dylX6CLa85cZgw2cfoklMVEuM
c6+QVNn6VKnh6weQ1j0Ufzn55WFT6peupI2N7isyrgVZHNoPrEKuVPnqt5GToqfQUZcQPSywabJd
NZZAU9EGme8o5/0cm54sD7W5cb0wkHg6JFOBRgN8SX1rDLq4/A21yTv6U/T+XP4JC/KgB8svAMWH
slkV1ktvYvVtDRq51+972lp5YKSC6u3BUacm39HGUfuGuibI0r6hbwjD5qsivN8+iqG/F2WskEav
Yqtvj9up+2GHfjFR9za/p+az1jFv/3JL/W7M8EqIN006kCKYCHLoR+b7wN0+9OYs26KqbxUQ4cED
2TAUiijM/1iVvHsHkp7s5npojhhes9auypaZ7gxBmKe1uZH856YynHME/1kdKcbwr8XFwh6BLTV1
2LVdoiDVR+b7z0w7LSuWsfHFPe2sU9Ot/zcoW30UEn76FpjM0WdeoLtYWTVmCA5AtlFr3KnQrLD2
uTchsB8Xc1pFCl9a+K7fJas0Wbg6jb2WoI2g6wegYppor6QWhE81VHdOPStcEvx4//vKigy4yKyE
dLQcbHnoVltfev2hAS/kEsxeFm6yxtBMvZrHvkNydDumsBvDK/9HbgFUWtWmuWOS6LMOWGEEYTux
4SoPIFpnmIcLw/LUqQ9xM4YMNPNXnFGZ3C6D3z4hQo7uOvl9A7oJf/QKxMM/yZBpcx/tkmE+c4SH
YUEevV4+29Uf6dNKs2US+1hUp1K5AbF6XYzl/fLpVprsCrSeZa/E6vRmHBHyaEEEnXcmndb+ScL4
GIgSpsgxbwBYrqZORjZKsd7AgiS5Qg4W1nodD6+HcpP6MkNGqxjzsqtdPtMleZ2KUCNQgb+QdSM4
GczAYE4r7o6N8Kc1rVQ4L+YW3BJF7CjhXk26p6JLbP5TyeCHeqzbAOP8+G5nXdIT17uuNX9ZOwmA
EieTgfysBx2qN3yzBfNOCs/j0M2EtnA5+EqkrMqFfpyIlSeBllIxdIC8I3urYLP7Z6/S3utu6Iq/
6EDhTnjRRG3fsln7/6yS4sknwV+0soYbaPQ9DAjquVpJoo2XTh6AQzQhwSBZaqKmGZEkEljTGN0O
XJi878jQ5Rl2p9JjAZ/NyBRqo+HxLjzSmupJTkY1An8SqZlie3vIKdWkqoeEta26ht9RGKxLbmIA
dvUiDjSNi/Bfw2CJa87PMYQYgM7iEZry8RmIoSU16m3ldvRJlYEc8n8wWmdI/ij/nNzsqGvJDnAj
9Vkm+MFe2URTBDU9obNR3apZPpxFEviSfKweI706HuaLHSQKjaUYzZlztORqd7WQspP1F6g4jjQH
xrYKGN6u58KjxgoY2gBgVP7J4KWz4nqpV8k+4nZ0V6vdCIFcDr6biN58FHsBMLkxm2fwjsuPuFJl
n3rE4w1lMsaFb0EkGYJ95Cn/Ilt9QSdbx9DqLARVxt72UnA/GyK/Qh5Iox43drG9AudRxrR8Me8B
7cU+jijZkjGIDl5wHUtroWqJMR+PepIgqXIKhiJ0eJMyTmxYhE5tdpLxh97Bjjx9tq8M4zJKFSD+
6B5AlQ+J+hH+1BrlDaB7t0HhLLRPp93preCteWFJFMpLan3zXXpWgESAPYPgqMJADdsL2Ah9C2+q
1v6mP677+EZBb0nKP0g6h63RO7sGqFr+7vW9TCqHMTXcF7EdzKtf1hPeTgzkKzxxEcYJ+BaM3aNI
sRpz4cI6Z/a4/J2q03i+UCztQ7dlydVrES3mAeVYZcgQ8VOVtVm1baXc4NrJRCTtAssnaDGe9yeT
OyBdbKPOEYnm2yU6qGfb4I8/r3Dft4awccNIh0aEPrNbz2s0PTZK2YyOqK0xEiim/dXxlUS/opQg
NTJRf4EBrOaZIidDkUo32qOcfEhXRFC7xC4xEMD0NjacAoJ97hROlEWVHH8EeBgMYVeNZKk9Gcdv
MGL0i/uziJXx1aEcAgCksfXtsb59DpSs2tP7EgaE/X1094O7+6g6nwOPdxiPHcacxm1mvZCjO3Bv
DtYI78hh93/qYDNDYtN3v5jF4n3+KPDjt7aA4+s1Xcfj0rah72W75MwhsAlsW8E0CsOjLOf1ZxB5
YSjW9v0EqJOuyq+W0ZJW7leBN7HPnFx24crbMyx+qwb5tq6ROfpTbU6T0xAky9Os6D+zdiTx0LOu
tUdgWoxkSJUpSaXUM2rBCevZ5s/nDtQPMU0uClJKYBgX/BdBfSLTjsFrg4dd9GMjEQ/UVWBl5Hge
yUMIf8h0F3kUogni0IdttaOx5ykRSVcXJbhxhIqh8fvvq9OuojWHnDan85Su9V12e+zSp9Xzx5vv
KWAMPC5TR086+YjtrjtCzkef2KZ8bTUhaiK0/MnhSxkan0xQn0nTsJzzj0AGmmmTuVDHkDbgk6c8
FtqZaPn7pHDJNpxpOphU3nUgpqXrTl0D/evufQkk9RBH/w2k3uREVkrzVdWraHEQk/Ob3CayzDg5
ZeR78ArBwyHwRbKfhTcQNhZrgkcVtlxW0Da/mPLq/+PGajyIisf1nuFtCwmABYR30SRcot07YS2j
Gr5S+y1gTG+V3E3D9s0/0j1mHK7gxUvOwrEjLcws/cc3iK29mVqTwwGGXHO3TtDfKfh7UYG00VMt
Rr+iiGsFtNHV+IKRNSWhxwqJFSSfalD/kiwr3NJd+EvQISc6oxDslK+4LU/40ieAhcKRHBoMSdmm
Ajp/2k4T1MDqVmeilr+0oqocK69OR2hqD/lim63b7luU2wdzRZxM6aePXBjvKY0aGQwqAzmmgcNJ
5eF/5vGKVEQjf10H3JhTDCcOVZEg8sReUHekF+Bbb0M4+rZZGMTKJxI598bdQEfRAJZEEG5yIEAZ
KukLjuWzdRNd5UFTnxKcQP9S2iV+VMjWNH87Rj0ydX0dML73TGacxyiwsprpGDCmE/5w9MDfl8v4
hK/WYsW5q0lUejm84Q1NhwdOLn9GUDjoAJH1upo9wxJotpEscw9UamQlfTgEwYw+1DaudtM26Mo3
KSfDILd/UWf/4acdt0DAh3n0OKtaelWtyu/Re+Jw3CkYuhzQG6QGVtRU2Piiy5gFoSfDB47QIFKc
svgJMzgSQqirclkKIqv2VZKHCX7E38vYqPlw9lWm9gBexE7SFAMuyhSlt7cndJyq/C+uYu/6+k7o
jThypcZ5vAk9rjJFen4xmKuGGQErif/yWKN1/1+gdo75T9LXIyf0aIMeItO5yjsapsxJb7r5q75D
cnGdlMH/eO8PINUPy9kB8CIJqIcu2CWMGnjVziaS8rbGLH/GKpu7lVIL9snLzTGKqlUAl5nI7UG6
LQcV6G988eeI7Bg3KiBEXeQ4XPbcxOL57BeZZICkQ58UoETZ77ECYXNyzffz0YlT7XSONjOCpKMz
lYXOM+tzrYxK9YwyW3lbakkbBcAk38S69D7QsF0quxArc6uULGpsNBZCLuBiM48Z0iwAWMYGisV6
PA4emGFynk6tJfnZAsUnMaOzecMu042GsuKITxwggvJ5lljpO4+Zr9+x9u9DkMi4Ie9UOPe1nU26
0cRx7tPWVb7ZoCI+ZmntrsOprOWN1RD75iFX8vEPQbkxLTx6k+Xdc5d//tZFKYIK9vOxlEXPY/IU
aDb+RVdHz7ieXBOg7G/uXcNMvmLJ3FU8eaChBgdkeUoLS82/1XFZx1jUrH4hkfDT2bZ/dKnMJGiP
Aik4BKYvRqYNsTTXksFooPz+C1gd476bWG1FB2zla4xBW1JVBKqiJu7G+hE82GMWRmiNuIpsft44
aQRIHd6O2SWdAH66ZiCfJMr/+GcTvmBjtN3FX9Lxp+m+qyxt/oPx0j5JOPejvtHWaz7yzBVwSZKE
YDqDxkBqsC5hmmNxEhTV0xBYKMiCi8EfqpdE0QvwYoZURt//63TXwqYCF2sWdzh8oJQVYeIKhG0z
ZJLsZwUx+Wg7FdjNeLCBn3Bv88llLCksUrAlIWAlXnSQK6VQa3E2pKIsIVkwll2YqnfVs5gEMGch
E+PBRV0pebSya35jZ15sJuulCTcUH5TsGtW8uykQ1G222UwhYF8Nrh/t+CFuAXF6cpxhLKEZMCa9
Jo5m8uB0EKoPPfd/AMoT28cVEJ/Te5w2ot8J8+JpHZjGQPJ/wWEmu9vNUMy9PVGs5yZ+JMe2Owfh
QYXUInRKtdnCDDxEZfj9aI/or7NpNCoTUg1QPn3JHluaoh+qqMfkPCbRGCTlV3Ev3yJIyStgX4uA
wyutmJkwO8/GhR6NgcNq92QHqOyHqLv45XXF/55n4YR6XVqg39Lm1PqEwcOQV8HR3LH2xcPMj/KL
xb/3liTS3c2Ms8GUntX0AmcEpBs0+icwjZkqGz9j8agF5Ta3c+wHqZ2PcQF45YQP56YdXyFLt+v9
oAVa7mzcdNjQy5h22rAo1jeRIqjHaeoSuxc+gM0WtPWF4QXD3UvPsCxwpEv4TeXPXlM/IHwFrW/Q
AF+c/WYZiLUe3d7QQ95yQClaTFwG0/T2XjVXgJmCTYOwHpAxLT+XeJbpoSKNwGyKBIm/xOQuwVvX
709sNMRc4SBD6rCnDYfXjrR81fzI9ehXCynz+qrMJFJHGuKPT3awYFDmhfxxqeBgGazAH0YbKY3K
L9LJbAcp58UwXtDms2/LCWjLfxCNlFGFu7S6KdL94k0GyS7mpNypKKzdUg8gJ9ttPLd5K1bWzms3
yjvpHDRek0Z+Zcgu8emy02/5wDMS81EzZLp7iH+yad2vpolwhSx9G2D2FbfsAhVo3RfN41/cvO1u
8ErRWjx1J2Ck0JtQftqMOTBJEGeEFcy9Vjk7FRmCJn5gk+ezAQIQOmZnD16SBQfttTU9fbkcmjUV
f9a1lpmiNXJLhzR8dIPzXbraXeCm5cHHeUhJAGzVm2xHAOL9fe92Pp9tOxO27nufNG7ZF5Dpyrdl
0FxKBExSv9MHvCQMHFgjvj889B23UGnc+se5HRJnSprRU9cH61LtiVVbtVpBA2zDsj/utjgFO38f
OjxxvS9PgZlE1HHSxGCYgEPCnGOyTugHVr7krKINmcK4YPPNWcNiBLw9uDTw6TnHFF9OXz96ctcM
jnhnblWMcol3zMVBp0RQdcH93sw1GntcCYMmESriaK+v8V+k+L4/7gOGDjy2pmay9QkgaEklNIXu
p2b+624SJcpR+LETqLLECy0igIgNbBT5ZwmNbmMR15KNWwxRY3DQ2kDEfzhXBcYcuUq6A6w+8c3n
rE8GoxjTX0VQFG7h2VGazuZF4Cye51Cl+2oNvmVRlrLBWz/06+p+U1E+BIIjm5GihI89VBpEAn7a
QmtFM2TKjRVesHgdvnMuSYI6k0Pvqu0WVFnQUZnQEhBQGwlZ2qt365/iWyneIUZLvdhbtvAO6WPL
8FfZq+AzKRZEXe6D95lA6Xi4IR5m85lkuDovyqbMbVY9jtubJXggjjIIuK/mvrQfpmMOU9oIhnpr
uGPgbncp3wiHCVp/SQX+LXTD7b6gTRapscvQdU53PHeosVvcPvNfQZmpg5nI992MCDk8hoPCMYYP
y/6dHFQBKrUrdKyb81eNQImMZ6E/C/FSRk2KB9nuZtXiobAsZZLgqWxvrC9+sFZkQYFApJ/vX/o0
iQDmGUQhr3LMMSk953vFr02mFAgq0QQ/+Pp+TMHr7+G9r/rWKJo8Zcq5HY3uyzRjfZYp6qdyZ8Bj
6mHTrNjSXarwN/VJfY/hQ9eG3p7UOJvbIPzZO0Sg569UvCqW/6L7ZaWlAPirz/sGbcHCtzbGsABr
Id5inWiuv516DAa7EB+kKcLuIhjvPO2YCPwtGsVWfl68vxrpZT506jREyIw8wOtiRpt8b3220G1g
CmO4BQCdYO+ZFyqlDIUMoaa6Ji+gGJ0D3/0tFTPTivhFshtjljviu8f5IF87qp36NVXF12O6v3Mf
8815KqDwYT/lgZS51Z7ZX2JbIwQPNsB0cRDLTZOSF4EoLRQLrOGR5r9/4PLb9kYNOgrhgNvzojV7
wkk+haUTO79kMqqaTrySOcjdvP+Zy3hZ/M6WPhmoeTB9C1/vDrkXasveExz+teSMkCpBvuYDcFBn
rMsqfL8/G4Ukrzf6RwdYEG8VErz1tZezUCbXeSEfETdgJi5wiVPg3KtBXdRJ/Aj7EI0IvAb3P+9C
VgnJsQ8TOoBVcZmEWRcgQlhKGiapy5OO8+7cbg0AQeTu1bwU70pmB3vJe4yrYo/hzjhr9sgrN0Qd
+oiQJSXU2W1R9/YA+RL3CSoOBk3/XLsUK16r7uMhXpjAJ3xIuHy/NsFlJSoitXVTvI1Garp7cJQW
RR2R/yNVQCm+V2hzh73Aig6JAe3TVN2Pzcj+NTkrCPBB0H3Pf4zpfG2UPjYouAs4XHI2LsZdDmNU
jwEMWtd6sz0e23daj6pWp1zDswowp+n+SMIFEBwFrgckoxSfFOEfufEYESLR+wqmQX60A6Po85fC
BuggIlYu8GjTpqPeqo8i8vgiWSbqL6Od865Des69+OXi1QmsGSa+sq3cnYf2Aajy5eeD4Ls4LE/J
XK1RR8Yu9xQ3v72Jyhwk2xjKWCLuomrSp9/2imsnyNzApFCns9xLWxIpbN/ec1bWKPz2/EUh54zK
NMhO7XXuffasuH0LljAGqpU/NdqvUbgBxAjtJKuMaJTU2LcRP+0w2hGpPdiLgnFoK+myG3tDTapd
/y6mW7mqqj2nKNkZ53EcGGvHnD1ZzJNAjfQUeDudh7IfgcURNuCLZn7lNJd1TO4fkAcULt+j9pjZ
bvRDyTm5ZQ0l6dPvfbJsFxNU6e+1gp60cyQQ+ZQ0b355c0le0R+2oaumuw5zCNjQHtZxqJLwob7E
Xu/09HY/wuteyOh4pK0PbXJh2gQIGPuwYFPA7PiSIkFiauKnKEmfzg7rtcs8mlsqj3p+9ZZiRlqo
72w0rTkt+A3JQgnjq/fP1t3/K2taJusrSzfP+9lpWS4SvR5/muDVJNP5Ff68qAaXj5QPFPNmNv3l
JFpQoWq1bD9zPcrFqwRBKJ2TtPNDkjWosPCqKpgJUq3TEZLtITvMH9iCmmhiK09jZzEjXbgYMVRQ
uihYkqStKEe56pKEiIgCzcGZH834L8Tp7LoxVkXauB3tP7eFp4Vn0Iok6cKwbpCB7m8hS3kNUGnE
U5rhcOpT04r8+IMSfM0DkH1SaJPfJC+a4TsQH8yC4WEZ05YYmkVVjbms+KTVqA3EOJVn+0GVVr2g
TeqBkrW6j7N8PzzB+EjJFyBKFeTez86TpMnqOa02v/ptAzM7FZQvfEcbLsxcUvYqh39EHTJBxVvU
+mTCrB0iLOX6IvKyUbqTg0pOgVddILMsI0WAJe3u4eS67AGaxVYdHdebLlakxa48LDTaUQHjb2CO
FdGx7kWstrAUEl7PEthWczI+wTPdbY0UcvTiMYMzVrkxdU6UjTMMUR73C2w+YAfxGNfgR2LwsO9J
E/F/Qdq9ZmCQn4DjQVa4rf8qIp5r2HzTy/rzReop6ttylBW7ZUlLCtYfJo4YQsCaCjw6drA+b2Y0
H2EGr6+4SE4JE/pjziWYQr8hYUecWlmDzCzsBRMLIlB/ghrFpD2u5BqrKerxfESunNU8Kx8PdrC5
rC0HCmehYaqlXrvKcyOU7mKRo5cMG6L8M0JgUVD5Yrgg/q3nCB6ytkoHN5jTtnqvfsoDdZ0z83sN
WqO1icP/UxXmBF0cSBAydLXL7Oo+ZgEuvE7Slt0rRD5mhBj1m8x2yHmKmzZFF6BAGhZJU+8pMwsv
coGgqPkjVqcJP3LbbfQ//qguBiNS653/7QL6f53jcKxgGiN6mlEiLbgXLGbUn9CkTUB1wKeV+vdE
mbzj51qFkPzRDd29tqzA57r4g0Lh8P4fIB4wVH3uvqdeTYCB0D3X5BUGG6e3PO6xga/8+pzsxdvW
90S/OQaNp/GmD67XpOm6uJksPRP52bKZFeTq+5kDk/c33u0r//LSR8S/2c/mVUVf21fzOJqGexsQ
vovDH4pQ+j5Lk2gFrJFDsrok29XkcQrBiX0OaYHl8gBQC5XT+yJbIiv1t9VfxEb6eZx1c12eyWpE
+hPEYTt8qZ+xU5yXXwfOkh+d0OQo6MaPXW49Zr5T1TNjNRjOTIMwWP/b+rO6bBmhW8S40hnU0Z6f
plOBEF67Mk/YV0KtKq7BZItywWatanu507+qPoKzTeoEsD0oqLVr/HiAjVCKtagCv4HWlHVXnkWo
Uuh0LLJFMl4erdAkCuK/aQQ1aT+kdugb1M4BM3Obq5LpEusgK+0fprSy/g9M/GucAo+bZWEPmnjz
ctVGS9j9twuXhW9uFCsuMK0tVlDaMOdKX6eF7Oyc9BpcHpFOFjohDXXh9Ua+OCsIM8ZGKVN5dkgB
Nm/vyHCb9nduEEWcaPblvcWITbLDGaJRECUYoRufX9HJtZ+snROM3wKGDDJxldwfSCW+uQlHJljQ
zhXBeX3jiSi9OTgDQgtNIr+MKqaMjeap5cG2XZyTcc3YhzjC4hhRTLwxAC1+gwgltdG/kG+gRvl6
NNuhyKetwyEHkOdZ73eR6+yNUvTR5UK6ps+9zs/KqBGdQOA/n90zEJHId3YNNbg4PqzetFzPM5qM
JdVzkqsB7nmsfdwUzY88YLR5h9r/hUw5VZ+fCREtHPNQJyN8VO2VuDwm3+iJ2iMrVfPlCy3s9e+Q
ggwsdoUooRV1wnppiZwavFmnk4gwZzSs/03UqZ+51z3bJL5woAOUX92i8lvInrsHSsgsmu8XqDTw
uuu8z4bkZHfGxCbx7UaTJnkRPJGpEV47ZzzhO59g31SgyHkybmQtvwDCO2AVg1stU7iJm0qHp59O
w+0e4pmDmmUc+RFDalsd38BQrr6G0SdddIbmhHoVWqRcG57hxz0D2ziOH698y5vDFId7Oo14dxCI
DYwmnimOWzRxgqtDmA8W/A97dAH9tG68jy01NkwXSDyvaxf1JR3gCm9ZrOkGogUxwha8jbVLG9+y
hBucfhZ4SoGXGfVWn264f8YISrf96Q9gQsPpTwGvx2YRct76dmqDlAdnIn3X22vh+aIaenMCPH3l
9mW0UOVJwzcpbkBU4mWhKuEj+IfamBwHHOeQnjM13XM538wqV3xSaXB5nNqleYXzHUWkOjz9UIr9
moFppOnTQAlheD2wjUpjhiULIHVanfLu//Gqd3Io0es66fjAVf7wCuej5cblWxvTovV+qK8LXZKF
aZHok0qbgXRDaRQLJnXnWeYBypoOcCQcnkmhwxFzp1+V8Vk/0knPXeef0nd0CtrCfYngO3FnHr1D
ZuaJ4qM0p+qFZp33pPMn6Cuf+kEez9UX2RPi/j6r1EkPvcGVAie9mEfvhAO554VMW5XAJzJksoom
jDzFxKYKr3UPbYGv5Wv4POSGhtHCWPLPKrFqRNd3VWzcJWUXVPdwUVLZR+qtx1r5youLQ+G9yBkB
yXobRMGt+ragohfCRa6qE7LyXkJ2YnS/F10QmcSmwXd4xsR4QysQYPwFTnYLqnpa9O8CMZFxRUGz
7pq80d1eLYl533pICQpCctebpvJCGoxG9w7AV9N6KH9N2TDL/UvtwVLTGG7s42YegX+jfMUR6XBs
DBpyYJnmiP9qv/56J6my/r5YSK7fApgPWymkkx1OZPKXUvRQuG519P3hwRy5OocLHROeUw+22aeX
RU/fisNfQsWePHN0GdLsfGcxnGca1yQ1coK/gGY7hCWO3rZ1cgIetx5OaClGLHhoU8en7Fjqss5j
6yV8gFV9NF/MiqHX9eE2AuHE03wCuTW3rnTrNZFo6p1D8kQiyGdhDrLmlRUyAnuyMzNTuwGv7ky7
ggyPhKR7iVOSBZUNEaG2HJpfhCxYEQVZate2siBPNcwW8wNe2P/a0JbbVebtb7hlK+UoCUoDB5wA
60oEi5nN0YHSm06s/CsNrcxlxTZvBD1PclTenjxErzNQyQY7pjWUXabfTxAwhpQRcecIlRdsfpZN
8++fHxLT8xInHXWuNIGydvQlPZ+k0XhCPFdWaF0jAGbqiRmLH/fX+kENqY8nxWIHaQ7AK4QGwepM
y4hpoudZLyTWoAQSQuVZ+wgIj2L6Z7gqXN7Wb2lcwV7huUkI0PR8y224PCSILCjp3Yj7O7ElCTLM
PKNkPYLjrCOe1ch9ZlbFkFTFlHYwcFe5dHN5rIVfKAAEt7bkPL5c1mT0DtMRMhoj4gTnL6xPNYaM
k2NdgPn6kD//eJdSmO+lhZF7lJ3Bu8qcBGfyK5URS6I1PCvi861KTdPU/jaJWqZjktuTjlUwHlqx
bxFTdT9kG7tolASj8O0TpAFkH75ynOQYhsrpGsbtalYnSL3TloDs9zF2ec64wUyU20sDkufwgXWf
rDYqphCPpue/JrUnD04Qkioaryl3ghYU+W2sNVum1z0IvABzAgE2CuLUptWOHNHu95P91hIflodr
7EPae+JqYUo+FWzFoyzs5qd9Bpnp6fdtF2XClHRYYU2J69wPK1my0wV5skJlVCuvJKdd/MSmUVxa
8oTtz2c0LTW3+N5mS7KgZE+xlWK8gnSvhQdrpDKW2agpHX5qTt363rJrcVQbci2Gj1jlnW4fU5LJ
iRrcXrbeQTKQ8zT2LYK5yaDY/NdZpf+H/Zki2qmT0L3lgw0NzZo1e0B+Hwrr7z6OD6Yqav3W+tV6
/nBXbGJUHzxIwxV8VgvAhjEnNVB50P7YoO/nE+nTuvDc6/GQ5SpISt32LTQHv2jNFaLxGzWl1XAs
AWeDA8gDmeGYU0ILJa4UK91WvfE0SDiG/32vQVRqMzgu6gp/+t/G2qfSAkseZFKObISBCElKSd3H
ymXnfuDTqaAhF2Ag7Hqm9u0G3VYRxJZPFFmJn4MslBe4onahy/a9D3OuL3wPyTj1dVC7SkSZ475m
UB5LVNutmftHxzaePYb9508OELirdoSrAs7nY86zksedYFyrLwHKt61/GCQqrCMO40NxUvsa0TiU
A9XBZbARqXr1Id85gtsWUC0VtbOG84/ZAUjHteeNh6N6OUlftCW5m0Aacbsx+kfCf7rUnLx2q+QY
J8ADFXHZcRLi+vmhEuQ51+6FZ1GkCjaczV3zoMamXiDQPiWGu3JNfDvzZmFFkBV4ZBZS4zVsSPy3
rCj3XMPk4lUyJBjF/CHjN7IsWfRk17XMV4Ij0WGEebp0KPe7KdHag4vVrvBu5AncO2pfdmssSu2o
sCXg19tetGUJdFYPmJV8qPvroMWfG9VfCaeyx3ceOwwoQLc5+/2AjBsvAxnKz2AkJKmPh5uDz1Z0
L4hfNEjOnbalndnrOdwBCVD+qnIZStcaLJgM6gkDNfJn6zqB+UeOMNV6w/v/wpDIhzGRWGtbir7W
0HlzyEPWfB/pM6ZlesJTUQHjDHq5DJFV/Pv8Eoh50wYnykR8ZpWUIXYIMWkBNm+YE9huMY8OgiAc
pe+0wqClFsn55JH4p3y+Z2O+O9SiwCvJI7v+pPNMRW3cnfZIl9oxU/cwKNjbA2Y3ewlTt65tS7vA
MOViQjCpbKMexJDu2ZKi8YtZ0s1/DnDa48Vd/TXthlE45omA5t63vlHdSEuNX6yvgMuEenrKVCU6
ldUarcLfwg0cO/6lZ8zeHOSUyjzb+oBtUxis6wLCVWmWFl/8ApwNxRYGclMsVXL98y5QqxPAtVQp
Iuv5WkTJYS41KVlSUd+cHWu+sjL5qv4nZmCFZVvjHrun5wCcv7pfWSLAXnJfIaCN0qpAD4r5gzrm
UvOOBZH2+167bkNNfqZ3BT3099hnAOrCblFFhw8Ji5GvvyrpXOeZX7UeRR6XiVEmmrcYZFhQaOnJ
CffQpLLCQ/VIw8b/dqwJhPdiKaqQzxNsPsaO4Ygyhym9325/By+h0ee+xUQXIoxmZPq0gOX/qn73
GmgzBOmtVP2Wj2cR5zb2CBhREnAEbuz0xgvJb6c6UVxuNlFfvasHNFFhQnfOBm07xr4bI8gGBef1
hCxoHCyQvG4Jslal4kLo+zHCHePCsuSb+xD5tHsZwQan7bJGR5Q6g+ndWQwIJ/3ZstMM7c/BPWoZ
j0PZBm77iR3rWSd4FLXii9C/rIpptXPaMNclM/QozntuxDBiSeoK+FbXMIUG1d9pVoZV5rXLVpqM
OSYIR61WJ+9UuLQZAjphqzU4DThwvYGAjT8aukqNyRJl13cCMt1qetIaAJ8+9oJHoJd43rghAljU
+dt4anQaMB/jZuqQqfEUFgHyU7n4cKXolF1h6QytzI2wnOM+XSjnlRRcMJxXvYFvfLBBq8co54IK
wWK/HpJkqPZxpkFVPUPGmgnb879nLOtgA6I0cPUAi93TodQS7iFDdlbV+YKEALCkjY7m/oGLNEWI
+rbwJ0aUqXHbiE9Dc/FUMWrNof7StXN3PU1y9cXJZVur6VFOWgJhXVkVgr2QzOcouZ0AU/d8TV0z
rSJnUDE02gGDy9O17As/5CbLJdRmc6ThrDaPUMFj/gMN3i/HUhUxOhnAYmUSgLLmj8LXJQ/6mbNU
O9Ovhi0IDm4BsyzFnmxjIqPyXem8TX61/UTHTXpkpwUqemyGIRGyqpzRTvS91CC9PSWTlp04Cznu
vlKIvbVGmfs5fq1P0GrQJBBdO0IOmP4z7cdF652pw3wQLzCgnkrqG+qN2fP0c0DDSuYePtN+mSjG
O3lxRcMmsZZ0TMe1Ti3ZGWICvrjW10nFa9X5Nb0ePxAqj7ssjilEdIwlBViNllxLVvyQoom0x1vm
psmWnA6NqhdLZO6DKdWHryfb6H6Pqqlx0gADhsyHjzRet3Lm8weQUNVznlyXPRI3YjYqgd4MvbwZ
XZauPDYyN7FG4wzWqyhb2ff9lKi1bZyhWDoPGREOZi0GCyrM4VCZ3w4Rbusxlxp6dfEvfFlDt2p0
zBxtL+SBQBeJajbtBo16YAkZGo4ITQc9MaZAqtq1PLOG0qBNPlKHYFuWxDjwCpMH5Ja59FFbXGjt
m4tEwAS54e9v5dN7f2s/DFcByudS05n50iYVi9to/NmgfiP4cT+zW33ZwnP7icuVHVA/omA1CFBp
xqFo1M2673e3uGqKWSuMzTf8aOmNLQaKbr8GXFVOaVdRN6Ziwa1mx6LnOMkXs5sz/YTdoYPna90h
mFYiVbn77dgcA9YLZBRFeX+XhTg9t52Ti+MJ3+ahEL9Fu+ew5D3zvdkMyR6Kc0U8YeZdwtqiEIGU
lj3abrmHc3jSWnLsIIO8ZVNswAlAsTknJB5fSii2T+6h81498CX0l5e2HqnwjY/hYGbXwsJ5Oz80
WIbfLwRIepl5IcG147OoC89ehpIekxl0RXTZLExGNBowKJ/QG/OP5Dls93OP88n52e4LN6SHjXsL
WucDLUkkXiXVpyX6bV1kA2MC5nlq+hpBM9tx43q2/7u4y2qSwYwBxqz5rrwUTdfCmPs0be1anYCV
/Pg46j0pqrvuQndDxPELO5NfCtyk0/PEWb1A8BCYGxsemZ+yzFuZAwynMM2noFlhfphQQVcbHIOw
U9MNTFjXjh/+v/KCBmzdWtzaDKgtL3Qf3MKOuy+4WyFtUQo8rc+rX9kr48gG+G8DXADy42ZvJ6Zy
ldWlHeM4Woyij0hkvtBFoSkT1MNTGAlKOnu3/gy5M4GuzIVIc+xF+7l0A7g3NOid2theiRp46Aqk
UgDbZ37L6jwrGv2ZBe+0Hpm1A1C9PgCa8wSKsZmcVkBVkSOVF1VeKF5lYT4gryX9ZgR6aDJHQ1eg
P9Z8J45bnmE0Ey4qaFoKGteX6aK3drV79qfhJQ0Fu4ciyzY/exV2aKsLfzoGAS6hYGUcMmC4Fn5g
tPzCkZiMfDac6OF+1bKg1xkZiUncGm7CLAtzx8rpVgLZQhRvgsfZuwYZCtojY8llXBhZH5sUsJ/s
0WfwIEjr0gx6AxnyJOdA4VFBXZHct9sRDTVn76QfkWY9OJze/quvXv2f6ZjZvu974uF+fh+BUpby
+xJeV4hCLNFVQyyX/ujU8Ii3gu2yHUJ53nr6YbMm23IXQOu/x37irr8h5R9tRPnd/7DIluvPVaAZ
ijF3+MHvm6fA9Arzjjx4ld/3MGSsWfKsQkowN/Psc2m7avRpoMO4VJ27T/kljH8vRfOWxq8+0X6J
SRLoZmrxlt3TqA/VzDAH9Kp4cfq5mBDDoA+4C8yiyKzPfPB2nHnPoH3c6R7sIqyg1m1bgHWcV7x3
/HP5Jh8fQSuV+BkhsTCEuHPUmFwULhoCYFLDy1cshN6L2EnqyThWOl0UdZ8i1V3zD/YxFSwVdKMC
hw2guT9YzcTW1Bpw54gOcaDbgRWrQIEyHQq/CQwU/mpxhw9vhx/1Q4mbBxYZaBFTYBNZnOgfoHc8
sSAfhpUuh5p2SpoMAIVpybue7jE9+o3+RonU/20ztEzySJ2Fz8r0yceABRv4MN+grBiaf4wXLsef
e/OB0Mtn52JKGoCF7psTonANGcAUE8/QFvijDWWaiFvkSicVQ2L0ypFMhjznkPrpAEjbAHNGUU0I
b3elbjo98lZeozg/PNTeud/GrW/DVSN5Xul7oKJWNY7jVFF/HrcBzRUt5waNBGQelGnNEKbItd1v
2oLs1AWLLzwGCxUcxI0EJf0eSYOLlTdi5MKsy1DswkyaaROLBuHLb3txnTEyMqkpdbQpe3Spez5Z
DDRMjdrQ6Ngx6XS7cfW9334biEquNDXfuaRrai6jgiS9Y0JueTlILBC6IdviI2HOW1IJMYbXWzOE
gtNxENjD3KR2felyA6Kxbod9SIVaggLTwbw3K7TQvcmeWULIK8tgpc99j+7QtFDPufyxvCz/6RZs
+FDANWTHyEvI0BE3qAdeNyROeIOaYp0xS66SCj3b4hRX10FHOlcbdl5MND92pmeV8AsyEfUa6T9h
qUXihPNoV7xfAtLDC6reVyjcpJ6fnc+S9qq79lAJ/nFanahzDioriONcYKqkCu6s5oP9hIUJ/JiJ
sA9HR3GMXyk5gO0AEb6SVyBD70aL0bPRxevfcNm9yQgepMYWg1ZbZWV+lVenpaImDZxasgxb70xQ
PPC1Im14qNWEPuIBgLB0PObkmxUxxts7cHsOFaMq6affLyz3JiM6jC6zKNlw+1NKGo5AqoX807FS
aXE5+JF/EylewcSUFMle9ZzOpmXK2a6RcK3+3vyUHlEObJyd1JfIU6ha1eUm0KPZYidTKbvgMGZp
onc65U/Iq5g2pqqwsvEZFB/M8I+hy6dpDsSVmokcxx8yLGmhh9wkLYRmk9n6rG1EQOWrYeJS2w5a
JEJ/vr6gcGghkN+BvNWgmSGN+raTBVmbGVEIFh/rvWqV+fBNxYAMlvWVI1db7qCMZJPqXkG81rrH
rvFNHW1yso5M6UhDGRmY8ZRfDObvBo79S7wy85S0hhVrp1LaU7SlaW/0DzqbKo5lwxLcSKiyuq9O
KewDrDQxxMUGFaTJRmJvY1ooM3TAVhDzxxktojdAdDUWOfAFfiBB4gcBU93cGkjxsRx0TUT3E5NN
hK47e8l1PRuSxAvdY/kWCk3VlCtI1DVFXQAz+XouZZSl+b/Oeus5iBI/RLiaB3IXkxAlNIAmGDZI
VEKoiq5qRu97P9oldppEXedxf6p9G1L0swN1Hqhl880lfau2axE2GPS3edzfp3l1j8UYhFTVwi1C
tF1828ErRmc8XNI/2FzX7/9fglb+GlQ4LDlccCrBCYgOhiHEAzKBI3JD5rdgLp+0kUcgESZW0tkj
0paakzqTRZLT0WeO/lQuqIvgh5tlzEJvDXP9kEBYb5AolXKeBLUOAmTrHrfxHXhAxuFzwCO8y9S6
H3RWZMiYId4iunBrnbnf1jttuzR8Q82scsz/yqRRfGxnszoUnrZaPlGZS0ZNi+eHkoLfXdI2T8XY
I2xYXBkgGpJS6P9Ol3T1tgocJ7F6EEg+fyhq7A1W0GWmJW/fAU1rQUaSeBsKu1sg0ROGLwL9uuoM
0ISFAdjQZAEF6yXjGD/+QGaD5jfd5zmaAFc0/wGKe/hrR+nf2f9WFO0hWKcZ3kenFtwyi8xaUV4V
lIkHZpvl0+RAS/EkCIvtQANsd3X5BuDGMDDydR+gbYosdQsEoqTwai/PBuUSkrUCjVNiDd5Dcw0v
3w/MP1eHk5GJnG9zxQatfIsx2GKvyWpgAzzstn3dBp8GFHU6PWUsOx8ZR9UdfvvKUcI0rSBrbLDS
SD/roiI0v0a7L1RGQ/iBjm3owL7FCuJiIT5sbvX9gAEV7nq1WzZytOa3bkboCMl6WPsP7go8DXwc
K1iwIz2MzdS7cM4LJbat0kfhGewLSa26PgBRYM0+gTED0CUAH9ZOXc8WJn675H++YfUoyl6ndf2Y
ySuzzrG+t+0ITYcZe4hWjj040dqV9vVtqilLlqKjPmWmeeuUn+JJPw/niLmw1nIUwDUZigwBPzr7
ywUxksCLT/JH2/CEo5fJyvX93QBUJY9SQhW2Xdwi6fWt5q/hiBtj9Qlb+STkmqYsPsIdhH4IpJ8T
Gop/PduYbCnqSkcYx9IXmebGSsVwjJ1eDWMmLMlySD0/IATScwxbO54RP6DUdN8zsMrylkqG/L7h
p/SKJJfOPPknY7YPKR4Y7VTMAluSzwit7lphR7kvvzTrhBNF5FSEhtq7S3hFME4A82gYd/J2po0B
ZqS5S42RhGJGi5G/MrgSWLAi6v9yiCU/0p5cKIc5+8YobVwIekUdoXfKq0hyQdjMbyyBQevfhx5Z
IASbF8hJIyk3TBmQYwANu+E/gKBmNkYC63hm00TXcOYW1G4j1vb5yclYFEMpBp3p0pjhJGIXJ5ve
Qbaxb8rlhCzmMI3Lzr/QkrE9scU1i37Vvaoi5Y2G2TpQ9GvRyUSrA93L4yMIphe4FIyg5EvcY5m/
LJp83QlNQpVIeaSSrLzKXi900OJQAQqeD+IM6P2kWDujGa8gJsmTwmZumjJlt1+am9YXxDaSpZ7m
IK4nGUeMh6BQV7eNbvmLDqY0BjInfB1fy4G4rs/B5aovOYeErmfrOeWY/C0a/FnB7AQAlo5w3XD1
EdecVaMOMeywMpdHwyASSkCCDApPjjmyg+TFsvG90RMSkRkApKlxhkaofDYTLUM8xYkvZMJAQBAk
UF9Jbr+jZxhRpFSLisW0ifRlbl6WcKlEoQgIw7eALHJyaEMktXY7SuiGprUoONzPqZJaN+ivUHF8
zC++r5KiuS+HDVrfnheDLlsc/yQA0GlqrL5YUDlJOnthJJxDLfXyFybVX6/BjZaSxlgjbtLQMz2y
OkGnMLg623tcyiotbKDGfME4ThxoguJFypLyz/T6mtKTrTF2kxyzbpbxsA1t3pwHdGPxtSumQQQx
VemkgpzoHFuUg+7+3lxzCw3rue4Ntn5Qjq1op2nB80D8/etiFfUyB7OinzJSebLkZ5IUPdUxyNKe
whwjOM7zKN+Z33gyQTya0CfYEYTsj95QrPfXtI3txmyT4q52rADthKMF7uqpeM2Ltoa+F5eBrIGU
c73yKMx7PTzhd5sSEWZUXT2XsZGTSj4hKQa41XDYecmn2Le0Z+jTYC7Z6ftSNaqMDrlPqMHGXewM
8bcXPqRZ8GGXhw6uMgQArwU4QQZ/ad7sqtAH/fhUz2N9nXhgsOW30/mbvzpX90LdElbTm+pXE48z
ItPEw5KY6dbteDTXE3n46U+3SMtMnprPQy3kly496znembz++VMTzDSwC03O8vqfnXvXtZVKeLXq
CG7FvcdeGEnne8nEYDuX+Etd6RDxNBJdW2RdDftL6XZsbSLs/WL/OACc3v1XuZarLA81DSMj538q
oaa9D0Oj2otCkyY4BgBzWHHR1dzpDZP+9HSjwi5t2gHA9Q7BYwKMGHizXVMhLd4xcuwuqutI3/EC
Jo1Q+0bl+hedYHDOAPYUrugSwhcFhmm1Y/2g5whpxFwOulxCSpQECBGOP7x9jt8U7TyHeVQg4MZn
TZa5RqimxfnF7DLN75IZFHggLcWv3dBeK9rEb3DpRrH+2P4yBXJf5IRUmkxYeGvl//Ge6ruqbl+O
1vkZw5q6o3ykhiK4Dg5i/js2DIM4ae4woT3HMk5KMDlYq4U5pt98i0Kv4reLuWGrlKhe40HkCt3M
fUBtQxJnSg1/eT56CbnkUvkduuCTtHwpGSMvuZkRp2ZZp0m8bBO2zJte0CeFJcBdfMNeZKU83dYH
4NANrBn3ARSPn1tGaJv3AgLR6hzaIYgQ1E33bMLlYhQ/Xe9nGSZrn/c1ZsBbYqylFB+nZB2LO82V
6EuADwSHfYmYsGtwbq8LXNg82T49VuKc+4ZDLxjWiXNKXB+VX0+fFp8Sdbhahr+DHKLtzSi9aJc1
BHyMxmBW+92uEOSPFcP/I7An0CmyiS5L6Z85QHQRRzHM5pMqHDVs/juOTVuUxfSRQtEYMlpyPpuQ
xyYnVAD+pXiz60EGFuhCAGTpENKIFVqsSpQoltS63p86QwT1TS4diUyZf2XyUIga2qcRisIclXMM
nRGkr+xvAeexgRTbDDPSaM3Uc1zcXSy1SnE3BPHVM2tppTWdbgmg4D2oUIiPTtLSzI2FJHRNnvo4
Ulvg0PJ5rxt1Z7IADCmNuhCuretLBxn+eiSIorCOVazHqZyjaGS3vixpoMCEfa+i+4ZEF9KCL7gQ
h4T+B5UtBENhj/XPbk/HPlG+CaNgGHWHWr+jB4wnuyTTaaq0cPTFwM0MVg0dtDikkbf06VbkCpJ8
tB7ftVf9gsm9HLZNwKnWRyuKq0muQed9NaOFL0FWldD9N5vxFbeaLaEv+8xQgsloIPcxG+s+RAL6
KdtVt7l/DpXe+RWxlA7y3AndV9C7lS6x7x8XAu44Mvq1uiiQtSSkuz7u+erl0waCXV4owL3iw1MW
ljcKaG67S0zcE4BUnncte1mDt6x3J1IFCXb3u69S0qTUwXpIPgqPrEaZt8AWWNvxha1GQYySRGpH
iHZ34TdhrlYCVmjIy2LXuWrpCvuywQmHzaQatIcN3t0Ri3eyTb5s7hZELJCOIHiKzKzv0DmfPHni
JO7yrKT/6yWmkqdbwkSaTv1OV9b62Twi2sT7oscJ2pfYVOOZGyQ/3KMXPEti4yl13tPfSKc2Ay9Z
GJHnnk5booUiQNNb+IseXwYXmo8zpPbNkMr5KDUH53pnDYb0km5OYpKtFjFOvYMIYcgCTiZKpnU8
Uy8MpwCge5LvF6gAHVArZEpQTOOPjX+LXDgN82BBAKYNsgpOWMBdC3fTFo/9I+MFrxsXxm28dYGI
B+UBCkro63jqBy4weCuB6X/aRTS/37mEtAXlWVFW0XWIJKir7UzyNxwjk9FSK84aLq4UHWrH0Di9
F4y1fMft4ear5AnaHArZMzymsCbYg0uLiB70nNSWGurK3gIcnbkHc4z6Uvzf7i/3w+vfn2Z7kapu
rJ6PK1GHAv4il6K8T1qSNlvE3y7d0uY9ed0AccYESCU5O/UEly2fB3qfu846vqG4JUGq4Y/pIjPJ
wEl0+xn9GXK/Q34hecblJ7cC94rsoYZsYu0gaOh7RlU5V0elLEfq6jXZ1posCj62X6+hnXg4SpGc
HIDZ9eSoW3JDxCr3k7v2fMu0p1J85KdE9OPNjY2EGVsLi1EG2i2m2vhQFOe7wm0/IEY31K6slc1U
vHTl9fI+EXAnUCQ/n3UyCdMG/7kZcrxF1Ovrvye63o7PjjLGuhbXWKa9+O+A6FyGfUX1bqX9CrZK
HeQRaRYc/2iIxJuw7NCA+B+0wfzr3qTv6jUSrRbWn3mwj1c3cCHB9HXoTKZjkiNMOvsSvdBv1Knk
uPETv50iTZ7JIg6Ndh2NPViXclSpZ52PDSSC/C7MB0WFovQD3Ruj9/E/ZmP8FoF7Db/6EF1QEi1T
XgzpJb4OZJPVa1ynkCXwFpo4MtC/IvudBeIUqjS71ZoiEBd73+xPybOt7QVTg4UQZmXMove37jlc
OazgmP8o9DTHXRU5pIIjE2RsFHFJ3/HqsvAlNddxV7rf/YD45jPqhRrEy+toeWJkqBBHC5ksWOFY
n5UIaQfo1hIJu8YAN8/sk7sFS/929Dwsjz8IqGn9svOvppTVlwEeDZijx/gRKk/822QFTwYkkvrz
YZHknSTLZShZw6vaiERQTMXsAVrZSX9vMVKRKbZVuX6oJqzEP4antcZhUUtfCT76U5f2/fmldftx
4DxpziKBJ+AqLWET7aO51hNT8+AJazCGIOq5xwsufAigDU7O11WNkzTeFCTu6aLRB1GJOdDefAs0
SacWIanWBaeGFEbtqkz8cuLNBpbq/US1UITJrVCFWaYaZXducW8+p8s4YdxRrXrr0VqMvOX47EnD
B2vTnB24Vg80Y5Ye1rsWVBE9vGYdZVR9YhrSj+kJFk+1+KNQVEQYkEDBywD66HEn2VjRwcTw9iVV
ZgNvEcvF5BIXyV1svtw808pT5brpWFk218FC5eXwe3RNi4pflrqxQuyXtXZzAV9e2vOaVA5kXHEx
LhkWiR20w7HN83PTvx6wUZRGMCJSNQ4NMWgjBO5k4ZGXlTQg0HFgbKq2Xpq734qzPUeobyY59RC6
TF/rbFEp+kSbU69SXxJzPR+fWIBJT2fCfWQvZNB7v5at6tafBDnwhscg4H0mELBtQ0sSCcTQmAKl
hw3UDEI8+zzEn0MNUiG+FScEHqbEph/78a3HU01BSwe92rW/+YlPlWPTgezeItI4UavBwFA3/ZEx
7+plz0QVZZ2i047dOnrsyTuzqiyfU3jwFpWjcpkVOOVNORuBj6GGxoJ1yo2FJQobYtUhqiq9WPmW
fOeQREE26AgmBAZT3abWoxRsXUlDoZkyO0XdQfMsbMFyTq/zLLAdQognCKI2Yv9I7yR8xN3+u2KU
a8QxHPXkATK9KHYrtTQYgCSrIPlx1TGeg8ILQzvcaWy5pNIKs+4Ti8u5Pn3GPv/5nZljfrbctmvA
dSeovYkaJ3UCN9iBHVTPL+DXeRgphFfCq6144I7OiVgkfwRIud8HiqxAZJ8DE2UpSbRe6vylM7SM
B3In/tsrXOh1681DZq57Kcs4rUFHEBKAcH/dQ1ccHdslSv9cM1Qi5jq2zkWspP/qzHZQa80UZdf3
ydUGchoWOcTV+o1gRt/PSrXC2lPSWq3gSQHs+rRyZOqoJnctIPM2BxG1fK00lddjJAW2fAwzQqSd
OEqNY+JLCmQxfNMyZtlO9eLtMEjjj68cL5k+5Ngd5v5uKON0ox4Rwr7rVeJVaAAyuJRL93L7Otrw
muYv8TXU4vW4AcdxmmMcu+37dq6PQrKLjNXHRxhmB5cniVGY8tTummEkJ6YmFy8VkCpRDtRXcL5e
npPI8wP35FNwEtM5rrbuQRh8gNXmsFnq+dDYm3Wp0HVB7J4vIfL98x9fFWN93l4QARi8AZMHHNaT
cN3OCk/yvLqUD/BfE68k+t3W3mtV0JXx1PtjUnzzDbvS0pv0NYjg/eK5KgGONU74kmhxe8CmPO5y
go3TCYZFAUHF0OrMQxzGAdlAohEqIo54MLG8yBEgWfNKqJ0Tu0SDoBidoTWuQglhz7jnvCECzReX
vXw4GzuMEJAcbKHtS7NjT+05qMLpITx9ebkkPRlaBu4DzAPydPD8uGbIsXDPep6Xdphw/9NbUElD
9S7lmltuzoL2d9//RHD+8m8/U+oE2TRkSu4oBdgEnzk7FYuXKtG8HHgB5H7KnRnQMXi3fXjcue9O
qHFVVEEfuHmFcGfojxvS7tZdJ7RjovWcYzoJ+LoiuWsJAKRLXzZdRgd9H/OubBXNHKMLQGam+v8v
zz/V6RPyhkmZ+kxI2MrvzjImb4GZ7HzJzFUGcT2890DrTFcFnDRNVri5gxTfGlHS9n/0Max1gTAJ
S+Ira29PO6Y+vbjy2a7gNiZE7vGLBjwT6cGFgBb2xCnoSxl/1wQB29MX10AglbALmxGVVe0C8ElW
2HPkMYOP/PTXuZORG27v/iZ0EtIwNumqBvkP7c4WZWJI0nXBaNO06lcKBu2V/EdpFLJQavzhoK9E
Eb9iLIGzecbFKiG/FtJNrC1t6bNN1RwytRLiWml4DsSQ/69IvbsYuEajIJez/yswC3Txi1L/hLaU
8C4DXqEqGMqfupjFXRY06ZB+eiVARCkuzP31hPTL4P77ipJ2w7kw91KSGa2jBFGB2zoKsRL12Ory
IlDMaC1MoetXhFeYOkVJJwOBsLM3HnE6Ba2C5lrwJa68o1cXxVIIIVc6b2ipBpvgckZL6jGqQFAF
XyWEXFSXdMeVJIyoB+8LLBzKq0JthLVSDuRnoJvLqE7ezm8XShCInnJDnfFUtWd0ocA40rSWLHDf
bI4QrSSqOwBv9X0dfzv8BQhcp6BFUZJLcDsjokUKH4lXJbqKCAe/E9eVb5AYhwPy6PSNFv8JujBo
6H0tQHrh2bA2PSH4WV1nAeoe9726xElTKmQQdLJttYv6LEyBJJWm8Pip4y+epTyrFSKsTcUKl+Dj
IBNFA3p16hsGi/QrUQtLq/Ywl4/hzuknHFQpEYjIEouPis1/xB7UAG+fQdXUmQcFedTyq2ZChig1
0WP3QInNVa6mEo81eTV1hlTZOyemiN0cwlflrVFLscRcgDCzLhYSnGnWkXH4D6INXIvNxSZ9bPSB
kpASAcUlN840m2UZnb7n982XtQRrZ2WpOP9LV6Ae+Gt/MgRMyBoOyYSJoY9GHallKc2XvSKbLRm/
84ukGoxZ0Pv/qkS64u7rcYPtPcNhsYfkhwMZE4AyIpdfowW+TAjSzP3v9Zg2rqm2uvtOdRhlSEcO
6QpSGpG2C8XdIAhsziHqIg0mv/mdZkWmoIhEtNdQ/pyYLiZa6/SWHZNgX22QXqCAOYnBc74zcRai
Ba5aOhBNVFw2GAQuLKmxcGh7si9pnnyJMxbMCtNlAuyg6VaeuZZMq1zOTwh5RhjwM/CAbZKNO4Kp
CBaJPsXZUChKr2olbS5ES4MTcuv1EEaL+llfIO1LT9yUF6ZI2AMVBTta1kpnhenKIKpusofQ7pDW
/2gFI67t0DNMlpXbLnTK9aKuHa5Ourhi1awChj8Zhk3qwJkvcJVUKYZOiSznQVM3++xyiSQ0RVBO
H0uA1jSlGy4mq9tN20gIWPBHGZZFnOifRIIRE7ao/GqeNWUgLhrlkyPCAOl6TYH4uKNcRuXGoT38
MnqVDmWt9fkDh7WdnL92OzYEZMT0BY+uhNxD/l9U774TaBZVWV5x/HdHhsADrZmb+QkIHZlaeIzx
dKAkgdkJBfn+piOcg8O+eyto71C6VA3AWRfuTy5h06rEAAdpPY0xah8WzCP6N0LEak1z7mUjseRR
b5qLtCV5lhZbnPmE9rMto426TYwogxHw3NXbsNvdCQYCYO3hmFD24LyqwA0CHV5nIy1QLaqv6vLz
n9LfKrcbwIbg8dsNzjsjBA6V89tJ9nSUlB/Zo37ZyXU3zi7ed62qrFRmfrFudeYzcAk3jfBNUXYq
MvvxwO/P74ZG/ByxU/vYKgVuzQI40PJvFJKsftwDJbPVc78eJG105vap3jWcc5OQm7TlyzVr1aMh
x1wVyNr5lImgHxZr7tzvHqs37k3w0rxlgElvk4NryjuZweiXE6aMr2d4yVCzFhdoc90DnYgMD7K7
12jMtRTomTd61+FitBVV9QLXF2FpkwFrMHUaKol5JMqwCutsirAERwQRes0PsoXFg91b8b2otPqJ
pesJeiRalXQJ8dXXxLFSaQZN1Wd/esIIDdolsBU7r9hEnSFRqfNj/UnP+zXSdHS+UHewVx4MmXMq
lhlu/Gtg2Zq8dDSkxiUJIZByqNlSGfpFNzeai0wBHDr7CO5ovWdSBtzr7MbrE4xOEdjxXeEu8m2m
9ajE53Y6mzHtXC7RXLdGQZd4kKwp5E32Xa8enl2lXcUW6mcou+esowNgomshy0TT5nrOwZ5sRWzp
KRjoUyjAJuBbGzzQWedOyhPQAutfPNPS0pLzHt4qTRo2cm/5H+BWhGJ/v3CVhe+OL17CeDai4gV9
LXRviUulaOYQgWzLKxLJknQw1Yn1S3EzjF4ATC+nLmmoGYXOtGPDCwe/1UF5biI2yBvK/HjAjk/x
L5WlWk0b1/dGUTpnrb9SH/LRG64EPdK5l6AMUhmfA72BIpp/3MKJN91PtLJASSKgfiA9DGstWvS1
Zc4vv42h/h4jnWJXukrL0HLCSd9Tlo1Sy5xJpkWH7Ed2oX73X8FIaiCcIluBZGii6snfF91KC60g
mXE36PUhr5gpJ+4cf5WRknmPNnn7NmR4OZhskrnO+5XPY+ZLLl/Pei8cRGwT8bM+LvWV5PawQeM1
UfUGVsGirI0CXoNBneBkHee5/gx6cwl6M5ocA0F7ioDdcht17sAxSwxAOcijv3da0Lgu1DZZbUFP
73Rg3J6QZrmf620tIm/b1V6k88DK2wC3h51uzoCFEpoF406+asWrTWkVKusUlKInyboZIbh+0ZGG
nirrILOUGWDoJT9Uncdn5JpxlRe1VlmZxECXmwe43qGesa0zgRyD/anhYB0Otf3CP8WJtGbWbSdU
4wpGLPi0OycI4sizFVqzPEqseC5Y8TKBeNO+lAUl9XvH+WhA9s0rcvDwiHdzJfHbvXUck7kA60dJ
ilzNpiZSDPbPXIO7mJWRso6F3Z84XVyjdJmB4OvJuOWmPEcaTBmGXf4zl3lxTEgt5i6nWPGfON8h
4WE1JxH76/AmOFfrpjwZOuiECvBSaeUlvHjRKhsTHMClZnjqk/gKcD2aD2qcTaqiZSov61ZIyF/f
qhrbQKoLb/rtQ8rpggew4x2zJMDtd6kSiSODvPx0bb9LeVrCjMgYFLK069q1o9DQArc2G1uyQL9k
fB9s22WqQORldDfHX9W1PCbKzZSiSdHvoxy1xLtkG6kyBMumU2LlVgjXw8pwkNRNd/p4fIJhYUsP
L7V/e2qTIPiY20zoZl00TPs3NgFWp76vgCtPm8shzTyWURFXcO0DajUCwKu+brhQuqBmz7MoLnxX
zSdEBDwmYEUfXWE723vYA30I55yxNa20R5Z/UlL10Pvp5x5uO6t+yF+wbbPEaSM4+ng02+vnqDh+
3bPbOJa6btbedMcU+lkmGPlAzYmFHycPuWgbAbA7SLHpi4PE8LGDXhoQTw/NneBlUXlGXHbM5AU2
Q8DIcBSkU0gK4nllKYPzU4Id28fLUQnmg2bkiy/r56B0R5HI69iFCTnYfcUkEfu1oDsNs/t0oau5
AfK5wYurnobxGPbd/VREy7wvmGkYVBz8STWgdt6VF0DbXGt1UbTaQaWMuukpqVmahQDwk3TJfSq/
xg9DZ3EQ0mb0yaxrwQic+oj0A6bOrQ7/neCM7MTg86IBndY9PGWcpjBqUmRi14c8cumdr6iiQec1
D0Xr9QOOLHtOT9Ksqsw1pYqHF0cuELBAu+TLoTAdn/4gF34g96pQgY5npXjHrnKY9xigNfBxFZPJ
KMKgKi+eQ60S/RoDHV8zQUTTdCwVEh8pzLHGYf+TZMxvkY07E5yMMygR/VKDzWObryjHT4behhCT
o74f8SZ+LJ6eqaKvx0PW6eSAGUBd+xDQqpuNSoCzde7u5YcRAd0wnOal5tn3ptdgSH1UCq4Ajuaf
JS9um6fG22uIWEmHHnhrYKdnRpbPsYs1d+HlqNDt1+JnGGOPcXaGQrGNpK1oHrMLLTg3zMjmk0tf
ARpfHtDme/gVzY2E44LiimEGeba8U2UYQ/3DFb5ZvzMrDIsqH04lRB2a3cDlewvJnzMUqpYWZF/M
/lAMzZSAlVCf9NNSqHMzfIWs0YAbhIW+CxZxPlqn2x2goFbNi/n/0ckilWUoK5BA2hBsqM/8ayYI
K+PtmNMOhc6vjV8pMRDcVXCifHpy4r09647N7yuWTcp/3t5mA3ighvFSBiEHvPvU9PBdrL4E+rho
O6VixpfYllV1cE+wt47xr+Z8E5D1zs3MENSEHM/lIKaw4YwimxO5Gs96AuX1i4rMY44FYBz4VAR9
JfCwbmudPH+rHGcltRAsFac79ytdtVePQeYKLgMV/VyUUqhnHw7PxHtH/09cO/OKYGfGnpanBsyD
ZzncmB1Bg58DfjADh7yyZ13dNKE77suNtLJjLlIt3PFjPCpjhqrIeFFNvVwOzCEo0U7HI91MTWlJ
/EJb2Sj4qTb5oNOfUfybdti7eu5nYEo1VwVbkyYfcNYBPqk7sIQH0o512JymPtvdgZUxWODqeguF
PwUB+XWdpKOmfVFaRcSfSvi8iu3L+QE4thZQakB++vAQI17u8EM3CytKc1NyBpUJB6Z7UJTsMFj8
JDjoEd4tsWQOC7qyJnyxvvzngYLfm4Lp9OlWrKfLLUID+8vLmG1e1SqZKFs/Keci4oXekxLoKX9d
/F1rXoAC2unBgO0pcsx7RlywvGo2Q0MEh6OKF3LlzLvIN8Yk9d5geC3z40L4WJz0b9iwSnT+ljIr
Mf1d0BuIPT7ghaejSBAViHGRrusYXMlIQ9cNHlcf6egzcFg1wnbyScFWJcjz1blmMIuIENLHu9G2
wlMbxM3nMnRDxWFfzF4JR89qHOWr59QfhvuaSXcvpfdSmTkyvFiIDvJD0NumpCGerlc0K0spMGef
Kdm8V5Ng9d8cMCQOTeO+R0xaGHvrSzs9jQPr/UuuKf+9QRlfmMoYJECqT0SbmDrRrXBVzAGtXMpE
IlQXomudQqGjMca17kkXpo+ch99542ZbUS/Mgg9zBkah4dd5rYp0FcicT4LsBh70F2bvxF9STANe
yz+/6RZBtU1+/vvFxOZ5JIrdpwHftz5diCcCK45g9U2lrhqz+MI2lD2QqTk7KFPedWbHNPiPVehj
v1s5Ev4YJLNHBT9S25W/da3BeKs2QJSKxCnSsKnjQEBM4Y0HpNq3Mva6WX64NOBEs/qVzA1I0XXV
98mORNokbIhggVYJvyDqSRjVg37NPehy9CTtut6jlN/cmk/7pNsa1kwIA74Q6+zT/OpOhXBE1jns
THq7PIsv69j7yJnmhTuDF6xfmC1p1yFTOkQFbVTRXqJArnGYONCMv0WywcFeWpsAQ6ITnT28OlVA
+XlU1/Rzhls3OV1WOeezHEZzLgpjlyDF094p0vYMzO+htjdOIcbOfBkQhlmpm0i9Z3ztaMXzdKOV
qfsQqQRY/zKlGpRA8sj2i8pUA8wzDMwt9DXxylBnKcwmi63RdPmJWaOt2+Go/OlZTKaIeR4wkvgW
KuMVEG3fxksdalBIWabBw/xOZreytW7MXWOi/4AJTCWxE7bEY3+nZQrxYrBdM+5EMxw3VYh85GOr
+2neYAWKgDtFyCUgdA282pSOP3o8IOGcBoLLpIIcjhi2nIWh7dcmaEu9tTrBWEVu/2fywQ8YjVLX
PvLsN7jiFothgZMw21r6jsAYMYFb512A3r4rflTja5Z1O062tKwOBwWW2DaEtu+0mdKK9WUrmZog
QgWs3oxi0F7vrCzUauAs4ra1IVjpzzaAwQeYlhRuNk9A2/TOjtGlGudo3gkzxPR+wWKWfU14sn0+
wVhca1hPht5bgeAxNeBzurtVz9BVX/XHqDdjDQgSqmdl1fHlhu4ChTY64wOtgJsK0jJXLuVZfLvq
UgTpz+TU1jqggYLALg+BbwjaDghyrsAgNv/AoSZXTb0zk8HaPQE6DO/4N6jEy+g+adV22lDNOPR9
w7m2H+wyMmD8iHk8gICTBuO0O80jHI8g6WcH5f+nXOX4mkRB311f5RGOYj8EkUAs2dG//E+006Hc
vU22VDDlSNHeu/NWrTHSNiRmLyLAInQJaC3s8wviR8ro3LQrYd6nIsMFTqM/5gEhNm/8/yRB0I58
L7Jnx0lFbY96pJgf/oPPsKdLJuYv1PG777lNe036ry2uwaTWDUwj3ncLSpdm58aL289rvCGzUFf+
G6h4scPsqQ0G/sqvFv4IYqC8hgyLKv8IcgDgs53Y/e/jZRnN/eh7WeW86PJd177ZK+o6XQ8/1WuZ
UbK/jZfW9dVbpWHpRm26YNK4ADFHvUOvSbL4OjuzGUPmY7Nigfir4jghO5bSG/N/n2plmUC2mSpX
GTSxkrq0S0XC69GHf6BOcdrY/nTm7Fcn4SIDJS6xJisw+UwjB3wwWURJguPr4CDSwdH96WOQ1Imo
4PgxLl1+vCjyyDX/ZK1ouXlr7VYkaccBUtVulZglVneLc7h3Q6S/rUWUBfh8sR0D/sX1Cn9B7lOJ
cbuT4G7eUlCgqvZ9MHWPE3mxLVJoAon89Y0Rmqz4voGvYaevjMOT9S2MsskQvoInfuX+sW6T6qhJ
v3Npe/cOk6OgnfmcWwRimX0C4ylVkAQhsyjxDqYLKpnpf2MSD9rPhk88uyWhGlSxKnLTBicVBB1S
m7O+gbVTAv11wKOIAQ3xS99iHX6vgE/MPIMByg/Sbj8iqThHK0fGcCEcqISXjbw0jDB6Cw8FJ02i
DgAWDkywsAtNaGJF/SxNSW6fTOUmm6QHn1e3X49HX/j0a6Ro/j1rMbgyHV2eHnPEF+dAsm4ZvWsi
bV1q81gqk1pSwYVwMSS6WaxMAnhkN/CTsXhmuoAe46183wZfjRF3EE8wCaR4zQyjxyIaNBcgoA3V
EeLQaSGlBf9X71kphSNUMTtiPW0f7c/e31xBRxqCN1yJxoW1751Y2oShH5Eqr13D5Gu/Uc/JlNTM
SvIFDB6XtYUF4iyNZKpMa0xHabLFQ/LKm0N/jYC1kN1nowoh+iJ/FpWzD+gmFIcrx2o6p6hZKcP+
1x24iI5/jBT/0XRe54J9a5cZMT1l0mQ3JiJVzCEWxYr9f4loloPRA3L+6iJB3oXoPrbj/0904rww
fD4TkfwF0JdwIC1I1axnr9sXv6H0XzEVeZ3SjfSLxxh2ULavq4ZipeBEUDskdKldUJJPVT33X8bY
uEtSwFp95dhwoWxgXJOIZDr8jafQ6TDTswSBx8cy9+kIbmwRgWPXdx/GaYIUEiH77Ofad7BylEOm
f/9IhHLLW9ay7OXFRXgKKlIHKeHTCeRvkTcVyN2UHrYnSH+O3hYW8fzoM4wXpgkKjWklBTYiGI4t
wCn0s9ZoiVXSdYzA03MIevWsCgSNZS5vvR12DmxS/aWEAvlbgYqaXucrkNymqRqqSwZMFPtGp4o3
aBFRxprl2WnJCPKt8m6vKtJ8zJTGbgHOv2w2CZUIVL+B9n8xppHzpy4c94pEHo2U0JNS3ik9fmLg
rYABfaefRqa2CJC7LPnQELSOCFlV2v3oqO0OEDhgyIf4RRchaogv8wYUewII/ADl9y5gSwyD54R8
uELSmEidbi5qDjbWjH+iQurhC28pH1xyND1K0K1RuRLD1mIBgjcWPRyDAYuySLWTTsjvoBPJ97tZ
CEU/OIHnoQOTmMknVGGt7SomZlO/O/3k836v3iwIXODXYGmnHWL8uqVMbg4xvW3EQDdU2lKPuDos
oAWUanp2D/+SgxyOh/NaZ2dV94p3aOASsMxPLz6jekTr3iw28ZkHZ7eMS+xdilujQGTaZ5TzTtn4
W0QzBS3IiWYOIHg+LIKPv830z1asaRRHNYDckAfTpPFgV0t3+qHeITKkR1EUdrYxKR3ryYuXxnpW
9pKklPq9jXL+Lzt9uhnxo+1gicUeAEEnrgQFrd87hg7uqHrKx1wbRevX/iidFxnNw2EUXHkt9RyZ
ysakk4RX9ZKIelZlbG8x7olAlof9itSKowP1QuKecJsjA9mnnyie8IufxcVDcdjgu3b2Xw4q2lF6
Ge3oYbg1zwQMWjst/myhPDhJ5NbGS24C0RCiEyry+GqF2JtteEPQ3tWXJTG9ITEbkLD/bDPxNjjQ
48C4FPA+lHvA+aXdgzgLhdbTksdZ5DabbX9X3NZDU1P79D4m9AXW/VrNEktvguioceBuY5MzLEQn
HMkXISGIPaf2UkLfHoylSrgvNQOdhzid8fmY8Wu8QGVE5+TbOyQ3lSMrhw/ATZvwjl2FVBwX8O8z
I0th40tj/UsJAkhkCTXCEMWLZg5FuuGvvLxIpRnit0wF1ZVfpUV4q/TFkIViYgoFv9ehkTbkI7xm
w3tkHoMkU9QVKoTIR13PkrK6mnmMwSN0TRHI0EQwVvCQ3zL4+2kJl370PKGwpWr/cHVGkDPIzYl0
oqFGHOJqlkW1AqNJ9E2Hm5w40TSt3EjEtu9pEq8hu1DWYtLIpqBP0fAEMGXxEskctKNocD/cArpn
y1N19fm/Ty6gg04JiApAX8XufuovOZcfbNt1RlHG4gqw9zn71UuBVloO5FJftowr2vwqdetA9D/8
T53iPZQgvo4J3kBflj3prWUcHzJlyDe3ugqKch2mKG0nxD683hP0/xmYFSfKZo5uGA6hgxsLHsNZ
zzKK11+FkhrlYxvOhcOSKUSK8KV0vr12q7hoUmG8m/4vM+E0dlCMHni50yG+el6ninbgDAjZWq51
ApqkAcyqR89U9pkDPb549e2VfLeWmQ809DMXjvvIU3iGj/c29f6rp0rL/QT9QBESW6YsIxG0nxU+
MwQ2D9nV+eH9Nl03uSStwQDG4EQaOdceqbVYoswA0b3wgVRD9QZR8JcAN8hOpOjwUxaBnw5yIrlN
INZhBf18TKehcEazCIAHQeuBNx6uo5gatO7uwQtmczN6gfsgLHSbVxNHl/6VN89tz3BONsmyUpyb
qjahsX4lTRKUFgyyGvcEOqQoIUcT851HOrBffUI4Xph+cFNKQzMMJr3gpixCEZQAxBt0uHU8qUAo
zfHcSIf0BnRE2dnSd44aTEyx9ANWmUnR4+mwbK2d3XWRM1KOiFrYoNya5gklaYX4/SFGuCr0w/bp
ApOxMRlUhTtp+ve342uFpsk4EzqytNcFDZ15GK17FeF2nbYuMVfFHJVC85/iNT2RxTkVq8Lk9zR4
IdncIXu0N6MTMVJEKaONqe8GsSvo/Z+wYP5w3MSfgCx+9JfnZ9GHekwtF8LGEGmZrDWwd/pjqHd1
O7Tu0NRBglkzHAL6qDhcNLZHxO5RqzGZTgaNicglQAgrSLhxWqw1cDZ3WDa3YWvApFZSGsWL4m62
SvwdrcDL/F9jzDnX1U28ZofcCn/7WMUqK8bLQRyij5S+c/lw/liqlOI52CS4QMD+wsl1qDBy4eem
PlL4DkSpyLoCEChZu0iBuyDViFH4nlM9vtzG2YZ1qpta6xhTxqGrhQ3+pqbOdLtAcHp+YDeKmg0h
VYFnMxYnDMzXtkaOb3Bh+2OZhXgMSdyifPHecNQWgMPQB3Sb4up5yvn6GdHB7EWwSxjwPB3MwtSY
03iHLa5sMerCqilrvfbJUcq1VoiwRKbnGnG15qaoL+C5QCONRi9JFGoQlFmRNHt90AunyWEzdvNu
FVJ1hyhH2gK+7V8Z/Upemh1lGSnByS5XPb2WpD/DytF5Ac0i0rdoRVeB305ro0cDwGZTu+yAy/rF
81NnIV39GTqSDQTX70xub1NDACGZlfBaSyqPEVp9/C2cSnnogULrCq9dZH3IfpwoSG/nSMhcG6Dq
VJ8bBQFwaYYNaaPMgCaz7Cb2I98Iy/Bu14kYdAAsZ+QiiV4mQtFBrrVpnx3g/FBN716pmjzynHjj
ohqkPGCxN2xutJxga2pfG12jpqrwiJoNDmfd4NHTfllFNky8DBcMq/kz3JzkvFx7JYCWsmWChCWe
hspS8eMAaVYpWIaF82UILYjei8wjzVdXiV8BCDwsUxX2/ETxZJsFa+lLuOzkUlSyCCifnIXrIISg
Ig8wWulUeKzftnDgzec9Q6EvAAAYFS7FtFM6J3WEm1LRUkMvla5M/IVpRnsg2Umz5J9qsf04+2P1
Gp6Rkc/WpWuv9PAcPCcEUgVKQdqcsDDyR5MESCesz8Q+TPzSQLWewOkeKgOqcsrtB5f1R0PnRwiV
tNifsl5crC1Uhk8eiKvL+Cg4lU+aDLGgJ9P6lnTd2Mh/pMGy02bqK348fugeACt9pUJjgoi85vJa
+U9vuWYe216xPh8WOHmpiFfW6Ey5jEs7+E/1AM4+pHFZly1tCOxCOoKhUqYyPalEv5DZvwPxPA2g
nYQTTTisM798iYcihrA2wls9StwUFiDUF2K3jwvlxgG8/jcvU7dJzIP6hPqVbZPzF48PnzTAy20l
wzY4s+EVs20KblAN6Kw/lCBko0rhuQCap4MepcCcGEmDBuooPEnASC+X3ysbeMDPCnj6Y0RSDwS7
C+bBxSWqs6Zb3+Qqew+D/p1QXvNn+a+YMQd9jheDGthj/eTi7j3mfQV8ANO1HY9mw81Y1L64WTb/
a61WH6lZjauV+VF/i2hHt36Bw7kDGNQQbzFeY/0U130H3ZmqKwVwEPFZmbox3DYnzsck5X+BhAYf
8HO23aQ8++fn/vlPOtEIQeT6K46hGSLqhrQ99xNixBA6J+kfjWjC2tGsuDmg/ptR0PgAYdBLa+8q
Xw4/xm8JImdKZgzMFUNV13bdLdv/ZWoVRAs2i7bv733dKncHNmHqYeX5NTxgBF+EIWIopBTxks4R
WKt0+FhVkxE51HZO85Slq8S9j3WlC9KT7iAOIWubBVONa6zSuem8ZD0HW6z0Kx4b5RVXg7pAhRZH
6iZ82PhwufIhZYTHOivbzGH8H2ohZTFAMemgO3kumlWYGeeWfm4/8hAL3y3zBu3RK2DbzXwksurB
yWLgkrNh+FRBPrXXPcRsEfVEdkQuirDbk0ZsbwcIAuwHLjzbFBD0iqcij+pWuVKHieN7gttWCu03
G3+ZEYKWrjLpjFswqsV0DEN2549dlrIRYJTEHn8Lr1916n4YTqABFGkOfz9T61uAupDdM2amHvPx
iVfijV8mMtH9ZAUeNGVdCT9U24axmnC3AbcLB8UGvMb2nwJZKdJLFTQO/EHYAfNy/xq31TL2eZWu
Dyx1PRExlk5oEuAjkl8fpF6WWj9YvmlEAkNtzaUuTv9rYqqhOvq/kPXbuGSIzb0SW8kM0sCJw61H
kO80l6NC7wRMEarum+MB+Fl9U7K54rl1kNvltRpazqnf3grwaIXl/OQtlF+Zspy/1z6c5OeHOiFn
GAiD2UyjOE+CV2Vz/vPQv6aazz7XT7OD4GHV4VpPXDiVZmdC8u218GAShz7qQiGbds2Cr61rK0Mt
c2J8Y/0w5bdzc1SYFQOFr1n1FksSNhSWl0uD7LbTqNJloF7lFMwlGajDm/YUKt8QK6BiF4TXuNox
jdqHXHeCK8Ni5Z0836V4uP3mDjZqLG1g9QtbHLkj/qxhYLfNZ41ztYnFc8g8oe6qaa5V95ixkFuV
V1xjdtK28/7fWEk0cwVpAF5HBtbVXwlkNEn8dMdwO8B9eRpjzdj708OZQsnXllTAjBtIketqeTCu
/nh+5kwKKVK1sw0EVSPW8JwBC5Dz1sH3dCM7Y/o1+GIkRrcWLb/tKJIgOyNbLjTCbGXelliuIq6f
Gs8ul0gs5wdnEpevPww+qSvaci9WiawEILUrXks2oMZJXQg7nQbZG1KWe1nHT+Kw5aiQ+RjyfyFq
Hss7eD5zMxltHmIcWgHKIXO9bqeqv8PvJHfDWmgAjWhNEgN/8QD5SmmqokSsRgb9xBbxDOp58MN8
e5aHDHMFIyEty0ZTzgIEFoBMh4JfBAXR1ItTuznmvw2hAv7TcJIb1Gw56PS0yBqU26+NmC/6PKpF
ygiBhFhgLZsyqCieaOSpkabYg6R8d+VTb0Rxpe/IGhtNNVRF44Rlv2asAcw8ElLCIGqBYgch0i4n
x40PMqtD8bCyFKuy7YB6EqD2wMofpTUdNWvtOvOc9YOk1P+hcAHNwd6I/jrCxW+a5SjMWlzGxvwK
n8CKEryhgMWne01O1M8bYSe830EiVsGoitX+OQCCRe1O4YYlHmmJq9nZg/pmVEFTgdoOOdogzi/O
7HpZeBQQoWCpBmCpRPgCpGLRnlayMcGJGudHSAGeb/Z4BN/CapC6yQzqO7hwW6ob33iBmHZoNXyb
Il3jWdUDQE5ZwQ97KABEIuIUuDndHW+nn5B85ZtNSBhEmUxT9p7y3CMV9dsUDJThNrAUBf59y41s
463r93EFrwUx+eDIq7BqjNiAM8lXjIwoQ/4ARMAGRStK4aDXedGUV/b5NDN2zMr2O6ahIKaVrY/D
DVcEYfW0THjgvkIEtdAMN4KBx7rLyY85o4JHRct0e/BHP352GBS2ESXrh2pgXLiemuaSJY2Nfb0+
5pexNrUnpVtpdfvw/UB8b2tIYKUw3hxTzZ6LbH0vm0FnZmjLkaURSukp1OCh55CppbcCHzt2Njgo
t8+jWdPtdHzZ5+gHvNRSbI01LA7h/8+jxN4zOO1jaAWf8bjqrxJTjr2Ga7nvHtzowP6ptrpymtXT
AOsQgpOuwwLE6KtMTzjprxYhm2W4lUHNh3LcU0HRcGSvYEq3Cqbfyql1XAuYegsPEQzpn1LPIo+M
8ivax9MRw3FSlsC61cMlj0QSPxfnkYf95b6HXMiqDC38anu1FBrAkIsWs6jHGLkGC/X6SIzyBdh4
24kBfv64+Aw+rnn1fopW0eQDTKdhs/IK7oiepVgG8eLA415FRL9FUbRMUSb4ZLp91LHO4QCbZAk3
dN1ELa+QLMmTaY7+84L5xcT4VxT9burjeGH7843H341VbKEDpXIU/QJ782eq/jvc57gD+2MAGGjO
sKc3iiX1mfgFVKC2pq4CHhN4axGuVMV1xKbbDDbeRw3m131vpSOFOigt/phGqllVHzA0R4+D2WW2
EgIe7kayRWsCnN0iVGNlm8ql+1DgwHb7svKdsNUId9UMHjeaRLKL3C4VhkhSbGfPEE2lyuJleB/x
loA+rq8nvd1ZxLUmHHn8SPm7cL9E3gAbioqcIrfvUShiBreSZodPj4XQSkMGI76t3eDEhBsyiUtG
V8akjMrJdlcjLGe0H6QushC0795eFrCRQYgXwyIUriIJzDjlvWzWpQ8V1mg7458tRLk18fQjRKBL
EB5ch8zLd3mpdauCRQJi1wd9V+Z72SyYQJe3BPrUxH1Mpshuv59fRcRATKBZtAC3cXpO8E8/56X2
8UnIPinOlutFwaGr+B+fNQi13PVBcEqEYFlJdzKbYkOrph6pkybNavgvLPxPuEtBlaLjGPH1v+g8
purme4lOpUzAS4+gGaoeC3evkvrlVKRlHPIChAq3HvziRlmE8aaT3Bri4QyKuDiRX/OYJFWayjWY
6/EhuXp+GcuCFEzqOIS2rks3aa//ym7ChuXpEpUSg7GPiZctlE6v8Av8WWY9dByA7WzVESPHU387
y4OEF7vw5+PG8GA44j79jfyuOsjIdX3/j/OeiNzWyBrFneiaCSbyn/ok7sJTld/4Mk9fnD48iyHG
Sd+7BL+jCAXckSFK9L3EYbbs8ht7ERKj7BEnvsIO1Di0o0UYRw69lSZOTzcLR+28DRysJaz4Ont9
TjLtFq8ki0kzqzzL8d9unvkdbreKuM6fOHowh+5WhHmx5D5JDjLCUSJk6VOSGywt+DE9iqvjjm+G
WKmdNWeIQ+lB01H7N7miUcI5RhRynT6t3JPlobfmfzDdS6053D+FefcHa3bPEGaonOp1R9xtqtII
K9vfSecMB9vbd897HSRvX1HbCMG/MhZZR7unXy2/M5L5+mg0afuFvSLHfADl7skorFOZ30W1xdFq
HD5Bxgxpw4h6mdDOT/fZdCdmKbnsjUuhLIBHXyHQ/+Hz4I0G6lemcbm7s/3L6GTM3WBn8SkwF4Pf
DYDQtjcatVEx94tZya/D0GFfgb96CMws8kxrLZCBjpsWMBamGkNDQxLi0ELRSgPQf3P2Pf5Nz5Q4
+83AsaBoKblVHG8EQ++QKnzR0JMwmPgcElwPyP6DiRo2T+O834AncTqMjpKYcolXnPjEdWzFJlmR
EcWEf97YemDrOqYzkv1MSWtHFEvqhzR/HS3xQODTSezqPuD8AqDDO0pvJOnFyvUnt3DnGQiaGJeQ
GUyCciYsSibBFhDUKd9zyDgOgRARZGJDWWc+nJ1N0J1oXwdNYd1M2X+VI4o4rMyIajUxaceOfiE0
q/Y757Zry6+8bmsAtBVESPbsi4twlK3op7S26LDaI0hLd//RXFfEyhzBwSqUinjLP7PagVLWg9ji
fH+H55My2Tn6jMs++kQHzvM0DUXkdblYYcNdCNj1Kr+NGc1mJe95bhRaDqZ0rr14KCAMOaASHsU0
Ne4ilOiOBlJtCmYeHmPl/tX7ZAwdlbXgEaKH3yhLiyi0nKLWmIHdsHO/OOQepeLeMXQwtMqfDqwx
dw1BvDpfaSZc/vhwg4wSVGRgomj4eUMJheDpUbK7ttiu1vdS/R60wtw0mt7kx/YGTEsbaVWPPI7j
yNMRL1Mu/4gVeIDsG+LLwN+WZ7D2RKejxX8fwnKNRmSRC15GRyCJAldmx54JxjYIGS8ly2L8AXCI
VYVHAYbp9f16w+FgnJY6a3N9YwbCq/A7MR6eiiF8ckQeTjd03uvPRKn2K92rR3LpwwAFyENZohMS
ndzx6j6zWnozNUWsf2fmen9txo0zJBkrRFp4QDRJO3/xmgxFRWAC0EIdYlD5nvcbEYhI18CITyyk
m7HZgBI5PJMNVdaM2tngQ/BMPSA4H7j7FAELTPhmQ1f3QaVJaxYH2pWm+Pz5nJAnt/va+uE9djTt
QnB1cbhP0c1fs4t7gGktDNkahDqtqA+iwL5MyMkmjm6DmBMQzKr5SrrR4bOWS+XFU8aWHI1V2J6j
oHM/a/U8vPsiW8PZEEeBR0d+g99d6S164xXaFqzbygiClcB6YVddCp1aWvDu5CGNRJ135M+isXxB
8VON0hBHGWReOMv/0qHHIE8StqleFgNhKgwQ+7DRRABzQJSQZy0H2fbSA9nfEEVIF2gyhWbPbxEz
P2awCsseRMtPUKYKtCaV5icpNGB6u6oYhz9y/151f4ZMYcfcBnykP+Jsj2O5ivgHSxFfJ0inLePr
V7OAxoD6vaOPLEycZ5edv4Nl8/NPq2EjZkhe9Wv3/Sb4lgjiTo8SSHEWVJrJNGElIcdks9tctF4g
9waqYxdm0psgv2lj1zbrhYkGOKr4PSOe1O9LxK2jhNt5nVlCQ29V/BH/MAAmMT2T7kD5gY0Hvh58
ai0oBnrsHfWPhmC12HRcBrEnHaXhMdcL98inKFLMg5IRMNnyYgY2B2Ae3VADwKfpzI6kAJjbi+3/
eo0JN/Wwv8LQwwNaiMQcemQ46K1pgS5Vxgf68Arg5TB61k03hSyQpGUoOAYBUreFw3e1dD2+aIci
2bNgGObjy6kRJFuoeyVgjXJh2Aa8eQx6EtLNfcXSzfYPQn+8gjbn/IiqxTwl3uciBbq0V86fFSTC
OT5DSXu9J1Vqc+rlJPde91xbg/D0BAI/WqLuxjj/CoOXsWy4/qDGEhARhVWsL/e2QKftCzdrb6VM
q9RcYqoscYbDGV0OAQKLXYcSvrBC14iJrXw6UCDVlRLDDKVC63EwtOALiWb6iwNj7kJeteVnaJ9q
4nhy2fy1yySmaMD/Xczy8WQFQgXl/UphRvAZ1cYlsmkNqk+OmtzHZ/3CY0qUb9EmiU8XFCVcZZxD
ubvxI0jfluKa0TVkwaj5p1+uXemsyZQLjpZpATkrsv1Dgxfda98xMAISxjPMerHmPR/Sp3MTWZ5y
EExNP4sZ/jAPVfvlmry4/EtGIyrkElJYoKTBIs90fmwXFfyjQsG5tZ2F1EhmRpcY8puFPGnRJjbm
18ftXH5ke6kM6YlRSRbbLeaODxKNskX7UUdwwAGFUXbkRAmM/qnJg2w7L6RK/HVyPCsyuw54qRwy
CLdtN6tUlggrYdkcuwgflZmKtbdS/Pn/OioGAKMUwH3V6fkIsRs7Nhw988UqTKcxXeTyDMcHNJML
2ihU8ZhtbPKs/9Nx65IZ6QzkztNw8HfSjI1D3ckBLdEtpN+D6aonim0tHQS9jDd5Gkizy5R7I4pN
1L5hthGwCSKgNR1squdt/HOSaw1xof0mOdU300RgrORwLmZhWzeoSpv33NdeENW0uEMFxW9aGotJ
Y2TkoMNeJDOqgAGAFTmQIz6IKI8dSBrLBAtOMlBtc7ajT64FBDZv8BNJtzew3F4banNncK/46bb6
TwW0clUNF8F12quaFRSti4qDS9toxufARsbaOLlOY3x21oHWjJ9BOnvF/jakrHXyvIrTAkRggik5
HxpWTNaj96w8wfQtvVW6NGlPl2ssqrTK1/wOqLsfeTeIGVZJGAhCSeZ4EHIrFIBHusyEykdo6cx+
07hvgsnNlk8nOxxE84qkraUel8ZMSnjeUJDZc69gE3emtW0Z7n1br03GqLUmHmHHasE3pjxez4xE
GpmPEcnU1cYZLGAB/JbIylVPCF2D+pAt3m19M0VogG+LH4Is3YXum41oE9TrNaDnIarPfIIeuRC7
XrKudZ3Bgl1LrGpKUVtIjRl1VGF8OVaSsvMEkoFp+DLyNK4ASucJfKkaAIwnIpd2ZPiuamEGDQ4S
nVWOs/DWIOBpz3UqPJyQUD5i/88k/m7TvkOWe//92pnNtZ5v1YUUAGMMmIv7V8NtTM5LvwcRkiQ5
npbBlYLZ8Lq1pmhMRD+aZd2aFyNMm5CDc+JG+iAFxmnEBOLQrWdnO6uQZlsI0qiADopVo1M3kqp1
odCwUULAiCd5ZpKkae+O/VFzQ3zCxEfZtlVdiaTlr9P6KIsnYmy+WDtvEaBHSqmQv77wjucE9vFb
EgsbfB1umY4Mo+MEs0r1rBCG7m8hFt4H8zzWi5tqKOhxYOyQ0y/fLwihr6TRnsNJ9XG2WL2C0FS9
Cr1xR0HVpschhKCOzFZFxmacXS7fHEvZO/SPSFFqpne+oONaAapk1hpe6Nvo9kF/uJz+Zwshex4T
m5bQOX2BHrpCE8h9XgnWbOWuBDEC7NRZshkhWvx4Pec+NaXBjS4MaPIMjLbXISHV98EX3Q4uY2kH
QfEUu5KbkH0WeZ8yIR4Fg/Bsp8O2PenWglIRAM5b7y8g89ZZQayL8Gz9fCjZceSlVZISF8GZQSkY
EovMj0JElEicIaQxmwsVqt99kGfljyrHed5U/IDdFx2V1f1kCwv8aOP5kkLMSjtsXrMKOoBe4DDe
svyCFVnPW02wBw0sDZkFgDLNwpuA4pJwRGLckKD69ASgsvC4z8tbwT7m/XEBrv4a1Fzm5wVgsVfL
qJEMogNFCYnYYt2t/R/0sFV5LtfdlJgkCqLPNL3uWwg8hl2yUiv/B6A8ifHkX5kbjlPBP92esgU9
tPgSeD/g9KsvQ1TPOCkdPEweG9Us2qV4k+mhpuKH0uOPma8mrYTYohXGqHGS+t7tdGIHQXUQ77Bi
5EnGQkNSPfPPal/RM7q4q+Agl5L8Vw1Ps+0HPDrHTQWSgCMlA4x+6/0tvsFHZ2nCqeh1pEBHay+3
zuyHAfgsUMKINGpcZSunTydO2YjbRnqd+WH6O70cDUUiJ/06abgWc+7DKvQNF/2wE0W31WIkUeGF
7+SiYgZVb5yQj7euY6cqCxW5ileYbnPigfcsbG4+4W5EhXQ1ZQDeoODrPrrTsKXEgkOn5aTweEf3
JX0a2vgripT1lmjJmMHLJ1tD8WFtCZ2fsk1cYyVC8ZVWZSBeDuqxRwmYt9TBRVsQeJ2Jcw2Zab5r
Yux/5Fr+uwpG29vAloYIiDDdknhc6umenYt/bHZQjiKvot9WLAhnELM5jw7zo3ubTSdTU5Lbg/w5
6cPgqCMskQqYvxlcKccn1LTu5Y97yke+5I/Gb5IBK5N+nvAQ8fGpnO5viU2j0JxLQL8Hiq6qKGD2
f2XxdVVBPLVV4fP+myl4whE7iaCVuKngKWke1njfID/SS24VYdETt5oDeaZjvKp0+BVNfWG2xwdr
Jion5wtQXnKR3VxeSogOvCbsi6aOhbh06QMNPyxFdm5gwXGr625tOrqYkCBYwH2FJ4gQzPt48kFm
mmPP64cTRufNqPN2J3S/8r/cucZA6M+0dlt6HNhPuFcDfcDiKO+UyAWWdD261EYccMZsQeiwM0ZT
pzp+IO3ompTYuWUDSjGbs6c1V8aQ5OIoIMhjoApgVN0GPA+m9+OT2m3xrHn9bbDCVpa+OxoHzggN
dcNd03HvfI629KKqPIcNxXOQB0hYezzj++2W1Vk2+9pc+/hVG+DZK3EQYDTXIZN0gDx3PTNv5dCC
7IsSeHPoVZl0tTrCwkjJHX8A48hMxIXGO6p/GEa73GxFsdM0zmW0s22oQPMQxNdnman6n2hiiWzN
FIQZgBcvK1/HsUJ0lmQCPtlwj1pYuB+zHr0pnejpVwNIYWhCmf28WoZkWz83STnGfmzbYcBfipYa
/aNAjK2fFQDhKxCvvG7RZ4ttMxyfboKPb7TW20HlO1UGQgwq5R+yXhRTlcP0iX0xbXSq8R0B2yd4
k/ahHokBIuKMOhCxzjTo3e3De1iz6vCLqca/cp2G3rRxdp1m1akn4G6GJNNaznJsoj2DSTgZBmuN
NUzkhH2HyF2A0j9LNaxOxmMckD95ngc5qfn7MWVrlgPUOMr+x9kXZnGbNO/QDsyqSkPSmRRSnf+Y
hnBfZfR3ijgRxltdiYbUG0LazYzGua0TbVn5QIRyNS1Bn6MxMGl3+s91tXiwlDJELN9804GlgF7G
6VbNtbbzquA3P6v2KqKU0Zv7qZNtQOgx/TiAmEf1qp4B6kQDaOWyNmIwncENDudewE+Fe+Nxp8z4
msw+teGV/inauDMPaxtTxyJn2Nu9TR4K6/todqL9FcvdoIdMFs1YiXujfTENCFlBfhI16KSBEP9F
8RwGIMMqWmXG2P0c3n4mIc2NzXV7b23u289W+pQH3StM607dSc78QPYpBGtk4sAQV0gzaxJATthk
jPwYH9aFr5igUNeq2iAmta1hdfAqmsNxkNnmPfsQPdjmdOlLpLqyRYXqm5HjfmSK09GofDvzJBnZ
G3nPMZghqtCOA04ZCp1+bpxYkOTpE0WaPVAsmaITUYY9ruxgb2JDPh/Xyh1YaUKeODgVaqdZ1NFi
UUmBjUK5gkGRcZbaz1WP84aG6KCxkOIJ6NJ7iDBlhL62TlcqPRVU7ln0pVqjx1F/X+qQAhuKQDzT
mkRleBkG9nCPcGRUtINA9G3K3VHMyUBRRfL0CwQv5xYZiexyuWQ5QLt/ZIOT1Vt6sHvE/RMnqhwD
ftJ9l7DaX4J+hVigvW6eQm5ncvh+8aK5SdvdlBz3BVQSad2AmMEtk7dQ4hGsg8soXAHXFUKDUnh4
B8AAToNw52PN7oAre/k2GFCcM2oK1/p8Vw7HYauuaRQP7rZmcQTKGVimZmRvmR6lnggHIPqiyaWr
84WDlFU4KWs+CCYgnP14j5YbedovOKqA1yZFrgvfRrgiDZblzIWb/W5PFPAeUFWAY+OHbSEKGQRp
1DS3mBtG0mVS5UH+2dAhAK3l1BdXK7JNtDI54xqU5cgwnqmmogZDfX3wVJ5IkSuT310FhSmOfzVP
ftS7cm2VSFh4KgBD+ZmC+2PvQ1qF2qqsPbSuOLjNN877JWmXzwM283XcYSPzozaDu5/huzibeZ7p
wZ4laB6yUgpZQsyDacsMM09UeQpozqvGoA4KNk/YVzFf2VG4IvQ5NnIs/OdjoShFOA22hIexsYik
777cck/DbRH8LjAJxDYaSDisW4QJdp+obMVZhQBTwEx4vhPIT00aQln+eEu+VA0G8ep8jfXMAlEc
RFy2XvrQwaCuJWU/Yrh5hJTGXR2x5PoZCacNXQWOv+xDuiRiCY/WWlOsFrvqXXmvrXwjWhX1raq8
ygIC0ad4YCUxSDyMA1xjmuFT3tRVB8Z/29bt9CxipIXWj0QzRZe55jKgAHYRxw4uJuzIwlAbTGAD
KCo2XRHbilhyD98vZLBKGVLZphMl0cc6BIcxpSzo27xwjkD1D5nsT4DvVRNqwKy74KQSAP7MUDmX
mKWOT3s25JqRr0ZciZXg7Z4WIDreVWbepXGkyU5EJy+vQwpe+cnxHX9KldJPchsKb84FAUpSzFSP
qlm8TzgDdCD0a+THhK8m/Q4zDS7UDGc+W/S/b6PaJoVD/0FAJAoBjBuoo+zrbVeqUrjkYe3DMtRc
251lfvdpORBox//ydfmmKmTOB/Gu0EJ544xkqsvhZhM9ToeN8bxNsd8c8HR92OEIY3CpJ6MZkp42
a5c+asm+1NRbxXL0f6J9g6FHnNXE97d8isLvG2Tl8KzEkTMInXklOcVka+j4G+VD6uy0K2hvhJS5
6YEejkWf0Ck0XTVnVofwx+ONO3q5Sj79vw4EJwmbrXqP5f3tBI58TZPr1x7YoWR1kgvQuN3j7Veu
jICZDZojPswEDWMaBPgSsQkZMKLqWpX+mNsJ/avjo5JphZcfA4ZM5/K9jXFH//RC9FcMp9+255EV
TuqTXYvMO480nKjOnk79G1nyLV09n2f9eeU9uKLxutV4z0RSDIi7Xn+1AkK9kKR6vauxffQPnHkK
dYQAqWItpHMmgSmA9idkecSWl3ReIE9CO9VE9OQaAaMqW67XKgeaIJNj1pqMa4DcQV7uPfGLJTm7
lmcHyxguARJiqXzvDL7GdOcMrRnupanV13XL7coN2mr40X6gyURwUZh2DKQ10em/lTntrFJV5Fak
zSYEGNPbdOZl0eAmNVgiNcH+AI0fkhGl1JO8s6tttIYy3ddmFEqg7QDkeDP5vfFJm9LbnkW46VAM
g9XZzdRkBuDJtpnQEFzxWgHTPSP+FH0lN26I20tufH0n/pX991I0l77O1Pd5Ht49z6Hfl+Md5g+1
l8QijxPO2ecePofStECjACiuOK+zDKr4TKVW67vRia2Ttmict7TEweaSn7gEId7eEcjGGLqo6EMQ
9hthszsTLCFUVj+QsGovb2kNlyJBBCxXowlCfswh1AjxL59CHr1K+4gbMZj2gN5wZJE3IA8obOL7
S8bDH0jHoeC2gOOwVEPwdy1WGAIuANEeCCtJyGb1Rs6fqBmnutOTgNxtLArU7et5YQwRRvfwhOfq
L+r0v2Ot/LIooEUR5gvK/5zWX8bQfbI4Oo62m154ZiIo/RgEPQzTMcxL/WhV/k5WkAuvVTG0nGcl
f/SHAVvRx2F8COoUDVUpeSLZIO+FsoFJlj8v50oIJrnWOHbkwl3UGeTQKKeVGp728Yz7KL5kDiCM
NoZoGKkidmdtoH4i4RM3dG8424AwuI7HsFY3BtQ1wZxZEF8tsVL2tHhItgt8YIVo+kle2UIPC+Ph
z9CptibU8xqJVmApDXRtQlepOIsklGS9TZoudy8kVcr+8VO4gKKhYA9Q6+9LDdj/fCv1TiToVkSt
G+CBPzGm/1Jr0o6Uu7D2hXBQcx8fBebUa71QVs6++CEGMPaUdbtbiJxrflj52VZlTB7iq4FnGrZx
EOZIzpukOjo0+xl4oxImOXWU7XOBHzII296wC+nic9L6pC4Cp81jqNzw7Y0uHHx895QIT9oVXqOu
gwY/POqGPh1oTczCCMR/aFlN/9ylP8ZL81E4QFY36/eWPKaJeAf35i332BZKK4yE1CtNjUtY2Lvp
Rar/hklw5lJ73Y0BDrI0Qc5UCO+RndvqWF6vAaRAiBY4uLEhqqKWa1pu6Xv2UdRUO5UrQYYj5Rna
oG4Z2/J1SMu2gpd4BzBWtznbjscFygtqotD73+HB6AL58h1EASNZYjTFXj1rbka1f2zNW3mhV0O+
QSUpCjBKefdRL7lNGQn/INfPYrDAqgcbg2OwYflqRRLizBU4GSS2m2fd9NaU1urQAFu+CduRGxBd
zKlxscRliMe52EFf71rBxvmHxpp/sCEJ1wTTSkuS4yajtykV835gpz8fQkxiRgqZ7TWSAjJN4U0B
O/7NBG7OgbTF5zkxiI/7lGoVEvE812eRxkyqTREDoE0hE5OCFPR5bR7lyNx54qIZIYGUctQ1b8g/
REdRlSP1+yUbAPAlAWhZaGoz6cTDmEsYCowF/r5B3XDNkvqJlo+J2Dd1tY9hXz3MUfC4B44ZiWba
F8q9VmqAjhvOONwwRSabgNCCobuBHJ64n8AflyGWV8gjsi1ojrUC0DIrU9qfzaHo8Q1zuKTjhHFx
g9b22T1ls0JNICqLc7HYbCl0++iOW0LW4UvvBI8CyKOjQHrIaPhQc6plmGjBJneqgAbsZbWwM36S
XKtQGSMkgJImSyUwyfFn7l1reCwLCNhXUd1sLSE20C+SN7v51CpX0HBABQurGefOhQ4xpc13nZy5
k8+DuYgSFUhs4vNsQSbc3lBrFO8Wul6oLCEX/MXOM2j1aAtv02uLgPfcnPOyGQZPTuIVXdvW+zLp
AdsYAiZihSzAi0gTdT54W0kKO/vUbf6OuBhuFLVsdXdojnn2Hlxx5qp3QLg1m22PKexBgi38/Y5Q
t3pNMrCqNYtDrx2daCA7gMwebIDky3i7R/m1joTnqdV7CbCKpoP8VyIeu/jE5gi3xCnM/WSdfWEM
6mI0QYHcJ6NrsQ+Glra+wY3IStAhbOK7A6grFuKff9k6vb3TSB+KEYhGvDkpAYeGLkREIvR7L+Ze
Z7LR9sgHSDrgmL5a7WkC69xhZ/imScrM21AzTuGj/49W4gME0K4eyQ4prgNC7TQjqEE7WeTBVASY
4xgjNolh9OsgSxLOcrF4eQVre2m9T3zsxh1C2bojb7E2jo9+LoghYgVSuAUrOedCeAaIN+SmYSpp
nz8Y/yf4vTY3fhuQfkz7AEqsPYX+gRdFVqFMeha32clZHeAbV7oGCPeIdlG2txX0SQDjvboQiqTw
soppY3QOjQ2gKduBBZBcR5ykbzWEwe+Z3Di2k7KmEiQzdHzCB66v3POEMUoHq5kQPsiuX7oJkNUX
79ouSoB87Tfup3wzx+DtrGPErhoVWiI+ROxmFEDgsR0VQjYu4BTUdlAdqfnUri4WX0REB2AzlRZN
xdlPZy/2pR9fO+vH2hlHPqZ92oZD4J5Jc6eXBay7iAFJ5Ivzpb39fdam8VcIf9Z5DxRN4kdHvXvI
Lzxaq2NqhC6XXq9J9XId6dB0VtCbTl9KkOhZMmk2IMfaKKr7B2Vr1hnAvMMw3caNekMZMbu2cPxo
1/rm//4Oj55K6PVX31YUwgxeChZin2vLRkPDOM9MFyLc9gZwm85wGD4rTUhv7K9tYCf7dcJtwmYX
sNu1vR7Ns6X5wvYtq01LV8vqlyyLkli0368yhnwKxgkEEKPcmNuOnomYqSx37HA6tRvISl15rmBQ
9NeBh9qGVjnYkakM+Gimt2fyxRz6xY5RQdKXuDqg8cScmgu8x3KR830FrhrmzaEFNN7QDlSJmujC
eWr1jY/cs/0q3lrPjrKDfCfYd4zhzhHkOPbEHzBy+1C9pStYZ28kZNK7MASsztwgmJem6xVW0fs6
YVVdi6ZBuDZ42A2iWbNb4iNmfD8hyfnS2NaLUC4BflCMjSO8PV3SWQtuj3bAqQCs4f7BrbI7YBCb
1Yan53bIwk8RlFJHgj137g85ypcjeehCd0ugpCKMc/cj5nc2U//pG8TTGaOsil3LOsEtC+Ey/+Xc
yOmZhMghw7vecz3XI0yb4PHEHdb+EDgnpJM3IdCdr6+ZenuZFQZbBDBm2HlwuRrQ6k6lPzYGD9Pm
Cwmg5fhVlgxppaJyHb1n/KUqX1bo9IVd/i4mFWpd6aFZXO+dVj8YfdwXZra16Ig0yfmK3tOFKTxe
g3GA1QtBGxdz7YrZIm90xoJ+17mUWQi1yBtBqMZ/l3+XTiE4/CL4KNaZCJb3l6u3/31IXau7HUjk
Gv4idkp3f0cdsAIsRxbyGKT3pmWRVeWg6IIABIFlECOof8s2JSv1I1JcvlA1zji7j81gWmc+76Z6
QLkDj9cgn9pBBLY5pAp6ox7h7PzMO5ySDgD2LEDDp97fm7Uq6/vDHXkDeO6TZq8NbcKugeZdLDxx
VeX31j+1HhaTtYGqU1Eju4ytHW5c5hrAemf4viwKYz5F0pItnva3/BJPh3X9OjLPW6ZdfYw2R8Ui
D7PDFVW3uP6TQigJOvzqTivDl8cP7ZGZs6L1GLh+Q0gOzk4TP/BvHAIius1xDfsVVX87CodTxA2m
8H3dZscv57ZxINOpupa91bBf6ePJuKkFic08VhLg3I2plBPhucS0VRWpWjnozKfiTkHJB5vf3Q/3
lO5GFRB6Zdc1Dfor1xp/pKzsDgQlHOnLgS25wDIYVridNwIBEclmhtwqK3XJJUOOl3CtDyRmsrtZ
9npVlzFaoSKwDMW5rmVa0TDQ03e9p+WW9EnNRNyu6hSbSUaud48mnapeQiG1F1FRN1ucplGRLDzb
0RHglCrozNM8ahNZuoWuBM0jfN/7MlvgVM1JJjLWqAGXfqPsQFPf/OSjQ7HMUben5bnv4zz7B2Hb
CzzQtXuVBjcMtcdStBvDWsSB54NYrB5qMRqmYKSWcynZMz1qPenLqCm4fUWj4dHmDGEaATqGe8ly
9dPNTi5aL1LAuynMxgFaHClJpIU8cJS2bIOVneANbpFym5YlZyye6HUP4pO3n+B016i5Sf1v/Ykz
IrY5+lX0XFGABUwwPRpI55oDOfUr1ZXChoGtMDaXt0mQQMX81tMxRY2yTrPYJ8TDUiRM0EzAGRjF
a8C84Tyh0NsB6WPYNT6rghLEia3MLTjFI8nZz5fxy8o0002ydzhGKK0CE3xCvdi0Jt26+dH6C/09
yozJ3LHFeBzpZo47tQnzBife80ilZc7VsiP0GydnneXjmD9XIeCQmn4IuNnnZM50O+0F/taewKRr
VC4WXDiLIfM9uO7d3/etg8PR8PKGA7V07Z6n+efksTd8rWP6C8MB0K72WUGM2zFav+2qjM+J/5Fb
gX/tdpr+UpXA+Gxa7ENIA0I42B0bgcgwnyKmRKD1Qbq2KZaYv4xtVFmr+Rhbg4pqMLZ66SuQvhok
CZAXX5EARj0k4Ay/xaXEaDJSgQ7l8OXEdgRVXmgm88hkYBMJnYYW+8Iyy4PwmeOldLGjjqyoO5DL
JCQ1IBJYHrRrIaVEU7I1IAll1RkqIJ2QN3UPUfvJ74qnakl16y7trccq3w9tJN+WHePImDUEW8Wx
fbpfFAps4yWcZwD2HuLWPmfwEavPIRNM/f/as1QrgbWhXEdcICWbs2+H7URB4cPnx09REL4mSwy1
5yL6hxRtWea8k2skXxjbHHYWEyhU5IcRWOUl0owJ3lDSueNdVFuhCdoXANW9xganUU5ylj/VKk7p
QOjFRHvazqkqORLkC8AHFaiW6XPYk+0wXWZyBVa1/YRYSL8wMx0XcWNVcwTr85ssWfFwlWVLKC1k
Pel419+S1p5Y+T2aBFGhoh6R8xrba2mDCyBX8Z3waGuAI/Ue4oYhotN2nBEkNUA9t48gODew/Jaw
SA38w0+B4aVoo/0uPvoFPeqyyZfxOd1fqA0zFbpWdWK6NDXDreSZXfBcy31CKvZ8H/+VyZeAONiR
I7qWiZEO4ZKjW+KL81ycTYQVjxGUhjLjdf78kkSZZkvSRYKQrkbL7Ec/pbujyTabNgMEzMRA9i81
sivL91ZtMAo4Q3GTit61SgY58pdOouYeIUdIjKqaQcpjspbOuE5ivYTCH9nipN4w/ndUiepzbpCe
T18srOzBF3OkoBckVIxHN/m46KZn4AKaJL3WzgXm4maghQlpsVmk7pnLT3HHH+84IWW+BD+PkZ6q
w1GrVUV9MDHRTRgA6I71/TcJGwS4KngO5FPN/xSsVLfjf+pv/8GLxlFxRnetfiqLwQZkLupqbbPD
7ys3mUHeVfHH2hykTPtZkx90lhwbXXSMzkMHoP6otMpM4YGBfj4GPS7JPzJiDhX7HLlRf3Nho/zQ
k6uFU6+rRalq9ZZmkNSCIcQATKu0kQB6PXHQDsjgf5f+dlpiaNZkPaxAxS2k3VcM3qi3WD7ZOfvM
Xtf7ql9/H/x+QgoVZvGSCzYPpj4pel3eBoSyFMnYcHe8TDnU6WWe/8+qgI5aBUaWwSCQVGttQU4M
7Df4Di89urmjom97Ss2/KUrXXEIjScl5fmpFr0a22JvTca7AhDAtwQkNbJ31Q0EnaED3TucJLRbn
8kq9L5mhBoPI9QV3rEtSETu1d7HBhj/m1Xlzm6lhy9eG+OE4eRqb87A5novXmeEmkSsldJ5bi7oP
56DJxDhSJi7a5LYNUuCUuOgBrdU/OGwczBhwQH+NJLeK6v1y3Ap7D4hyML9La0CUfz9XxKuyuZc0
4EJMS5v5JPf0zJhcF+Bvy2gIHpSMQ4qVyD0SvA6Rmtyx28si9aqa6zcuom+nlEHYW5buI055NEP+
ZvLNVoULN/3iOMMd8hOb+2l4GaOP6dC8rhCzKRlEOf7LAgxBT4CMf97NkCqz4xjdWZ4oG53U5HIF
/xb8FW34qsrpG8bwOm77nK6Ii5980jKGLVzzFQq/pSJr3m8lV7RRy5f3wAUvs7bL1kQF/dA5Td4P
U3n1le/vdOEYcxQm9wIIkb9AiQgSiGxjELf2xTxtF1PeVFpn7zm7mTVpA5c7007gy7bOgCjdw+Ec
KGlSUIt7IGBfBZON21zj+95YI9oS0J8cFUOJWMfVcV9roGlO0mbbBw6SZNxWrBjIJ+VLeBL9WRmj
evExaTo1jaRH8/EiNhIy/C5VBM3xm/jpo7mOU7U0KKS5y1KlfaN0MteuoOI+0OSwBUlt95I/vPtm
RdBc1kyO4snZEPNJbqoDwxNs6JAbAeaQq6MJdQfeFESfHSrSNnPanGNKZs/pa0rZDt3U3Gx6XiwC
PMj3EeQ5krOH954Iq/ip6JaIvtM2/bAyR1yvypfbBRvDljE0RT/I+S80ElBQ0JU7ETrH2831rsww
D7ifGOsO5g+A2x3JIYrgtbrgLICwzerECw/HAdomyMW070AQ0lB/NK15Al60mwa6JFkvF3h010tF
sjQLGvAhAgaS8WUcfloZB1Kov0ObuGPgoOjKeSHAdix5ik3ybaSZa9Mw5bIr32safgsgMgFGUDmW
gZLqHddgTYK58Jxktzt+1fbhEtRgvkfPT8CI+ipE+Ghim2dAyBLjAUbZlxJzxz75zoxILNsnleRQ
f+nD0vD1j3uqw5rn6Xdl3oEdkF7y6ozA0HapXB2iRfZAlu26KPsOeg0URgx8sdx1/di+x3kJsMSc
yGfGMleWQjh/RKXfUL/p2SXUSLinkwF5gZ8ytvPk6JwiURwGaXMs+8wZJcMpki690lTy2IiBNg2T
3xqwxyi8CoJNutz7YOavCYkdj9Pe9mMQloyLhj7IJ8vPYxYdQFKPGf7bls99rvt0D2d3JvDumE12
G4UI5T1r9UpbeepKi0DnpEnKtbS0PeLpcw1bxbM3Q75TyjB/hYk4MlcfiBRRLN4nPrlMce9Jnl82
KD4b5qmSEy9TPpespR0E1F2NJHWy2GbfIXF3jw7jbRHceBVw/trvsorCSAZ1lJgsZMRRo1rcdO6n
zruzCpR0vof0LYJ4BhNf0mqJUJIc5g7zd/W6538dUqTDnW/lu+aJQKuLCmiruY42QYH1vCrMKr7d
O+UvIk0L6KzBRBRet5X4UItBI/ypnLQslEinKDqCQjfOv2H7BFP68iYqvSh4JT1CdpFyzeygNsbe
N4zQq3tdggxdRVtcCwNmW4/q2z0YbtrrxmPCdU+XNuryGeEYA8UrAHPNEvwm2lWTdWlui8U9YRMQ
uru0ounaqL//nJ3GmfBV0K2vZ64GRJ0tmMVePL5x5NgHwvGXq3UfDsitC2FyxqLifJMWNHvZVpRM
44yICtA33fT21PQrVi/O5DH3E9bRuz1bD9+tl4tLeC3UbfBrBP9tCemprsUX2diWFP4lfYeELreG
l9MBVSny3EBPQc/vowOOfzRs5lT6OjAYr3A/IaQzthk94tOrMbkYuHx80cPXY2TREm/WPsQ/L5Nz
VGoNoD0e4w51vy1H50ua3zDKzhXyJ2ZUTefKRpKqKRKGttNOaOc7KZMS61xEhWDEng5fcgv7JEfm
XsIZ3cujyxMAi2jQE9+fIdrKjRbRMIYdI3WAYeuFCuxGRUFB+rfZgv30+zsDwOWTPoOEQJYuIRKr
Fq86VBivE9nMJ4gydhZzQmsxIv8gDrLRw7WU+Ncr+pASfTEdDmLRiV26PL6hH0Ibx3NO/Y9d1miJ
Z85KVkK2o714Oux9oX8QobmNUO4Y0pWlHmXzFe5Hbhy5zjgA1dFMb5oyUv8hgOHTsil/2BnPoZ+X
/gsyS8spf427pLKZNnZPoysjWbOM0Jw6ciuE7Lto/TUf9px977YdC71w2TpvXnip39wl3xHfbPVR
7GLgyJfbhZyuSuj21LG5DdzgKe+ia5SdKvpjGw5D1aOhAHvT6D1DOkVVoQ5lqEBUWvlhuhF1TcqU
WvvRR+uF7buWKRG5nx6gZL0G1gP18XvBwgt7DM/XbEHx4dEmfv8grSvaS53eSR+ToGle+ri84APT
E9+91OUtxLDOqIDFKqr5LfjGv4Ry8msEFYj05xyYillP/QWMYPm1sFl4WCdmXfzwQ29a3v9bW5aW
cTDDNQM0qox7u5O0ugSjBq0ZvmlNkr2evV3jcXDRsPGyw8pmZydiOT/YxmhEhvko0XzuYor8wDg9
qYztJ5bEsUoVIbhzrJrbWYRHQJZqYtqe4L36qnUpbEl6IPnO/vXiq8cMbSB1+fVsSGg7JqldEfzB
dNuvT/td2EzgsIUyWYaK8txuBsm48S7ld25i31+KYCKtC/+T+N8KXfqiaAZAmFTl4WOasG0qHXOa
C98pSCE4Itxsxgp+nboA05JgvV5bKneoFuOJjpYo8fQ5WJivmuCN+icMUbTyQbeDnZX6EncPTMpS
VyhkdHGvQV8nyNdZryE8ruw/NPIOCkUgByN8pJDEAAZkpBceIUUwwQ0v7+fmw2lSoPzZyV5q1InU
1FntDxYQzcJiPlKGtVfV/x9okpJrK7u+s1TINxRfXvyTlpeWNaiS/w3ID/FMjISAYQ2zapTCZmOw
jkqz+5i8jZ14UviB5kALD6EJ9QqKmSlHkCtVT9v6av3FFagkjaU2VKSz5EjkFLHLx+uYlHx5o6wG
I+JSOAH0JkqiDw3kOwQjtaQTVNops+C4BJtZ8PvbpiiiNRRxDsHoNEbmqWfzPKrdalaq3wvFEJNC
LKbcd3CTnV1mVBNaKHTa4YrLKEEWiJraMlUEPKCvIfUIZ4Vm+7JaPOlIQEf1yQJ434fmMpMf8iU3
OXFiooNbI15RKfyEilEWtg2HT7zKMt+ZBYc+h6WBdlw4CCbWQ7AJx37pHvOZ74RGQgt0avz3vXnY
fvawAwhJNoHALsairijGLAhcr6QL+zov2156Nn4E0bel4BuOEWt/pLrBLPO3dwr+j+XEI2ucn5ce
j5XfrdcUuSZZMYtYmgu/q6U0NlObb58gFCKL2OTea2e2ccP4R//qTVj20ND8syXyIgnCBZgOIgX0
gNd02k2X9FECJnkxH80+7ZAXg4ARwBXrmuW4fLI/PHFknPBGTEErJ3kHnFwDKRNjfGfQH59I08J5
sZXShwk7FFWJxRmzPmlMMrEiJFwfDmIDHaTpTOm0WEMIgsdMyltd7LafP0hVeasXkkH8xMPD1zbR
ekPX6jrfjk1zRrflhTP5wzP9kEMlk4XbAOHbjKxHkiNj25MFbxkFhTJ7AaI4LDKW3nR++0o6JILr
cmR3MnU0qfh9+w35hwxDO+9KX7WqvBzpx4na61o4VPSwm+xHpMzwJ/YIzhVbGCQdtbE+n3YcWHan
50llURdS+BdLkypDRIRwz50wkMApH32lZOhgfhswjVcPOXkrjZuzp6W97nNjo84/8Bnb7DGJgUR6
we0kvl5fcUnZ2TAIf5rAcEE/RYIw5rPbqmWafWRP3lB9kDGHFs6ylFOv/SRSiHN+xqtELTp2UDMG
sR3+IC/zJFOgukbpYuEmFVpjAtI9kk7F663X2SCJHifbi+y3nxu34D3eAaOqibIH03H6JWbsi00u
xHRZebwQ3KHFEEgXpCCLIq3y2MqWyY6fpKo68/LGyymFOKzLFfADVk1BwqiRyRUr2OeUn3ijR6WS
Y68LM7GLgthq7XyWkA5HMziZ3wB0VlkhegYMFbiWPQI0P1rrPWbOZ1YVn2/OPdApaQhQJOlOtUT4
AD83mVXwH+HCzoFBwGik2M63snt5Pw0zCa63W/VPcJdtAuOJ+xutmPKbCMyEHrXGyFzsj444n770
vo23nCVenKQPLE4JiIxYooQkT8ch/2+eQUOAi/6xEhjnIW4zfqgVjFGIG79tloXtFDR4eizvBWik
NmBrgBv62yvqkbh5J/e1qhIEKHuFDVFMN0V1rHC5JeeV+Fbcz3wPjYdIRhaSmBHTTwDyTRSBgzPp
LEEXwJvLD67AelQTNFc8GOy2NC5+HVBjRxQ1fPDwvPObMzQUsXFiR9XY+smzJwH1OHCh7sngki/L
XJN3iRnNgWTIga710kOvp566k447FXcZuSOKgqXhUD4g7xiAoodrFWZHcSPruCY0066iI1WbXRQh
fYMv9Mxw9J1ABUj9Ok4ed38TAjBT489CYQJod4pQNENA1NIe6SGzXOD1RNhKWenuUMrgoSW8keXl
EqMzz/oYQiE2XEHbcBBaY53Xj/Nju+T6BbO+rgGwp1sgKoo2Mj/yYYUSksGL7DMzhVGX2Hiwczys
GmxpqwdbDbOCAtLVjc8KNajW8bBEGhO4DsR5ABX4WzP24h6zg9jtlyuRBMlRxTHpSbAi3vICIrWg
dXOMj5oHPPF+AmI70fJeyw9WslxeV4dpZlj33yzlaakufhv/1UGtQO52UwmXQcAcM8Uwz3yVcKIH
3YH49dTXmeoCB8j3ZjUVX0+EOynE2XSgPou+YN7n4JJT98UOZ2JU+Khf7jrkCT7L7B0Zp5orYZRp
u5dKv6nV/6GRNeRcNhXx5GJoMI1C/LsCWyLU3A+qHcD5/v1NTNnT7KABg7dSEsIRupqzbGOzx6TX
nixKIttm5yPd45DDV5FdTxXdjUwBo70xW4dRwFed308PMY9QFyYTqekNAxoDwiNL3/V8JNDg06lg
WxYxo7uAYy40vTe9dWituKlMOeVjZ2Wg1+s7kUtqm9qWBuEkmk8dd7BzniAS6ULOOBb9vDsvOVWY
SyFbluWc/+C3vKpTApouqc9RD5g8a/Sf7/OIhDVD44TBUepKkRVH9npaniM3YJuushbOF6yDpo5A
TYa8IMXLXFz9AdS8cFV11uL6rNhLMc6JZ2zIdJ/rC/j77/VWWs0M4uqSTYxChwB1fkkE8kZ0qzG8
Rp4jJShdau7SIDHIsIpQv9oCXaemdtHP1pqfDqxw7j5IwQqxotOmXEdrVUMubm3NxMQM8BYFU48r
tKImASy9kofq0/pO8XKWacnnp4H4CDPQZPmZtCSAJ9EHSI/J0CUMv8YIUQ4SlteJCfOTY2z0wvl1
igQn1gj09zqOQtYuADrLqnXATw86NnWbaRBie4fqS0UH50nAUzUNeZjydGHYn7f9Anx5XcItIgYT
kqcLh8wvN1wBVv4i6cha2rMBtZl/bq9lt4WthuYHdwcZ+e1hpKqsxvdLOR5ybINFE2UKtA3w+c5Q
WWwcENC7ahBZ53qfi2iuiw3D8j/rf+mB7F3TZ2W1q3uIke4U3vMiyElPApU4yCvs5qsYSVNRQrkX
4jRYDugutAFjxjIGPDODomeKHyPZrqlkASngLcpLdMSWO5FBZChH1MnCn7RY0dS/3nFfmnj07hN2
LVMOAb1PkZ4iY8fttwjfYhg7BxBYH1QlMOSOaiGDV5kVMzXs5NLJdlzWWN8fkIm92lIwEuXlr0QT
keE2+gfw1jxAMNSyrBTTuDazdT+NUN/0im20iBWMVI+EQzjHsmAJhNQ8mBK1GmeAgwwG7/Hp3yP9
7J6fPW/1FbZBcezLw9pzCSSraLz18B3O15adjMuA/dNuSNaHyWdiPQkC0+F2NOVtGxJxScn0RN7t
kAF7jBogmVOxywdpFowtYwNX11VuFe6EzWgP3QfeCHmlI5b/tTDSWUy1+2nPXHDn/rL80w4RcxPA
0guIclvid4SwF92VGIHqOL10N/He+yXVbofuCO1pT5DfbqVztWty0qu0XRktB7/VMDGt87Tv2vgo
dYcmpA+sHb0OOMLdczGzSGkSPEyYNPR2HmmWjhGZ1ZnPBKp1GbTA6x7tKj3dXrapAwYMjGJU95oc
LCRSyNVR6lMMcluLcXYvaqn6ffAm/gqWfJu168S9AlYCjWOZ5OAJBx/sfxY2YpMwM8Kg3+xpGOvq
kqwFVBEFzfwvpxrkySHj6iXfLKsLHZSwQ2VrD1trYT6zG/TGGojpoyN0TGavYJqlZ4rS1gb9IpXI
7r1FXLTNremCKxPZlRWQyRBZgHpcRqp8xQFJm8W9g5qaY6cOrPoCNCSa1RAtIRRNZ6BBEsT8jRoG
IfdlyADq2N2exOp2qMk/k3uoxPbFwIkPm3RgeylfX5TilhYoh+swb4AGBHFomqKByGe5xb0DtnbS
6mijOhBPU75pfpU0MgCarlarxpoQUH1DtneVbGZBdeqsLTdLFfnKTiM5SRL6ToWqcZn2N+LzaQ1c
Lp/4TYhZ5TjTZqPfyy0ZkBJFIlYAjq2rMAwqqKRlQUefdm++jDIvTEpw4gT94LJYE1k5Z7zqTVIp
xjSJDHvXeYeYz+mc0TOsCwWwcdYvB3o2PCx/AIog6bEhwzjwqe/bEDBSPDIoouzQryJ7GhNVqpnv
WoOgWVs2FIifJn7HeEClpvkrbbsIFpvFbfxEoRYdhViscJ/gtdrxrq2xhfygTijR+3yiB/Aoi44n
QKnzvkvw7y1fLPAXanXqJYBX3ARB37o4qlCdZEmDrInvgn5QTdMmAlNTSRbwbv++LnSCyq6Lqhw6
zieD4c/mRIO6jczTwHGX1NS6EFL7nPKIqoI+vbqVbZfG/I7+9Eo1tMLoXPQKYAG5D6nRLnrvQe52
r+M+N8+ccgD+OK0RMaxfAvcir2hDsEDiwZnANVr9nCR6453sXX80L+GwlgrY2+q+1PfUUUqQ3+BU
+KE2Kb+CQfgrxwPcw+84/coaL1eWjVWcKgV5h/YFsAkq+z6i6ToY1G9lkfG2feDbhHBGBTbSgnaD
3lZxSEzMr0oZ9xlTsrJqhEcgsK1VjN5g7dLg8iJ3ZvTvrAg5TrS1VBK6YweM9WcAcRGbZwYuDRM2
ZHdmKIiWbqI+nVPI52urSUk61e+PDQeL4XNGs8XH0PPI9hG/PgAnZgMWlcyklRCPA7/s0WlNded8
LM0zzjRwI+TQMjTv5jQ1sOsQuEeHsI4OsmNzv/SxBCrrIMNjtnVWIDzALG143wD5mUJIC5WvKLsa
aBq+UHCJ7tt21qunO3Bd+UvQWeKnJnmSaXqLFdw3Zvc7IuSs1z1rRs5GnJcH8yCG9PwpgWDSl4FF
YBiKDndtcGTlaZLe2UsJxQzZtbA/I07Mn7boNoOXXu67vwQKcT1HEfpfd5qNFbq5o4a+12mkCf1k
xvysC91eD7aUNnzYFoRxYA2UfYP1k+/bdFoudM8Xgo6VR7oGGfF2OgNprF287PAt9/asO037RJUk
FUo4Y4ZaODTLhLKYc88LMt3Y0fTHNVlAeceHFe6SMIYyeWYhbuVLX+PKMzP+b5ZG6PDqMHWlyfNz
qin2Z2CbIQ4wvZRJj/JVXPc9aG2ZHUYfxejeGvWHfZM9ZH1Z8C62b9XcYHTolnVfCpaalsmTXlPL
7zM3RMleXBLwYS1G/DzlQAPTB325ptJi2oYwm432qXSE7e3xZa7V5QvmxkIaRabLB6FwwZ/KKGIl
WW2xqxKZvO+zjB7nRMZz254Fwa9nRMcJcbCD5jnKr9PhA4qCnR/W25915NE0Ww/NHC86XYXL70C8
S6QtryKhD32Xc5581fMtNooQQAbfjjkZt8zfl7xUST3Q0Z/ZRNob03G/EvrLbwYNqztesGz+qb33
SBMZ3upDJoa6Mxq/VgJtthZCfSRjeD6Hi49oekDxW4C80DM3dHBEPLqMjIQkvcg+HoYBdKsANJZG
mffUoO6FD50RtQyGSdbfThHdFm47lRXE9j3nidmJKUYr0C/Wd0qAf/WytmcXXguzTVDgTtVR2E0q
VDxnx81kktneUkn6ZkkxlD+qQ1gDXVlmGjryGB7ol8DeGwjqEzh6I+A0fiMMclDo99rQPY7XCT0K
YEchv/wjhRpcK9xOEpvUxRa0quvVx0AWCVcW6TQojLZPEwwgeO2iklen8kMhLrh+qUbzbFppHOph
W272A6S1zpecQxjOGyCFL6g6MO0heYAl92/PMb51rASTLyqK2uij99jfPHcvWtrcfeNQoH1quig1
W8zuEYnAFdu56qVp/nKTNwYTGUGAAVTohyRThyYtio5D+1EgqsVi12mGLo0JKnFNnAL89YbsHYj+
y1gRwmDPjyNQv6uiSa4KkfA6QpPVUATZbvE3u3VXkXASgqZlWic/EZGxLH1HPoqk4aWir/sOGNFH
YCbW5mslLKN0Jaj1NeaOl9zwbuEb3RsV6pp7V4o6xjGywwlrGUqRjOeMAderB6xjN6dmYOC5ZTXC
bUCJSMRCHSE1DQj9el4c3EitEg1tazXhzmUQfKbG3gfWiTWqY6UCsWtfDLT0TUpb7TVoqddDmCtj
HNyNwB/hijQwujs7/yVDatX8g7mC9MZjPKIK8CRLs4ehn6CS4JIpSjWn2jDQQm2OJygBN2NBI9Ae
I54uTerDOA/fmGzpdd5Ghn4rQizkhD4GGP0v5cwdXouaSH6yxaML4k2zB3/wYPqvomwWpxUcR6oZ
mt9LkqhvqfogB7Pqrbd70zKBF/XGFPsdltbdlYRd4tUrhfUO6uqESquL1kz57hs1Zr5J9hS+9rrK
Ynn3AIr2644nyEFUjqe6Nlll17mUcz6pWMEEYCrcwb9Id0AId48WEcibgHmI9HxlvvjPgaVhoBiN
KiLFYcL4mU2uM/xJG3Y/FvtX6CYdvajZa2A4oZf4XqWX891C1EfMB2OVHJThnz4A4uSMAvqmPxOt
fefwIjzNWwip/ciC3B89RJ50gq1qTijrT7pMdRsB+tNIuewgkmu/0+dfni3+4Z8yPhoGw5xqxj7P
9A2MkYnuCDo4M85HtQ6bN3aUpwxY/979JyyQhet56070hhrhFLv3IwvCezkFoXOG6NI6mCBY2GJD
Hg/xIhKrSHEsJFsFF+DeHPQh4sWTQJ3kqkfDBI5d6SEWl6s98vf5NaGQYnuoIwWmx7/mIHDHBMk4
smIlEkZm+A6FMKWfXrFc9dgxj9JU4CHOuefaurZZNXyFeuS578WKa8+50fEMiN0sCL9GXseq/ycL
DI396NJaol0MEGQRngHmgEsXHH+Wlt3WD8GjSyEmKP8pTxsv2IRMx3MXska/9YDPUYyiUi+gy4uo
5XMYRg7C9IK5MuGYzUU+SJljxKDFaejVD0T83sHf4TwBFJGCILn5/uRcaH4HTb3IW9qa9kF2Tp9x
fHnH61BBT32kLc7R1kisUGGWUaSlPB081Cz/PLKqQAWN9iHJlQJY6Vgm8TJmt9JxBakK3JgA3IJc
AiNiGSk0F04kGy/nFfaYDyCqDUX3YbhbP7hijwKgo7i3n41+ovWrYbleC2DX/kXCeKzIxoiRBDsp
Ks3ejpJwPfYMg1FJwVbW/istybq/LwOebbaqcZ2ichq8YmGLd0qLOwcDkTePdFE3ULjTies9k/Yk
8wG5i6/3/EvfsOpdtiQ+KVm1hMlO+WE8wM21uEv4eUyesH6ErFRfEwSgQY6Jr19xqKHtyuZYVkv1
2GC/yOXraxlB4b/l/rUUbfphQxXTvDXcvMXaTvCRwY1Z2EIYhUUapmR2aOhAEPgZux0HriTl04wm
3sLcVYdFgjmRmjIBQlvlrE4ouQbULyVcPku7+SlXVAbgvfTvTgiB/LiN/oDTYQ0tWOHZ2KGQSki0
4ehGESd/1e1dPxCpmSwX/I9sjaEs6aj+1OJ7IwuiKskoAeYfDdSwJ8ImF/PkUKuDhCgbauHnz9I6
lWnTZ1louJW8yUXr5hF3i9UgKRI6R1kg9Oe5p+H1MjuXQmdFGXFWv3db7oebsBLdfw3O8AwTpRg4
0iCc6HL38bNctsSIEw/LzIgSyJhgM1LIp+FRyoTtDHzBt7CPD1Rs+4gQd938prTPMBxwqKyeMxSx
Yf1CrI9wbwCzozMMA4xHpftp9rWfg78EJTPM1wy/SePr2RvVxLMsgNkEnZWnIOdBk5fk3pgGoPoC
FEHITl0p50+EVOYX1RzKDZDOFkiuBObN+Wnmxu+4V3yX2GdKPJVuOmv/T4wOUowMdm+tGINVzQoN
IjinvdNp0SBN/3QqD4Vyr2OjRf+30CkypqJ4fUC6XUxUEPPZIC4eymwiwRUlHVZmUqNOwfwJuBV6
4mKWXKrgyFXyJ0tZTyaong+rn6jUkacsl5kuVNIkNRuzH7mQHuxnrJvptfI4jgFThUmAyvYQakCo
cWE6qGUxcNUh9F6m4CP4cRSDpw21Iq+mlaomTdhrbsjSdHMe1fxEAwaVzrQRsYIZPwjfzgDlQlbM
Ej6E9hF+y/lL6IuSwWXH9sdz72ajm2FHRxI9j6xBV5PPTkqf/K60XzkHIbuHJy8S2YE14HG1S0dM
Rh8QmG8uGl8wuqo22Mj1ZJH9s1NCAfZcwkoIWoxV6HB85+66rw68Ykq4NxgVfBKSCjeL1gjQRBeD
ZGCAU5csrW7mnLugnKj5lVyHbu+X4HNddWNi3dMGlY2i6o1zDTgIUFrUeDt29THO3iP79+OUXoFH
ByJOi33nEQKblJp81UNIFips4VgiOnCGIFl1O+qujWDvhLBpnZKprVmcqXCgtjy3Oqo8edj2HDUw
F8EK6/GMFhllDHYIAlLLPRfQt+AQE+k4pGXElUgp8EhKEnVJAVCowtoHj7/AnJHewUg4b8/phVNq
wuofmiRL6TTFiYeMUwFYsgsLy3J0RLJbkh2xyz+lelcU/wVn06Tu08nESOD/KtGPDL7C+csVtnT5
wpILYyKhtiP4eSUdfyzmFJV/BzPtX3gJUoQuu+4p3tppARc9/HIid7R4f/QfS5i79K32MzpVVJNM
rUkINwhsnK+2bd13WjOwm53xtjBf7H+pexB1Lyo6PyXrHqi8/UGqnriZhI5ebxxGHx/1pTxYJAB4
Am0jJA40aqY4J5H814ZHiaz/lZfqlxDcSFSrvJjqYfLwo315Opuok+AjI3QlZNfuacqPjAVgBw4l
4ktLJcPbrNMwsrndX7q8Ra3p+1qiDasC4RdwpXcKHMayEZSnj6R+AsDmXuOiVaTA4sl8m6JPZjyM
Wh1eHITwQJvkOiBd1JGT4ynl1L5ij3s+ke1B4wGyUK6oVRloMPee4inffRBytlODS9ntVS+NvLEa
KV+1dZeLpq0YlnX+pLFP0QSmrlhKsZSiPFc/CKkNEKuNWV9AGVnXstbwfwmGdaRZ6WpqbFh0xKKE
u23e2lkMRLnswcuOvxdUdnA5ajZrmSSb6xq3/z1PI7o5ESzVVBgJan9sYeWBPUXMFFMNhUtHm+Yq
1O0bhMDj4f0yr9FAYGQPWFqO0pTduhGFopGQHuwMWdJs4aC3G7nJ2jIDI4weTpDbpc0Yh3+YLynh
OEf4T9TlbPe/gn4eQ6G7itts0clA2dpxQ7R91QdMs7/GqqbnDfDTzhJ4n3eq/RbPRYLwS8Og/VT4
H0lp85a0LtFisRU4218KZlc1YHY0rP6KzR8D/dfGWIyICXRyq5c0Hc1WA1FN1ntv2azqE58PoxeF
m8hKD+d9Q/IxRiUT0DwqDQ+Bob4QDkOJV94OUWDR4I2dP+9qcXQUGm0yD7w61TptOfwiwD3Utz72
0Dh4MtFXCHM6ATD4SQE+h6n/IB8GA1LyfC7/4x8vso53NEPV0b/e3JCY6biNITRNYmWwJcQBTFHb
Lyf/efrbTZnh9MsXeSsXwftWygenydWXjBhP4+Derq0Mml1VAZfWALWAtjIuhu/N034RPYYsioT7
Gi/tCkN7kKlakc2dUvjc9VqORrWI5/y8QfC2UjWP+u0BbqeHu9Ctd+dXpY8HPQpU3Sw7KydS+XNF
Z5ujplmeCQWQfEwR4JFvOfuzMa34N6N2cTdZh1bhOcBxDbLkg2x5l5n9GpFNa3Zwsr9hGJBiS1CT
nvRxuj6OG1C3exQ6k+QLbafI42kkY7Yy07thgufxokVI+MmxHDExyA5dPlZ29NEgSvO0pPRf++tv
FZ2ul08lQiTktN9Okdx+X3+U9cwxN0hlOEku3gVkcMq3Yq/SqukDf9gdKtzWW24MA+VGfxajcUhv
79kinKckCPr9L3GvrB+pFnLCMp2wk4C4znWybMQWk7QIVU52x7zOjceCPlJ9bvoDzZ9Im00sKLJ5
0ehdHzInBMUO0p/vXpiaAuKL4hW7RWz86Mh93fstOPO2EtYyLsAdysoGAGBDFop/RwdRegtSwGAp
okokIWnf7Mp3XVbk3gjHK1RLdh0vmQdstbas2iyPLMx50lHLF9x8V5/v3K6oqTIAYoRJRGA0AM9Z
vV7JeAUVnv9b9bLTKFz2urwAYY9Dg6BkvPDvTCww3mtZ9GI0siu2a+9uQ9RC+1mfzegy0n0NzGME
wHh9TNFb2CpihLJaYrxW2ELy6/KGuloPNvgNt2IzRTldeHVm386CbK/GqAL4LrH22rrf9Hs/642v
D1U7EL75wsOnbTW52d34T34wZe+rE/xoiZ8Yau7jy9bdanulbO26MzRCQpZgN1zJumsK5cYubuV9
p2V+4kXtQ04KAvfoLzevYpb8ZLf8dhVnmlqdc/1Kzrak8omCxJQrz3i5xHVG9ZhHsAFViRquBwcH
FJnMp/A2wV5EzK3pczyqA2pGL5siwrsvY1etUBzyV3KjfcrFQ7SZju4WYW/OqVTbZNyzX11Nini1
IXnBCrM53693FoO7ttnwBYUbQG7pKi1DTiLLRyVAGLdY2K0P0HYNj1rc4DvvpSG837lU4Kmgiy+J
W24+Eygh1c39Nchnk1zN53rNpSU+spGoTIZPEYYwTiOFYw5RPDAnm3arD5wdbZ65e3Vzcc3Lgrtl
obOA2RRz6qM/KrjqicT2sTpmf9kN0iVkaa0Eq+MzmzpEn4RwsKFxbYYpTkgcB9xpW4k3Dqf8u/TA
ayg5qbtYOrwfnsc5WlZcZ5yLVfdisHi/zauZPNWEHTZ0bHg1WdL4P6he1nPjXdyksEB4Gwcin5dU
yarGeTHkE+Mef+ZHwRzAC1QOsNhC5FSC68ijIXcte83QnPgrdgZd+cQW9BqY1X+Ol68Zyd5fNKNX
zakA1DmQ0k73xifHHKFjqr1eGCX/friOyvE/90r5uCSmTK2jo/cBJauz5t/eDpIjwEWa8eGRtotG
AJI881ec0NqUXHps6C6GhsbKxy0oCvTumOQCuLO/JhMpJijq22fg9mYYBA9WQrmbjekmQqBuj+zI
/xjEls3OQAjJYP+OPkPBuOY8VWftI+hAoKmTSAbkS8XUHXsdbYwZVus4RRAPMYduzYV/vX0gqkFd
0rsuRjo1PH33rAqQ+3EKR5nnMrwBdme8PXJdQSIXY4ZmGFxE3rRaIEGa7FnoPEdC2BquBJTCHQzi
e9dXmXea9q4SEQnnh6NQXCKuzb+QwehIA1uk9vl59d+VuzAnre8JlJi2JGLYSehYnT+4buNz4ue8
fcgOKNvdMBy8gAaEfnWmhrCVjViR4wS58909oqNLidDtywT9i2Vm/skhDbKq1u5gCoOaIjF/NoSC
rQTcYJKIfaBd+4ehJzR/Fb0OjxCIcU8mSKiY2z0ueS3fCJwD6i1SpXmp1iCEStvnW8KT2us8PJtQ
jS6YM0UUujBvpMim5xnVaIywVQGM1FzFrtLg9JmiVFxXlLKs0U5e2BiIl485BFcd7IX+tpUE8/h0
q/7cJ1/kxQoCasF5gj945qvUUkdX3DR8jsVYCeeVS/e6yzbCQVphN6nbRSw+EL9Wcr+6Em0COf+n
MjWQ4zuwy5InJqTvKEfVm4KByUhjgXni8fG/mK48seevgW1jJJtAzDVXlDMDp5g4TfIQsbMB/Vfk
ZNQMlrfI4cwmcRyKInOYnzdnXem4O55kKvbKTOc6xsnkCys1US5hI1S+X1GAH4C/yno+VJzVfEx2
ajaAOefDIVojXgeMta0ZXrkbfeLgpE0qrCJqiePyht1WoMX9R/2cIo9sw0je2R/mgyC66JUtzIpk
hdbdwXT27yw08hJl9Ga99UIXshea+WjAgSoIJVBRM7UkeLsagfbDorFkZs2BoNwn/jLr6A5XYdXM
Qpv0UiKgsI7lKTNuMpfhcZJcOd09y6dnA+AAC8h5hqQ1q3Lro7XpEo8YCNSELYnd1Fj3zgEQDosr
H9ZUqXrpFZ3l1Jw+KuToV3Ic1msp0wI4qox8D0Nq7dipwpOcby84moHUEk4q0QcGf4c8+9MAYld0
b2pisv3/xc/TD+j4gyYNVLFYW/B3QYlZnZUTMi6TLXz80wg2lblwLf4ohgij/MdYKKX7rK2REWKS
FMRvzOcRj0BKWWKalnSx35G/pIxqmk1v0Bb47RMxyIpPjRVZlrfbB+vgrVIP3RER6N1BK98fCCcp
t9ZCrI8KHbzB8+QtxaJKCj36FickH+y6YSbCjvHOkLu+uciXTEUFmsCfSQojMoO5oDCH7c4xfDqj
luH93PZsbYWxZl0bvlwlEmfEg4ihwOgGhmv8TveaDKF2qjlCYz7AASPqxOXjUT/ZRH2izMTM61wq
SZBNt34hZEHR/2E6scYtWqLE6YNh2S36KKBIoWZ/WxakvKSTrjOkQKGpVF1emLoFDjD06vEvmKW/
umk2BLcmEww6BkemrMV+IbUP8FsQ5FnBX18Zu7X0B94TyJnUwpaoe1aNVT57gDcJWFB632KMQU7o
ryRm94K9w46kJQixwEUCMW2D9AoD/AuILv2NAzKn1TgiSkINUyski+9BKyTgf+d7g0Ec/11J4qgY
qSly2Ly4ncrMR/jFPc+7+Ue158PTmzogvn8CFZxDncwbE1uBp2qpiKXDUL+ywlod+PoZpVW1H0PD
d7wYbD7O4tTu9wsijgjYDrLq2lnx7XLUwZNpiIQ6t/VL7oJJkcr7I+HVdrcDtz/ApN7b3Z2b0XYi
SpFPZyMGLKE6w/Fr6ulcNCTyRL7/3+dD4853VmyEBUEpp/24yos65fdcQtd5fKm8z0JNRsCqyCKJ
Q6wq2rg7lBZ9mniaCnAH6n+iioEoo6P5zN4qMRs1kD+VbzJmUMoMqK1eA3fJVRw2cCiPmRgVrhku
gtRyrPgODUjIQRTLTrPJLNzDvxY6JIImqyfxbM4nAp4YehAeuoi0aKn0BxJavFSvWRbgmhO02bMe
OT6fl9lFqGArQ7EXMUNwN/KZRcK7+x/HOoD9IfvJG59D7BQNG4LlNRkn+XAJ6IONCQ9OJSv4vcls
91jZyQ9O3o30XT14xUtJrb88n+sn0lM99AFjy+fWlpTeIvgU5VEqQNep3CN6sypwQYNaCCVqVXYc
fmpr4dpBJ/nH+nlKxM8139naHISB5Do+7KlQF9pAQ6YzM+LCRUbamNSB8R9XmcH9ZBDKNTwIGDe6
PJNZKn/9zB7+RHsNSA81cF7gphmw8sLoDN4oPTYw6VtGVTPuQcyFDqkdOmf0bAXhYxNXTUn6HBvN
90ngzXMiYbwIifwlo8KxCtjgIZGXdu4uz+xba4hlLwhMIg+9u8QWkyab1xswoTeJJmeC7iCgGvmI
9ggBO3x25E46BnLjddyWpc+TeY4zjJ9Abo1oG94ytTKNDxfuTYzjIlUvMT/8CmkdjweX3W+3NHpK
lJRIPC1dp91hh2o8kUoB/ptModH759N9JukQS5pIFjIuldO5UDqhMuFEnlsHUt3VcnkLmMs06G/G
/odBULPD/knez+FCeewlCwbhhIKi75KD77PrtqQ8RROMBmAtouORjMC5uJuchIInrqEM/T1DXcv8
SJNHdjk66jsMh4C7RJukz4W0SG9Q2JRmQdji0U+6QaDfcTaJE8f6VbFpZX01tyZ6zR+EI/nsv7MV
OWf5VgAUu4i8wIG9hleobANfkQXkz4GjPiAi1wEeAIQ4CpMigmS87lhE6pauJyAnEz8+xw/KGEVo
fT6x+V+V4jrmdpuSTxdw0vlZwo/mUxgokqINxj0Cq0Cx2RcSqOX2XdMK73RYhrjQbXCzr5LPxI6l
YftxI3AHsOYU/12OVDFa2A+8GS3tUNXF6f8e8ibIWTHWZ1o+8apnXoQxl/uPj0NvOQg8Oza10Fs7
PEsUZxFO7ysgDu+SyQIaiKoyAI543rtyCNv6ERXf8zJ1TUTp3LMa/jWmGEoriTPQKeuxDDcxeT8M
Mvb0+0/a+tqOuobrP0PnPJU0eVXspgpvz8b2BP4B1PzuS3DWQJoejvEMOhLJ0MlNT1WdG4gPKxnQ
DsSGAl26JeI/HbEDerEUohq+wqVb2RdRircVCJh3G/5cZRmJMIJ0jVC2RwC1gRVElJQDRQUHWngE
iAw8VZOmcVbVGBSAP+WExw4tpPXmAXNPOdYVrXCqpSD0W4wBaB6RinYwFbwPoefyFd+807EvMZlY
HV8kIbLwLOZnv+QkDXQZj1C0yoHyV+9uPS9j4mqkJ9YJ+H0B+HzPYnpYep5WrZPdmGe46FKah6Mt
mzF65VtDNn6qcLbrT4cGSfII0iKh0HiY4gI6gY9S2zMBjdDsW+XRGZWs0Dv7H0vjTTUXid73b3ZL
mZ4evyEVwN1bd8E3izLJ9eljLNiCMF490HqaWqanYnfuqCT6tR3CevocSaqyUULUgmO1hMOKDNiT
2dt60UN9QD/q2wtgHOC+/lt23AB19R4KTqXr1U2l1nPouLKfDHRh819/u+Yo52DiYBq7Js1cbL+y
sU873K0pVCtd9Uv2ItsAQ+BeHVvHSQslnqZPniVzd7wIgTdp5DvoeOud0f5dMcJA2SXkvd7Ev+Eh
ZQnFDhFVVrUZzRic3Qvdbov+GeNGPtihVMHNEB98MDA/oP9bN8JRGcVCC7TPQEOlk/0SFx3yIDjN
Jj6fmbkiG+mwZ3Urg6D4AuVljjSGp9IypXc2EDnB9lx52/50gY6mdCB7Ne249vtOaaAxBIlcvQFx
sHrLjKAPRDKY1RfElOqNLg3TfZBdAp6sgK/mRoNFTs1BRGv/uvItM3nomC+U9Zzp2v17a2Clo1nY
xLum5TOhMXbVbAFBgxvVTTP/w14ZSIqKujb39wuSO8Uttqiio2rh8YmU6VGkXfQtfXVjnD9D0UAL
jMLpeQtTUTJdWTMJqqZyeRlagGjzR3qYpgq8Af2NwPjeowqLKS2mFPSlUaBkH4NZGO7w08LOhwNw
fZCwP3rkXtaF/IOxL6KqB1A5CgPD55NN93Swa+g44cI7ifX4ri/DcJaZXh9ZiEz5rVE9wqK3T3xN
eU+NGtF1ROFDSkmiWu3vNsgfjr3oARnzuM3qUqp0H7Jg23zMr/uURkxBB1Bv6M/UYUVOtzKxhyeG
vLNjXDrM+EYgtjYnYG/3TPpTrV8VmX+94AVQ8ICKj4aKQ8M3ko2L5M9zRpPspQ2TIoVXIL1MgvTe
PfWLGZxxn+ayRnfdSzHWi4TyrZla07VNs3pU2vOEpMNXZmVh8T49eQ5s3UW2+sd/x9ctbx6EuNqJ
b0Ti/44pKVGurs3oIEGqxAXn+MG3bGK9SzgvzIxAWBTIKcdgO32d8wIlqBfGVV6rqgnBiipQ0beD
3Vb1Wy+iOc9ITnPB7rbSbrKQsBKQGWgdb2MoJSGiQTv8wIOkZzp5Hf5xiZz041z5BIyUY26knCcg
X9d6lUjHMTFhuxR72dqoOmFs7UxeXO/emeETgbOi5jv0SdD8+0OZqJGidHPHpWjJzfab/ALCRskf
r2RNjp8Uq+vGxlXolFIlzh9KSKRC19nBnN4sVpSbjmk0QB9tg0B0CxOzDVH+sRzj822Jzu6zpIvm
n29DyBQ3XkHozHbTpRGmU0023QEhnXr3MybA03GMj4PTs+VM3bwctM5OEsNZSfecSA4oe2lLfynd
7mIXmHeA3RX1UNIcjVKDDpEx/T0hOxNrtQJ+oeo49UqnmZ+oDc2kNz+SJ7pre+/DeWTcdKpdvvtL
y368Ldr0vqhpFN3d0lw32TsIyEcdek5SFNPB2wMZ12h356E3PPuhXQsWpKNTb7n4hO2bNT8YWw9W
52ouc8hnRP9mK69US9Wkte0Bm1cJWhXJ6t3aL7rxb7mexyHevbB3Bl9iSe40YlekAoVaQe0jJnYs
NCeI8dzT7o9snVLEajfbJpJIYZ6gtdZt8R0DNZJC0xCcAObJdlztiNyvjT4tNw8FwIW9N3ZJLFto
4Oumwdud5oSgSASeuOZZhSG08JbCU8gB6njN69D0BySpzJbsehmtGSP7OLhdkYUQLvX78yS81/8+
X3jhoJkRl3wIaBP5NusI5+M/nCeinw/TPCDaPWqjhjK4KMqjH6FgkN1ran9S+Vlu+HoQkiZwG1BQ
6IsfszLJNKLh2NLry7xyX622lhLzWRYfMBEFc6ebudFWpdvy/Pw/NEWlHquKxj9KQeUbRZdVhUbh
T0GbcXeZuGSpXjrWUj7clA+vqJCtuSX0HexaVnNUIObVZbh1wADk5UaUczQPgJ2R/QN5HjcTQWIX
GOZdVXbcOaus0E9NFMfuS0JuS1D9nwT6Ybb6o8kgDHspt9gtNlI5n87FgR8szgNF/e/70BboBFqf
MgTa5UA9sSzSZ0X6NiltfXCb90T/DfIDlD0HZByC5u6fsuWVoWc++leM5NKfXSc/E07l9rHV7sc0
s8+d2TdGsVEVmnU/yCVSbAJEHGP332OOb5DBuTswfh7RoU5O68Lz6KIk5SUNJ/tBahzLCCADVcbg
arRjDdkHzINSdGfPH8yx25PVXU1f02GucwPny1Y/B7zO098VO0Q6q9CoUeGc2++tgAboDw7RfQXg
pVUbIWo5aIG614f4IOgxaWS4nx/IKievarv8RBbUD9BX+ALU701xu8nKsR2xq0hjHPEmtnq7pTIW
QkGQSgR4rEUJlg52cR/Zy01+Ydk2fWzhdNzU2g56W2V8EoDaLPQo/lY3gdwSLIMjG8dplARhpzJh
nq2KafltM8HNaBn2TU9HaQSFmmHJMdhJAUSzYkpFL5GWbaK/3r8IlVCQn/yLr9M3P1KbWf+e5K46
oGsFFa0MGxg7HZZXIij/ztZ1haq8TPAN+fUJ4BNLELyti8MxGbjKXFZms8Qpnd3M1+cgLS1vTqTa
MW8QCqZ44qr+93tgCOs0/Oy3hYvXU+yHHsMRFtKOyWgDdxsSn9hxwf24zbxDnSJOlFWJSzThibY2
tPRvP344npGQE4iq09pol1x6WBdkXHVlf9GwGlMPIofsuN3Hb4KXh7mkNNqjtH0iifKJe9SWat4o
YKlalF2T6MNzI8a+NrxoyU2Ih8RtwE5yNPZUlhQE5NYKc08PM6LslFdf+VnBYbumwUgfJgBtxkUS
apIPesmLVc6TjzF9seHzWF7F8UWIfk5MuTB8uN1Pdz5rUSWEDI0q56eOkqSwbYotmczFfJHc16ln
Q4iEEGQvWJYCPhxAE5G1oIVxaAN5JLt5dPM8sv7lyS1AP4EIFAM4OfslaMu7X8SKuWuo4G5FFEn5
sR5N/7CYwi1VSi3Nvop9pxLgM+iQ95At2482zkqwnX6IVoWUqteaWNUBN5DSSbH8Ykb5DruqHnjX
8up59pPGYP2CIskT5Y/B30oACsjDZt/1FvsLPUqqTwrdtAJVH9hbCheWSob/zFkv3MxuLoy+fHuD
WH6FZJQGSW8TymFbcc1w+buzmWMeXp/cu/iRT/i6W1yioDrAMvN+MCy09fRdNR6u92GmNB6C5Qy4
WNiX+WfZ7nCHoRMtUIn21V3rveBZu0Bi6OG1UME0KjWbRX1bUzj4oCBicpegAhnB+b5nGyVSAB0c
xs7LEAkIIfVVk16/zBwafvyR8hyMsGu6Ln6D35haUmz61RCHcKOKTwcGNQwTOgJS/0fbZXIjlvaj
dX2A1Id5NeHdr2Uf4e6ZS+eEdzPAPqhaLRXfz80SziUrBNUMKMLKASz+yS57fAIyGqASZrI1Ib1g
ZOlPp67V5o4Q5IOG5BFjHJLiR8wtrmeNsKPgmuGm6hM7ANiW04QurWUpM5Yzrg0nXNeUz/LghjGJ
2v/h1DNjBpBY5b+62rupCKxaq1c5IPbBz7IVwKD6bZGvuKgCFWTgXTfqYnc+HTgNus7jDnSKSuQb
HsWvR7N+1Rj72qkP+yB1IIS6jSvh2KxkDdNZgBQADipwQCYOfxp7I6tzH3NSFGisF358+NfGRPRd
cTQjUEboqsKNXFK3AlnpYMz0hZbxVgJrrx79SYVTkVG9oo32/TD7YGiB5sKprlJ9rWMigiYSoEIm
5UqsggVFj6SiPeCfWU/9Euo1GwU/9h5sQqTJtVyBJNAqMNVy3NIr+5VX5Jw5YUkjdR4QYxk/6FGz
zqgstFY4lG+uh5rWdwHC8IFhcSCYgIBxs+x7aC9bFnrCSDPVPB8jpow+A6+h3YTmwVKPlItSmaNA
iKVIzETRVA8z0/mMslJB7GsXqBAa5V12s5oUkW8ljKMvyf6EANqlFlOMseFuXEs4rKfibC2xQi2a
gIq+gr8eUT5ojg+gfgucEHBUUsDdRwp+zGYBl8FPYsXMk7V+pB+jMh/cntsjBtLZ0Taoajs7y84r
zGAX0NrDTmoGuxMjBDLXidtqWNHLzalM1IbdQ16NqknIJIevqXpRd6sen+Fqp8EOsnEj5fEMZ9q2
qLl4KiDeGxcDGu+u23NTFZukYI2bOp9a8evLa3FdQWZtnWUJEqZF0rBDVN2afRZGMtiiPCkln7ws
CQazvm4NDKS2QKKRD8JDuwbmVVxOuMnBekEpV02VIgImLdYD0oQ3FxYzokSmUTGUIW1uAuZuEjWb
F7XKTOF2NSRtYEOyVn51McHCbNSZW+LyxHT0bzG/8tmfS3lLxorwVfxO7ewcCqwB84/ceGu1Pm8Y
+uMbidIsBeFC9PjyD2E4M6yUrE7lVSzzcuaUPkbVoEiNR8uVNd4Jiug2/TczV0EsnvW+DE0Gea+F
vCOG53/wKsq05QbhlXxGFR/2vLPPKuSYJbO9wluDRaOzS4owwmB7IFiI89kGLSJIhoK25gdMNW4s
dtwTYk2NuT89qwrtF64HoFQMJOEUgXTfU/yw2iNSEH0fyXE+IogAwWkF9a3G01Xm1OpVCFEXCCm9
mIhUqBPAecsdZ1pTkGYd4H6pgBkRv1SVVfJcHPJMokjNl+ct6zaQ0IRbmvejvK2YPU18n+lL2lYm
UAB4MMLQO1z1ndOHCyPzcnkro+RVsEci59C8BKLnoH6lHQsCDtlaQJI6Q09iSj2/mAhHsJ65iZwP
I4F71s59PKfisEiawnHQAMpw8tVIszxURQUFz+xfB1cQj8lR9C1gnh3Ln0wkP/IJMghopIf2XVl7
KOjWnYmE7Y+IAlslyJKMLsmfRoF4svo444BTF41ub9j8pSvqYp5XVczS8vKVvN4czjX6QEXoOuFc
5E0ZZcPwuvgh3yCpRPTtkdgNOWc+Jn9uWKUIsRGzp2vuCIPqkr9q/i7wnLWLHTaosGPOsmMz0i49
HmQGZHpMHmbf/C5hiQ3eQqBcR/jggx4fmEcNQoTLFFQBQ4f6uTDbNldx0MJAaO4ejqetuxwvKun7
e5O7fbnzf/RrHvNcXEFIStoB15/pbG8vVw9cc9Dwu14OLhMLmRjGE82ZNJz2FMUHopt/FaaVhbYw
tUAS8hT1Hyk+xCQhj8+Itm2HIQzeIDRpGzbHmyqttc+seH2/C2YjR3Dr3O/QMeM7xqp6PczkiW0+
figTc8W76vaEOJtvNPU/re3yXMFnV98hL2iFKd1124yfYP8vvZnV/BoHeQR9RFDn/s0MLGLnzvMe
wN6dM5nOsyo3RThfIclGiUt0zaagdP8P3aDalIsydAZd2ApD1bQsvYQBQNpcD22COadKshhzzNYh
1SloyItWysy8eQ+imvOKHZXuiIdypw/86rpNsDWnHFy4tJQIGb/uUEnoqjlV6EWac0FiHZh5mE9+
NfeA4yBZc7rje4nKNTQhFY/1vSVPxYOOFrLnc7UMu/luNUI8hEpk9Z8YeW5Hgk2/KDk9jakN1jv2
T9iTsSud1x9uBqPc1heJBhzIdOW+x6sg7nA2pdF3VZ/p2gyE4e3bwNcqIy6mfgymlWiwyrC3DqE1
eH5O71p5JYCwFM1LZbmwrVDQUNsDtxZWIiFs9bzJrVohSZ6qWfXkHHpVKrqcOs6+VvjU2OUsb5XA
sXFdhdSgyswqc4eN7iQ2cBOEW8ebJqZSE1s6s6glbUJOW2f6o1nadRf4K/k237jDVAYV9zsEm22Z
IfXGBp8/rolyGX8l/iCuXiq35JsVyFVmXHsQvN9gr+KxFme/JCNjNVZKl6Xm90ufRx2TCr745u5i
QkPsiOvUJSuu9g7/BJ9r7MUDdTj95TMfSAiBZROLNNHVBfTHTWYOYPcXue8GB/5/8JB/+PVm40j1
1EItBdebv+QuO+BrYKfYXiRd7ISQZ6uhKykJ+ONarnI8JcbEIKQEX7MjQMjitEO4ebhtOUd3hFx1
D/HnH+ek8ZaR5vh4bvimYio3QCWPAXrJSjtURUWjMLZRWtJ7svRkhIXov1Y5PY6MSDX04t3/1k43
tHuYXp1+yMHgyXBXxAOBAJehz8pHiPAC2lTbMwERUUGk7eSZ/NNQfJM3wcmA/rpVtnWSjK0ttmWq
dUtk2giMYgOCqH9Ba3TeaPp8hud3rv9TNjsr585aodPAl8q4cPuK29byI83jGUu7g0mYBRu2zGqH
rHfReGifwg14VerHvFZAxBWU4GRdw7NudE6fuslxAgX5uiMAzsJnmlWQFgeHahSj655HlTRpr+rH
MUKA0Qekt1xOAbKH74mcB93l+vTH3W1RUDGFR5zwLS2dhmDzDYEwp6Duoq0kFX7DMTS9KQ7COTCC
V548tcuGTf5ANocfNrF9FnZdR3Ak4h31XP/plmBKgO0RbL7hh9Z3mwSGPuaQ5M4Nf+VzMMaub8S4
/+e3xrBIycmOvYsGvGWpU6uNGAVolKB0AYP5OkveRWkFu9j8H6XFZwgV7VJ5iuuEbBJ6m7yN4xnu
QlOx4Kr0hgLAOUegTDWqD7oCkOc9YRPjJ0Ay7JD410DZTlE4r7joOksDc96ykGevklVp5Y39km1G
ErvTafPbsMli2eD32Qklz/IWU+T/Zf2pvgyTvBzU/8yo8bZAxqfq+g1u0TS0hazSEDL1/I1Yukdc
A/fhEj2CR+GfJbNq/u78qVL1x66ahWDf0I9UCPjyfgDxaP6v2Nw3mmnHGDSBC4FC/R7dfAlW96Y5
tNnUHDael0dSRtpANFCQbR7v5nLHsTcfYJV5A4UNtXJrVyzgfRxQKHkmS5nHTbcCvEG1gjfi0w81
muErQ77wf3c/k7KFPjwOKwcRkEdV9a2+GDCR0EEJ/x5BI2mROdyIFe2psSnyw6bxZfYXYt2tqdak
ThHE2frxkVuyOx40gHTsdaYiHXYqn68BfeYDdTVVDevipBqeNmEoBbKB/1xnDgVM68w4URa2Qsfl
WBSo9cYEZTOvoGlneNdrmzZiEuWaO0ttWhgvquiJF785/RD5/4AjmgXbjt8qRTKdYjnuZvd8rXsb
0+gRBVLwI25l6eMEXe872f8KbEC3noBrjqOz041GDEZxQgy66t6WjXr+vgBhQFWMP3iZVJljKvl3
wu0z+YGuk9+bq2siehVgHM4m8qNzptyojiv4LLyJ1uqXkl8/EaqLc2J+tA140dtzcMsFBlA1Ujzz
63U1CvtKpXSWfEMqSDyn6qezZyh4Amv7HubRQ8fBtiRFX71Wci4KQWwmrEmznGHTa1HvjASHlAXl
n/6QLbbrZJewCFBAtBpkH+X8HIaPry2opoMw4Aoq7M6mt23f7uVc9vM46bUKKGlm9lK1V+Si0Qcd
aj+SKn1eENVV3NV4vHslsPnGFbNwbVSbjIdnVRQd08WRaOO5tQ3ooYF+/EpVNpvIZ/3gYjmg7IFV
rDc+xjj3HbWrKJsJQDC6zRE/2kd0hOmv755fpe70ZEyC+jt6N2oOK4BdZFRE0CHmhJr8WVvxyzLh
b43Ol9HUEXODfH4Xfu4BJeYelTx41EP4cSHiwTb48kr0fdfub3QIPJmInkRwoM0DLYLIFUUGG9yS
oKD1gGr8rt79kGYpsNTp+mhS9C+rXGyXGEK+JSe+Y3NBePsPohJRfM6V1I2yWsK9wgDMjOxDbwKT
kpeM01tObYq+++iCHC5jIE9gdHUCXhDhHOqOpnJKvqlOQY8Jo9UkKgWtDq8Zm0F1wxpnVAuCx9Kk
OloMB4uxLCY5A+FGo/6C3M/ZDY7W1yEcQwRV/MqGLE41KvsuSA80HQr2E9vMcOI9wD+TxywLLMfa
2GSzfqK8mvobd/46bMHN3TT1AylDyCFc4Ev04CGBMcw47fO2gJ4Ekdb9ViWW2YnOssAEKG3FQJbl
L4xVOce+CiBqvTRmY4HD+rLwoQCnOlgmiILEbzc9FQDliaiKvV+6d3ufTSulnCIjTjXJxvdUYowG
VA4c+zC+YH/ucxAsFIs19wB7AieiVuA8iVLhJ0eMd9r6K+RPeg/uCy0HSv74jxCmL7fvhUhkpRqT
WoX9xR8MZbaL6b+EOVdLEdhFdAO56xDOmYIlFw864BOvUa5PiTcm0HEWtwPlky9UEpQP6kmiX+2s
qb0b6qICMGkjN2yCz2dZG5hXAyGOHV95phqZ04J+9ZZGl+tYkat4BolJpmbfHnkB75KvOFI0zAGP
YHwSZU8aRX2gDtohJHdDP5ttXZ5UBNwmSFrTl3n66f9zNsfTgPSbfE1njDjjWk+U5KLOcZpiX94O
VoO9IU9/K2xK5Au8YhnSOzHE0m2BIPO8UKvKOg5QvmAWRcPaoLIWWlb+kR33b+Xw5klxnTrGrUK1
t/JoBrQJHAxnzxqizzNiGc4IKvHOZ9LXMO2VKOyoGd5oqBmwlTrCueZk+9n9T5AiQa3uY+KiKx9I
azvS25YcEaXhykzcxRMnioZwsqB0ORH6oIsQ/5YUtUBJHaWuJZyzSgEQzM94GZPyN6GKnuLdJsR5
8I8udFA9hylayY5KFKUC4hzdYbT3aQkpMv2zlX0YNYviKbGnrMRgMHj8z/ZP/7/YpJHKzFMTR4Mz
Hx4Kvn/cHM3wRjozc5hM9KRxr5FjBz23p9yroljBKg4BMqNpt4q+bfTSoXLW+CsLIeOGubZtPgoj
uxWmfEStIXrgLnAerOAa9JLDGvk2hjFd50QtPxV7I2f2DNlJ0+wQph50VihbWUrhPDWyLE+NtzaH
QzXaIFf25VxQx7hHwkgiiYfkyhw7cz3+UPJcdF5mwGJTHE8RXC42lQMtHqF2yQlgmU0mpNfGGajS
8KjT1roWhhku0u/iyc+qv0Q36JULyF1a7ubtCAXaLCekUTecKP1bYYFQ89hJg1ONgz5i+4BrbgYs
jrXFi+wVAzsYh0fdUR7elSD0vsobZowMq1fEhP07DdC2Y2GM0xqBFAKZUMdxaP5uK66OCL7LnCWH
Fe34YQNLv7SaXevVGjV+p/RR6M8vLmViaQ4L43z72xU3NJ8SfyGnvU5vQOWXwxBrxUO/Y0a4SYXR
MX9xsM2CsHBRsM8XaEhc09FeK1QG2saBBJKaD2WDW5X2peiu7b+Mv/tNqSbMuCGGG37R7XAUHEjs
HYUnxbbQikcEQIRDMUSyedNPErclZpb3oGCD0AHMNQiceXsSgPwp/Xa2Fu4BuVfzEsjNgsvFo6Pq
n26VQ5id/NrCYFvjTJugPv+SPIH0OeMxMxivXfZEeeLQCeYeeVLb1l1pNBPPwo29jnHI2Y62KzeC
Obxs8kIQCtCeLq9paayAv/NkXdjMSc++oRMSLQLBlGJNM9mBe/kNHxtg3MPya4GALfWml+wU8n2y
7Wyrj6HoK9wdHSsDpiQ4KsaFL0LfydWUmYi1VPo7NvoQVNVCtnla2GqjDQh8R0o9MfftgavslptT
ZZ/CPT6HWNFNSn+KAK6dbI5FGSKQgV5iXUsy/vDfQ6XvDC2e80r7G66LIR68GCvHZVZQae05zjkz
lLljg7F1bepR+NAxZotHPTwazhV5MkyI2BwNG/51CbN0BsEnwwAOWlrdPlRPRoVFXgz+nXzkqpmJ
Iyn7nx3ClyqZX+9deExFk9Y92DN+Zr8gZm7r2HUe0YDR0odcydqlUYR56DlnHT7HiKstNicxkvEt
NHkIh/WPIZh5aHesGfxZZCRkxkJ3MaCXpOBxAlIJ5tKL3SNrJ6sxf6jeVCvU3BCL2OihuI1by45P
fCN/jNiaNdA69UYDP8FQWUpO0DZOGQx7TmMh8eRrL6EXG9rJFXEbfysV/ALNv13dKO7MbiaV/QbP
QwpmwwMCtEc+ldyvIR/HJuZBjlfvIaKMfh06HYy32LlPENSOWBSCd+4QbRtAb0v2FX5xnrqThpsJ
rxeTUM/iQdgRWSJX3LPx9F0aU1AIsQAVYOIR2k3PjgoiHgBEPmpfb5mQ6ZCcnO3qNRYpjUY2sSEu
0QjBHpQyznOq2BjEJTEEMlHgNBhKO47tMN+TapUxo4eTHNaYRFg7Um73XK3sQUU+qh9bS4dyvzDX
AfjGLNVh8YMvcatEc/N/TKTC0GcYlfSU1Q65why/rq1jR+qLCUPsNVHGcyDujciiNUZvuVsj31jK
BxQrtPtUFuKL8CFnR/1/9yGYmTtNJS0V6ynN2iWWUR5yYPxm50Ugt1ZC3xBe4wgJkvbZJB0Gmsed
tTpHYF1MIf2CjGl50y85s9J7AbVSgyycrIZkspqVOe8T2VhmYn79Ti6IKhljU4YdPQ0L8QE/qJOo
XEqAttBjbmPzD7P4q7Ukx61vAS3Pn5PcJHqft5XSet6KXx/BTtb4i4sD0Hil3x3COCd2O8lBoo7P
VOxWuAS5GGGfVxW4p5Lk0nNmbnNLrxHIwR+7RzXYwCuf+/H8Xo0obxjH5Zx9yYqNxiTGlQLPXdOA
rMu/KT7R3HUxc09Toh1b/H6E8UkD9UH4xSacyWiHttF1zVQDNux9NNSbfuO3yf+lmpvjiHNoP9XG
DKgRJikyMPobbM8b3nHXpJXoF5Rcmc0QED6hSuhIuBh8cZGjQellXXAiGYcaF5qW05hfKmxEUGk0
YYwP4pLTcJhSjUU8qSahKO2QFpYwl6TjF83DlzMHlYd2VCLT9fVPVr0xrUexkqwirb0u3gnNcGyV
is1w3AMqfAFoBy+RuOYqd4MIE32Y3WEAFwY/OgdQZm9c0pA3jUv3PEZ+g4myOIcHaAeVKD5o+4Wt
JhQsfCFrFEfNmcmTqPPYBL4vNyPgodPbug3sCqFeZbFspdGSMmFzJo4AGiJVIWEkVlGqezK31BMd
ufJTfpKA98ANw1jRCKMpTZz0XN2eQxcHIamV/oYD+hGc5RqLeFmXZPH8K2+2KOWu2PC7FWzUCnmf
lHS0pieqrpHar6vgBNHlwIgGTdh7gXVI3cv+/ZxlVnGMdnMgBtgaMyPg+9a7Tk1M6ih1+tFtZx44
s3ZU9Or3McuDPaw0ih7XG3t2O6wfN+3yv2UOR1AW6TGUv2l3m9zlVvnRHOQdcfF/OM7RMSsNvI6k
RuiGF+g1UJErRNN3EkOL1ewjFQx9SU04etHOPnwz6A5WFBG3mxwrFU1l8P5/b/DzJMONDdm7aatO
YdHo/+EP+lXS0lI1zKIgSY1H9DbC1Co1TwUPiGPE4BjB6n+y/70l3f2YebK6yypDmXYHZMcERuZ0
BBgok3VKgGYrFMpDoOHzo26hCi49Qq5+ij1PZhOYXNgw6XNglzC/VznEk3K0Drrj41TYZlt1MPSf
l8dl0ARkkg5T0SCaX/TKXSMudOpW8q9qBnXPjzR5GB7SNFjTwsjVc837fKnDMx2pOuspjkdnEwON
nl/S8NIzucS4bHLrQ75q8D6NWULWC0/mY05ydlYCRjXY5/2Q+/WzsQLnMdel78jlR7HEaCyM7h3Z
jVZ9D6mGm5u2l6gmyiF+G9Fi+2baSOlzBL2uMgvjHcfBoOKglYgUt4rFuwoP6f6LjQVBhtTIpAKU
Ppq2Ft7rzOObss8KlwDWa+YnQXX8dTSC3fYRWZQKGxCW+6K7Hjt5wZxeYHV5fMkAUnV8b9t24lcZ
D4hV/jOkOA14orYV2mG1xcTiqFKxMCFWZeaHOXbs1IiK8P0UhxVCoQDlMMiQBBYUupTuoGSbThol
FZM+K4Ul0cIWEvW5fvXPTd6LLyfcD20wK3d9hUNfV/DaJd5eh/L/929iSoThw1LP8eyVJxQ0rsec
NG8jdo7MyWLlMqBtRY69m108TllU9vd/bNIpFOfqduMJcOtNj3kHMYvO4RSW4/0GAPP3TxAustp3
x+uxndMuOV7FD1/Ux2WP5385BFPmv+kxxZRCBit82+V7qrg323LXbND+s52NkImtCnnebn9PuNH8
JCDW2gaFTqs71Okl6gjb2L5w4C1I9GvRGA62ziOEWzGPv5JF+Yka31JhionU42g3sveX/f0HIp1M
4sMALkkMFLZvGJy2Ol5NUQKqE2vPvbil2IoT4GsJU2cYq5ZhLjxl2FCtbs0fOYGjeRFpgxtnP4hN
GGtYIUPwF7PNRYrRYJRuIYtk8n56LvLabqtdDymP5gL71EG1FWuLUaOnkxthHeqCDiB8DqsVI85U
CG6wNMun/lhbvZmu/bxjRsLtQme+IWQDw10gA/9pEZ0xIBofzs+pN6YFTqQEN/+MVguAc50jCl8F
gWtPwLZwCRi4MfqpLFq4FixvvkXUuANAM5L336kjMJS/mzUaNaVy0fLcW0ZHke/1ikoZYs1/oDNj
dnvx6xLFXzfDZ8rFxS9waoPj2E7ZAOS3yJgdYlgwQgupYsvyz95fuuFwV9HNvlh7ogNWKdutAPmO
+5TGtZkMBdkp4MIQcUVVHjZmcKBkSJ4kavZ1k876v2sNxC75ia6+aYIuJQTELU2f+2D1oBRgZ4Be
4HxguwIXEgMrlcoLjzxsDnAzrT3zFC3axuFPJTNspTF7PjccAwmPSro3KBlRvUFG128WecMuYZNM
9Tolnr3otBfDOPd2LeD0kbfqt4VZgc/7ZvrerqjloETOB699GwB/eC33fTmIgiK6m20xr3g6JFLO
/gCoB0sS49StRsfXZY+QNpazyaUfkO85/7JVgdkZAL35WjnS4Z3MrpMefW5j7VIFmbI6C5CdNveU
RsYCrgCsOqbrJVErHKMBkdKfmw5ybVgRJuSC6h4zOfjgbDqgZABPGAAomCIGRs/SQfsbMKcbHa1b
Sdfc1fm2sib8Tk+vS6v0qnzNsoTOG4z6JEDhV6IiUtZpkCoS/ZiV5qTvDEIeBk9C47mPaFZEdiSy
jYhLjb3phwdIayeewkU30nnauUN9lyz9d+6EGWHwc9J3cNJoD5nBCY/Iwpec0NBWeiFqXkl08ARj
OjyMtM3TK5nmAaedKFF+oW1C5TaYwV8RwiMmsFXNDniEQZ0Ob7BKkF1rR8Cs6FHB6BUo+rx2jbC8
vGuPLoJR/87Ax/9knprYDqn1JB/fRdeSs9yFZ4ahiGKnhablShU6zXggGjpAqJzXqF2mQgWnu64n
xIXUA19K6WIu//qpq6ALYO7ckM9eqCHLyMEI8sZsvLHOIyc61triz34oGSqzEZ+CzVexh4++kY2W
BuLalH76AclWRZSaZ+XSFsKhuoE6Xm4m3nIaOoR/GtZMjeui/thrt0lbjg6cbYKAueqzcM9SVzD1
6YWW+66MAGr0TQmwjKiv06J63a3ek27KkAyDolTOI2JyDedNWe/CntpbqNPB8jlmYOD1rbwM4NwA
WjWgvBOsDWMD52VlxvuL6XJ4mBpdwRvaNf8UE1uMC/OKkIqayTajEiKWZD5q5geHsVXgJSnL04t2
rOW+VFBMktGndoQRhJiSX7nFqyZYaNcVnTRM0Bixw1EsXWWc0WTjB3raVd6l7X2UWx2pXypkhQ04
ybSBjNHqU3fsGnvet8awBN/Gp/2nI3EHG64y0HKiQ5tu8Yr14ieacFyA/mXnNuYVlmQrIRkj6Ofh
NJ4bC2nQzaQ6gJ8ndB0sBqo6LegJD+4H4fc9QWbBsps2jZ8VqIQinHEvZhq5KBiMpTf5TqOS7+o7
+yyPlakyf2bAVP5+jrMtA13WIBsvb5gS58wS0m2zx+N7JWNMz1tWtk5MTvnVynUrY1GL9djAW3xB
LpZp/zTrXuAAO5I1erD7r7gyp2NiBlJHeDM6CmJXqOkGhZNH9VPiWkDheEiZ8L/O6n5pSCJK5Qxr
xEEppSvlw3WVhvt3E57DQEAiZpmOG4+RuBtaRG4wQTD1S9tdElGKhCXPlVb17YTW7ZgyqHQ+Yncb
Y+/yqamzWL5oJGp4ynXt3NksuTZmdJHY9BekasFqAWJwqRafTO4mb0QG6ibQEtK9KwXikKmH7YZS
eeAGxLkhzt7yDZ4h5LYb8Smp/Hi/TSLaU5PISGVCZCrR1/3szfcPe6LnSOJe5cUoAfSv0e9GlnoB
+TY2zuTlyKZw7QkimhjoZI7EaL9CjrKUlrUYnnyiGOW/CBEawoYV5lHAtB8/F5kJ3R6dOi55doYj
Sp7AMtmMc55RuedDavDcgAGRSaj49QY9Y6dr4DsKqCtgd415fPgFn5ewpD8CTEjuaJDh3KvBgUqE
cUsY3TMOcWnnWw3v2/e3+c1hRmZjM/HrrGUPyW35KFRGqV//cXvPaXqrGzOGMwTkVeMYD8FzrP0J
gJPL768tIjbE0eMyGDdwxIW3vfPOM0uZ8w7X3sqQEKry/GBMsctdhUgi4RSbhkW37duRszHAe3Eg
ciykd96/lBwL/h+YgChkLQee8wASgnAzBABKPrIN+QbznJex+JzgZ6gzQLYRwxiNMLOG+GhYPYe9
m2lUUCA6PP7RhOVaqaR+HhGui0pj3YZNMzGyDhnJBTySasKeevRE2ZZoVSum4S5SsNFFzHVVOXNC
kmlx8h2s2680G3YX3cTm3OW/3eJeKnbyB+eTGQmGs1iy6O9hynqHO9k/OVhEp6sWYaxJTSVn0ZQz
SvR+BG11cfdKDaxG+fdVJ8TwYPznLc3hg4/F9wa8q0FszUVkDRGe298BbqgOQNG8lmkKcIfMizEb
r+Oob4+1PYaiqfrFRT0m6IIUlVjHtYU2ZR49vdIii3qXegKVE7Vf2ilmBuVXRQc1P5+Garh/020q
ioUX5QdY1lWoHGogub0yBT76yNetiHP4qqVKknUiReyG7A+Wyxfk1pdFPIruUMaYbwGPOr6wCGop
1uRb9L9u+bYynPsDEAvbqjwW1lCM6L/mSfXjI41/UQCf0lR8YElqGZKUvZ3nEjIGryoajH1xrZCB
YNMwtieGNfmb3m9jnxDJhxpRolpbxxZe279IfN+q5L6manT08JKiRMC/JACxE2AMWeEQtOIX5HXI
AdzNz5AaHoKTYvOOuBcWV41n/mq2gQWf2zN4Q+I8f/lpcNzh/Vehkyzfwf6zbAcJdBQrvW2xkmtB
wBMxEBRZMPSGGiTUYT6O4A0fgJkA23r2oNYw9RjH6Vk41/G/zrXdgyoBX+SikwKS3AqxVsClvPJM
HldjEiiU36WJKY86RFGyZyXWx2C4g52vm4bs5WOV4dOIxZbhpH/kVA4QaPwuYjTWTzHgUpEqgajN
+RjzsHLXQJqAVjnjWAyw4Eost1WJuePPZqAkSjjO3iMjcqT1jnzICYYXgpKgIB14N5aYc6cwFKqm
L9WcXDIaLLAGex58FU+Yk0KQ0vl6LmiPBNMmf6ywOnbr2/VLmxDheYV3fr2GSxHaxylYh6EKiDgO
WnQvzWbjwo8VM2+HM4cs9pderShalFcOr7YLz35xNyXw1EW7if18GCwestaWolCLA5Hv81eabXC1
aGGoSr/ER6MoSPLxIcGB+Vc+XtQAEb7NIAE+QufUY9ryv1mZv74oowxCYIK2ZxGGU4L/sbvRKQFh
v45c7nf5P/tou2f+b6G/m8Rk3AuKfEFa8xyJkI+kp5oP84H//OuK4HitZWvewLzspCOS6UMCspS7
eDl6Q+bOs9QIfEyqUJDrE8Sl4KZHVcS5+Zzr9q/S0zqJTQZXTlTN0fwN/TmS/2CTO1CNvmp3jgw4
1A2VG2ntX8cfaAtWYpcpDSbC/QLMnoSmEZPzdJ6dhw42fYS3RV9ZKt3cwQwxt+bYtlr9iu19RV5r
LO/t6VX9pHFjU5u9sq+g/nkTaffNnioXCL3rhtfBYpdbFnMdmjrscahGLv2bu83NmBE90FzV5X2I
OPEgmg6kMMrizJMUE2Tfs963EdDDrq2nmeHt16I7iOfQR+4JHLcaYHoP5N/Q6p8tdultxG55rho7
w2e/fydT8c6utF4dajv3j3nRXzvKwA2Ry67KCnXXHgj2J2lrmZeYbjAiFRYh39eVES71yvCEDWZD
wzC8BVh4iMfZ4M3oRkwQhTbU+jbhiwRMRlQVP0a80BhZP+41sVTm/5dHo3JqCSPuA9a9sY4YynUE
fr+8AQVHRGeSlsFdzcruL860n8aucQIphWPft4b8LT2Bsbb2WBcXPhIVy+tYkmEBSWClBleksgmk
vXdLRYvIKQT/GYw4ZlwhooeATf6lddXl9p4iQ3IgNAeuwa0OIkGiJcib6phXzuLd4MsUZESClt1g
qyMpTeOriOgq83K+6rhf6R2Dwk/T3qeeyhw3M7tN4R1QEKdPi55lKUvLB4/4mpvl6jn1TWeFbHeq
xx8HOEk0Z5SgJWgMLkf0WUlTUzZo68tGVK4pzk/CYo7TEpBCz1xeNs5NvsSX6BYPrcOr64evh5eT
2qSbW0BEc1SCRAfw5QQBp9JONKERLsDTi83tgdLVeQvz/q23e7oX36x+004z/ElarSf5VkPr+p/u
UYir2J09ApPXjAe9CVVckoX2vemDZiLBod9wY6Z5H3SPzDFBTRU3QfuR65rZm/1AsEjGoXHHo7uc
M9ZUAAjehMloYHUZUU7zm0HOCZD96NsR9RcIsYtOgdmWyXB0dTDH521uTXni5zNi9RPf9GC/+u/7
OR2TVKoQtvOvWC2g77+tZbCnB/liPyIImKMXP1G722e13fgGY3G2Df4reoa49k1hq5LN5khdHmnW
Qk4HIF/K+wz6G2BXIYEfi3FEVtXxgElGdGmi/ymM+0R7jXDX1dsCaAqFbXg0xm1qak0iitzvUzmQ
/zrjx+jgnz1w8h0gSLms+dz68SvzlR01LnryiJYNbk8v/6x7KsMkndhljwevJitvXBRaxJV7qZti
1yNyssR3D+E1EAwEabePYCWZ9xcQUpWHZ1QK13zHTxRzY/75I/9zGUjTLvZYx6TmPCHMzyEOjSZk
ZTvB6c7S08RFP/lU4wXw/NhRZopTh8QWBxrYZ7Xp/YUweJGUToucf8iba5rFAYbtxpqd6fDxVNoi
ORiQdTfdEZDowoa2lSq7s2pftTei9aZoZzKiEDheehyBxtTa1rnxUIB2rvVo9n3Jr6VI2xIgjCOL
qQd/qW9m9ZeDPXBuqQX/FFtdDlPKbjLmsfXWKMEB41txzfI4aywt8n4Hhd4P2yGXg+3jgstOmyH6
tEpMOzJ8H921vLyXmNnU7seBLfquPbRRS9zIPm6I5Y6xYrLAp1IR31CgmlMhpUnxp+UFrlj77bUw
aIZfmwL3n8+iG9NutaKZWeOL+jWjUFROaRkZ9ODlquNvGAHATq8SWA1ePML/xGxSVaMQu/GbcIT1
T6qEmXX5El4/HwKeTUU0wNEGHY32Zs6ru22kK2DtfL24Ckf7s7Kzo+mE3JSyzFBHX6/aoqgDovbD
vD8HrM4fjUyngZx8HdoHJiNr7TYP3OnmI+3eOUB41XCTAvsAW6tBTNVKKIHq/Arcq2L1PGgGdwdr
8QBF14xs5RTpmA5yZBP1hrKmM1JSA++J2d7S6jo9cXmlNdVbrFRSrUBlwcBmfVoncEaZnaeOq6ty
Od2Eg/YP94LjBL83ljRpiOl+m1WrW0f7kB8VBdlV657Lj8GY9yI2rXD1rLJtPOXYgQdiKr1K+l+s
8fgeUbUVV02owZkPY0H042mav4WHpTKjj2C4iqA+fXpUh+sW5vuxp5KKbejoCH7CYjig7+niAXRz
WfNMTUrs6qt2VfCLX8gwxASE8eZwim8/D0VY7FdDnwb2BE1xAVJaRU7DL8E7MK8CsciQckDGtrJQ
ZXY3PlXMdlWfzKunIMlWoIJtchTFPQr2QUpQz1O6BMX7lsWJSCoEhLsSklq5++KKItwKzzkyuDcU
btMSU4trocEEyYxY1VRtMpIgSmYyzTwm6EpaMJmnWOXzwlcKPSchJdmrZhwIwbjxRy811x93KPOr
ljBPA5u8WHP9Id5Ua2TAsfiyPJjfQLmw8PprNK2YMsosj+DvW4oDw5fpDFT94KeHgBxQzBCb+uQX
XwVeAsjWEgmonFXc3vyE5WVKZeYHcOsSeXqUDzGDT3SaJ4yo37c+vzv7oRdPgdK52xaDLzJ2Q/wH
WRzGZZnas6lG5lbcdViz+Ii3Td+PMPoXUnTsm3/b9Th7ddSe6MzIrZkzdCmb3yrmv930lRnQsSk5
T4ZrEQVYAmCVJGLrDJDpdLU3gr5nki2qp2w9v/14D2B402qdHw3Q4TyTSqPMJqc8sHbt+nttdwld
1/+B8TucE+pR4oe+2rAmRfzNzsOQ0LrzugiLlA6aZVKAM3ML6Y0nfFws9a0LSj7tE1uvZenTFmSu
XS2s1SPV7Aiv5oelTXNmJkhN0KuCO17FQCAg9fiCvCysAAAXp564t3DkM1inRMxz9yzVoBG9IjkU
vmou0aXERfyrpqhI9RoTewOP4ohbtl9mniijXvcDXoGfqXWofLKFgKoRvYACDEeUimo5ybH+Rvc6
5UQwqih8sW5R+l8LrtvRBXXPgWRYV8jJ0E3swYpgxFSrSZm748tYWre5ybvPAKYFw40P4Pbl/GrC
z4eYav6NCegtr6OmOoHrxPRCtnuNi05rFH1nTQTys0FiqSwkQ5q3XPDFCwwPMP8uO7CBMApkyQmA
oEIzyXS7undlaMGCOcVxli16bNtveamRmU/YmcXdrZEuri26tMtQX33ZD7cbfVk/W7pzc4UQQ6pX
/LEc+88t//8PcDw4gLddmbwjnNgk6CG+noRrc/KjHs+zOkT1GKw1xoBwTLlrZkbn+EeDN5T3V5xJ
jUgzHnHphHDmsr0kh1Z580UhjLGRMTg+E3ql7isECMM5F2yHd/ackQSgaDw6807fL2bxaxGn1Kty
OEqdwpQPpzPsON6tjZSYnkf8/KHbT47fRDM0LyUmqNmsgFFtsuBCsHin2CTEs+iXhlbDpe2hIRym
72IxSQaoUSKM8Sp2FjHdJiNKuHJ5uu6QqcMfa2zh3Xm8NrWYn1r0SFTuRhGwexxL1zf4JW1lt4NU
00HISie5BMgIL8eNgCXKo1k2CBLxd8FDU4y7DXLd4VHb77Bm2p+ZTsWeqdT4LNEnbRJIgiOeINq3
ZBUjwHN58Ox5eP5u3eYI8eGsE9Y4nRjnk3QpQj8SIE9qy6P+jjjvdWhxkkKEDE/XzFXa27zRDDyd
UKXTaEqJtu1N6NdoU0HgSZysht8lNZ+3S1ZYWX9/LBzFd1JXohn+mq3BP9CcYfPG5GTZH4vFyS7h
LbEJTVKnFd/MCd7EexkPnUilCvE+9j1RxepTdNXQnrE4UMWYuJN7vqxGykauzeLZv0tAnHXhQ8f4
/ZYGt+8907C2yA3lPC0ARu6cVP4yEi830dLlnyNPEnjuMhQM/W1gk/EZ9Fx8Nib+S4DDjYszxV1e
A7hYC3DUtzgYnIyx8jJhwSd2p20S5KvgKQchwwVDvGcpZxATStp8eAIPyGzg0ybWAeGmGtTA31mG
C6Ig1jsZhcpvm6/kcOi7HFB1OsGrqlRk7NGDbrMO5GanWEmJjmuSRy09ZfM0fh1mr/t7xvdlELWT
PM4qaXmfy1xqXhu76EbeNmfvzPzl+fpVjZLhEDtBzvxlLPZcrRGj0wRZodaah8XJFOlPrTeiJF7i
u1RRrslyT/m10gvDjOINpRd3D2sfvmHY/biYJa9vq5rtdG8Rsvrli8DkW8urRcjR6hSp8AGJn2IB
tN8LoqFgCd5eaDBJ1ORWQURGOgoEdGCKmRy2ttkL6AlX2HCxbwonK4itUF67yQ/xgKbVrY0LebkB
iab+eXQGOyoornSf1bBTyHYrhaqF8GZsRh9V4fAFNKwHqxNEnq4knus9OVfZ+BAQ0TaCq1KSi5OU
oXbEie1iEFHEirSpF0zaz3G1hiLxQmwNQZvd8iK1A+PL0UZ79QyAJYU7l/ukHDFeUkhJHssxLGbB
4OO5dWHAgH9/A18D6pBZQVCzFjAC/HH4C7QsckhW70JTA74Oa1QpTgxXujZqlIJBRAau/CO3vNij
M/iVjo4l8NHpWRjcTmFiO60+k2c9iOyu1TSfB0tkU460rG0NhrZC6o9jXzhDOcoZprq8R9ajOZnB
A2/FbXH7Z2vzQcq9/A4uKZnwEyOqMBxwsxwbKd+aIBkGm6MueMHSSTB5B1CKHIsrTx6WYzTyKL+i
JgZi9qAFNhoDYqVUy/GwC/Bc63dc7pK5Wh334VGtg3GOwoO9TMuZ6eO9DUPkiG3YaCBNbzKa19Ho
hZvr2wjpWGLVfuvXQVqlSuqEHn3GSBlXSU2bJT7P4K4ZOCsVnW71JoT0Mh9Xj2782D0Fx/pVgcug
Umc1NcIMuMxtbxOf6lINyobZ+O0BhohS8ZGj4a+kM2V7giaxQNKuJdspCxockotzOuEkZUxYjaWb
9zpTz7OxXKEmNHMQRfL3FjSvrtg7DNRQf8s7eYpsiQlgug8f3dE1NKFGgmf1w9KUVbhMDMpQjoOv
1K4MM8A1JXJ7hELXbsiFrfeIMa8hRXvH0LSJUMjL4bZv4BGl/9maFeCrltGgUy7owhU/PCyLyqPD
/tlrd3RBhh8t/Sgbcz1X7m/Td+49KkUAPqWZ+/05F2IFdC/wHtSqxnj5bc5iDm4SzmxCwBpsljh3
SSrS3ccKLEfAgCJu5lE3JRhMedGEU994FulP9y8ekEI7aIb6mnUNKx/qsjkcmi058ApX9GGo3s1+
4U28nWEzBBu6KCnSFNmASIAHnhRX3CJ1mg/PnCgMkfBat4+gmCYCh8+Z2dWSAIjtB8r4Iy8L8rWn
ZwBM/7BUvRsoO63pEogmdrhrruBmGYR1j2Yz9J9wZgbCDllKzrq/whAJC1vyl89wQKhC/V7pQIAa
zEEwqKcdW7Sm/fR7E3T8eMiB/ladje9oVunPkCrjhl6Dwc75uw2QNxk+4M0rblRplp3QQMJq5j/+
SRDYP+cnRyBAcjFEZVYn1EIF380ARe10FJGlUy7jWbtBvLFszbyC27SJvaqkk493eGNQ3GTBKEah
ro8l8DKnwZ93SmpTLp32qPHGeRdXuU98BnbfBYZjk2z88u9jMhSY0/5GkKTwZsfk0AoKkq/DyRAr
z/Q1FxDNCcS+5ISdkT8SPkrVWfYNoo8Qem+unWbcTuvzxdSH7ujHJ925VbB41tqGC6fG2kJQ7L4d
BFYDBDIt5xV8GXCnomFoUwBabSsr7CjaSKzddJ2pGtEUHGccPMudVRCxz303/PJpUwBT86+PPgto
XuIHY1FSCMjHyb0KJaoM1xYnJWnxOZiY8gwA2HBA71c9RetdcsS5W6bmWWmpXhyRqP+C45lO8u/k
o6wZR7eOhL/4fOu7V1ITmGG+a5jE9nmGbpSZSJlpxar1Ng1QSbJNQ1wsCn3yRiHRrW0j9QeARKI0
HbFMMWHlby1nxac6e/5LHp2QQHaqelGFOoHyhY0HDaaMEWktW2iQ02A7Go9cW6EdUxQRJ8HGGPyI
l8vhuHeoKvvdmITG1+a4vFLgopkTzj0dhaSdSB5tp9IjYVT8MNExMiX+at2a/CYHbKdwhGGl7zz4
5eZ+F4pMPtZEtqWPX7YetTXYdcPUglAEZjlmmpYEQOwkzBksbYhX4keDnUKawYzblgapq6W3kc5Q
ae0GYtkU9WHiyNaPZA8Cp1D6u9P7LKN0aLgi+xehNbajQOqJmTVe2MCM6I2VgZvWRsynRvPhiSCR
+0vgZsM+c7BhZioPFP4UvHf1KjXv60aAFVK1jfvm4kjxh+DsmKDIrh9eCHBGit6ZCDRCpyqSzV2E
JainmWDNvY9MjUiXHWNgehf71qAGTSN1qUwFFH2fgEyG8d5STg8QCf5BaRQ1+/CPbnZI245Ayvis
VLJR+UFolFO9EVGc9qaSiB7uitEnDgGNJpDs299YPBiWum+DhQqN/chbxHT/3VwUYel5dDcgrRwv
HBF4IwuBoJxX/lbWAG2LNZFj62UMrwSeMwC++ImqIRptUQerD8RuK1lrE7Ibh5yeYtiqbfsk5AA5
VaAaTgaPZJQKRI1BuFItlDCufge1Ij0DBxb/WEWJAUpREI645Im3KPAiO9R/lKSXIAvijjJcu9iX
HfZ0NvVAUtHSSx/URr2+FUUjgMZXQ1Pz4K92yFIktZq4F6eqxrqfFL8jEWblFxiKBMINGmxr7l2p
WQd+Dun9olZ1D522DhZpEhesdfTnTgg8psFMZh8xw63zLSha9romz7WFQRKbBnoCpmCtGpXDphqt
Mi/xmn2qQIXkSfGWbWnT2syDF0vFmrWXLFFchYLVj4yRisspifjk7OBozu3kYpiWE258cgVd6mew
h674deXLLI+iYI+0yXtrrfXedq7i6v0L1snCu/hxOEfe09pLA5MWucPPpD7yddTjcj6l8t/uebxL
WEbEEq3lYxihyg5DLXpClZsogdj2kxLVNgPE1SuRHsDxhR4HE9d04LC2/cdfLNWjMm3OI10C26n1
xDdyDQC72oohWRfySrV6UGzkpL9zxV9O4izyCAcJ2b3Femo0m694SjoOR36uPkq7HPhtixmVqYPk
IZDeqjfOUxa2paO7fq7tc/O6YFnVl+SmHUXny7baG2R9cy8yehpVWYfBYyzzzLpsngsaFEgbGXeF
65xMI+WQUYsimtYVhONOXzTa92srEXfHMsdE1GuU8QwPzcJQRZw3v9/WeeP3igS7fAQUsSPFzqPk
y+ENPGYZAx+ulqEtAhWr6IzVPG99hFTIAdJ04OfZYV4bQQ2GKAqV4h7qFJyvJ6s6O8k1KBRBzgqm
VEQ/jvU/HIGkeGEblSXaj7rjhreMU+H0j4Hq7NXPNt5wl7v6t/M7vhvRZGG6R+VyguG6O3dnxwaT
WlVTY3d4SSVaSdKWNOnwcl09cK1xdJdIr3+a4bp/p9mrrNpWHsacbuqM10A4YrVpsldhBXQLiN+P
x6XT1kJgifRCJfq+VdmZJRz2SezT5ykNjve24/+pDizy66gM5lS/mracNHA7cZ8bSBX4vdUklxYP
IkM/i9S/TtJsvHniFjpdwtPSxavu+dyaIGEQIbgY4EP0MEjr5YPqmBJiiPJnOpI3C8lmvysQUkBP
mfD/R8D3wjUpYBXQ31Q8K+280Tz8Dhw2QUCsRwO5aXKpkM/uH0i5ieBa7U3KW8IeVPRynf/nIoa2
d7BQekmvFuizqwaSKIPMDvdTwyPX+TFZy2+LMALuV2gp8tZ32VTRwnJZwnE1Jqq/2ABLy6Jb71oK
qD7xg2qw0tN0WLYMWmNw2YPmnuvOR1uKK8Tk/F1ArT/Owvby+yZlCfMQyXKphX48QICFM1h9fzIZ
zv3HJ4KgYg8FuXVr1TDkn7ECzaZlGIMIaBvt8O0JR3oopA357akPFIT5tcxpP4cPc/XwwejdsbXi
uRkoZOth5zbIM3copGXhAn+kIwaqj90f7D6SEA6hqvZrgLKGjRYegP2ZsvjjnsgWNU/LG+UWD0Kl
QM/QsUsXD09gO8mCf6ufSOIqTP9qUlxKVwvFHH9sszIxt68SkQXTOnS9YKqxqy65bTZxe/hZIDUF
QZgDCHHLGJ8zPtg0gJVoNeqFeKcWEsys9QE4qTnNdBNCRxua00RyBuTHUCQYcyBpTeKATcWnu7rt
21EtnUhOhzF3oBwvrD4sLYGabfeoQTJkBps2R/pRtGlOrWCc0gcthPPnvZWM5woUEs+wpkMTJfEI
aZ9FWRZH3yZoEp1/KTmR4xViwwG7AkeLjqre80+T/Uz5RbLx/EEN1H5uedl33jfvDZCebNOStBbJ
JNFYPCC3ivMtuPMMSVv21isXiaPQNdcDAqR60yvGh1FQBlPHZODQslNOSDH7jSkt8OzipNkHr5/f
DcntusYuMJI9h+ry9LlBuzIhhY2aeqajuWAXXU+GNgsXp9dpaS4qBAtFfULA65VWT7MzJx22uAzB
f4VVBLFTGTCQxuLu3H6uU8U/7Ehc4M4vckKrjTN71uqQ/D5xFlpCzhdHM0fRgPZ9tw7RtTyuhxn6
BThgV4oCYRkr162iC4CWbHXhyu/KmEqNERb9/39m0DCYTHWVkMlF30FhVym1rQmT8XWj9IYJRLOn
jaJ8lZp6P7+EBMkPnETH4o/DUNUhYKtQPqcjEkpj6iE7g+YTrrv/zxuHdkhB3EXsH9zzotCnm9qb
oF84edMNCizoLZ+D2KuSTZR+PxqQCO7iJCHvdkPNS5L82Ae34soYtok2bVuIcEYXU0fnFLrBPqF6
TMt7YLlxoUe1yJ9tXU1rHDP7DOGuavHT5Acee8HMDwIm4o28XONY1BPsSMuIKxC7UAC7uc11HHXO
dSbKHj4KT8uq8MnFUEnFO+DlMiVeF+fT4lUIoh2oSvJs6nhsLrXKbEsAOm0AkQOpJQrMyEs/PONj
xh0qRYLOZdAFsDj2JkBi8T6oRbe/sVTZcMgHvxNAsG37BdNtkNjE+ss8WH/kxoLY6OgVZSVxlCJI
kC3Lsu/1TV8I0S88TU69IUF3VhbgilqLJ2/b9j16tigoYLoeypHmqrM5hAOawKQ2AoQDVzqpWaX3
DZBXj8UuuVYOijQDZh2uq5CJgkbClINqp/9Xq8mE5ALNdGu3N1v7KQ6iQPW1uqR5gBHloZ6bBDyX
BBHrNjCJ9gutbj9casGkwLSzI8kSpRb41EWJdt1vuZhTNkIKTy5RY5WmQlCnphgqYgn/6Cx+Vwcz
4XYIDPnULuxeM+eomLFRqDooU4L4prg/blbosLGpPwNjb5cWWzNAookx2w+NVMGcwb5qHzSyETlu
LaULkT9iI3EcAtE65WtDwSbMuF//V7CtPAo9rlvJwtAgq8JCdirJ/63K+UdGwSs4RMHHAxxY7IG7
jSkWzNTttShlJISDW3npBwSRACLgePq0MrbHYRJhjcnVXKqo61kMfewuq8+Ti87iep7a0tBzLbMY
OOC0SSh8oW2NesxRbiyrrMx4RAaqYADdL4d472+tJiR96aJ0QtjhvcoviHCRIRLQjWVGT+e1YBhl
Jkvu0ENTtv2ly4tTDFPdfD343M3NH1CzfKGT4H2fyDNVLlinV9OismYGMgfL690ugAQwQFeU57M0
E21tpcqAtKn7bMKVX+besJ8ImmsFzSAzbaPC4OIympvNP8KEsPYqqZU1Sr2GdgFe7fz+M5dltj+2
JR9XqsFpyXUYdJFXZQ6Q4Yd3c4PW3NtkL1GtflZlqmq7RUgYj2UpOVbYn+AOGaPFaxL6dKcpMf8o
e8xhWlfzRdCB5xtLDYlpUub4+OUtRaeHNAlHDRgv8OFQmlkDnTZrKgo4xwVlj96uv7FINmbEVLFS
F/EJXXLx5VPYAXQTEj4NIfLrysNXsC9xIma4i6Qif8ss8B8L6oASSqJ93KeiI1ARLrEUQ2SCfd7b
QxKluISyN2far+pIzdZVHQ7cs6QNdSAZ1xBXpPtVaWT+RP+JICSy/xL5zjqyusfhibVRYmfmgz1t
oP0HtTdDgm31u/tFS+BsJCh0wQh2IWUXCR6k65KPakRRHvhw3xUC0+4mkW+PMfTReQbuXQGjT5Iu
hT86qvCf5Z8RHsZ7cUpZkoEEPnB5yM7oXKmcSkcRoIFPKNbYKwsIbSghpTCy1yw3FuSbqsBVXZKf
6ISichsjUdJGHGiL2o6y/bdrgTHeVsHLqOkTpYdejvZuFp4XJxj5R53wHPwhYQP1iCFDJ0S6Cef7
35RXpSrpG5Wc3JTFxjNpzNUWvIbquI4hHl+3nlHAf2HFaCTY7/ZtyjRh5TWy5aRBJOgCT3gzzFl9
DXBrIkcR3JK3iqzT9kEA5uu/oF25f8fjTd3ZzdjMOwxnz3gwZe/C0JuhQxv+00NVrHer7H61dB3Y
JeHTA4ReLm2ZjH3Ujjx8bAF7vH5sgyuNkDNthp7BlIkvwVJJ9Cf1z+L1CiCOMbh4whVzydLjDGH6
4xFPaLfME3Y7TmVbNuI3yzkWwVuVETvkrvD/S0dF+53zuQs/fxetal69DEDRS/+NuYW3VpBp2q8y
wcEyf3zTMpVUIorW8RpG9iCxaGlfRc97K4N4G/HkAj4PS/R6AUQc8vf5yOMXONPU7JhD1/+2IMrC
i1cFqkfjKZcukTP8nhlTz3aIRhHjCiMCzBQ+Jy+7VIcY3/ai6jAuxJLo1Q6RTaJK1VbeH0rFU8Xm
oLj15skMaJqDiA2PD1GHc6+euUn7rVlc2d7mMzn/pIYB7swQo3/C00b23rhuI3UxbeqHHuCrmb/v
BL1vSBahLA9WLV51PZ5qTVNlmse/xjCC11vnxr6ENT8Qv1No99OntUzm7zBMqIAHhhwURLoIZhvZ
3zZXYQEiLb2RnbQsQyILBAYGRCiX4ziuR42duiMp5RFr20GLPSSgrqutkACelSzE5ZmRjJprR8hU
ZMCn1Ud6p08nt5JL0kTl4TlwyVmunKYRlz5jwS4s5v7tIekSa2VPFvunaXUzzKLYU9hriCa3eeRR
QP+Z7tuVSs0ci7ynKtQRq4dbo7O16OxyNL0rv6oKE8YtxvIFCQnpj/I0jt2qtk0Nu3pEX389jpAl
9pRu0yzPRi/MAGHBCKRsxRDz23SsP0svlaw9e2sllX93i/FObaIgakF/AErWqtipE/P+X/xqSxYg
SCwO2QVBe2Z/d4xCFcTjVdJe+aXZfrsHMbQssaYnjru47LrFwubxzi7yIW7mt6KapAwb21KKDJkR
zJh2NUe4SQetfYv+XzNn0m//7TBRxMotqYR6bq3UZoEhMVNBKxS6Qm9vgnnUab79yY0vn+mG7Aal
GEquQxNsviq2QEGF7hhUSQU4xwoJuqPxIkC4FTk/bijxBKeFqQPsW1xAD4EJyEIrkCwDq9pVHwzr
oaGD5Rg6062btX43idB0hAQjetF20dXT8k7A3K/Kmz+mnGUosYJoDgkyG7fhOcePXFYd2ceV7MWc
CNRb2dXdquZFv69NhfJZhlDClk6fvI7aG676VAiR1nvFCqndqJXhPreqNAIJGwYHybCQF6fd531l
BK45z4c5HN9JPLMWM6U4WgoozRni5HzdOSM/ClZoa462GRtT8h4XoDp8QpmXEFqTQT95J6/szniR
l32LWTDfnKB0Z1Lt3qqS5MfaQqRiWzr3Vtl07vAMMzqcALYJ6wttjBuimNFKUHruLIqgmLQxrbnf
2wbpR/1utdpnwkRHHQ2qj/sdE/7LsghRVPMrcFC7BUMNn25ygTEmgYr4QCHQTBVrGCkXfIOSWOXW
YmXEzE6RTzz5Ow6p/X5vqwshzwHDbWFXoyipifg8tLdc+vKQX7fDjPRNnOaDc6EJzJsei9ZmcDl3
pGp/ofEayt2txyUvJaCXufgObE/pZ7rtPmKd6ElxLuY9IwIPXQc0AUuV51T/qowXHarUYIACrMeA
IvirQzb2QdRQ+cJNJxCxO6LjUpeILpGqVGUm3Ah+OSDy00cfZr4/8hTGBP6ar1Xwi5Z7kEmBpxs1
oH65z5R02u+I0Jc/FuZjhzDZGMb4/JVbArOArsZDOiL+3zF93KftMQAr/izBWGpqFnvr3zUHPOIh
jxCirD1s3lBG9vTPf4sHx9RKIN4U8ixSxR4qQ+BflJqF+AnNak8H35mXnio9rVNWy77xGBBA4AW1
YKdB8dtijvp1P3SgUA5/9gB0nXmI1K6O61P+h0QsVaVFTZ0xpNMDWJ8dn0MqjoIg3oNOH3lvwOOj
aINRYmUM89vYY87aIJ6GW6OYGYxmJbOzSL/K8T3eZ6Xxe+bQ4Hs0+bYyC4lWNT0YPwUniCqVtdgP
14gPe8adyZid+EGLA5a7Av48WYkrkTCBmt//9kQ4eOfimIiH5eICId7V7MI6UYSGd5uMV36xiEB/
HKHGY0RS8aftfke+YYkidddnZnrfEC32e9Im8Wg7q8d9R0LCEEJwFI/c0b0CvN8osMuB0DXNxwFx
mWs7LhYxlSbY/IRa7P8+cMBIlYVb/LnxTyAHMrG2rgXU/WA/yfABemjgxA/Q6KClZgOp2/XPqWte
/dcANcNybvm8PkQeEqZIT6iFP9MzWijbNEek8HSpc9dYMIP0ELcG/JJpe6uZON1+/hqV2IAfhm19
CzZKp3DYLLY6pz641Fcd909Byj0Rc9HyxnEvlObXhzef8r/p42hwdDC1uRs9Zltvp9HkGZqTQHiD
qWhQ/H0EZLEjg99tOgxPb2kCID8msIQhpsijiOEaeYwxGJon60jhCVxC4f3XxsWzK2B6nI3M2s05
08S3xR1l+K+UWOwNvp82t6BmoUAlvQ9f1HTdnpgiOsJ1NtGa4X0uFMQr5HfmDbQES5/oCmKVJBki
EVFr9d2JgmcjNtxcN4fH5rXrHvtJE2+LNjq31o8Ii/u/e7mzEgecA8Xg3WmhD6hFGR+OT/b1kkTb
jvzQqIOowj1EYX66yEB3rQRdhY9n8QXHnz5iKK9+6kJURfdgAYGdYG12YM449HM+MxrWYdYLxE+q
+R1fq/OhW1Q+NQvT+Ablp5mdJy1U3if7aa/QuQPWcioc+MrXydcBphSLG74WXxtuaTrMtzxhICuU
g0DRJzciXSmk8KRr+HLYP+DI9azkV8M+Jza8rMPzEpqg4pbEAuCRVtncTWiXssCUI2AIKrC6dk5G
aVKkzeG1J6W9NQ+DqsdXlJA5j0i1xn3SHhlCKL8ith4mVJxEelrHcMGE+xv6pda7EZ97p3yIuwAF
7l9vYfCiycQK44y0ky2XavWlAwielL7cvbr+vGsZ2yWfe5zcZWo2NpsrXvtsxaxwRmJXcS1SzGHc
0uZYXghAm4YuLpTY/c85dOTg9UV9+D8U+CDoyDUI2mkQVBSPQtjMclrxUeczjTqsCIsWapGwqR6c
804pyw1jg2jh9EYlx9fKCJTSZP8+BChQyKk7Z+UdsulS7Qzk322lDjoMFKsUtfNC7pa06go/Pmqd
qniqSQ2CuUHi34orc66kGm2zIdIOpCHLq13P7fCLgyUYj9vkWrwCzYWxn2sNTjdDkEP4n5wBQJfM
iWtzZFmJXAIkfS7wJaHJSegbENuvCZHM7c4spVow0aXqc55PauBcn5PUNG1PzFW3ZfTz5ZJLAPrm
Y55R/iNn9fPNrU/VhXHsJ6BabeYwh0oZJbXcbjhT4ADelIf349ECtmPcT1oRoSILvWq4sR4Fb4ZZ
885q5LvIFMsSwJZP5e19ZiITvDjU/VqtFu3Su9mPZHkhdzKEKznckjansBJX5sIUDQHJo/s6qtds
2l5kdDHPZLiVM43svXQPZdV3vUKDzI74VwKer5Q/qMy3sZ1+w3x7xqC4VD0PrGjWfrA4zTc6RPDZ
v68As7vbaXZ/gunnIx4CKqt0FXhOihGzTxMFcfQRugeyX3vQcM+T3D0Cn1GVrpjI470BSces+4M5
aRbCnMdKArIipFx/95KYtQdhDTSzi9KJ3R6NkYJkCCCtGbU1FhBYYYIt93ENcbydzpMSMX+wNbQM
1D1ih8GQtFgRMhPDjdN2rK26M36mww4FODRhXYJdKY0II5Fd/xcetqHMST/BpT4yLgU2AnFSYuNl
Nxfuxy1QaCp8NA6A8XX88O4Qu5q7qyN90FvaUChiw/A/YhMDjiJEhh7CpoA0gLHe9/zgXAcT3qj0
Ftoo2RtggdkKyJqkfudOoj9lgG8azJQNm4T5ifMfilVkmAaaASQ+5zcodmiPOhHU1Hb5uvic2CN6
uQEys6GWWirRX0XtLOA7Wo9Nt4tNxJm2K+qkYekyKk+3DdGDQKpoqfBncTzE8D4yIDdo3tjhp0BT
0+yUWnDfiAHbAGgvSq7airC+EHyvyRsa3BAmr0iaO0NyAYJTVTtZHAAunaSe/6xBNoBcWUsDC82E
hdt9REBghHZKW5jmYFWOhyBdKYpMZRtEleThxTKW/qFhBZPt5wfBBl78lI/0cCkTPXx1eLwA21mh
01ORNBAu+2JRGoF5ACvWeBKicwlaxa/xlxkG1EbJCoWH1W92voVulLbrWyXMeflLlD3EcuHiyMhG
ojnsiHDpZTxf8tdX5dFpkAMBTh62BrS72bhHofZ2BKRdV2b4LI15gyaL6kPDfz8pwSWG9n9YH0J6
ErqqsVwyBV7M6eXbmJHkMMPgasR0F/rWmN7vnS+LPKy+CZFhuG6tXgQp9K8fyJyp1eZInmwwd/oo
NlboiQWZ7AFn0IYXSpI/kAzEna2wfMTnUrabOivPj/SqpBXwL+oFKDzKITvbcu7w4oCJ+jDuwtRT
7rKl9UQbkem50JDhjr7oydojh/Nz5T9JGEDTSqelmedoGgWP4yW086Go3NRqHUlY8Es+u5vx5Ghy
ILgLc8j0lJiI9NEomr1qiAkR0UdALS40FaIFHQAGfFid2Ix33E6JhngaZrEXzxTpyp0hOw1FjgKM
vEhfGM3MWq3B9eTXAY2Xn9Q6ViX3I0v34+GE5rYVq93R0ulz2llIMAfUfBwfY6wZt93BtK2Pr5Dx
K/14rkrvU10lugsunuU+EJdysuDb02dTP+R5mXgsCgCTj5wM0s8V8bxLPEo2fDTrAAlYrOkYbo3z
H6Dyvy0vOvuXiX1ocTGlsZ/2K0FMb+U32wRto4pB+ezn2YFa/meB/wiCeaW1nq1XtasiVz73Nkkc
SZrdQOfBg135lgrTGxc7mGf9ZoNbbv7Rnj3KavzSaZGoWpFeUDXVjV56d1CkIqJzws5d5ZOBpkGQ
keOsaqMA/YrT4jmSdPRr63KPODqSE/hPVep9qXxZ27DtcK90zp4DeqH/KHkqwGf0HH+B3BE09KPs
sgg8s1XFbj+TVQ1I0JSyhYCM+EwBgEZgBZWC8pIkMoe49WwKXoKretn+1+vxpFqDMWnyrs7kMa+T
DfxAJktjtY8fRKcnhqnLfhPCeyHIba3OwaNYsWPvxUxirnNu8nHv1X1z6rg4Us64Jd4S4DM72Ts0
dU619T6u4XYj048/MvF2LuTOmUzT64c8d2auYMZcxdKrk7Tt/kRy2RNfhnC++BdoheRxGD6O5mBz
1d1EdTKzvIUYf2tsqdYxa5Z1AEVe+Lvu39w5lCmt2r7XLiSUjitqbAC6JaW2ZR1+wg7xVNDr78cK
oHrvuqsf9UygOtd0HzchZybHNPrAaj6qa8KWjNetXrROqG6MrkCuV2nCEswH5J+2Ln1jHCNZ7bgd
BPmCbs/vbP1NdVSxWg6GKZN/kqpsmYNQm3jmFrHqS0sWcnsNkfLU4CDdqwL9IW2za58e8G3qosb7
CZAorcnAT7YBpFSNtn40mxHQnad6CG1Mduz0HYEvjmeH00vsGf1UVTgKt9k7pq2va4YkChyMWnQm
zL25RERNYr0jHH5r9Dk/8eorLP9c9tqQx02hoPMLX6zdcBF0QpQfopppl5x1RJQkdTzkxwfTBnuV
wTQ6cdOM2ApBrmmEl9HriHAt4gOykTE0HK/PF3TU4FsNu9VdQkxLzsKDgZ9gSItHpDlYc+8ptSpy
bMuj5e5190Qi7NvTgP3j5PMIkSyRMbvg+HSUdk4MBLhCjVGvpUBg25VtJidGtQOfCrd7TA4fjUJo
wctWU5D6xVsfcd7e+JRW2aX2U6f83/STV+lLqnH6ilJ+52FWUGIp+3rL5dYMj/PGEODQCnKrqnxR
aCstkIIVAAE23U6GVLnIPfHN2gF9+W6zYCKDBGgIdaN4Dp+SQI7tDM12BoAFPjCILqQQilWqRyVG
OpjQcrFpF2Alxv58d9P2n7j0wpZb7q8wNjwlFz3YDISo33zif3rqARPtlyAD3c54zw+iBtbcayCo
RPYB2ZdRvywQd2vS1qWaCRfqOWukEPLwulEMFSfIMBXLn9lVzD1KsHteyA/aHvpjnO48Sy7I0nbO
bO3J/aS28+JMtAHAjaIHIeLzZ7DuYcHLsPFAHYq+zC2Q+9b9uhpw4mpQ4HHI5zF0/LCVZY18ZyCq
nUNTxsetyIml54BcNlwS5J8NGZyVeOsPN/jxt3AhIC+5wApiduUkvXr3+2bLTe/ZVH6KTApBOMcW
CAeL1A6SHYBsUxjCdaxmK3KPbBZ7k8oYjnItlPu+26qJVTw2ZkFZHe+5+O3kKGp3o0jrv5jyS1gj
xGM5T1ZPxQn0hKQLAnLOER49XkkkMCS0eEiox60UTenDE8V8pm1SuLRDHfJ33aHdXyRyEdlKhgAI
1ToY7GjHtkri6Itv0nDuBH+d0pmFgu7sqtwDz+4Vgy1IPnKpn0cnuAjo+HbfDu5y37Gl+yDfdOe3
CMvZcoun0L/hX+SiJNTR5YqOnWNW34WUuuQ+RljocER28EHzH4PR97NjboMsYV/Q0xUnEYk9nGw2
WSgwG0NK69QO6e5OfxkCopHKNWogPsyKuGOuFKOZGghj4o0WMLQvO1N5V6aITT9OPBWouCD7Udw5
yjbQydjrxIy6F5YeO0Vjzz9FXz9jtTp9xnCci0/O77HlUzNNob+rSgX7NKmy73tLSGdFcgqHwdyf
2KCgzlzdjya3GnYAwRFLqHriJQMoDIiSyzls1xGlsA9OEE0uXoCvZr21hTxy7j6JBUVBhy1jUJ7A
A/uZvJSOvbSQth/6v4zsbBqGm7uJaLW7f6FDOmN5YJ14jzOaxdNj/qaXmXXILv3w+6/Iixutwahi
voGKcquaC1r/5IiY41f3VHI4SvTpUFAe5qd7V0JchTJqgSGR8Ku+dIdRWC05fE8TA3GKcIWGB04g
bVrPMeS4QbCfmUVpjlkUPsqbby79nmfRlF7NVSz/vdpOwXCIV2HI0xMrHUA5cocObvaO0V8MOfq1
NqSY47/END3BherbTI+2cPZhhjcD+7PnnnYE5siOYkLRuii5wTgebf2hk1P7052PscJpB0/uGBDe
wx9yl0/X9uGUC9CYgP8HytYu+kbDCwg9MOPUxFnMeWFPofNZ2iNT9y4rJSZWXlV3l8u5aP8ImYtr
CRJSchBrkWGG13IJdYOIfksPIsZOkoaxt+x74cP7Q+vQ2GppAVJKUDUAS6xy2SU0AA2pqsk0HJUs
5V72Mlo1ZhyFBva35wn2piJB8fTejwd0iUnqBANgP0xLjYw+JRnJR9PfBaPqdGUtYw50nSNv7ohj
J/poJRIcDattRQT2HHQH1oP8yj8AlpfYa4A4GM+cXBzV/XfvMrvogwkQD/8/N5+2atupLSjWo9kU
yQv9p4TeYF04qCEL/pZZE6VsrXKCNDA+VpP8x5jyNNB8ZDEIWwFP+eDBtkps3UBJDpaBB+g4rjxn
lHqgdxRVbEiriE/fiIO3zYgqNMxyt/HAMKXZ89tz6UANZE0cJQ+O3m7MUtbfjBcHGR+zTHNnPFXa
Gt3znIb5aiWM8spXxHCyyvVzXmcegcofWsCz+92ku+tQcIY6MT3AgRzAm0xIa5JH4ReTds//8C0e
ac9/9IGyC9Mz9nteRGO6SKEGJHQJL4uY4Kyx3fkdj3hcAdVwxoWczjatLcIa194uOzSINBomiRhe
Vjmklrd3ysSAuGG0Ce3EnbvmpDljPLwjj6k54OxW8Pm4moyAz7/k10HsLfFYB6oLuocLOM6B7KG+
2fqX/Rpr2NCZpcClRujhmGdo6i8GyWIqYhCu4JxxWI/9Gt9RsB1DnSR6lKZQJgqi5rsu5ghdvHnl
Iz0m5TIOEc/UVPumDq/QgAtJCqPRzXydFPw6oRLsnwh5mGrEgDSGEZBW8fRtDGT4hkW1AodbI/kX
n28giTEefaM+M5AAeYeq6y6t2JmTxlPRwjex40Xtu9Np7IKE9VkIA47oiTkoFFT2uMLhs1C1EQBo
IR4+fSvINi4z3Ql9lt+K+puBzEBAe0aiBZnpUylFKYLkl0NQfgiz1ckZvlTjNkuBI9pUlFraxSw+
FcJnos5rUU9L9AX6g3iKg5FnycO80voJZG/c1Yb6FPQ6nweW5KhhJVHQCyon0YVoHgQBWi/1Y/bN
JwaExXE7YS2vj+qH0O8EYJLn/dCM3fdRN6mtbyov+WZEuSGcTy69ymK9RS8EwHVtdsXr4pEts22X
Xf//IuD3w/LspJjCO/pr74BzMNBTnl/dhGVEZasySbIWykGSqgYvUc3k/Mw1XJyxTcZsDNcp7xew
Fce58ofNvYfZ97xiFWKkfUGCkggmLcSi3OdLbBcUANCVFrEI8JALgbi/4V7Id4aDTMhClZEgsK6Y
zIsJIl3XbI5L4rlWTFnSR8nUCf8IhSatKHnHGMKIGIvXGoZkSWfDfNgky4qoUHeDC587Z/+5dO6q
oDKiyI9qinVV8UF+bD8UxicWPaNtFZNapaDwU/JxiB8fNrFBydn5BXnlYqjydb7KIoRaUAcwCOgL
ymzMov0jMPNpkkh+uYUs4m0gqz0NDE61COlllbndEbqfZ3goL0foHq/FHRZddPHmtmUEjf0uccBp
9YhbokM5+N11NCCAyFgKEFrpKU/WaCaolOQfKveDdT57Ygr6BuzSopK0KD6QtMfNrER7/3grDwcu
l7R0j3aMjzTYe7MUuFQ7xf7mngYAirMmvEwbf5RnioANf9cEpoIh+VmqIFoQA5hCG3iVY6if/1sv
HsnK901BgVDb4JPFayICUNr8e8Kp/YEXJW+wmMSTwp5caxwFlH9lZjx8xPxi6Y0MhWWBE2lCEFPM
1o8qUETTmt76HQytlbusoj7dT9miAaoURZPeQIYVLm+YnKOO1DYNkSdTeo27INBCh+pz+0S+QZFP
ovUDuiTvQgFZ/ThWtma4Rf+ivBbDCFl+yKG+t03+RCNc86Qs+PBpDAa0Hm+XolhMGx5wwdLhHh17
CNouz2U0IDi5heMtcRJjcF7RLm1Sx25yRq1VDXCrt7RwUfdOtIUe+luHYKOyzLR1B4ooKjZ0T3Fi
y3qfqnvoHlNFaYpQ5Rhgqh855NfTyiygvDSYCE7lcSgFnq44TtwQfjDkwfaQT8dZ1+kXLFcvWAwM
E9odFHeFqpTJEfe+eDkDI8rlMRhXnFLsUrvIulkkVa/zi2x5+zy7NmfqA+22DdkSYQLcPiIM7eU2
jO4l2ra8E3xeRyCE01I9RhS+u1KC5XJRnBpgtb/K4LzbXApsMWJSrvYVKL8ZxyryTHRD9tXEdn+O
gU6qvqUqL4Ens0EwnobBSz6LiX0RFqknF3S4lzTULyW0XDbfsAwvJAQcYMfV5hDa3Mia77tC9NdZ
yCsfAtd03Kb7nuIKtPuG3Z/AlUGRh+61KbmTbGHqViCc4aNSzBDFMcGKWU6jI80qglHjUdlTqjOW
qeuz1f6zmj4PYwntrdU+YZu/3JBkYzPPN2jKiPrEPKgbFsxkm7H7hCe/Amf59u067SoFiovg2pya
XMGORGoB21FOKbc1cmdei+A56CZWDkvZVA2A8DQw6Qm3jrmq5BjeYZW11gF+KugV3bsH8wxcAE7W
aVbGi0Zv0lKOWiPovWt3h1eS1z02+UdmMBtyeqERFTmi2v+oTiA8Hcze0cWdyPkXI9Rubd2MjxCc
iD3UDbwgKdw83QGUAWquEOqt/qWP6qSHXK2uTCRNwg9A2YSGVlGLMbxY9i9ZFv4k1+3fS/Tk/Oby
s6RRBiKGav8XNx4KLozRGb0na3+i/mzS2aaN0djuw+8Pwjl3fOjcLE/SU7+NtDGR8s+vhSWSk3zl
vccre+YVqJVd7ONoyL2UISgczEX9Gz9TgETkAFUXJmQUCWE4bwuozyedUFGCVDY1l0U3QGHmvGeO
zkPPgK+AeRjDKvCTuLSjEwsCHT0qHqhNrf6nawsugbm6asZNqkOYtsi2DQVKwbNmFNb8F/3Z0Xdy
czTVHA1ODhjBZFDtT1D5+VIXWK5/i6BHtITDJDmM4qGXOTE8qKpjq+ZYGCgWya3oyOcKUcFSUO4K
x1JR7vXjBNvFpss9xEX8DrNqEzOSAHBdT5DWFkZXCYiI0bFxXbiiqtT3DWG2S5xSxSkj8u1BOmC1
0z/x9Xbc47U+r4ciWkpa5iSyWC9UHqgmljjSSN+ijWcE4XxqvB5k8jGQm3UTL+at1L0KdvocHli1
QPBtIZ2ar8IarlVYx8oc+CN5kTkqtj5aVC8U03dCVLE2BNDeTUTgLjhnYrEoQJ5Db97jLFT0UhU0
hCJLQKoYlNox/NPqdw7fcuRxj2+N9cygEa82gLj9dlQudirLVJfR9M43zlEsEgsZXl7B+pwT9aNZ
ukx/VTFTVyhLd6a0t2GSLfj759FY6W1m+5QeOMKL6Fc86y9PWFGaacVmEYUL7E6oDZ966mkQk5DY
PLyYZHq1wxAgHKfblfIvPk2/AxxnCVjHENt2cv4NBQJP4P0XXs9j/zgDPHjmQqIaeQcMZmaWBlGA
XKGQD1KjwFMtcHc9E3uRNWzCW/Dp3749cJE3km5QzBREV6TcuLR6stQvk5boaZlqcz0VO5jEEnyD
4V3puOvSovg/awp+wL4KKCQRf6hYxcyC7LVspClhWvJVSADqISDp+Yn0uoCyTFxFEY3E0olZzDho
iqVSRlH+vgFaR3uSoOBrOPWVpWJRPVmd1VDq5PziRIwGZvFiUJNUqQxhdvGyA55qOtjtPjn2zqR+
fDYCoJ/HsKE7BMy9N5wLTMSfwfShPEmxhBgwGVSYIIENv0Ej4QEN1QibmiqA+MfcFUt5vHQIKcup
Dm8E1oEsUssIIej/j8k7Pv9GxlEZv/Qh6YNoLILXPPJp1fyPSVg/W5HZ+lZ9vqpVgmDcMG+jYssD
Yy3zqovWNaEXCaWb0rVG4PfS7JU4tRGyZGRhfsnJ/AfaxJn2fvHWF5ouKT6kQz+ZQcw9IpieFGSc
mAkSJGu1I1B2LopllzzUoM1ZaZoq9royJxHQ+FAmxHv/ITjOKSGv8aJOMkRKz2j21FmvTtrOm8Wn
bqjJqkn7nB6D3V/1F1jzLCIHvtKvmlOuqLh7ZlTSEFSwwd6qu+M07ztuyZAFokdcbfIeJSYckD2l
tDjhczLIW2qWI4D9ZK0R7TMREpfEhawjvm+mnlvqQiWxURNlEcZx4YWiEZ0al/gqwFtlIMhUetaV
qiGLMfeGP/LzSm44x9yDic7fyR5TcjpBZgDovVhV4b7lTzIM4YdhfPqdG3qYMrTfSEs/92KcPOsi
fPCeB/2Wy/Spggl9YpoOa3m84GAFQ+tycr4rTFE4Q6mAOMg5U26Jk+eoYa3Am1VdFy7nl7BcQQmX
39e7ro+k+6KuonHZi65kkzYjd+XkQpBQo9ZlwLUnFreo6r7n6SjS4LSyRHAeQkDn+NVDJ3o4XnWL
rpns3TaKL+wTBXYdWykmSiaaki7+2aPA3wBIfS2A/qrrL+SmpJhaCQ6qicdyWvEZDS6vYcKqWUKr
Bgqi6PLzveiYr1MVCilemMUuB/TxFF6U8lupjIWJ0SOxUJADLsiIGWJq4rF4IqqbvXCUtra2LbM+
Cbv2Rilj1YrnAjEgzZXZIxizYBVK5ZMtgqspQUbVMYZe52f5dSPbWh0jC0Zf3fO00HWUtSoR0V6v
7a478IczGCw9acx4DuBgQ6wXViMgh2L4DNOdfB3vR/lkfV30+tUg3YpIBAUOvnQXQS7//mej1+Ns
t+qT6UTxQMmGaVqKNnt6ONa/9fpRobEq8f/6sVMYfMaVmPsXC+drAMs02pk5iBWL8DtZig9iDsQE
D5rouUP6/h0ws+Y//LBK8PrmfdrmAkpdZJ44iWZDPe8SDGZrmnYiupBeBJTpEBO0dEM/6z2X1Oa7
aEQGY5jmFoHjmgmK7px0wHPUZDN2FHOo0xcoBAJay/HHX6aHI1Cw3zffQb07PTJaqorVOWiJuxQT
Fy0/wvFRutymOomSEzXtVj+eJDnOnr27zjNaCUD4ICe8DX8RPD6DD9NWCMi13hwUPoSmZ7vtMbVn
PnSs6QRu82BlL1SZq7yiKUTi6E0rH1JTlbhPmASgc5EQwInLUY0BqchOoFkKUFk9xDXAdJphpokh
PMWsk5jZLq4ZBeJ8c+SISQ3ulYZwu2k37cotDcT7de/3xK95plwk6onUntl3WutaIZmkg8vMbs88
+Rzu6woBNMX/ttiXI512ZGIudvwdCZJqeeLKXyOC8ChhX/miABkn6VwAteN22Sn1oWX3DhilnlrR
JHty05n6Jlmnh047U9ODkknrjGtbtwyaXFL6ywuKc7DKb35n5PATpeIwJvAgHGhTp86bI3MFLNml
VQvsc0ef6IqICgfJRKoYEwCZZ8B0sHcEK8CFfGNxaKCnPHliqyHXh2ptnKr9/kh8HDwPAUX0m7Ju
RJHLTAz+NbhAQe3DSxLtSfiVurdnpIdTbeNGjtBBsWkSC5fbcxsuZprUWJXhFABBg884OkDrF7/J
E0wJTIQ6jJFDBzo69pgjr3fytZCca2TJXCSyrRGr6sPKEqRv2DqUSWXNaHZ1gWrWxoyq8jkLQxxl
ZoO1BCv2373aDYDe866/ZNXXmE6w1aMVrYXZ3sDUMrQzSszUwry8jiI7dLpAqSa4RXUbPnbHobiZ
Vh63lL/aGNCzKyJqPG2YAbSw99Scp0sKjr6XebVtTMCLaahKEc8LOpVZE8MGKGq6UDSNkUrmNr9r
cj4BJntFl69LBlJC1HU1e/bc6HseXcv50bVxXvXjMU9FMWO1/PLRHnvenE6dINqZvYfCb5H8fTOb
Ndml5OmHXTIv2pzAHC/BYIsl5FOfXihGqLAzSMAmr7A+eu0IiT2VN0NKAueyA/lBg2ESKKZj6PGN
umjHmXD54A2xuCQzesHP6Ziw2fZBb2MNu7tBvPpUyUxiMRj2pqzA2sAdM+5gDf5/dtT8WPlSG6Rp
kqdZEyVLK8xGWcIYQbLiHmPJnlE/R34Im+ageGJRbFyP3lhVXLCr7McAHW0g+CtxPEmnP0Wh97vm
DLAqa0V8uJ8LEqvGd72gKkn5QMRHvbyXLtNqJY2Y8MBbfiXJf/+gKUDHQE5LGjcLV9mpDauMUrMJ
yTfN7gXOND4O9ng6RylmmGAWhRG4pxT45f6DJWNsLCyjzh6deN7sKMrnETl6JNa6NFWKKkOnXOjy
6UOMRvrzgm6P7OUxEXNcR9DgZx65ntZQHZYGsEcas6qfuZQvTDCe5R6pKScPy26ef8ouWexQ63sW
50tKYgpSJwIE6Y1u4Aafzo3iyJR+nCFuXhdGWkdOWP7qpMvQjr7mrHiKbeBDynH6ekjXM6TXb0TI
Yg8/qqcF9jKwQ4+cUbWewTLHfODBkDBdNFFhky8aW97NVo8lYAxZB647NPs+fkaRIYKli/EB+2YB
GOeQ3TZJcjoQeCbqGXzkJ3D5qLnITMSPG0phWw9krFWdtQf1fTAVDcF9zN7pq/2+anq9CoIwY12h
Pwyq7meNL/HNGBGmn8IIfsT38MVHA6vdj0r9CaLBqH2oVyZaX1lErYql9A260cVubj3gmOacwrAp
dL6kPIeKv0Tc3pU0F4FPb6HzD2MqHlbTNLshkNlnx17FcBp/ZoIjwlVuTsznA7dE/6f92dwfJ9aE
wV8fgldtLBOJAPBWRlP0ABbQcNln9A06vdKbn8D1O+wh40gsicgG5tqGPJtnhtQaCqUHIQtF5aHN
0okxBCuiEMlbFE35qfO7w0qy8QGew8KIez/KQAwhB+ReypxFhhzXOx9rWw1fR/SlxweJGN3MqluS
NeqUMbN1VGbEIU5IkI2/AAj/zkIPgU81XYra6OcodlZ67jWDfdc73yGf5JuXorAsr42XZNDEkS09
IBAyXg9WTmIDZXnm80JMU2vHwqYWD0URqTIE/YNvvyd4W2Ye0f4VXrkGLn8Xt7DOk+we2fzJLxnx
Wm6YGbCYB7UZI2E0+emyPrBRIAJBQ8QbSq41L+Hm3Eu9F+niyugtg3bEQlIfi1uL21PwZu4iVe0c
1XDijKa48CNghIT1aecUoxwMF3/zFCcla/p1gTcIHwkQV6SIp1lpPbcguuzi/F80w9ysCXyVVRfM
49cS0uRfI4YC7itkAv9Z8r8AW4TJkz2UhvVBW7gyHTYTmZYW79EKEOeyPhk+C0jBywqwnQkDxRw6
81F1P4iIW5kc1+KvE4g/TFESyg7s/xGNU30oabmrNqqEYi7mSX2FAFh8SFWnsgO9mPHJV1Ujs4XE
3B1Kh+nTi1N26O695hWco++8dxZBP03cv3jxT+GJA0ZijMilydgjmWSdVOZe+M8oYzE02taGiwiq
2BLiXKam9xaE5ZaHD+Fig9cuct2RRQ3WYMYfkbSQcU9dMg65MGFi4kdTSDEOUWTf2UC3DiO++jdq
LhujerWKVsaqmSiod2njwDfCSPI4Ui9/5VR0zbFCejySB2VMpzEHUwI5vVE9TNXDLqyCkAnw7ahN
uaZKfn2NcsqnD3Sy1DZXmj+cbDaJW0kLTGW9dDuhgeCjsYlv28uH7BkAWEI1RYpVzsWeVwxRQ05E
Q460a51W/QZEGswWjkRpTX2ZbJ9o8t30z4VPvjjObaHmAWY1LOi8Nvqxv6yDESC/ESHOw3A2NR4q
EwFA2UVPXVfBuYlBp2FzVjlsgCxA8RrzBP00PBUlV7O4ARUMbgSQBYrrm+2Ba9VknmBxlP0IJf1y
N2/76BsOcOibPQd1kNITpU1IXRI9phCLZveEbKw9NHNTjwiAKRLgO8EwGE2UZsIGMBKD9Sa4XhpU
30Vj9ZOATajWsZnk45+WXuRMqb+AVRHEt24TFOm3ZA+ddBkHGYUYMiabEWnVgoGqtZuCvtUI7Ny0
hssT8pr+qu3FO6PUwM8GrLPHQEzF5GuovjJ30zk2Ps7hL8izrck65JgRAJ+clsuIV2cKl6JIYt93
B2NYqpfFkZ2FlSDbnak+wfEA+5L1Xj2fgoILW+N8p0j1mnnPycCbXRGq32NM5288x9IxA0Y8YGQL
IFUqPay/9OP/Ew4vtZbZCzH+ps0yIQ4vSEKNqGHZ8ybmX2NNWKn01OfQ1/pH62/eU9fgkrHdJuji
9vJGQNKC/J/J7nFyxgsZB9m3c6kYWTZoVM9iz5A555EBVPPbFgG2cxKWlNvSTk0qve8EQHkWH3fo
u+LYcQGT6alzkd9iYlZtiTrG1b9VEBE/dAuGOjQ3HGffhWso7VSLPo+X4cI98djcbrrCFVmyHqIY
UL++erBwepfJwKwwi5XxT3syG1ec/R3KvfFVeFuh5Aq+pU682a3PF3YsrUqMZYxQpa+CmBgK7n2g
FhCHJPkHzEgLD3jQVUWzkg1IR5pJ11gfplcro4AgOTEGMPR3suRN36N7sqzoAoXgzT2MpH+ZObYc
ENypfxDQ7M4IoNaPA9ueiKr2TTMlCfl5Bp739ilhme4u8KkyG/kEFoJmDHrBSHWewQyzdSZNjHoh
IunQ9+JS2ycuWyyHZ7eed1v04jzKli3cbIiSLMBBH84oa2+pFOFEF3BAIdxIM/dVtujPqblnYG4g
My5AS7Sp+bZWBIPQ8YPAFR930cNKHN+xuDYBNwrcm9iire8/pJjk5Lixh1l7r66H1ut8zDlMWF4F
LpBbe8kF6cYmL9eHt4xtl30sAvTtVpcKCEo5XGio4AetFTxY5UrgbS1mG+GKn+kBqz864UTm1Yip
DWCRsCAWGIUuhU2JCqUi/q2hDYC6QahbI5XZeGvUT0Pg3AoiJMd43jZFLr5iuXVD+7tySKZH23nv
LxIQfVNMdud91+oAAZ0Vc1SPtTiil/1fe8+ZOLzfmOlUkkX1AcpYoXg+TnwPOW4OUN5w+JayHAe0
0RwB9ljNdlCJKgNj5ENxu/0VZluPcANrClTA1eLjvwLVBfQm4pgKRhhf0bh8sZmL2tsxupEa/7sd
MoUQs0xdartX4fgjIV4OntQaByyck165pspSNbIH9r6+esx2q87dlovIRnQJYitNRBYvgbC8dN8c
4CGDE1uK0sIe/1IP/4dV3STd9J8qC3SimcK93KFHl1u8SckiWqMKG/H8Nc/dlvMyU+u+RiYvXPcz
O1kgPvpJ8JQjyG+yzCLLb9DkpwGQ209h/CJn1oYMsQVeRNDGSBcwBxg7OEnaQ6kCQpoKQ0Xw/t9e
RrorfYnFaZKWgql068e+kyVrTxCVN2UmZBpCOEG7EwZvE8ephlugQZxq0nDbcOyUCR8XurYWxU1g
Rfz2Z7ZcgpNn9p1+u07+IDNTEno0oAl4xU30pjfHTuf+QeStdsKv836QlMLC0kjxO+hGtN0E9+TW
DcNWBXe2kihOE6bTdqe0V8Lrb4h0u1RLMSpbDBY+E/yda2C/J5D3Uo8wfYYnmNz5Cobq/7/zTAV2
wAApYv4GpuQC340aKu7V5ysOUeVDXDkdwWWsEoXPGYXd2Blih3lL0qyurntrj3YFk+nAz4KrBJpa
zq41CiPhIcGEFKCposcuZLGcBc3KcDKrE+hqRVdvela8CFF3oEKgLnBVaLXfOom94Qn/SqfJrdMk
9uN6GgzQVRYLobRnTjVYc/yV2cX9xzUoW2lcA5JmY26snAh7wUSE+cnFwTmzekY3UH++dJTdrB/+
aYSV9sGBYZ00IxdPThsWuVNYVN78ptpB/DoUkCwLALkBthxky/lZp9js51Q4kwDuAUbfc5HXUj+S
fkxjGwt+Bsz0oJ8xo7a6/wyF2HoOD7LTaGesq4OH+3iyDtAlYbLw9/WaRSfzZINtoL7qJTV7/9NI
DU14MGKrmbFiLuJJqLDcb/eE8/iCwh5nKNSiiiF4HkXALsNPRlKbJwulEhFysMCrMFP4IdKKxcyn
Noztqtvd/FVmOao4DxN/yoMGy62FtGnGINhuIRzpotNFHi993BXRPnFzPAdPG3Y/RcLvPuPyxrE3
z/R8BnwaVWNgRroy6GzxQkpsvbGVY51I451RmvK8QTRNFjBKpm2q+0Yv0hJExl+rJODVEBYq9xRn
agwNE74b/c0VcRQ1gM9MnvLzaIr6K3YivmTiOlWxLH0HU6DIc62mW/OS+p98Il/A/T1gDsMLhBD9
xsM9JScoSgPfveZonLrN+Pi7PSJq6rEvLzvodENswbLswfqBaixF/H4TYb9juD7Q6JS6/Hl+vofk
cBiEkAM6ZAWNyOmGb//FjfpMOxSvtHRZiVVvOIJEdI0b2BEkkda0yGGn+5QCbhRm0RsK+TRRMq7N
Drq+i0IA5vgIb/xA4nSQkZBPFkvKoHG0+f86bk+P7APHymrIPRP7gvZuQxCI6R+JLCX2QpC+IY2x
Zi6b6PYp1vanWupwQUkTjVcP9LDxwKJeOObp6X7pYpMtnQZxBGacsfRzR7YIrit4zUmDvqkj1JLi
fGU8L2neE0SNX7WfYV5hBgFwWQvg91F0TUO3iFL5dHPtR4cvdqzUXIYgSPQMCE9+e3q0Sih45/l9
2NPlhPHuqGSK7XlO9VmpGmXvaSGtiuvA0c8J+Gv2ywMe9sI9/YATna6yb7HWDRgom2rMjZrxNkL9
yNmBgYJO/2pfmgN8GnA7rTABR+2Eol4bWi3DECg+H7uI6WZkimzPWBVCsaSv+HT0gJVhHR29st06
hYLt9LTGoa1XfNydxwcej0+A04WqTw/qDl9SjB9vjl1t4JV4r5WmEZqsmVX0uQA0y4Jx8u5OPpbD
A+wet6F96cfjpT8IOFFeHHJir3v6gEXF1AWrUuHrC2U9qz41YZvXtLrHUQDPDhFEzITrVFZ791CY
JH/VT/BXlA1XrObqG5Gfn6Cw3k4VLJHxvkTN3APQOjNzV16I5G8P4How2ckDxtRcRj0SWqM4ssBL
XOZKveqv5Agiy/YKl+1Wb9MyiYNNz7Do4rqeJDZMhg6SCJbcoMgBWrfFcYA5yfsEEqcrL1Dmsj0r
RPe9cK55uPdd/S/4aXjw662/JLD26JHTx3i/VU+DFES70Ey9N+sU7nqEAgn27LaROvfTEVekiMfQ
fVUQCD6vwG/FJQoJ8JhRSVp8pPVtcnm55ns+3ybg5c1mFhi6mEB/w9FLhaW+WWyHRMjYbXVsjdxF
tcsbN0ox2+XRan+wdIt6CFpoanlfZPyJfVMIQ1FGSWOXZ1dha5+UDXbYwtjeK6U/gm+6jp+kDw2y
IPEpxfX0yIIP6yzyVrzHyWWwSKQlECycrXqXViWPQp9/j7+Uro8ejqJ3riX5TJViMvO5xarJqheK
ncObm6+dfMxe3PWqWAsWTsDIEQpOfBubsK1fks0rMqtyjOoNQkbKy4BmgvIM3aB1yjh7cGCaGDti
IBQPkMq/tzcG/ryOoQWY5jPAozGGj/CwTqInncyYSl+Kyl8EdNFd75g/C1m6vcUjY99YyCI+lXAP
qHDzYehYilE2m1q98KuZoOVkuNly2fIHzfRLk9xjkQuawFfovyuV/HyLEl8cd3F2K2nP8E/kjH1w
oFSuWmj4FAJW1NhqNDC8T1hAl99mqZDpUR7q4YI65r/P5eEDVUNx8iz1uby6lxikhGGyQAQ4y7AK
Ro9LakAaByO2/3ZlGiC1wqvLF0AWX+Rq622TaKbSIP6IDYmC2lq01cpZ42hnSTPcmaO23tWTJjQU
FisoR6LiqwyQvQcUq1g+6rFERb9seq4swmN3dObx/FGv+i9AMOsLs6weo6WkC8esu9eUO86st0k+
pjtZFLXvGsWPgwDCpAINNoFOaEp2OVfar0M7IZxqNPeU/E2J41OxEqwInJNEVem4gr72X42Xc78w
usLN+3iH/AVknIBEfbcvTNEYS2/IUEyFxKQ8GK8fk7UAkaW7mst6+3m+qTukxYrdDw5cCmbJWONS
JR8n0EkACtSiK7knIHX3QoBH0XnhvUdscOXill7dqU1s1arcnezF1I9SRBnUBxaZmShe3udw17MJ
GIBD5VredbemhOeGx4fMPcDj7myr3G7XcmcZjSwsD5XI1FFZaLf8l0mznWEycDLbZGpIk0tQaJIm
TL0Qcv/7pux00HBfp3bYGWF1JMiX9w+HDUm63J/WxKI8p9oz+BnndK95BiGLTKbasB7NE+evi7yu
5sV6twyv3fWPPg3lss+0jrbHGjymu1y1UnGYLxIDUyXvYMW9ehHz4f2g73ileKWCDbv4H9aEvNxz
FXLzW84BnP1DAryxdW5U4XLd14biYCmGY6AnqO8LZvFcqe/VSWsDjZjjy3gQIYIRo7m/bSnULFnS
i1INrPRZUvergOl4bM/hbllBOwmpqVMKhGsLsbbLk8fCyMToxeO640nYu/apMsAeR9L6KktWkwQ3
s0oY2vREDpSd5gNxkTXvJHAG15gqshB3vcDu0Xf74jtgAhH42NR24wuKeLeG0ObVx2A7XkslZczV
4m23COwgaIX50Nz13rrcAJDSrNn5neRbyHfwUgi2ZmP6On2dQyJkSNrs41VDw94HVDb4d8hTViQq
BWuyWFsuV/LGCZAV+cwsTl8UmOTI1gPR4ba6ZgRCDamhg4BDr8KHGagIE37AhZNyFISTBIgCc9cv
aU0TeUybgy7htxtm8r/fL7193Q+tvlftGmLywTJmvBOszVAjb7HSXN2UNJdK/9kjk6COUrZNBlAC
iIUCgfMvvJXh4o9iByxa1A5stLvHLPUYmkkDOYfimbeiiyBE0J1gAf3VUZSrsYH5Gh7MPoB6r1Ih
eRn4JJ0hNshZ+YXWcjoD3/IYnheDKZ0lNy3RkvZoy+ysHHqs4G70OdT8DxHHrDSp7750Dm6u92Jf
6p239tSnQFNcnL0lFpkuSk5+AoMJaqbWuNPZKuCOSMXsXyah3N93CuzspvqnVrITUsv3nv/tycKl
IQJUhjbdaZgdIho+xrs4Xv8X3kSa7tW7Tti/y0j9HhaWTJeKlvU8RaxL36vJ4lsZ+h7GPcC9lHLX
7dkME2zbCuItF9S3gJ1H11qY6VIF/eyx31eCejJphLoL+2P9QONMzRcWFXeR7C+XMnFSKymA3D2N
7vFgUnNqMJNdixwdfbZfDUuoiYGu+WkIiAKsHJynZSDRbCpUhyH08qf+Tj8WvYGcmtHC9QoJUmE/
JSF6OoOZjYQrm+n/4SwOrRMDYIo1YUbe52hdNn9Uezt8+xdSTQ66oLthfAMIdhEfZ8Papr+8wi7x
yZ07D9rBShGZ7q0miCChMMcSZX+EMbbDXoUc6a/Dtq+ZJZSuQ5dOUyDP7nRCwEkQx96yEPCqIF+o
A9p9WajGaVWZjVCFcLJf/k9ld4FQJMIvDHbNdOaR8ZVo6upc17FbSlSOqJcu3tW7Swjf0cxJa2j7
28UpAyw67eY9rgzDFZtab8OjEqR3d20D/kOUtqde8+5BM3dqKb/c13FE7KvJ4tO6OWrk/sK5xYFi
3/PncXUjo2dZOouZxNnxfNl/axjHyA+8S1ZN8MLqLJ7brG25XO9CmwwZvlahHkG6Y2PCholC4hpp
6uArBLL5tj9V1sTuEb5cYjsIYcvJlWVmQ28whYwod4nxPkfHTbm7PyZ0fXwOeMcmbddCHAzKq7rC
oxi6oW+t6Db2shWg5rAsZYCAHwaoadKZgMVojaS+WGaK2uRdGWgSZrNuSZmL+gyNfDtGA1pFESaT
1caufwEH8a8xyqnpilLDGeU+JJQpYq7z/cmJWHhC1qNOHyJLwcigaMTaJSHnrRJMeeM+nTQaBWg+
5HlPcaTP/zS4JMKnejI4/plAeFjOSZmHv1YHBRJmWPnN3YpovMdXOieI9N2l4J2IRidI7oDtuYkx
KL9nT7f1RSMWtJYY3lVtMwF1d8fV/zMOEhl+6S7rM8qWlL+7/1v+j/Oa7CK52LVV1pUt1AbezLcU
/u+XUoZ+V/thwIFl7/8gAwJrITG1XaxIsb8RO6sfQHRg4BN4FGlEenicSFFv34xAtbSEo6R6sJMV
LFXX7BhawEY12JLlqdoY/UV6TzFSsIqXKFqSblNbH7i9R4/YvrhMEXtUCphmL5cn/KiSqeooPrQ6
1h5m1QcV+tClnMNLY4WkCgXqtevLb8tkYN8Gq6xKk5sCIPWqqCRSIL2NAYFcfhrv+mtkc7wRuev5
Fnv9tvisdaxC0wKi5D3yi5ucMPwgUyapx4cNTTO9kGoAnJJsVV54yWWfWofmGB9VIUBZa6SL/043
tfzNWn6dN1xzVpV0XRIit8KWK9aFNLmHzwTFOv33SfadILi4efUmOaSgTAc3RsX9NFbr3kwLIRnZ
KFiP9qUkX/lBDuTnwM3AWZ7UMrXNNwf6hdfmr7CQ1yBECR4vqI9U/c2YG0bw9F8AEnhK4UGpR5RO
MBYb6cRBIfmum789ituz4MTBrzobEGKiyGoSkK+djPze0rGWWe/3WYJA/b35aa5EEzgGKqGc/LeY
VeOPTo6+audgyXIknU7tP+n69n5Za11cvbLrE6oDt51qshndFQmchYy53Y0YK0xVLoCWXOVgl8Cl
DI74DQBfpBkbKCpfRU0xKCAxF/wHOZ4JAPH4bDha5z/YsFE1zIDy5O9yXTOAR5xBSUZP9V80xOiT
1xZjIKxiZu02VvvFPs57/y0+NXat5aVAL7zeE1ZLkFrkpW3pY2/0N/+5LIn7JwEMwCaJBlrFxi03
08GaAtQCgBuErHuWHnqljEpwBQlmYoPAzOzlWbEcW7J10foCLO8wZ7NXTgOOOcWbzgg+WFdwW3gn
OokY6R22jjvG/vc/pbLCjjOmWzO/M85tfMGLY3sqFcn4X8e5vcbWGl09U0I10m8IixbHv1fKSDd8
Sx7oKePB2kcvYg947Wk71onQ11FIv18ZCwn8usRLxqv4HdL3hcVpeJiWZrmkbzHnLPHwNm8I+f+z
Va03erhEfCznLnXWReFOzq/jGTg5z0JPGzfKdcuLI4htP4YPNKInriao0syymp4fDW2amkxunbjW
gsLY8WMnipYZfpuM1INm4c0v/wazfiJ5o8GcnZJL0njzrKHAj+CjaPYvI9mCa1VR/5syEQiSJdGA
zmK6/S3wt14DvGf61rofCELO2QvPd3gEyGzW6kCX25lLJohwMI/bFbczKwa/RJXrCQTqCiPjpzWI
04Q9QaT8LcdEp/gj47IaAowcVi9WQpJPakP98jBFNYvppqhut4x+CfwATZhbSBfoxC6YEVW7rDTl
AZT58upB14mXLXUtwiwjMpoBr7vEF6ggExzKfL3r9E2kXQNiLsmXJzniimHkoaExjxW4vbO0MpjV
0v+iYblXB2L2A6YDiqdZ42yvEeWXlmEQPQ/WApzaqN9yLfCmzt+Pe5RYelRbAoCObgcM/wjlwEg6
/pfuHriWOyicDu7sOp5QYU3th7tYRFg6+9GoRG0riT4EjlaXiATRn3Wt+IKvYEU5/GShUdrk9jk3
256VNuJcGiLgyIzWvP7ZCmVMgkD5TrnhgQq+kesmtekzUMSSglT4KybKAV+Da52+nvAU3zpntWsU
scfrptOOCRLmZelVwvLf9tfbznAJS+tZbH5z15vb8bG8Yc/bgj+kO5swU6BSCOVPQJtDukwFtBKe
mQn8uOYbJ4OCdnjr9Ovdx7rWwhTxO90dH0ME/xCLFKvjIQRXTD79Vdi8fm15vEy3oR7IiRbIudXa
IiH5X2zgnZksUtJrefSGaJt5WgbSqL59DQ2K6qXW5FZMCHQJDbgdKDUzUg0HutT9VWxsuh55SOzC
N7EIV4Pt2QkhW51Oho+SOOQ+CVBPK0+p9JTscwceO5mro3Lx6DbSyEVlCrLwbu6YKrPFYLkuSkoK
yW96wB23GIlKyjCDYti2D7JD3d0w2z7vG/384Ed4YA9cuNrueDG8i0p3NJxpVsPjAwrJpHh55nlG
V/kOJZpmrBfmadk8vEOnV5fdgq7IKkmyUG0F40qg7NGTXIXhWS2pa58ClOyIb9Nlyci6gjUv/99m
st6tOknJTCxbUTQFd8va4CNHnAP9KfGd9qlDEBAYxzZvS9N8jotxBmgUsJNVN/hbrIT85su1y5TL
SjrHYWXbEdaHc0atMOIa/JxIJ+7iFkKy3e8mmf1N40joBOXULmuA1MhdChZKNacdio0tnF1Fj3Vj
pCjKX9WOljd/k9qJW/MPkUvKZ3HBwl7rYRlCGBnH7uBuOI3joHrhAKGIJlfSVDEFASav/J3MrESj
D+ySKKCVXwyQivTmENjyC8pyCPPAxVU2ppSOVkPAnihnZbgJ46VhVFWtlM6WbPBIGmtzlYOkoHU6
MwuPlry+yoD1pv8+08C4llqYlzs5Hk8ZczV2fr5j5TEBbEvcyfXzMTeGGPv7CeA1tjK3N3L1mHoZ
ABWZDR2HoK+axFFx+WDYsCtTrIVyUUYaIlTvqpec7oIjoKG8P7MsSY6Q7T0qE5nQqHDWe3FvGjVw
lRF+EY6ft9ND63quhvWbmNlGnhxtbzLgg8GR5a9Fsdl/Pt4IzW7MulE8DRdY0Hc2QCdZ2UrbK1Yk
1HQGf8CRktDR/RSf6w5OvHWY5SC51ZEt7JDvDAvs1AyEWu3o9ZpN9ew4VhIAGl0ka1COn/PZUf5k
vwW6WvEf7ePCRxbGh3fOXslecTMtemtEiEPPLHa5L/HZhEPeiDfx09a8bdbNULiX8wC1xKCFhCom
unyM4ikEji8ZqssFYfvshwBStGyIzDzbhvWCRF9pS2DxAgHKhcEddsI2pCxkzQOAsdqkuXb0Tb2C
Se6768rpb9VltpugQ0sMoGreaRQdCFWrVE7icWIP4X9X7WbPe3nQXOdy33uTeC6/c/cb8LE9bRe7
mQ2L0qQzGrEJ0+FYV31GlFAXX+nuZjThVjaQe53caH/i9TMjJfH79RGAitpEv5c5vvVHZRIAeVfz
GaG/hNEvaQfQkeW3kr0AUwy2+O/eUnjhRdJlZKvK05IIDG9KXgk4TUeGWZSPO+PvykdktfhSCR8h
xPnRg1tkCBKmlT5+oKcRt4kFZGK+JscUKuxdDz58LD6tvNnrl39jntLv9u1s7gqbs0pOdbGDAl9P
4NdK8aiQ+i2Zh7x3GDf2SCCkK63mH14jhZWnF8WM6xXl/61/ShxMaZGkt2hbjagFfW5r4ufWz7KE
RqAgQ+XvgUO/G1olUORQE4OwzwDgvychLzwY9mtAdA4Gmnf7mpeingBQXkn8MDA7s4XT/PkBo1X4
NLRaOtCajqU03r2GxSCJtjZynzQpBXjn6lAfoW6clBY+Y8yUnxsB9lB/87ylips5FXCQFsYykX9u
qKywbZ+Wum1I5GoDVjqyhmM2Sc/pU9ZuaxCXchqLUFwtAxrIQf79uMSEeiP7zeBiN7lPyq7Yibf3
LkvtFegy5RVVNfGEP63CB8C+pIAZtdjdi2dK8AHZfA7vEKO+AkxGDwBZiMoMFhHCcs2Am4N3XJHm
qhgxpOS1hZaaIo+TAMI99FmMdIGJyLF3mGb1VRm8f49W7b4e1WHlF0JyMT0fBz+5bdH1qlOmQjIf
SWJL07sKUIs/nCqQO58bIiAgqG63t+RXyjP0SOEyvv5FnvOI4iIs4n0h9CJfUP9HMkzhAtYpB31a
kalAiGf0mEVfGN0Lqgnk5bEXq34zA18NQZUO6mKUyq+qm19cGJgxvjiykluF7n6EI4kW+tzZUxwF
WZayT+yrc3sXIMqDKSUMXSIs51IzRGMnH9mcaNV5XQl0LtgDcwf0ovmtq4lMPQFfWz0Ojbr8I/g3
ymCNWe0LLwGxT8MSQhb6jlBYbumgvHYfr3IbP6y4Fes6BE2GFNVVBM5JgVtY/tRUNPxo0Hhi20UA
RnMc5cFUpa5gBxpDp6MYH5iUXIsDTAE07dm/qBXryg6ELxwmUZ/XRpcQWraWWDV0B6Xm/aoW+q9L
BSfctddykVKsiSdkJk23YUvrVduLaOII3vBxtXiV+x+1OATpV+Xw1sZF5IggoZijOf2l2zFm+W/0
LzraVvw/7YdMOuWOipaOATC4IFPzUA75RoTN35UUpNxHW3bBrD0CI2+d2i4F4MuTmrT+tYSnkHv9
4JkAUpVz2f525napvonHmNwsxwp0fg+AIPmr3ox1ADbaGPHcikhGzCkHfmwkvvWPB4f+jpjSUJxT
Lg/6/e79X7F6BsvA/Eagwt/77ngjVzxFo7A0YLnDrSxLyKCvJWM2uy9bcMWRCMlYcuHLE0sU1nnG
eeRHmK8RBDmVqOvpizD0psxap+upSqRF+Fasnsavr+8TIuz5uQC9mb11UsC/W7nAYiZa9e23+hhR
y2VFWsHPV9nlKkQsFq3EHHerd5gu9lAKb7VOUmyLfA0ldczr74XdCGrAGh3mZITAf4dCTGhPahDw
FZAbzT11zImGh4naFXkzmC6NmGD90tu3mr+Q49/z+Iy4SKiO2Zk+ivA73NGUYi50mazJSqPzc99N
dP3zDmeosKE/+to/HfL0/pdqQSU1QcT2e0lh80K7l3NBw10d0Sj7KirsW+Q0qYLvzOyIEqyGarSl
T7clblKnsmDRATFkvHRp9vKvM+lTQW4WClWJDdT1BwNzXUUXV1NQC58ALjMULS49VQI554Gp1f3Z
5lm8PR81Er5xr9VAd4391XjSc6zTuQI1NMuS1wq3TkHswIy+yyIMS7tyjqQOxDkJeFP0dbh5tU/p
XuLfFuC1lt/Bn51o6eQsz3iuXane3R8NJ8DrlvE9ni2ORbaSmZM10Ds7v4R4KN9Bh5P1ZHu1oo0+
9QnVCb2Skk5R5XQ2NZh9MahTUzQ2IMgFl//jshssOM6BKndaRIAQikH1FaAN5NNI5c+jqKG7moGj
rnnadoA/DGr+9cXrqAYHv91wmKNjTbN5Pan+9Sq+MJcIzuNF4YBLYRCKrQ9AUokOiKzxDcgnkrPG
M73l+NBLxncBFQAhSmmGgucsgxkSzl+2XBe85tlYfeaU9il9hmPiLT3NkgnUWO4m4CrcLPDNc+HJ
GHKSpVCGCBRp1Xci9ZKHXKuyygZFZgPo+VtgdiT1ZLOzQfp5RzEy0pPfe1cZ6/qaZJaLBkzW/+0T
YtizM/Oq+Z9tJEopvLX5viIeBUZkzdCtmJXy7Snmy58EV3FnTVbXPnJcaIe2w6j+XGFfIjkT/PHz
4hhqo+4XUFmm6g0qMfkCYqTyz4H/1Fkoxr1VV4jKFBgzvmcqY9Nd+HqLJ90nKU/pLZx3Y2cRsQ96
RxK4LNs6FjvEGMfglKxdFC4gS7V9i+TC8D4XuEo+4yGg2Dzrtzl5vWJ3Tep7UAVBgeZ1qhhCb0wY
Qd5Ad1Gp2UUQh8/mrbmGPFdyKFg86J3wSUjwGLVlnyhM7lOv4PbT+iLRsWOmGdx8FVL4MpFMkkz1
M745lo9ui/rqz1kAuuPUe4pO/QKPJpDNiQh95goF7wHrxt7zz2FPVPXl2iNAJlazuJacMeMma/A+
Hr03Cr+XkjHNjHhVCXZ2crqIgFnIWbLDNE8hFB9JH0y6k2CLq4hgOzRlY5/9NvHIqDsDaeyZKngS
32OMDzZVjKlotWEb6cvk1FdMLGjO4M9PddM8lL+m5Hu1RrbVESk8TKjhfJDVqR2uI/jIgoJA/UMB
mwvROi5XT/+Y8QDGEbciyHk6pTVlI5B478lgnMJX+XCw454y8xQjOpcJqEzDYUDtp40USeVlN/zn
Qe1tNsdDJq/66JYtb48E8qRWl/cGkepf783+HLV/yP2ls3kLAUxNiQddohuLa4wzAYVoq2PB3AwO
bchHkLi67bi+ZLvZqwI5QyiTeUT39FQDLW5D/E0l8q+4D8ME5BRXBfX/c3lnYczngM0u++fCsbFy
UiV9dW5WHfONTwFHTcRuNqX4JZaeGtErJ1X2ty05y1WEuBX/D5DTJTV5Q/WUFt5nhCxYVyP6r0fS
yN8kz/rJhLo02SF25YpZsqiZugo1MvK6cZtbSoxvH26WPgX6gc0IruCR1+Uegi4PJhJF8PtoxYml
/8kyH3w6rpK7ff9cheAqJCvpbyjoB5XgOVi2tlf/nWQkqAksH0qZ20ps5KKgWy6K9mVQyXFB+RWt
4Ja8mKTpTMPGWjXbBYD9WILWQes+glMG991Y+W1j4c3BF5rLuvPQMcEncR6LrwbPI1K+2IlUfRs6
TNWf0YzNbVvoaVKXUUTyHCtPLN/ssuQpWauYGeeO4T8orlagUVp5A2Z+YL+t1yJzxHyg54FsMbKg
EerC45VxFDFfIl7NZd4zW//rl/zZkanEylqFXUVYzlqg+bSyLANGPXl3t3DtxzfWbguNjR4z+xSH
qJD4eZNNCuTQVCxxFjhoE2PzrVEi0K5ZgussaPLpIsGq9Sigbgsau5SNBIyX49pT9ZIIFHwkPvhs
m8j8Iie2MXvzFjnEtPXuWVlZwr6UOnLvMoF/QxkiNwGAKBUbGu9P+lChAGkdUnQZqfW95E7rMs5H
lUHf5e1xMUGDCEJVCACUK6lAEASm/SMlvLqwJkOkNOLdXCG7yLBPlAe0y9uh7jm070jHnAaQXTUT
MtWqTZafRSZ/yi4Ac8aRKcrrXexi9TzS1H+X5JMYUjsbgVv+4zOTaQsDokJPbsTQb5qTVkQCYf1t
LzxX/qYrM3Qn2tw36dZQ/aKnL/wM4nzdOWqBZ8H0DcTqY4SvUpokZIMMgw+269BhlMT/fvIgSO8M
RYw32dJUpnD0VI4XGeEqdICvOu7skHBuItVJUb1UxSw+KK8V9VOJnkcZKwDln55vxhRDcHgMb4EJ
1tm3BTC39RFpHMA19uLhuXYU+wBkBU+9q9eYsugmm0tAzOKXCJ2AyYGyXaPopowHBWm8c0O+I24R
cs7jWrcRQlF+Sj6fE6KgopNL8DcSzbt2NWjxRCtLqpBa9Ad2lsIOsbte+qJBd2NCgtlC/a/kxj5w
whKOlgB/B+I8aL4LCLzynVHBwre5B5Fty48LNB//5uoSOvOo6VCRlRkEGZwWNisobGoXV5V+Vkfy
Oi42qfVw87hHdlqQAkgaUHcQwVw91bR8VlkxYjGQbKGHA2wjCV3d7WK6IGHFZ0nRjxQ6S2mgSLzz
h3RXh3AcmTLT9IXFNsRIzVElWEWaTfvDUX27Lro5T36KKddqkeE0at99hBTmGpa1dWh3mK3+pHCO
aYw/ONDZGNSmkkdW4MuOMZuutp1AtvqCMHE1gZg3Do0ZJTbTchTJ7ZxVN9i8xKKF0WFKhaGXWkvn
nesICWoV2hQZv8kU+azPkL5PgjGjQnigu3CBm7caZHEYGmk8oeZEyDsYCMyz8w+MZ999HBlqUd59
egoOtrW0o9jcu8HhaKoQe3jfZykEl9gIKLi15M4bgs12MFn2eYurbr5QfBSNP10VD8iHTntNUqcY
HiaBpte6z+p62qG8hMu9i1Kr1ibrvR0tBKnVDdwiUOnMNjwbZO40qXqYDE+zhl99LIqzWO3oWP/C
TKDLUNvrJaikzJrzziQd3gvSWOOCvBzQX1LrNqVYwS3N4bfjSRjSRRUX9USO0Zqv83QwqF0aLEI4
Gd3QwJYqyoZ7isfWv0z7sREDbUbFdmf+ceINF1f7D/gjH1DBgDRjqSxxSK6UodMyfAS1Sg5ODulz
C9AXC71O3fErGIUCP1F8S5FyIkeIMc4Gs+1tCyqkyjsr97cYp0i04aH3sYGYNFny0lW70muCNwwR
SHZTnf9g2cr8XqjkeWTqVmTPUIlbYahwkmJI1rJYxeulkbmkxd8zuibIlXE8WDsWa76XV6AU1401
7OI5o52O27mN5QTT5B77HCR4tQh7vOTaUtZulPvPgzy48d08LF7LLnJPKixxndwq2gNrxTuL/F5T
kDV9DbjjMdjQsfPxtP3WPTEn+oUXPUhgdiMbumOArZzXzK8kX/Wwz5o9M9edfmRp2+3vWzLM7a5X
2pl732oVY5s3jCnu+g/ErLgdRVN+/I07swMvN3IM8nVVFgpm+YsiqHHWdlcI+NNWSv+0g2HzZRd0
F8dbmURRV7ZHgIAfBCFL6awEIi0E1SqDytDxCLH816/EpiMyoWqwl9DB9taSVVOa95SF3U3XFgFv
/RmG82qF+29hhZRogMaK+mQd/+VtgiWamHb7v1IZ67lDyG/is5mSvl+vgoUtRV6jmRzuaQlwnmd+
3cmSQnchRdsIuw9u1PQ+ABfkwuHHJ1aYix6W6cqAJaHF6h4mw3XMjhF2ZjDGw3PEQJo4f+URiyFX
Fu4AhrDWzYMIAj0dWpjLlzLJajBXNJjg3paeK6UIG1Nyo5Xn8zaWTj6+bAqp+CdXfUzLOPvANhfs
TiGGvU9bwW5WYkTVSCdWv9oYCco/x9Uy/s01QiLAPvQ9nLRqHWZgETxdVNPcB6upMjdsW0Eegfhz
yBjOFVAIyJF3rxADoBIbmS1s640I/ji5n+I1vCa0iMNV2rgmfmP/me2185xvuwdO2WmjUVZkxSFd
EYfBuLZiXBNFmZ5F/kDi1vLrpBA/DbY0oaDS9x7ArXBExe9pPLhuWsA5GVEYGJKj+d38grFx/7ol
s5rASL/3i+QktPBfFEwR3ZX7iVwtqgO/qBUr3JKjE806Ma0T8uoe7QylIlxIdlv2w97n8i0ax0xT
GYkLPoW8U4Aqrsr9ghHVftPCsWddvzLsxtgojvh7nKhBC98rturwZlx8Q6vydMctVcHvdMq7oBwD
44mfntk4pSWnxpqWbEyWkVslRi13c8fdwhRM1S15pyYhUVKXLmKPugnbQabuPGC9txz16bny4NYZ
5VNcRVVIR3L2GWCACKEy2O3zD0AxOWInhivyH/fi4FTe4E3pJztZX4kQROfLPj3xkwH+GvbDui/l
cHjBbgXK0puAzg7H5LGg1M+Zo0sud77N+26qeQgUjQhd0iezQlCadb0fFmJDoWe0snRv6uBPFrWZ
H1PtgyLDJZy7hhQWQitiVR/Inr7Uyvrhpka8CVih2GrjZA//u5RRtpPDIjVtQxoONEpZ4W1ZrTYD
5owKCNlsWnjjkLadCPZnsGRFuyQBBkfwqnYd3hooqdscXNGPLiGTtRQbLyF0Huk6XXa3z60XY2zB
7xgUOqdWyKd4qOUmx2ym69E5KGILX6TQeOJ1/nKxUND74igUyk3YZ4yzKyRC7rD/O+BL5O2wHDcL
y14ERjbM76itoASmvpo5Y5j9AQJOqeNlDd/ABno14q8DEnuLFdqvu0FjnG5ijkaPodCfQE3hm2sW
J5y/mXxuAxDZW3KHxykMR0wrK3uo02gj6KnzLGyuYVzlqVwaqphyWsgYTUI/w+LX6H5SNZ8mS77p
49Q+ZC5BE28Xb/jGvs2z4LqeHjzAP4igF/UgxCEicWMu/z3OZJnonzfNpadmwhQ/Oz3WvGoyyXde
/37ESpz7oHGToAN7m0T8KIw4biV4AZxESb5oZZv1Qa4nG0mJ6NL268Zjj6pA7hY4E16F5shVWaUV
3x90yTV3TbAXFzojbJ8NxNLZOPgl9AuWXtKFDhUIYlcymLqQYWRyGFpiVQM9JTTST2TwL3WsqxW9
SjVUKugRT/HxhIlUAFxtUxdfHKHouU/H4pnEBfUFHuiM1bA8y5HxoVOvV9/yxVP8rwpNwHXqUi9W
H/j5UGPPCrPpjvEmYjko/VS91Fyc80AHEQcctCh/z9j/491GfXkd/Dp4PFq1wagoFlEctbCIaZp5
YVa+eT/DELBPHB8xdoPobyf4CwlXgzeYkPyafPS6OaWz8sn8Ii5VhT5lWUJmvUS6C2fs3d65f5ek
jCIQUKBkIEkQJQLHe1pgRpo6W7dPHOjwQ/3NBKf+1Z1eqemqvEu7XmuF+Yd87qffaL6g+4aJyRX6
k2yEttBuHokhnP7DFjHZdniU+hvTaRV44+27mMH2QwL3m7af1h5cfbrjvZoF2nBuF1tIkMNe/UIv
tS+BLXoXKRGX0CSU4V8epQ8z+54N+kNECde21YRpdOgFM5llj25SDsOi47bvjq0mM0eolajWVEAm
hNCYEhguvo0mvlaMBIJ5Oif5jUf4LfKNsC1oayzfy+VDzS2oyHrL+BkVUd1NY/6+s627Ebw6LvFa
GLLymrN1NabB3QWTlKTSgABpRmgtxp/u1PaZxH964NkJZkgSOAu+PkkmSZm74izoHGbc9rV6HeRG
W/yBVTp3XAmQLNDqOoUy+aDVQbSvbvKDKjGEorEZ/5xhEfq130GrhFENMfuC8drd87aRyaV45Z7w
fsRxmJ36nZFvo8u/OFUXuZ+ORIDx5t3Z9cL4f0yzqIl5d48nKzHUNJzSn0VXhu2Or2OWS94LltIy
enkLL/DUUqPfw09abWbGTz2dYIKxRQLO0N2CUQbz7pYhPzmkW7V0bybyTn6VoM2OvpnEZdXK5dKl
fnWlixRQ74qx76nuQ+zcgf0lYvQe0GGVdHKvW02xvnfdyLIFDb5oTk2hWP056ZlokpQ7P/X0rv63
X4g2MpUwmbiy+dGuNBkbL/ICnGEfbZlpsO8auY39sSde5nVJ37oVE+NN8g8RTDHFlSdQTTFjYLqC
k4DWW+BKf4uhpVozB6oh+YXhX+WhQZxE9FcllMxIhb+xTLHqNUKeXaqd/mN/uc/5E/jTGaoaTu8y
H5du5r4zzB6v4H8h2qtZEieuV7zZcIkikHC/ikHy02Vxrcvs9u57qui8b9J++N2JPmSTrSGs9Lqx
vntt9UjS34UDeiCRflDt2WsZV+LsRyKUNrzMpr4rwFlHktFGBtYe8vBmfW2auzhisaQDXXBSo+rR
aGRGc70FhJDOK86PQD8AeX+LjIcOzsFf8+FIJuXY+our0xTBqRbIQoZzO3L9YKd1kK3M0RQ2tdLV
PoEe0OT6APLs48H41ZOVACcFO3PQXi0lTnSTRgSrCqQNshqtBYIffqLD51HuOtSCQ+pvWtBjvYfb
+X5sNH23Fb6cRgox4U53cvb3GtR+1H0jYulMY43HNCF1vo7QwuIN65KLRsWP6rkibn1ngRWkqq0C
an4kAy9oh2oKBofk8LEuX4H0+jewBN7AoZzuZiQdOVo6h3D7GnDWhv9p2gkKQI+8Ujb8tOJ92nhI
XkCBYO+aSFSFUIWmOxqXn7glD024jdyTCS/uSHzfaAkPMhVe45HU62G1gZ32j943gsRIZKX1FAyr
00ZCsUWTDWyr8QXSJzfH8VIvjiyttJOlY1yyqVn1IS/KC54aQaDjs6Wls6SrgNJXNpMcTNDI4VU/
Po4pyYasdYnS5HPRIyjAIAyFDDDdSb/jKOFM1hmHlgE92k2qu4Rlehxv3nc5mVNFAy6NOi1gqwYz
lMqJ2T1IQ/y2ey9jGOxNtPuv/ioo+pNaCaXmAaB1y/nclK8YNFfwd2OErgK5mdGxIpfMmORYr9r5
utMT+Offsutgw+uCXuWNHISi0PK9hgtpZf069zMTt0T/sfDNTmHPAy/ZShvX68pD1uJT+KVg8TnT
fXA+VyxzPjgpNIzOgvy9SJlhivkyJ/HU33sZLewXX9886Wbi6370C/7PO6Pa4Jk3yBfxmu42/dtu
LrfyguFYI+EG1qUwskqYu/f+aWkJ+acRgQj+Nfx9QDgKf6hjQ3/10+73aCUXi/U0m4X2U56e2hHc
WZC9P5WEzEfyq4O4wsnXmz7RjddVEoyHSwUUppML95z7vMyHnDSa440B2go6G4IymSEJMueYfwuC
DjJCo6PmpHbwpWwf1n6IjEnaqsj4QlP2gR3WFQLC7nx3u2OxMvBFmkgb29lxKan/czO4VYS7+kZ2
mdd+DwzkvI8nsQBE45jFjdwxd/m6wBclSTEBtHQ4rpz5OE8B78fRAoAAnPVpvWR71/hPekl8YkAi
ZNEwHVPKvo5kTc9e478fJ4GimBg/vjNXU9INjHQ40z8nHpAICthlDt74VlbtjpZ0y4I2vSkN/x6Q
rqGvIc3uuN2sg7181Hr3CoXrE4KZu2q1mNLfBdRysYU9vvsR4YrtsMOHr5Tfig5Vt+ph22IIzJlB
Tmjl0/OBlD9fHcaOKrDFfffNXGoC7OKNRafqlqP7khAQq7tYo0JhcRNNp6wOaIbQv4yjLXvPabWI
dgqHLyIGI2zy7Hq6/RMVGychRumvryDdeICrmZAmN7R1/LG5CRpD1Hg5FotRwf0GwUEXCWqFtzoK
1Gr1eztGuepAFrO9wF9KWKyeAAzOrowSPfTLE0O2c2HiLlJxKLZpH8Y8+hog66VHjwyhnsjcJPng
U7I93vdKY6L2kcUgYRHz81LadyduDj1kqGAZMWhadA9rg8DS+CxQgrXBn+pOnEoLRsqCo/dOJo9A
fnHy5zcIHABS7SzN/jGN2vH7IFk+NapD8xod9xuS2uLKCMy4o1y1JJUJuVqT8POvcjBq+HLMVDi9
lER79QWWFtdqha9Lf0VqBjFlpMKxY/38w2MYffEDtIWb/nbwsoPzrtGJlbvQqrR3zmGGDub3rYhB
5xsdDJNzjCn/cBgOZ+AkF3IeZd3rop49DE12G1Q/CcFE+acKgw4ftmzck7xbW2YtFZ3Nr5VXoax/
g0piBQ/Vm13M61Lvo83JUo/H+/2i5CSB/AwLhRHDdIHqyadk0MurKwYCbHV5q59F11IYqwwAVOAY
kOIG4Juv9Z/N+VCYJU831jHttWIlk05jMA57rz7b4tx4Cf1q1zYEIysAm3IIxBsOTCJ48In6v8WQ
c+aeW7/gZKvdP0a25KtYso5wbsgf7E2D2x6/gMqTF3p/JQRNAH8jzW42jIMeft0hYM+Djzwl5xWR
CmRrF8Pvdn6L+g7gf1XTBEIliChomlb5rFNGONvPZykF0cCJ8A44wQgZK2a7i3deS3Yy84pqQ4gR
f6o7wpcF1yZHAuFrkBt4W/x9rnhegxSwtF/tJ+HH6/TJ7ZQZQojotI+TUphDgIT6GnC/V4IbE59I
BRbMf15h7oog6iunOJM9S8CDePhXwV9PgHPzI2PblDCSbVhkRlAoJPEzSmx5zQO5zuXkzBTL/MI0
i9MOVLwnbmgbVOraxdkE6hMOXq+cdRL8yAKtYy1miRwAPtnMGCkqGxqzV/Pd0EnKcYchjCjlD7CM
PcxLOx8aCKaMvf3WJg5QFOH98c3zhg1m+I652yNvM7wwOSNrkymkE/D6RlVlp8Aj5RJmPgmSg/WS
wQ+qSmNFxYOacePdgb0T644rgfVQLODo0RDZXarl/LfSq/e7JgDWUW3xmDr/pfA7tywqAJp519e3
omjnrvhib/KZb6sdWeYFRJ8kYXw1hfZmnMthZUsbfdD8AZfHoUEId+EVUaikv5YGwwqXdow93y3D
ZETVfJO0W3vbsPrI9NVCfEanzdH2XywaHO6fGvr2t5fqjOb1LQzev6mqeRLY2qRQ5PmjHnM1BuXB
Juys+aXvE+o6LfYWiDaLQLvAhHqlZTPLyJ+CvJ819kKp1IWAJvoPoanDI9yONM+431rKD0uqbB54
ujNhqQK3n/dxjgtzej1qOE3bAD/Mvixe24ttj+Ft4WnUkEwFzTHR3ToRWLXEkavAT8Jo0BvxNqBQ
NCLDK7p9LuSh8ZadJuCKKMY8Wm/AKv1mCUwQ8EBxJ7ZDbT/8UqZkIZ3FrEL3o2Bwi4TY/1wq0Ul5
Okp86ru6wotoi3UjJKLTBrgXHb8UeyDGn2OsAdlsNAjiwymo90fNKfBVAKqsIVOEyf8EsMcMIbpq
SMX3F+dWPNcbSa4j8/Kft237FF8MiqyTRznrMvf+BuaETzH2J6gXe7Ujlh1ILGQGMaAPZrWVVoIL
JG2u08WhHPx323Va61wTzXjH2os8kr5p9RMqh511Sf6dmbC4rQx5dDmj+wXARyk2kHmC/KgVEj02
r+Dqb2pMI7YUV8tCcunADP1dbDQOkPdiOKHi84s13LXOvACVz3jnC5kH57lz5G9gTA0gZUT74MGl
L1pVVVckuPaYNozuDPKaLItudnpZmVXjm5TfgVcu1C6c5G06kz2OSIsZMR/AE1xzmZ4Jlyvrtn+G
awEExAu/d9oTDksfapQ1nVxNBAUHDik/h2NIQOAWsGArQAH7DFerPSraRB3wiT/bOjSfEiBMK1p9
6lZiKkqIwblmncapBsA440SiWYm3kRRFo9W8t0DvD84lrhclLPuQTF2OoOQ9W3jF3fC/va6ORBrA
vIu5zALkh8W9/NGReAef3NFRA+GuA2Kqe9tuQ+Z8mp3JMc3+Im2oDoL7Ad+nnM0r/0OKSHhY9q6a
UtoYJO6xoaDAClGOpW8GChT7TFJbhu2zldF1sJ1uYDXQ6X/fDYqx1KQqs0RaDIR0AgAUfjZ185c/
T+S9sDK9jzmi2qZYDTL0NtbTI+iBmEJaPh1utmXwpRoS6zlZtwWFPpIsZVky8683N3YUtCJbniEZ
nUa1ycgIfuqrJyaJHG/1zJB3404WnyrWZAjZpC7N/HxIqAl2OhQFbkMhQCIsK8YUCRGYVeDkyV7V
ljf/btKqQMl/2iTa1v7T0wR+mJsVMzFfdRt3gwQj2xlkYZv5ABtNCf4/remGKy3jW8dYPFZGWTOq
7VBZ8ElaoilVeCp6wSP9c5kdMGiojNypL0KyepRCoLtsdVPcQLe/3JKXS1PKI9djjVfdmdD4/lap
TkmToY3+SOoH35Kt1ooHCYXNNxhMaDT/eJGNXVXYx27n7iCy/P7XVsptBPN0/xBdS+ahADbQx4cN
xhkWEGSglJzeOhrSHMJOEmI7ThlqVA2yNsMKg5GaeujwWMjeIwqs57+eLiQ/OkICsui/wfGz5KaF
mhxetOmtzix+F90H5qOtrqTIUnInPlnmFRDIo3G6qpIcD+DgjzsDyEbDrJkL1BOYN0hdgvquuQ8z
Ksiq4OEnofUrrornL+UVar6xBuz1zh9CXLZsShuGooXT+wSD9JTg6i6qziw5yfHc48WUXYqA2Oq8
Qy5F5ljbmM1vFFxxZzm13WtynkHsIfy+i+MuedTWC2Q89hwNJxovd8kyViecpFjP2wkURX74YXn6
qwndUnn+hVraOHOoSSRlt9upj2vXjuQDrJ52x4Q0UKojY8M/UwL3wpIpFdfWYv72DLYUNcIpKI6V
FM95Tk2vCQvPDKpdmWGK8zeB6ueO3T6Qhrfwz8KsVFZjSLkky33EVDsFoHFZNOabkB9sfXgTvrIt
8JC97DS2ackZw2lDJiDOgU0Y7niyZLk0jSfbMi8PmRQD4Aq/c5W8gP5GPvIrRvqQFLb6Lc95uAds
1SzitY8pSFR7CBgYadifaf9ftwDFPYLtfQ2qrfg8zOSQL3rB4Sn6t2TwJR00bQ0SJy/iUUAI7eWY
056FtQioJfCvDyALKp3dYGhjJ90pHKC+P7WQRfmGgX8R5V/YP41xscbxyNbwCFqxlm2OpPnsYglE
Kh8sn45o3pUlAU4tmettR8q8/J9hFBCRBxzfO0TSQ39Gw+9Zwr0f1VRQB7oCCHkwd0kpd4KClW6L
RL5aNFgZFJOuuX5IU2c/zoeCk3/QiIfQyp8rOoZJMT/thRE2sVROffHr8nfrR7U/HjDAbZTWB7E/
/LKCkjOute9lFB8hYtLS7Lt7A21R51S23dni9e1UivasmqKq9rAReQ6M+W5S09suyJA4qjw4g3zg
cJzbQLIxGehx3SUQM2okV7mnmgHD9VKA+VuCnPZvxwB5GjFYwFDNrj3BlSof5/SyyorcY9LO0kqM
sjgf4opxx5ybtyq25I5DYkAAJbzI82ZZvdje1vCGH+M0h47Oz5Cj/bmhakO6rhpVkSh2sY0QyzHd
PR/7pRD9IVorJeucHGUWg783juOcwdBPny9meu0OYrDT4eYnc4ddPG5VhWZhY0AYqspzLxcEZ0ZQ
biCNlky4QjZcETOuYYxIjznq2YDLyzN5Ju410q5M5mNShuKzfuP5yiPI7Jls7lkOWLUnnacHM/8V
Hl8AYMY/+AMph1RQozUputgrQjFisAb3WuNVvoH8LHUk5jSVZ9d3+s7rZZ3zH50dGCMW4Nq2qUWZ
yrPeIK7+MhB/odHrzAwvVZA/Llcs/KEpoGXPP5l1usmAdiFb1uri1mVVxUQNNaflK0tHlotwarxy
JkMWUMWsYgwWBR2I6wblOtDvc5sFxsSOX9tD1IbSLVsY5Xcv9ljmw4Gr2zRl42FSXriFao58ZlB1
YsHJAc0m5nmVaXth5NEoK9X5rlFurzN8PfnSxarMVzBaX+UEGGtEYLpa+gjk9MVIrvHfVNzFEKK9
S2/1Kif8Hyp71Q1tX2lbt3MtSOiwmkrZSQr/pcxDOgfkWRafqOcpI/QonohgtSDORcyeowxxF+g3
NbWBeFpzOEjOM29+/7cAeStDYV401wK4efHEuAhri/ZV4HkEi9Dib8p/YkseCtpwktB9ng7V2lt4
6o6XnlYBe1779EZ6hzbhO28e3968SrAhdRQe/5noK7WE5Ik33AKGLkE7LpUcOf0LnmDXU/avUibu
ppk4Ntq0/1EP4Czv26JsPuAih5fbJDGtKYuCEo6X/WFt2qRdqs3LT+JPeg/96jaJXCbwpHzu8vN9
ZS5LDMq0PjERchVuDXXSkodaJQjltaLu72SHKM81AvZshX9/f3wgAzKY2i+vu4Z3DebAzcNIJ945
RURWhh0L/3SwoVfnjPeEEPnAl5PQpHqIm4BbEF8FgM+zZ2ccE/zJFYpMgTKur1S2fM2TFGWTxpOq
D3fzKjfl2k0dbdyakB5cuuaMr1rBDff02rt9qPazCPwvuiNXXg6y9c7o/fKrhHtJy5Z+o8cOXmzk
dFpZYj11G7Ba3B1IGwrQnfhPTJuWLD/LAJBpMVnntb+jQPC5iAuoK4H/IMXT9wG1R4pdNPPQaDf8
gTFkPEaaNwVVIvzbbiAK8vsMuexriOngcP/NidP39BqlYYdxgfW3+0XXM05RnazWEGcvg8VlMjGL
yBV9puCEJra9aCGCJsze5Dq8HuSceRfAA8LYjo/eqyeTFUXYoqO+1KZCa988OhoYG4DiqEAk7wqA
qxsJy1NB+IMK3WgFlz2VDd4H6cIYw7LL/YoJxdeOuRyhXL1LS6QhuDNf56JToVVGDIqjfTL4fKv7
2qQ2ua6ZqMB1ejSJ+VSXwiGwPHyl/OD2DkIoV1ppZca0C+EHdds++lhyI/VT/mS5RBU1vfO21ha7
zSyzFs3kYOgiw4gRx2klVp8vE6gw9hayponPjCmZJrBzZ+spbCwGnt+4Fz/YQ6GSNMMzF3qyx9Fo
2nj5yL9sY0NhFk/bdZ85+cK2+ZrsWIQKa8upbXqsDasUYWTae8WTdgEmCvJudS3dSeAG6/U9GcnL
OZkafRZi5QNNt63Kk/HjvStHDNICSU7t36GsNBwX94b6NxBhS/dEy4QnZOAp3B7rvEKSBw3rBtHm
JQ+1BdFivvLzObuWlUa2KpLAsYHzVmP1ca7RWCtNSJAkWzwpnJA1o+hghFUE27K6R1vtEelztt4G
mx2OSQEf32dY3YNkEzJLmwcrzZjZt4fqoTD0ii4VJBBjRAk5u0nPt2DHV2Jllqb2+YPIl1Rqg+Cv
uR7rju7L/EHWStNzKzPx8RB/2nEQR/5e05LXLuz9Egocsh3JDKAVmuYDth+yC/May/uTKjCe1X4f
ojblj9nkgFzR52FYzabHsV+CA5iXy76EC0Un3P8uTtyzB1up380Filp7K+CilFb7rOLcN4i0ldJX
QKmp5aiMr0zaBhVfHEIemOYqJ9GOl5MH1RAwfhtX7pbGqWWNdjIlYxmBX4b8mEguV6jA/1BC8Y3P
dR93iR7PeN9x/2wxgj98NaZScB4AjXapMpqhhb9tJKMw+hLEfD4lnFgkUb5FyEjXaOB4avSgZnQ4
HlcjCiLY4oCjMZ7lrGL5MX7p+9Y9DUVjUjy7PUIseZap1QTzSTlRljEE0aaWQ3o3Sal80rAs2y5R
G4txmn5sTac16qkxak5SjT0YX+OLmiBde3ZvrzjkkXgJzo4Pi/+V1YwJdq+yaEuY2xU31OtdnvWG
KGULHQ43IWakMzEaGfZQXNrh2QUqA+YnHPoSL4w18ZCOuPozTUM+cFleYvyMkDqK2jmROHX43TJu
kJxNAFFGQCKetZpwM+vpdI80ONWHlcdvVEzfBSwji2ekBSIi/5NkR+7Feu3/rFAuF77flmsWFyrS
GwE8YKdobEaiAo7phg1eEmHelcSFN5A/jr/m8xzt/S4j+RwRpTa/jCOyLx4tACnbruwDOic0Qcl6
VJFxjNXT7FBKXLwKGez6z31R0d2mTdxxkcPhs6Dr/wwTimTjfTafpU9yvzGc8IzcfZ7o2FN5c3n1
HCrqzU33Eyev8MsLisuTEqOOUTWAS5bDndAbr51BGqk3szZoNNCEFj71H+vL7EATEUihKY1M+thw
nUR5/5Xg51BCn1XzdUkhuoHHbjIGccbcwvbzHb/Oxok9Thr0bC/x5m/5SXZ39gFNQI1reOCkXmYJ
eBZh5biqUVdGvGISK11bW53Znq9Dv2bjxpOC/67DkZjF74OvRDQT76WisMdzwT12+MViR2Q3nHBa
NNTfym/xjVh5dBh8gwPCPj6GdfL2MSW8X1UeJ+JeAHD78Q3rprMGYwXWc3Yd5U8xwDNIx0cZDRVG
xQ0eNJ+0FP3LEhD7hWmfKlS4/DDfNyujIwildaq4HQMLTgnoAPQtGlzRmFLQuousKs2ala9dUDkg
Mn8Ve4np+5crAZspxB3bcC2ZOxF8t7H9M8tnyDja6adJMlVzyUX0/FHnAYxA4xq2ymcY/B16WKwg
JN+0ZrpBVh9UF3P7bBDEnxkJFxbmRIS05rz1ud0cr3jg9gOkR37UeLHEQYiiJqpCVBxckA1Mr5Bm
yVF8S2T0oVudu//WTl2QU7sxmDgUYiPjeheR8hKKjl0du5/EIG+MZt9aVL/Lw2iMWPtaords3hUx
XjjPS2S5dSMV3gJaKpdIzXH/x4fWrPPn4b2WUgZCOPoPimbY/HPDlrBwQD93wYY/oEp4ImT+wO9j
DyFXgd6sxc0/nllySpxXhSdXd4OiJOFaFGU9ZtdGMvtJrs8orFIJOcUaB/KZZzERE8hVjBY6G1v7
7CdP7CPGFcOC8vPwwTvvJUbSOTthaWiqWP1RXM5NiKeVG0qOhWmkXrHbPp9IwiC1+t0E5/hUbUFt
N758+Z6nJH9Dg8mQ5v9sWJ9Tj57gRoJn5QjWpp/rc4Smu7rWFS2E4AHmAgVkBtkUybMi0I9+xYki
+lzaUn43omnqv98rv8qL1zs7BHFzRtUtUyinGrAGlTub4uenym5BIQt4TfjfuGAryh9EEErdlaeB
KPrj/ht8iKOF3N5BzT6szR/iyJUwA7F/e3E3JoJA65q+Y7jHXe3PQd0CowXZHveyHL2E8cd3twm6
efdRX9Zaoh73a9xMNCm/Lqamv4Eh3VADCXut/sSe+p4F7xa3Rr7+jvFBTwpQ2fm0Li8IImjIDrg+
o2mnjlRO7AYYsoxxJ9idr0ZUu9LZoxyjQXow/UqwQbmiV6PAagogjah/O7XvKizBCOG1FeN2OHmq
wv2pnMKMIlfBm265iia9OY2M2lnIKm9knaYNXh/eCj2lmPaD0THRX+IC8KCIAPn5Y7PT1XV1bCCy
wW91U1MF3MUreXE4m4ty2wLsfU1U3cMylUfNLomlNL8vcCvPdopFkzgNR9c6BP2I9lgm3jnKxJKl
N2l57Zi7VK7ESr4wV2ARG2XWG/d0uY2Ab0mrXI8Z6HpVGJqSeBPvOonTpN33X4/tul8hcvZvHE91
8BKD2jy6WJRAwK4HRphIsMRweDoHSGnZfG6KfLO0B5J3YDH8r3CPxnAi/sazlaTSszMIEKIaT1nz
rX2vhT8JBoi1JMQfJKOvq+UTYpTzj3ty9VfsTnrddJPi4GubrFSgm3dGu+Bi2rFOp1fjRrYzJjns
KqIGoUv08TeDVcTZRUrMDfQZJCoBspHUdBQntOo9tNvbAKNallyaWN4Mcuvm9ZbfXjL3uVzTB8tA
PiKAi/gGnw2472rrPWBFkVicE+2tOYcEuO6IeWmSqPS3L+8P5SJjZLifpx6vAi6zBINPQrNyaGoP
4JzqKOk+J2e8qmalOdGMYWookWV9qlobvmqETFHMYz3B36wlhfUMsAcf2ldfsu0aTJnB8vKdbCxH
B2fpPXxq++lEdoJHy6sQ3iQCFDzW+O768zMPY9MsFv6Y3kVJX1UXknbJOLSHqeQ3EftZkObH8Oy1
Zq/FOBbXXBTfxfFO3wUMTaVR20l1DynjnLYPwLQuUgn86Cf9dKiOp9AyVz3Q2miKx1xteVDxArbO
WTCTboDLWpHq63gBFBE4357b04F5SDHEYygOcjYnK6dwTZ+xw9bqsN8YqD4RJwR4AiPz8Z3FxF2v
506hPCVxtxBPKX53yfQB2EDcQEXozDUqBAbaQJ7d90vPzzAqFfI2+NVpAd7yP5HztgpbyBaXvhhs
XIC8+NjNfbGhInm2Wui7QFuBrbPNRKWCOwK29W0NtsBqC69AgFz0nWJj7uCUfDgzx10qTj7rcVPB
DaU/aeJorBmxfWwJ32XokqOEHKdskJiC5NP8lhPk/zWsF5Q31olMIT5a26isjuQlHBZvx3onrSqt
FXj+aQxHvBjnQdELbrGIaiBu7gJUNgFM4Q0+vlZJrtsfNJEiyBQEB2XricX+DMNMgpNj4caDmoDs
eA5LOnFXDMw1D0LbYKSNnu6n3pd96oEaLcOkglKdMpWpAeO1AtbPS9Nw0RIRUK/hAXtaNGSGOtdQ
ZEYlAbKRX6EUXZ2yeLe3aU+aZCP/J1AGGyFZ6MYVLz7KOdOoD+pFzDR1L+qpO9oskoOjdyWK5c+A
cSc1mTXn1AapU9P/jL387Wh/ddJQxHUB0L+FpqbUszyoDPJJcR8YDQjpGWzhgOZ2nWIUzZiPDeGo
szyW+6/pinJOgmA6EKWik2soLfdxpsEiwqfM283gy9pRN2VWsdzxVO24evtBWYMiPLm8fsZwLjIY
Ahyyyj/QzIChRDtLv6Op6sBHe+ECmKPYI0zNGRrJR0uwQpLM0Gix+nVcTKZvPv0R0u97IBy/UpDt
Z7cUjlggYczwUdjmo2WjKJryfyehzOE0yvmuleSrzWxA1LhKqr4+N4eYnIbh1ab0hwmJM+NCC1Tt
pJvCtCveLgGo2oTGF6JM2E1NdvddNPDDbsewL2Od63EWlGrkIE2QeDMbrTdbUs72Lmfam2mny1nq
0ZQlpGESeQO0dTaFYqtBJL55s0pUZYMEHZxjnRSINxDXNdb82Z7ghCfEhZUVJPGnZaoD5z8mnaz3
EabThYVToFB728rhrdWHwjOCZykMRpr4edAV9OFvZtqKsw44ANAjrn57dAo6cjdAz3NYYFt9bpJ7
Blc12cN+IkAwgMk1SnAOwFo6pQg8kirYNJR2BzrGmuxydSYUy1VOs2oWU29fZI5baNrevO66HsmO
uE8/kuibwoEfxItRgkGi/DZWp+a7RiLC3qxCmnNOn6qsNxriusTUs6BaYHpML3fLSfWQfY2kwaBo
eyVCJFg6N+5qfLGMJdESJFotRHKISC6j4kNzKC85ukN2uVTnt++b7UfXj6/l5DUc2W3SeMykLB9q
rrdaajWCe4RPEtopRTgx0Ve2dmCtApYBAy6VxXFMsDnpPlD1DR7/rFpZg2uC3EkS0Oh75IHW1f2A
utt6h1sUmqSOZjDS32nQoMvquMwO3qEHABzd1NHdMgWnkg0hw+r3sDlcluQ3Z2hdaDgDB+ARPkQg
N3ikKyVvyJuqqRhz07UmA86Fcb41/AiM1CTXJEp6aLgtrjDC5O5fu4EQLd4r9k3ysnSVU4Yvc1PF
Di4b8hj/eykj7SrSo2Oo5Hvko9KoZTyEZJXrNj3WsluyrWvykDkFT/LJvtOEfHR/1kPXBx7JnAbo
0nJWS75as2gLTMdFcLz1kFcnypxlU0SlTAoTEo0AlHXA0dewH/F+36qNJbBTlSwOA6Bs9AEEW7hT
vpkaGQuNfd0VcGWzCl7QPN2WILL9+so0l+QWtH47i57J34ica7KuMS1ZhPk61aUPPEKQePem3xUt
agegzU1wMRvJ0DIpy+GgRD9l1JpGIc4xgkaVdNy4PhO/6Ku46b07fAqWCLwgKOKHwZXnCI4quhHM
v2tOzdC5Pwv1hzMS8nO/dnO1LkQGe/o4yiuM3DYJUUfFJOPzT0woB2JrJRNolu96oe9kqlX4DRE3
5MDNca49TwIptFz+4xbhlUypag1h5YFm3RwNnKPYaPrlF9xY9wCgkb/mWifG4eo7il/52pepmXBy
5mVkfNlSvctxBRDhm2wXFbn8g/+SWc8N9lxGsecW5oB3Z2Cg00WXX8a+pDwXEjqjJgcM5Qx78DAf
iL0fQsubpepm9eHmoVDgDF8B/BAcYQGMU4EMgVSNiX7Hb1NkHslhYZz6a+qamJvBRQGAzWudRSYQ
4yul2FdmCUER3OXYzOQT2b/L9hU78Fx8gG7c3sAtotdy8yx1k/1YLB1RyoPK+CvnHxKrWwjkWsOG
nCrUVZZ3k9PpoiQ35/7Usargqb5KOu1pGP7WEgxTsEZOuQnqVs3CYmxyPAXaJ+AzM9JOV/CZGN02
/D0qi3RTvi9/oJ0GcSg4lgd5+4ZBJVZUpO54zsz2Yu1h4YWgBlP1uubHC7vwsW4FigsRYksKBh+l
0QJ7suKbHtfbLWOeJTl3V+vuP3jJU1paN46Dy57dOO/434S3eNLLPuKxly5mbgfpF5JrXoaPXYa/
B+CNXGPKVxJEjL7Axe4eQKNnJvoitYr1oJioOy7TYKICuc/LIufdM9AdIbQClNOGJ79cYgJLV9B0
7r5zwztWI4Te/zqdHh4adqYj3vHcZJ0x06HxL7UeGm9dircB/RCVucv9yed+Ve/+i0rCXkG+rNZS
LFu9iJUzo1fwZtGz4QzGXIUmNxnNoIveJ2MOfCmCaP/dBTrvcPl7PIxqYSVYln4TUy2oaTN//+BT
EaL8kaTUjHNblauaSWj/XzEY3IbenB0Z/+kg+Oyp20SIFbo97wuAgJv3vLxsIgIxwmvLKGlDZA5N
y+ltBtWItNXLEnz7iblYJp6DDL7PvG/gVXvde6cLWWUjJeQShApf+qil0gIOLo34q6iQpo7errHF
8/eZoTXUtn9eLHAOlilk8GYumiCL8KdbQwZJp4wt8tt4cvumwNxkHhnXxQJK1VNvpEoONhkBuImf
6IF6kKyu+0KhrWj/I+DQRfp9axKTzKWhi3b+kMWUWvJz0VoNyo/vdfnByxCpcMaYBuk3nUZe0N6p
CM0MfjvfpGZBvi0ObhY5qHcvs9TEnp5Xp4dwbVZCCUDW466oA9tlbXAilDcmNMhT6rdEQr+6WuEM
59QJMiyo/Wxn3g+FMwG87l4vh0I4jLNxRnI9h3FJWt7xcZE4W6T8yANQxPxUh/XlKaCtZrgiCk7o
ks11K3eF+aKvFtsO+KsgIr/3ib9aR21WvIV3PDp6FpxqkUbW6swyg6HffUsA4t95W+OyaH2XCK8Q
3JjB4R/CeZZpFTFP+QBfUFG6UDDd9896r/gn9GM/fkAocDAwiQXsiZOvQW/H8O6nCv+P78QmXgab
oDt0VuV/p1wctLkWlB5fZ12gyzFoD1YigxBujODG1WAU/8cEOpVnTnn/CzjFD6J2IulHwJ8snx1a
sGe9Z2fhorGnmg21apCPyO3kfoziUEMHO0YND/wRQq8L66lnbJ0kem8hpT6FTAxfe8vqENMeli5C
ldRfJUd0JLNqlUc2HunQugDy7lSfEcl3x5ZiaWYxGaPec30t8wSsqaojWXRaqb/DK6E0N3FlzpbN
RFzOi8g2+jxSfguGhimBpwZ8D4uWUIjQx9WJ7XQxtVPSbcbLuRrJEgDjc6HMVxkzszhdzd8bAL9X
WqWI9nph+lJSDhs9x8RzUBzVlKm7byMMC+oa/wd4hfl9eI+SpYpg6EEZzYtt4JLeByz7b4kgyIuB
zwqAufNadyUzU5tm3VoMKQetfAhEM3OI5shxqQgH6tSToROS/2CMzI+FRunZJtEm7fPR72pOW3mp
O0vAtr3XGnjaBaGXVdo4uy+Cs3zEVNZlR2KfKVWp+s8VCuOs6HYVSWVRs0G9yS42LIrQVzTugRO7
zRI9PoWYXIDmumGW+R44bw9lJqsWKoTnTKy85wne48lxgpu4XSbj6N6qvAK900Am21pL7KjQdqSp
A6nPGIwgMt0U4yhN4LbFqss1F7CxnZ7C8xNf5DU7O9q39PR5JeItgD9cDewAe7b6rTTiFarajaQ6
NwnA/NvDs1D/lFAhU910suYAtGakhlD3WLwRxUDfQwIbcWgcBmg4rS0fykhchsl/8LMAZH2vHlZi
i7HHkzrEnb5RS9B+YgkeTUWCYIxQtDY1yEzb4pX1WTYer5f5EgOtoPt7S1U54jRtja3J9gBzCsQC
bO9qry7iWNpQvSUEiS1/GvYO0Mi+cqrMbRUOxitW9mNhvum240O1tSGXpoOrrmwSHwM+E9+Y9cV7
SqYq9JgUoNKUlBeC2emjg5eZ8Y2DVNGccSjjCkcm/cGtIAm+TkoSdivvWz1y3n/tZdOWaruqoXEM
0Hmae7ZC5m1+/YxH+7d3LqOIhwPDzyND1YaehyYR8ErFOgn82ql31HanW1JHoySByDzcqjdRqdhV
lnpZFohO+Cuj3kZKzuZJfs8gvYeMHvi45Nh/9Z5OjQbYpvOiL94Y5O8H2X8q6yq4sSzoe4cJ691x
LparO4rxhPL89DmP7Jm8in57OIftJO1/iIvWa9YWEwXln9FMc9mVSHrrVaO+/K5nF5iRUL8U285t
HKkbfWRIbmsupSnBLBgXIJRVR2lCp5rdHu1NuO/1YKBYY7tkW9LaR0ZD/8UtLdw4m8aM0ZzxxHEA
fwudmJzInAQSYhnBXWCOq6773yHbilPzwcqCwySuziHdz/HJno0e/73olZi2lyjIY5zRyx2+ENGx
e2sI5+cT3IN3SI+H2ppljxPlXeH5+JGxqarVwKkpbyUhm2uvT6CQVIW8b2xNZd/mwnG9xu3XDsFO
4EejW14wtxxQGbT60nR75w6X9HbHJvDAlOSHmPIjBMOGWMlik7lCNKOuoIdu7r94gKtg5K86eXj4
VX3XSN5ijvqmKY9y5A84hgWE4NIEv2Sk6IiEsukgGZAgmEiIuQ1I5U4lLcMKEcw4Bid6U4VilMYa
5ptJwm+MkRumHxHLyKakddjNhWOumvUsSY3SlWQ1AQ3aWVzKV4zLr8wSvyOK3jUeGtQpg2gcYVht
6Yfn9gvUM5Q0/UIv02XcrtcyoPeXZoKSJDTAUZgR1wFh3xtJ7pivsDncAZXQ1bElSiscsOCxZpfO
2yxhC/w6BZo5AFZDqN3H1+kp0BbuCeUnEMbW453ihP2LVL/MhK9BWmmURCXUh8UcxcuXtFH+yoOO
EiTQXAyfTzIRBYGjNgFiL6uDgdSBa6i7pZpChv71IVfDRvxP8TqwoHpkCvAyCWuLZr39eV9Er3Ko
RYBwup85soTU6lo4w6yvMsh8DOPbiJXes9tG/Eeb5GgtIHKKl+2gNQvCNoEBzJWtax/dTNWhwh0O
zgjx1uROKj2T001TzMcH0hGRystBuHBeJ2ZFgHERRRMM0QbxqC4i9P5bNCjOJzczR595dYpEi816
ugi1cYGzTNRvVM28iXfEaLBMz2kMMr1GY6WpaOzd8y6m813y0z5p+DGdUMfWkP2bS3eooNfvwRhg
DcBEGjGD2mIBCn7nuh2iOdFRfg2jj/mboFmMc0ZbsTROB8kP7mw1sJp9vqquiou+W0bWbuaY7f0L
aVBePP6nmUmexHT9BkUn8p5BL4aRjLcFFjP86IbGOjNbuGdTyI3lBa1wlhSgGXBEsS3GgeNznbv4
58goozkNDYccZS9NylLwyugbYhacfdQDAO4mtq7jdv0Qaef7Y0qVihFR6vAUEz1SAcIRU0FSk30q
3HTsiV6exmVJH/UaXC56WZYZXYallZ+TaW+Dv5sNf4Sdq23bukAzKveEoeSGv8UYLJpX1WHe74df
MHDj1zspiYGW8yry5EVCfiGjK9Tz9JAuBE7nWq1ADpp4jCxjeLMzoXVtrYz2Bs1d7k7QMBSmxh71
y0glJCo9gOP0PvQWLdCogbNwvK9w6dmb5mpaYWZPrXhqAV7SyuXm6T59ID/SqfBfZNpGjGjIl5B9
eogk0UfAlRkkb9zqKxEPvMbDB0r4g2FIzbx4TpJZdGXr7Dm5qw0KDIT9wHYY13FYXRqQXDXyiih3
GkTfY7kaZ6EspyfU1qCCnNlnNURl1Ped+Ogw4Si0q574h+4ALswGat//Nb8NuExEnPTGJKKp2pKp
XoFFvVjhF0ksalWjv/z5DJyITUosADZEh8RVIxdKRkqP60tKSiLhBh7SMolo6Lm7VSnc+QPyhOUJ
guGSN9p5rRg+6iWBisNeqUF0YtAwqT1Y4jWqa91vaDsigkNNyTXtmm16Dq/FP/2wXpueMgegBxAV
fTGPsBxeQtuC7fjJN3p5jbZcdI9xpvgfrYfUy+i9ziD5KN0WXLQvFs3N17OHteOtBCdFWJ1iC/gl
A97roDJucGA7Mw9AC6jj/IW/mNW0Ia+Z6fvvludmh8/KYa7b65z0KNPlSnKI94mYN4ERL7klYlHo
znfI9YB+sMinS8OQQjO4R72U9Y7ttUdoLciEZexLey/XllvNQjP82cJybZsL767cQmt9XlwE/0Bi
HVGxcJ0ugzr4oC1eyREQAeD++SLhP5JY2AAU7tTOw73xrJREhn25m7KcI+L9rVAqMet3I5RJUgxH
QiKtMvvjWbxXztsXo36iQCqwt+EZwcsWZzkrWcMr+WSzh/wHKlrMBfCxmbE+38syfoJsDjHHbWdj
D+2G3Tibksa3jZnAqmRbgwWLH6EUYY6Bq3mifr4jjixBty4W7XqvwgrQLFNl3tOpmTQgG9x3gS6h
6AokmNvUbxGLpbz/2z4aufWCERb7QJcZkR34FN0hrN83hmHFuKgyyQFy0LEuqpZYbfG3HeHtOaGQ
Me1QIVsKHHx5e3tkD4x2vNmBJpVyD2xqe0IVY9W0wszahDho5CLUK+MI4CfTMmHOLFF0irOAzYEW
ueMNUN12Y7pqeM88oNxATXHWIbKJX/wxvcFoKPe2yg3XVfJGY5y9mJ693jxjGVJiznquOE5jjqMi
+3KlYX7f7ZMSk24SrB6hG4rvNzeLjhbC8kJrQeRkDVF6INrRqXPyfGLljzB8wh6GMS81rvpqIsvN
Dcx+ChlxdNcIYGjCxqBbRqDYX7TMNZTdVPvb8iu3C8ctrwLkXLtyY6P7aeWBO5boKjTfUwxP8ZVh
X0DjcmnOSWhuxD8aMeTxnk9AF8v/t4N6dvaznV6AGRb5PoFgVF8+o+sJT/BOT1itKTTUQL/ttb4h
/ZszgF3wxxD3tqiN+25GpnIQBpnldWqu00u5cHBrh+7e42tJaXv64R+dsP+Dl+HVFbdcepd4VrSB
i57XOYr0sanSd5u6f2tZadqsFMtIB0qPHPtp6VxIbmZITxaI0h6OXN9Dg0X4i5kqRmkIPkXDLkyV
kdpoiWMmNsEXntw4w8d1UGCG0kN4uOYKskmtBrcnLxg0qfkyQx9UiASCzyGzFU5EatJMfAierzei
OGkwJCoP0dL4fesaMN+g/5RtAQ9vf4W8equTLuQuaEbgp9W6lunjNd1jW3Pk6xP/gplhdSDNygpk
DO7S4L4dsfcgzwXHp9shfFdXvC0Lu7GnqKptcFH1uIEst33rbVsTRuKi2ZNKrUahHQtxLxoTQsnm
1ICtQ7DLOTWc2O140mzHHa+8k2/I8xHCrYtpqHzZYfHPlzfeqTML49U7W0mC0oviTefP1sEzgM22
Lb80jiFfUjiZQpUMAq0ddhWbvfPBTjMtrf+bPI/nCsBpH3q43zl1AWSizE9yveZ/CKS/cV9b8pxE
ogl2yLpvBj3DtApxhkHVoROiOdL8udaJqo8S7Ac6BpZq4AIzdTN1skcussKQzKGke8ssLrsVQRys
tBbMy4IXRwXEiPbIxpgCHXqjyycyCgA1SsCkz1FZmfEnzCdnKPMohwcWWsncB6KG809ZTQo5TXLv
xt7iMgsvVNJKH2smN0X7DehWIqzZALj/j6yIhSJEljJOlqh/vZHV8N726AiffGHeQcHH9kJg0Uvw
e5W2ecIgIYN3XgkItclwU+B06oABVYgib0xh7odkvm9qP9Vtwi0d6eeqYW/xNWuT9hFCd3/MpvmK
/lfrLggQz+wtuFewHOlH8u4U1SgIaFNt8IFmcmnGO0n3+ypqVkilIlPzPHbbzmdkl9NiEeqOXTEN
T71RifMjEj2sCmOCw+1ti7+QhD/6NGyGhLxMk9BSHIQHzJdSZeDOA3EBRcLhWTe4+/DJUOyr/or9
sKNq+ugMe6l4C1aDqXMgAWMyqjO+iUdj5yQkQrwRjg7ZDHDPfR3uTbsZZq2zriiswkJg+OoEYET0
eCGj1HQi9FEDrSaeWVOHj7fEJ6t4nlIupxXLpu9BJYgsZcyE6dKdERrHRMAgsnLhRNdsEbaR2XpU
Or2syefFLWXLCwLhdUrmsTfn7140lFxhZoZk1eQMRsJyQySnN3OB/TTF8m1RvOWQ8IGz5YMUBBYU
dYwnkjIFmTEOW2HD5QUYdgwJ87NuhpEAJinrs7jtqRNAbExrjcnD9R57kdh9e1Lc4x0lqAZvov3r
6vx8Z72eaJVY0a8bRxRvvhmnuO+0QFf0+Ib0hkgKGathHx5hQ3iqlGSdoKKbn34CD8Isgg3LGZrB
6FOOl1efgCTiDSnOqQVwl2vHi9rBVwMSRtnhVoREVgRbH+5zF/Ef5HqRmFEQxa81sEMITvB+0ijP
F1/Ll/TT2e5r4fn/zBixK5DIddF3voNQtumJe+X/IQ8/1VDZRITGVTcHMKMUOYk1bteoYjdbOgMH
KwSMS5HV+LK6cVMngRDHaf8MSGSS9HJcMzuxiEw73/GWq3qu5rUHNhFVyLWcRIwjzkxUwqzIRIff
geYLF2KRY6Ux+4pYg/65nVnuHeFv57vbFZIgEv9PDtR1ySWIdr+MvDRX14k1RjEy+6PTkQh6OYir
xsgwS8B9YznhyJyPMYE7lSxm9NNrUEYkEn2/EVyACL3hi6TEWtK6fObkiJnUlX+sr83ReMptn7Fp
xnjrSA2RVZGeCKiujFdi3ghpl6A7fiOwzmHWlGF853OcCQqY0NpoYZ4bXjwuBhsJLldPGuUTzzFv
tNQtiQXPrDUKz4Lh89J3f41PYjz6+Cxll1GUa7UsMTGtXMulhk/QthpgNJ9Txm209GJFawE+GLYx
e0L2lZp7UiJ/NRbgkTAyYcG+AeufiQ93lA3TCk4izAVBJZiYGThTJvs6HUrWQrlN4bwFPY362sZJ
8aS/x4YX41Z1WqnFzqFgXQCUxpnKoFu1O8TqxocZzD3iK0sxhEptK0rxOXxjIer9pR1Iv2kFXHDU
vQ9bUyjcSoOg1rZBXPLeUN1yWAlgGKLzJ2+NUhZLQOIez4hoPcO1QlC3WtluKuHQQZYV8MyB9ks+
Ge2z1x1veiY8Iw3DzWKplIfNZTfEOpp6H6bMckJhVhZ3oK1zBo/lviQ2J8tx54k9kZxielRzTRKE
nD65i6aEgDbQyH0Qtqn2QdZLzgdGJLIvYt8rkqtG76bzKNlRPpGzws3uFGGEf1YqF9r+ay00brZf
L29gJfcJKxibYjWYgMdsLBwU69kcfX8dGR2i1ncocbANTWVVJhjZUZfVzp/WhxoDCWHsgndtA6xI
qBT9DkCDJzcmmPT4C1RnXFKC63e6XJpw1Mx2lhorPuMuDWud8rQlCuqoNmdAT0zMiQ2XpxpVKs0b
1WuaeTbgllOeE0jMJfcfNjXXIaT3bkIGb34vvIzg58wzeQWL72acwBvss/xWlSbeSr5bHXDW3ZNS
JF7qzzNrawn7IWwAhlcZ0Ctv7Y362aPfX3AKfOibCZgnI/AmCdlygmZ5or3CG0BF+ADQGyQVLx1+
w4l+NuEM+EpGRi1blOhSy6xNP0CNY277r8tluUKAbrP/fNB1SiAhkuOwvWf5Vh9QVyk3q0mv2iSu
ZrZmD5PmDngVTflgM9eMwVFgKI9b4Q4Agd88oFXllfKSm4lyj8aQdXIEY+31BeVulpVgGqs2xm4Q
6P2JJvhSq2PqUb8gT2KYjEePXm6wrt8tnvF3TtzJB8EFTq8A2FcG3umqkKmdbI1vEGqvuK1H0K/b
uB2k8ym1X6wiPbDugU0CTi1+dJM0ORSabK9OIdY3B2Km4xbDaEfgn0C1I7V1oGWD+viaMsIYHUho
rMGksxtOsa0dYcMkXCzBZA234jrl0Nau3tUxztUvLtWbj0pb15iY1bHr0p9OQH1737h/wFWU7CjF
sGdxP3SP23yJJBm7Y2xBVSMD2b0sK7ajQB4B3s63WOhYpEqWXrtefALNCs7MA/G0ge8wi2Hpm8r1
eZYMHbFjynOPwOdwklGTj66XsgbsbUq3bpa1594JEHTHQ8cVJLd4UETpamivp7aQy21lWAMtAHUk
WJHjc/O2hFLHlzOQXnxD3J+3cpp4aLcqNkBfVXzbWjc0NsqstfDcKnYp4MFa0UnanGb8wLa3NAzy
zj5SfTVOtwZ9HkGWpd9QdrUfmsI6Dik/oT1vhHKbjaHI/qSkyVVX2XkzBT+hFsA5/xWcsSx1pt7d
nE1lzV172Qq8qjefOvSU9NVlSqd35Ckh+fWWbp47W1gSu9iOgCtvZYVz3xQuOOXG+rqS1AIn0uxG
gIWRuajJpicKZhWKoQkQmhRvy6DzTdMEVCptXz973Z7QF1TMkDBeZi/wfRcy5MIct/ZlofXqXsiS
6RCTA3JpbpiqPK35xYuBu87T8q56QGKcwkHJID9YHmvSjaLfCJk0IGoDwUq5NbvwfZsGT+hV64ue
WHXwBNhvNP9BRwahf4dYCCo5o6KX6sFa9B0HUSmzOgK8H/K0DUqiY9x//npmlz82X//35Khk6Ms4
naofImmQozjGiG9CcLTZ3NhgJTjnvMlcfHWw/IKh9Mp3bcUbEX6t7zkPJvbLuyBNyzq671JkR1Np
//MvusLoEyjtm20if0kb2v7ieUknMf+vPnZeIS07PMHWeTZRiCjUsL3rzn+pICsKBr4nurWXfceF
konNLXx8mhJfqNMTro6VlV4TXZrLI+ysZzaJKfYYxl4IbOzR3/L6mvl/5nbzZLOdskHJJ8CxSciU
X3+7rqJEmsZ3vcNHSjSNBNGZ/wWoVB9BX7fT/SoebB9GXeDq47eyVzrcup1vt9Hb7iWehGp7W12i
+Uvj5KRVFXczCjOoeQJcxFhIOSkXkk37JV8xxtmUuxgXs2G0O6s31l4XP9Gc4Zc+SggxvnaGA/7o
IqKMkwURmwr8xBR4bnNpI/2Ytk9Kas2k5DF8wAHhMNUQhpKb21OPkdRZNKDR2jtLtLRQ2Jv1t5bI
qFKUygRmS8O4Q6Oy2IqYpqGT/G3TldQ9ufHZl8VSHD3AxVvujjLDLmD3FrVe6c8Yy6tMuXcy8dFd
YIe5015PdsVsrhRgXZL5gzuWnYZaR148jtD2bYT/dhO0t+4WHBHd5ERNWD2YL/qH9qKCqcw3mCs2
y+vz1J2Bzw5BkKGnkaQ5tF42l/ZNpVpTL3kuQbPZY941lCWOI6dmjPi2R8ORrG6AnIyZ/f5R1EO7
0NWaFo+szu/jOQuD5wHyLfk1RHSM5GrcO1KrtpLLRWD59k2Tq61vSFPXIua8tcvQCYqPUTbM0cYp
BASUcClUFk+HLjjZ8zHjH+eLPf5ybmRwdo+QVVHR6Pe3irMx/HzrAWKjQlL5m1dfkMwav3bX3wOi
m0s42lZE3V8y5+OG2eZEfrVkxnv8vvNDQJSY9Pv8gm3mVs76vZrugd8jCEkxNc5OOZnASgwzSlO5
WTG3hQEcT7T9WaGT6ER+WUkP7qPScXAy91JoD5OoNR6/cpqk5RDsB34wiwda/0PZafnvjHUY2aTj
qHt7QMY2ZzUC1DqLB+PKchL/x8ZFKsLUxAtoAKHy/+3Y5FeMEc7TiCNCsSkINquCATG84cJSaL0d
9Eu5WAPo2zQiWvVQWxiXY1wU+9kSS7b+SLbTA49aX5k32nriBVC6cTbrgVT2EWS8un0lRpBB3pkw
/dwGTg3ydx6gMC0nY6ltmfUkC71a2vpVjSFqqV1Hja3WyUQViRstmC8XbOp5SajyX991UV5y+NmH
nTg8UNE/N5386koT0mPeB9CMEJX3XHx/PuBxnXduCiR+mhp90AGs5dG4vnrgPbUd8wHrwbxBHKdC
OC6tGcyf1F0Z4o6LaEMDDAVbIaOVavxzTAEoOGtyYLREs8I5VSq0KUiil8zQT0ELdZV61Ihb/rto
QAEgcD3uuTSFbn1y3bZuxyAAAJnYSQq2J60M0dwFFcnepHE7nSIMoaeuoQndxW9njhdPHw8U8OW7
pzip0C3XPjo+ppdwjNltZUMVPagZkBgRS8uHvpCA1vDidRY08J9jn0tokIrz2NH32zpVfn/afZOU
AdzAhqy25ZHuKw6CefkyWQ5Q70xScacPZzJsPy97CZ0MmTFiH7LdSnBZfhfl/MUb2WyP5xVCqfe0
zpALhxk4k2TMhtrCdklZl/m+CxnxDN42H6CyUU+RlF8wZL74jUQ4HT1mkTfm8CbWJhTY8F68DUnx
ENO502h2jWNHOZK8P0LYBtt8LDILtMCIQdtXdAnUvytIZy9us9ezyA8N3G7Vo3WYPo4JpWoDXef3
0LHX4LCTQbn+T74OXbsoe4WQNE1h1EVtRuB0MBO4C9z4hvwrN+/yqY1cK38GVMVhxmL5hy9g/ooK
BNuVjufipkipvbrpixvVELWH5HV1rZQP4UXJXxPcQzk7hy+n5lpQZ08mFvRMXFCVt5yQsGn3GHOg
V7E2thZZz6sctdpHigAOMqMAQ+srgtmPxlQqIL67LeTVjZWNcxD3qrTewyZiQzpCMxIAArp6pG86
vE/oj1jNr9VAhpO5LruMK8RQ9T4jBX6MT6imN25oAefLggyN3IH4bKuIprYTL2749xPHO3mLPnsT
UKN3NbE4bJfD67+Alw0p8pPTe4M7dJaw1iFrW0YrxtDCGsrR19uDJqeoh0Us65+Ts/miXH4qVcUL
Yer/DPX7vMdAMpqHhYjJlQM+/p0Icrzqg4TpO0FuwWXxXajJwrcGnnv/yYOGFs/bTCjFu9rC+l51
Pbh7C2sVZtga3pTruLUXSbcoKJBWeny0IgTfytoOaaeZPsBxa1REKMHxsMB6mlGtH9UZUAZm/Tgt
JfOPMgwWLemvCAlLHO2lYyCFd8BZaTXicF0JS2uoi/4YmsykHEgkh601zcMGbDIQ33mbmdNxJ5BK
GxrXpFaWA2Wd2Yn3gI/ikZmLhOH/5npQ6Rh2UBijWmzrWf+wfc9dNE/UqCkRxZNyss1+tpzxSKoG
Ze2v4n+vwdh8UWOtzrDenFSHdCID4mwE1IlJIc6Ur6PCz1Q06PehLVhJuu1/k4MmBrZSS1bigNQ5
8VEsTx5hAjMKwh56H3Hcu8rXN+p5wz3998SR09wBkcRoPI0LB6E+Vycy/QE9kl1rGLYsXx4dxVyj
eRWBvfOqXInIvGlHw6afYOgLLTVN2BSlzupX1xYIZObDhO/QcPniRgI3/9kN+SNJAqMl2lqKIJAS
TDyORXJPpoZRgP5saV+dIil37jB+cBWzRhbuBmpDTD6Fuhg8rDOqYkhFkjCIJlE9X+E0nyDXRBv7
ZDHu0x1zgeOMY8abRu1GpNAQ1Rep6gF8zj+yQGEV5eOHO0GRaxPD8T8ne6Zq7f98Rl9keSmpHHzr
3VJ9pGXh7IKhxSoGMsyxfK90SrrfrWTqptBvVKg3x+2TCTdS5IQiy2L44I74M+G8QC3Vo6wDMWH2
PR8N/HrU6L47J/54dsOkgURn2RluvXme/f6nU7BqMX+gB2RsmIGXVLWEpj/bUuE/lrpJiMYqmjbp
gg71EMyP0dBJwuqCgjkHwMNGEWEMlKe5wGe1OxEQEqhX1OmTgzeDSOKWtpvOxRx+MYCchxwYttx5
Jq2aHQS2U/AyefF7fWTNz1+uQeRETENhTD7ZEwnVvYjz0A2uk3Q/jQIuzRzLr+Le87aoafl5OflY
Mu2z3MURnN4+5wiD7+HuExMEx/4jCph1ZZjYjEnmVRpD8+rZPN5n6m5mlFb8vdx8w3USnwaKJ4zY
apXkHaZQrdzi2riS1Yu69ZHjxvtF2ByTQCkzQtCvVP7sgOyr/gAoCBazfMC6cQkgn7kBYF46tSkS
Bj1C5OUuDvhGMkv3Q98mZhm0CLzf6K7ETWzagNTsVjNNrogZxqzTIRD8pLdbKwrkVvBeTcXiHlaO
OyxuY8qWha/K2vlAM2y3EKlAsoyU9WCVmVClodJnYG7ytRGWhjXwG4W3aEszxmd1DX84g90Shb50
pyGlJM6+TQRs9TYWjLqLjbGva8rvXcIUOotAEXrDPJv5ZlM7XFy/op6tGCUe9KBUusBgs7WXwQ9L
mKlL24032JCUbpUNLWvFYW9MOicWtLNS4lmPUVF1zHmH/XBQIIxnne3dkLxp0SlF76qhEU+NIZiE
jCBkCxT9mFF3hMRUkm5iUvZuSn713FuJaHTA4e99aKxDgHrQp8xal48+GA+ch2H0VaEJfsAipN/b
jPNG/qq2llLGERLF6TkVielRJGk1R1BSUVTQJPjcTtJzcII8evWljIG8bRP8FDOvesaxG+O1GQQ6
1Y5E/AgjxBaicpSV1i4QAWonwr/UXJApb6watJHmNlvx43nB2wzoDglPoafDn/0jWFyNY7jX297c
Hw9lsh3TqyANDf1XU/B6FudoRNmHKFMBmF87wf3fhpuLfqaHU7EkekSWKKRfNe8MOlkUYO9ZClBA
x59AnDtun3KSZ44+U9xPB2sUeNoBNi95qNXi8RRDi6Ek3H9gajxKFU5qZgtpmMWY3Ag5XZhE2D2P
iC36NZTQcQa72fsg7qOzJQItO0sik0X8zfLaxDll63KUev2S/5esmZtwc3uOMwpSa9HXOcFRZCPr
Va/0q7IZZTXlXkLNsuC1LMoMKuhBwTY0Q9BUpMaDwzzjtIW5Yjcg2ITRPt/bChZEKRyiLdUTTbut
qrMsCih9hJDIyt1TWzmW8k6zGoMJMmCefq3w7bKgt2GYwhM2jg3fc6AJjYIpr7JoXNEPcWHw0rB3
VUAXtLpzEIEKEXDIx4Gd8QU1GhhcWNrrbQ1L8Kacx9/R8qT6ascY9rnqUF7EBgieKceU0lg72pvK
FqXVSzozEPznYs5u4MJPwjMN03oX/49dbly36Lz0zy39Mn+LvgfJdeo/kmWd1jyzRjV8fF92/tKj
w3X15pARc2JLO2omukV6zX3Pvp9SwxobMUS5kdeJrQg18KJZrGHA1kZcu2bWO7B1vrhNyhTHcNAk
eUN0hqQFE2kOQncflXMrMGC8Vzl9L+YUAbVlWNQSW5+HZdoGW+ua4HOO8Ew+5SkrHrSJWTYizjXd
in2oYFv2638ldpOJt+oEG8A0w52W5MLvArBPayMnjBe4MmzL8bePyynVHM5dEeNmzihy1WehkTPi
eIF83w3iZNGAKOTpWa5t7ze4otTKd/hdcaCnrgglV2IZpQMkSbv2dslxWZjDjwfEunUKKekCr/q2
qldoySH4TVkFZUjA5NkGWxwME2Kc7dmuZ4KACefEj77Pkx/3wpNt+pKyqDoy+SmemCMiWUVdc3jp
2QjuN36BzbKvRTVxz4r4C+BQ8EDt5Kp6XELjDqvBEy7jB+ZOH9kRNalojkuQ/rsN/ca5qp1g6r8e
S/exeXXSIm0B6fGNK4yKcKk7pAc8x+OJsKvAHq/4J236d6YjmQ9nqUnWMeHy4rhKNbXv/+QH44Xf
k1y1YKWxPW2U2D9A77FRtF023iw3IgRjX6QFpbPoGEzr8fIJO3Bbft1U6Y0AiWhlzxV8tC8+LNfz
7q7BE6P5rtORFicyMeNuh5aGYOCNnMj7r55rA6grWY2sOzg8i/ntBmcTkHt8S1sBwUF4mfH+PL+b
/DxhSMGa+StL/Y3zt6lvCwoNXqaH0ujoYQQksUinJNlw6sV3+8niKkj332uaxKGzN46t+tlJ1qE1
NILjwDON48iQbfWUM7QLZGHdwwZnAd5vCpaqD2y1TbIPAklVA4vTxiboOgi+KhLUJfswcVg9XbsZ
geh70ly3IknlLd6lW3boFPxqu4RjoC4nPDqVMesGzZqkeD5vNzaFInkBmKE5gFA/cxZd9ASrW5xR
Fulc2CptpgyQXfQcA3ndRTwR39urchijMbvyEsMvQqT8lTALquJXXeSa1Q+Vk1gw/41Y/kA6Xv9k
knSUxLxIfPDpDZ1uH7yTLhlpjPRnRhnjRFh1QtfXzvoR/U6D6J5AOS2MbbcVbojy3JOUS/K4ajH4
chDvMYvIInJjritmPTqln3nojsjPc+WrtOTpPN87iiiWyq5E9REcTmszriKLN0t1QURWWWk9dH4R
lXroAIVeCxttAwa2GK49B592grCYlDvVaO6gJlMUbLYmi/DDnnoWcI5Y+CI6iYNG1MboFhNj8kdy
UA6HoXkXiKMx0G9dYVFO4ONcAeaiGcX8xXRIKntyudbLaL7imfh4VbDapECmuGE5pNnxLUKbB2/U
HN+RfODobTJX0bSQT25hJXwpO26bOdqAYzvAgQbdQyU5RzfEAGeTY7akotG4VmW0hKzUM2K+xqYi
Ss9do/1NU/ApEt9q0xZWQG2jO53ItyaKp/CGKc4g8TxiuiZRkD1Ai98hrO7bWXr24Tz9R2BX3eMW
A5IT0K3fjEDiyoDiLcFebO8oVaoShBO7QIj1egEAxVLXJky+wmp46a8s9XnJoA5PNC/IVujgkBaD
CHLOSnmpGd6d5w6U/zmWIaKBwPqpAuUGXCIkDfw0R0rxfKSg08pc6qY++WNAOfChyiMPmFDoHnMb
y7yqloFYvC8Nrd3W3qhaLbSa+X8O0VBaOyfNrbtJvFz3Hk83IgnNG7RQmthIqfLkU2ynfvPxhed5
oMt+iuZC6CS7uDO9ziTaamROmnT7YKiKfjb5CyaA8i8+nHpR6VZz+FKaac08r2WKyfUax5AS5geR
0d44J2LZkD0HqHPILDndra0gX5JStlCwH9+7SncV3U/GbXuh8pfSMYyUUzYq15Vddh7EKF+e3eLm
X8AxaDMji1iHVM8jaERD+J3qcgChoEFjqD+8Wl5n22UceKDIF9LWFVc+lcJtsWhCSYuLexwRuY5v
2acecGagfXY4iECx2Rnf4o9iXdTs+rL8N/SLMLZiZ9WKBNEfYyXMMlo0vAMqCuLrDlq9+ajANdtD
DCOYOMRYOuT8b+kom9Q6gm89bA4GFjZ5m0IvMCXcMoBuBkwEb99NTRbZkVIpsKLQtkZpmvtGM/as
axou91Zuv9U1A2/YkFLnFsJ1JCaUt4dnAHR8sSBBHrPpqyi2u/qSchdaaROrOGxhwT4nRPjLjeIZ
47prKBPqG4V9S6FFLczjCESBGX5gdg9mNZJUgPBkszKn/OPj3GUSPiq6xNDnyX8VAB5Ftk5SkGCI
Pj7iWxfUNN/l7EVhV1aYIALXrIduXHZ7X69Tip57Fk/ce6WjkrYO88rfDs57w57iyEM2Of76xkpc
Gf/uO87N9MSi6bki4DSLEJLe5xEk92rixXIB4gpk5WnfokCRl/AwvPH5OEpzkvFZa/TaBZreZmUM
fZuPJ9+zQVN8U9/V8rRIgheeWMe6j3ewZriJDVWKJumrbOfy0Vc/PIu22Qj1bxJDJ3ptcU+7UId/
0qfZ1sXigPRdRtINU1mvUfKuuALy++ifgw/h8E5Gue65kTTOIaQ1A6b0PCBKAchzeopbUJb6RJcb
Qd3u280odm3AnsAdPb46rlmg3QyjftXZSi1LFm38xM+8z9o0xlYcJ9twAnoy1mlxtUBjHmbQWiSX
AGiPiqffyBs+UdbjPEE4lwOBJKMjakpNHMFE+vfZdQw8aTDqFd2TzNiPLEurS4BPpv2vK6+8bH+i
FmdM3dT3YNJ9FSCvmhiDx2p0gMXJaYNFx6VJnY9ToswrIX1WGZEFBHkM5/La0QlnwZJ2DyxK7Isl
uBPuQu5jltdKHTuSjRNyxHrNAi8S4ZYCZisxjinLPNGiT6uI3utyuZ+ZYhwDtbUJY3z/aYRMFx1F
pNqxd8XFvNVd/mmBrQebHBmqoGDPfz6on9g/lFqbaEBjsc/sdMB84LTawYKU+4G4hVsCtYhHXice
aj7SjmOIHAf1nVMiieSvFtO89Br36uWEkXBOxEabAcnlnKfS9VI1O8ITH3ovvzXeNqzf0qFqQabf
JOUD2Dn8awlSRh2Gcm2+I0+JRa3JNuJyWEE3mNlHX4AmyoImiWW95ila8nGbkYnKSkKw49t1cLjC
7zZfx0NSY92eeI/Fjf6aNvRQIJxPyyXn0BFAtNqrj2e3yUbIZq1EJYXvoLBKDiQpVun6ZHMXjPNB
OPiyN28alYae52CLYPu+GfhBViL+LNL7Bh0QKwn+ECSRznpjTTRHRAyvE5MLnH9XXsl2oEaxuLmI
jKlwMijD1LGOBYLJcaXniWZIDbhPzi2gXvY4J/BxtHGA8ufpi1aOEc35MlRcHq0NvJ1Oyj/BfYC7
poN5zUtTRrsouQYsc4G2WBu9B2836cPKKfuNtKyNr1eP1leBT6+FLO/L7wn3Ngxc+n9o1sLDU60O
gxQu7LbEtG1AFNXkJ6t44PT+VzhsQfLmwFhhmK7XhLIA30fvxACVgE/8/5lmBKmZ8GKkdujT9sDJ
/XQFGA4nvixh0V4h4M6PqYvv1Gxm+pRLJ/HRUqsNtrhOwlxVv+u3MRGn5PuG8SwAbFdsclCyEfmC
p90LReWJpJ9uJv6KlTwFAmHO19SW2BhE54q4ePvM6rqSUWHB/0bR+QPt0M/sI1FN7idRewuxy9zu
UVmwAX02DvODxNKTFGs2VvvQKNPtowdSZcqNJR5KEQ3dph8GImoHFbb3NU2e6qmHImuT/jQtvqT7
bTxBI5NQ8zYFIan/2CZJnagzhiuP8pZVV4FxrcQ4HGIhH3Pr2TuCDNT0M8HUMEryrBs1ZTnkHZJD
xdBzf1RLT++k8va8Ixiep3AapKHKZjQK95VRA9fwaPaBF0YUsJgzZpZVfuW/AiUssPCZeDpcJ1Ri
YU4ZPC+seoQvpuNZcRLW2vqCn3yymHOZR8cC+YlpKqa4RBcD5qDLqVN99JL2u3ckJUZE63Hl5eL1
ou9f49uIrsXCNU5MZppazTgooWMbpCOLlKg2eKI5fjWUT4mg3lgn4NexiDML92enFlTmrTRv5aCf
jqBjtINQCQrK06BVvyIpLjvH6ZgzRGPLgwi3IDzJOgN2/Yt/+atA0zeDTLUSBwSgy2GHYaCuHrI+
m7trs7ZIbWcuVGWGCOpiLMFenoWgJgwXHvoZpbc6Hv3bWNH8uQtCXMzf5Yql4p56qyAkDBkJmcz0
ohfHufaNymR+7+I7aQtAJB0D8ieeHd2DRzD19IClzkXKvcD7EMYckDiYelkiwXk/yRMyjFxYhbut
HfWdENayqg+VazDl5FWM+ldcxjOar9gxjJj6f+B5xZc+KhRHsB/HgZkGmjpa/yWkPOStKAci944f
DMy1fwaDeRvJ7cri3KaL/UJ1+FexLhshKNqSb5pP52WlUUs2rmUjCfKDZnZLjBc475h3pctdyplN
RMRQkqGR3qySCXldDBFZwRd4FBqUitT7uTLKETc8wDVQqiEvMkPnLmWrtW8eLfWNqswbH7jlPdIS
b/ohGCDecczfJMGwLbhP+5LFHzNaOJ/ng31eXMnYWmi4C8BjMkoRT9HUlq0ZH5JFHAkk35kBLYmP
IIvwqJqNmyueaFG+ezfmHP9u98n01w+UjEXdE+CW6Lpcrip3eQ9Mj5WIx2oI6vffxqDjRjb4r4Dh
VD0OxVXwIERY+ExcMGQ6zLqVs4tB9O2cZtXWrVbGDRE3Kus7WJ13PXyeYRf3q4yvO7cnp5ZqAukW
15wiGI5sa78wOC6yKfQvYWZyiywGg4P9ORmSdGHEA8X8XicwosfCin0y97mF/VriJjCZRz/R+2+P
aE/yrJmmbMPlHG5ERbnDc6x4oAqdTemMYQPRWIe6/kcmiwcsrE/D32Ul/Ib5yxiEFqXdM59fMzIE
DFdevz9A76W7SsVpAEOBAvv57jQ5+tIvC/G186XhjvT8BYX9VKc+vWjFkyJyQlT+9ZcGAj33RSp9
FtUBkFQ1bTHOhkVluWFhf7nGWRNIksVBzR4G2bgYLwHxOfrn1ai9+0cPnJOd+DW4n4tRz74Fw+Wq
I8cnTO3Aq4jR0MV65UTB9wpQ2rHHK2/KWj81fsFkBYY3YE50lzpQ9C7kdawGixEN+T13ghLHdzyg
2S+muCeXBPKSFqHifAPHm5nKk26lfcl/9sAs7OVrqZiWQ8KHufkcQ/W8DKMCV1dHnFBfP1qeAMeD
VFjPX3JtPkQaM0gmjTFs6gAJjv/SMYqdZEaG+ZqEc/xoB3lcKWFDbb62+e/skYbIHVCy04w4UPqM
NUoX3QjIrDRtg8jJRNtDGAec4KWHo/imYyEU+yw626kaXIzeSPqh03Ot/C7KtFMrppngaHFq3uwt
RSeSc+uKNC6thSSgRwwBJqE4neULTGSw2WssFRXweR63ZjvFYhTr9WCuKVe+59ag9hFm0+ngFiN6
1/QHAal7hJ4zL6TikfWOXPSjv8otJ267bRmSeDnLoEYNWW/BaV1bCLUaJniZJmM968PGdOZpsJRQ
x86TW6iXUhO9vqCEKLUlp3roTg7r94GkRKENablDQXNIqW/APfmBaXxtxDxNF3/XZ7sRfq/LZiBv
a55LtY232PM9sXuyS9EcV/PSl8i7+oMveWx7oPPMmp+kOia4KU/xwwYCRjgqJt0LBVEVELqMba7T
pKHA6yh3Yi3GGU5qvJeD17SlG+dt+1AGY28eS3vMmIB+PgOZ+kVcn1usMs65t3ym2BcCCPwV/j1L
3jR0OCpaO7QSs/iBuPrzl2irpJod2fGLnNLyBQa3pmKYKj9kDLf3ciFb+kSvOd1Fas0xQYIaf2ss
bML79cjskCyT1jcnmm9Bg6V3Sr+Gu8yvF5adiXR/pulGlcyeWa4fj5mjh4hiV+ybvmgkuFdgio8N
ZcT3AlGhRVyxDQgFD2HEnNXyWVghMzVY2rQqgb9hMH8ZXRLzgmHTecc4SdRslgAsLK9anzNtd+mS
rJdfGjM6244o8J4iRWs4HBZKJZkSLkX/kLfoG3S0uIOMMutSkpDYL+sT7IM8R9H2uJ6286P18Z3P
K7ZkGI4t1swrE5nQJhhZwIQyNqrxqdz7mEAY+bxSsk7rGexQYNoieqf43VBpCVhTgFPJWUlpVCCC
DG4X+JHnLSTQnHP0gJnauNl7pwjvPHKsYPMoZksFdcibUPfixk7cjUlQwmg8xTw/b28lb3lqJ1jE
+aBgja88E6xYodUmGnIHW0pdlv3keXZbC2sVUG4Az/AS0DnMt6srcv6KMvtFkaXpt9CRB6vY2PUe
1OZuYG3/x4oxw8eCbmROMLeNvNR37yIpWaC6eK9dNYElDhmNshADtw5xL84gvgAfAkDzb2si1fd1
X+pdNIx+9kqd3/ZzmaibGIAbB6U5uEFya/0f8wCHIledMcblzBMlk0tcq8UNSL+maVJ/FzdJwhqM
XP8c7+ULNkMwtAF1pfJ/tt0nudZ2o6g+qAuYab4LCBFmUFx0l/OETxqmOEqIqlmiANuEW4hn4efX
bXIJsR5xNILnG9j57HULG2sbxZ8fLAFwL6BuenP+KPiwxL0GdK8XIgCCt9GpYNOkHrFD3nN89pUS
wBdFZkdTJ5RwdfHHicbHeMvBbINTeiUCg5NE7Ta/71t7796HK7npdnCsa0WbyhAg9J92ZzMVJ77w
JrMt5fOHEZXC2ugg77wQc2Rm06CEdzebRxIITtDsXPQy89SK9go0sNt2NocL8myC9kACwRcgl1vg
D+iUkUo4dDhM3eUyZws8nHx335nL6DoekhUZpduRjRz9FSBu3L7zIQ4AeVwqsO3kuBh4nzBH5WZ2
uF/dCU3fKRGunQPl8FeJttofe4A9wHwf2kj7DpIrMoL3Hj/IZxwiQ0Rzlx+lYSY2MSZGcJOIlcBq
LeLqt2I4OcqtoPwHr5qCcNVIj/ayVAragw1QV3y7oX6JBHAyxcByz3rmMuoIOzt5nZFJKLCTcMvv
OAkMOE3rbifIyenEbSEVbupLK4gF5CcggMRh0r7f+SCJJR8darrKhP9mGnwaWHLetZKVhKNUQKfN
KSmih2QZkoykt3qUb+UCe3epmYAmYDBEGQ13+Ge2YeeurpNvxb3yWif/pr6icYx9ISvZg563Hbqd
xDivx+P6eb5nf7SbhSBAzwVEVvJ+WuzrtzLYIfJYMobb4kuc3IHTmgHNi2WVZ78DHTT/l57b5cm8
aZDeSVEv/CtIaW7EFvJzZmJaeMs3mWjbPDRCVBPzwIJzb+P3X9IzkXGtxxz7B1PtE1AKuDqWLxSd
+rp3Gh0j1H8YFWuIVMTwnOoVZaEvrEJIVOb97h7XeZKAE/0pz79JaMTFZ9bQp1pt/goBRFCxkRpC
Hq7vJRvCTUEOp848d5Nke5YU0X6nj1cwn+Ut7FERcoLtiXaguds2oZBUUPwmuyQLVMn18zv7DuSc
PN/2lBJonxWU6Mr5Wermpc1W91os0nvCs9OIh+BcK0PADxL/wyeAx1jnzW6AvNpv+bLQkZN3yoKG
kHaBV/cTCOHExj2Z4a7nagalPqXXRvA17X+gt0PAalmpIKnXUNTLL4dUO5ViaZfqitfUZwVEw+xX
ho9Yf3mNmZSS5ZLcSX/Ar/ffT+F5hrhQzqBjmY7X8gWQVPdbcLDFa6Qn57WW0ccrlIUPG+4ntrU0
2cX2O0kxK89zUo8Chm25JC+xmWaDhxHyWqWizVjH+oxeSOa9BJz2M8T7iK8D1Z7rvBQ/vOCKGalU
IIZdwWvsF2T7Uwvx+4j2qjWAH6bSZAOWMb/jJRjfLi8vQmfdkfau3moYC+zU+7bleQ1LBEmhHs+i
n0iKPsVvApJze9YBmueX7CPRHDBdn3mrpftdHUfawAafiLll45i/ubgY9ch9xmO/8oyp0lG1PSv6
qioVpeJFrs/it8gIHau8xANDbFAQGI/6cZeQMwBegGpN8RyHNnQgbHiUb+nsJWWtM4Ra4yedp7k7
w57puTJNamkn2DZdz2HXGP6XpFgvpZVcARk0JTciFA91+A6ebqaX6KZfFUVeNt/UUMauxBzGGpcY
niOysED7oDngs6Lw2lKii/SdOBviKK6AY2oUL3j/PuXCPE3wrDkdnWtZk3dm0I1/TMF9Nbz0EzTd
inrVvRPFkJiqMI/aO+Tlb5wgZaDMxaPn3Z4HB8o56NvxSF3M24DkWlfMXXmCMTdrtlNC2k9UWKu/
nSOI30E9S08NPhE6Thfzv2d3nkIzw1513O11w0atE/9bNf6pzTiWq9as7W85aKDJxSOZ1kLYyca/
eVXgESl/r9VUxXHcSnHad91r/xQFwM89Wa9lctprlWk+8VO0bw/MP1Npy5aQb3CYAniy01vd6QJ0
pt6ZUqLr4HUdqBaA8OQRBgUb7csWoIcCbRsrCecUeRW4YNsgY8hJ8EviaAIuZaXtMf+haxdC2D6p
2LQZ6XT5cxCxfj0FJvvaikzU8BGbjNg39HKXpzG2jj3RapinW/wNPEu32J8rJUCQiPjK7Y3wXWpZ
P5U7Q95WEDpbOlzpbDltDz+G+n5iIjFXHVMzSo4R42oWLSsxjzbRYPeuEWE274uVqqm1cTCu2JG7
hVjuXAW3qtuxBSmEsDN3Baaz0jZCxP1J2Ufm+ue514NL5ZaJbSoP/xWefBcJjPKiMLO9hDBQxHdc
7VJ0LPBSFmroQqe1bfQAsWOz11zycr8Qo+Q8CYSmPcnNmXXj/8FDvh4hFF6OpUx8cvwB69ESLdR2
U0VJsdsC+97ZLPMawD/R2PA4t/Jhx9XZSwOY5+LxMMvhiKWgXgzjsq10Wp04Ik2pekAX+sW/hWmp
mI04mHFkFLJBV79kYd4BBpLskZoORR5oOFNd4tbcrJRy5AV0l7kMuiJIZFehIRblIbmPyntEWjuv
HfcxXbChVNeE8O0uZ4u16RILBsfyC/UOVK/Tl6M1EaQ4A9fNLYqkWJ6ulBsOkG+hO5R/0NZI61gU
KEp/iHIR6cCb8EQWhYtKz+TXWsiLGC+z+pHOQ7aIPanZeNHz3XkG5K2uaCpZwJtCcfEuhjRXXXTu
Cq4GTMKUy1Lz7xKOT/+RKrqCTQh7KWyWAEGBPBPFXH4ID55UNlFkEKLLf++42ZUdQZPWiWFO8D1n
kR7fZDjfwZgiuGdyw+gbJaBohwfY1Lte94xPXH5ldUyKjquGTqX6r6q+dmBBs25psYoIWdxaTzHV
BMFW0bJjFQaV4r/3Oj1dUghDmY1SqVdeOWYOVHMgU89yNz5ovmNaYSUCdb8RyDUTHY4360FhDMGQ
FJ9Ruda0RRoogCzA1P9n5I5NzgLeskt1g7to4veb0OePC7V+PJ6QC9GkLkECg0x4Nd2avztLyv74
EfJf0DCmyBCUKMgle5ec4KnFmi7LGeD+FXLmU7lYD6MdI/UpACUo+IH1Bd6FJ0mHhTSyh9thJdbu
Fx5yUfAMXLp4h/Hzr9aJT9J9vXBuVQkGmSRRXTqZQKJw7yPz4yujMpURz+2oq0UKHPPflMKvcXhx
KJyp8QwXnvnWG3np+7u/V5T00iZiRdqXzynkahznGcte9rFNjdIkV26lNeeP3B8eiYl6bNksCWjo
ucdeOukmi2yQ70wEnZ/yEJ8ahbWL6epJWwyOub9g62ek6kjftVs2Aw7y95ZCaZ5XdopWqyrMH5VF
foq7iheMG34Avu/1RtdxuiWoDym1C5I8jKEDnUVwD0Q+jWNEeg5O/bNtjL7jqPiAoAES0l+giRu4
f1KKuSw4N+6oqM8JAnJYhCxO3gFu+Gyw7Ohzm+V9FOJPbNJLPEyNt2YsHeU8/iUORGjaVAWQ/zH8
HYxqh4K3KyYo5IqYIAiTHrSy8/r0kxd908PZJZ01nj2vPAyBiCJTQ0dWs12t9bVHuXljHlrjmPfJ
ALrffb+dxqE+SdADd5pyFqogdImTC3ICzxOe9/OH7ssMlKKjm7OWz7nM7u1bvoXyVP7hRzxnrurX
ySqhqpJJQNoj+tmMv9nFZWg4TjgF52zVUpNgUrnJ2f8bxy351V0nQaiE0dox93KyYaC4v/hIdJmo
YK7pH6Ek5jcxob6uBp33Dv2qWfChPDbMMarh1tSG+R9ctcjtZLy+x0icQwxOHKaR5Ow5FGCpZegG
/6oNZ2SiBRgKGL0Is46WiI7an4WKHE5KiFO44EaIllptLVvM+g0M7RbOneHYebDahLOBcPB5r8kp
GXccer5+8bZAja6wvA1mq8gY9HG6kxSJJvm1qbfNytCmaMKPiZj4to2NpHfy9jXaI1pJS9jbT+5P
b0M+EDi0UNoMc6N+XduFEHKS0aS+IEBVtfqdiC4VIX9RQ1SRcYRIrT69SaXrK/jSIl9n8UvZVUxb
gifUX5uTf4OqgGFe64dn8X9nbQDsLny5MTZbBDyKM+gOG2HColr9EhABvKRjL2AlPMxKbVgMqC3l
a/XtCtdLwK4n8ltOATNfCOxZxdF8g+4je2dppPzIOMtDSzzqVJE+OVdoT4OTQmaxkhYjJ75WVykS
peRAi4qPbT2TGvW3BbQiOsHTcM2JL34SQzQ3Cc9lZYV321bOQBWcNWyfoGYtpzQOYBetOJWPE8G/
F1idy7fGsGZ9Cw+aLsIElSYPGx9gbs/ORt6gadzcFnDnFRWUt1AiycZ8+QsBg/5AsdxxFVuabyfi
IwjulMIMDPqPyifjKGy78sj4w+8fffOkwspTuij8/628shazBntQSBNu1YTyCQQLNN+hjTGnyuEC
0ZcrvG6oqQRELqPsXQnv/IH2GSFlBAAMLspHw3MRnRetf9jPxIdeMTsYLWtalqcioUAukiO7Ja0W
/S9nnpHDCyZDQ3gIGZNRVjwJ/HC742bprChLpT0qRSxLXaBP006ZImaIOPOe4ml+OZ2X5NhVH9Jy
K4GzPCIAehOUiXugPcukxshlRgOLY6h00C+J9Sg+DMUU4fc38T1A8zMpib0JH8Whs9ktTF74za/3
MwmIgUU6VET5lY1uqIvpC6pCJ24+1ufWZAgWnSAsG6SwhwKYX54aDOPWbp9QtK9au66A9MQwB3Wr
iudoBi54i9BxnuAFSd2AhgGaqyCpDCbXZ2SmX4AotTOg/BuIi3S7GLEs4w4CCpTii+rpyzJkD2zY
q3fSp9SodwwNXMUBEV1xsXzEL1Db7obx71SE4TkeHEPZXwznUyQ2KoixSmLhQaYDjpDrin36Sqm4
yGSjdA9M/yAjqwrCTiNMsDJxV+vWYYWnlSCyXYomtT0bkvTInQ1ffuyjj9aa1KpHdnPOzUH3fSF4
nSx+nJ+nspxgCkRpxBFcZiOS0aXIjMthkpj8oBv26yPSGo9Mv8U/15suwrAPm2MzB6Anx5qm+UQL
z3JAgbyokPd9zc+3EaGR/I1AADiOKY88e7x9k5o+GM1Ylo/AxPRC2Vkcas5gj+oebD5CWjdJZKUV
5Q35sizffX15p3dC0vsZ+UCfA9WNZGZGY2YqhWXius03qRBMoIJ/9iZ7PS9OIfXAmR728yvjNtC+
mLwnVML2h1zyavZOKcuXMBPvTk8VRkypjRbA+zhGOLwZM7ozUn5DHAQPgxdFHODXyFaCLSowNL6K
MvUJKvFmfDJZ5gr/qZnDMDun9mWmrTbTiEDvP/YjIJuE5denoqg84H3cT9y6vkPRcYiRD6vLngcb
Mlv+vQmM5y2bV0NZ4Le32I2Gn9UHiwLzYkPkweSVE0zMjm/nZgkfoK1hCnarXYjJi4TOEaza5v7O
r2QygdUGSo5jxxiZsa6kcNZGU1MZnqHIQVh4VteCgY6SuF/0OtoJW6kQvpk2eabdfb8NekgsyLjM
DGwRVTOzzPR8MKjeZ8nco+pkFeQpHJj9MMUPYM4zdCRJuy6dIKbphyGKOmDpHnx+FQoxAI1QU+Od
Hw0tU7Kg6hsY0kWZErD6GaNjZYgZpYT5HPkeCPIlfDirnGm5AbZLdMOyObrXbA+BuG+2aFAoY0SW
/eikwq5x46PPgAJtEjvoNY/3Uxpz+L6EhkIFA0VwUK0CAPymUYUGtYDVManqZUG1vtdj+xc+N/07
cEMbXDS4pHTgm9nWRuRfMK98Cep6uE9tlRI3yilg/3wnrs+767w0kgkR6a+ZcYTvfSjV/IbgXKYM
1c/dL67CxsGECxovilG1rOAAdTnc00xz/iQzd9mSNgtELp5SBkY4m4pCZ8Vb81HhtPBP3yxmh26V
HuhMalJsVKyhx38G6BG9HKOw00odf25BoABHU4/WWQqzIssD1N89i3z4NbjJAJiJZraozKrKf/88
ffh2+sX13jsE4jib1acgx4Tz9nqntzipb9a0l1GzIugN5rhF3wFQsdmmJAXngy4vXGQS9jWmZhpr
+hRzL7/aVzDbHk1VH2rj40mHP35kGbDwP5hRWqSLcnnz6xGSs/w12Nor2xqEhqcwQdHH6VFs2/S1
e3Eh1Kka+8YUJeCZZ/aLkpbgNgYm+vH+2NLOC9mlsfCHBQ6drL9tYmXDsGwNuDrX3M0d1Dtib6Mk
IWUBUTlwCHZE/kaDrMvczueev6gvNNcnK5OZ7zSaZwMb4LhWwMQSYRwSd3WosO1KMpsam61GeVX5
++rOQt03b4gc9GuszHaXMLpKyZjuQ+bpztBPwmK97LsYI+H+LSiIVY6LrtwJnrOiLwVe4850JJpT
6pJ/K1y/WI/qq8ph1ZusY6x9Kqsz9hgJ7rnsApgSxhfTPOhbrh+bep1eqZ+i3TwxJgcGA0BtJfhm
XnX8XdlueDp8uyaVMsDB9qie5U8ADjcFyWLHQjFN2h1SrmiWpH5k62NnO2tuQRlvO0s40hJwjeCy
PveqUm/g6GVAoRhhhrqbubFDzksgMgOcHmm3qefD+1saH3MvIEM80oL3dK4Hvg9gvmMU6RBxNQPH
YUI2P88DYopCdFaPCENPh8w9UIRH/m+awdYTUSnXJmpiQsfKs+BQ83lMX2osqudK2qJj7u8fYs45
z+Uu1adXk1s1Sl25w7yuRwUqdm8GROjvuIBkJR2zbCd5gH4i/QdNqroygs7gx+/LYXMCMOzn7sqx
u1nJLSQONc89m/IQBMeSd2+em6CWikaDJ2Ps2BFuRFd7rlUNJSeER2+8LYkFkoYwzvbity+HCenh
vhxpntrtxFmzpajWjUAVZMBKOuQfoAfpJ9QK9mYuQtu3yTF6KhnfDnbblBqD/pMMwM6nXRtZ6V2Z
Gzg87zDSckYBGUcGdUN9YYdmLEqR0T6tyGXAOf2blbXUczgwkeRB+sHUmBQGiVGMUqBaMgJ/szDh
bNXqua7xyJR8A8YPbh+SB7k0y05BgtF5QYdRxpTeczYe+ZNfsYQG+YkOLd1KUJPiwYGNWdogteUc
5HSKJIDr4IOQz4DeA6oqoeCdDQpYRhI+qsJHwfmYuD3aPSshfi2tJT5TdaJnfXLODgD8u9IKIYiP
AKNBWcy4QF9NXu2l2E+f6v/yrubwDu+r2+0Lww7sUXfnGqeWHmcgne+fC5Y4mX0k4qjNUV7WFp+L
p/vVR62IfotGhkrgTtTTwW5C56jnuZxouDUUn4YFGF3zchTd1/9aIVtmwXEyD9R8hCAvlKYdYOKj
e7++8ed/k78naPMODQaYQn96ZjgsCxygXNFqiIaHu5UG+ZJ7Yj5z495mlkyDTrY0Qkc18oXNdCK9
cCUpGJsSVZJEiMtRTck9iGGMYpkLWB7exqL2lMuv35d6BAvM69TbZE9jJxDeBa3j0B0IDW+/Y/+t
twGYq02Sq+x4J3SFsGtqHNE6LuDePBkfSlX/R4hJcbaO/AfgQuAg6pTqelquCilLLnNEak1EG2Ep
EENCiUAZ4OD7/nFzgv0FF7G0DwGlEyeEsP5chB6W34KHwohzqdTkmmGdEANA5EhMRkro797bYG5Y
1KnexJc/UkiGNwnhrUFnR0IN5wEO0hCZmpkkmTQ+ojdKXPYorl9QYjASJORg5vBZJuVZ09XkajTm
CGciz2/9bUT1R0WrDxq1rES/Zc0dhQPXbuyvBUSktKV5653wiphs17Q09JrdC2IyF6Eiu1FK7yHC
FJd5ks90aBNMNDW/dw5gy47Uy0KLxyQVKRs4XQO+cqa8dJvMnX9ogOquGqumwy9+ZrSOsilw6D40
nyh8PwDjcWOGj8FTvmWPKk3i5sQL3ZY5GRKpFjuQwz/77/oF1JfdflZSI6muy5+JU1CnpMZsGy/P
D/9u8wPieSpSxsigJCSQLevlj8e3yHx4oBI5aQ44GbwBlaZL/n5a5bWyyv6YA5tp7LGkZqXfKpFC
/sJYs14MRgeLK91HLPilk4Jv+gmGOMxBN14v2xAUwDdLOZN/SYVuPVbw2XxL5GtC98WW0gTTZS6F
umEYb3RV5GoilRbgqbDtCWOS0p2gc+ijf+g07hOKRBEKqqbYm8wW5mF98RDt6jOGbCu9cWsPqIS5
XITP3BlL+2KpD9mP0BbKRnIEa6LIha/7MWbAuUvvvn8I++E1C6SANG0HSn0M8oELPYUfmHyyF6LU
C01Dc10g9+B1ebiN5zyPPIZV3V2YVl/Yxyo2HwtUS6FWoNKaEavAauemQFftc8JycUe4SWpqrn/6
RoAwNeN6VEywKHvE14RlX0blpOjNqSYtK8D1dFyspQE8fQj/DGyCKL56e9NyiiBj+75boPua5LZw
13mdRarIYbAN1Y08HFWrAg7CVurTILge/HkHOCWbrkYLCWtui2C9UQz7mV2hwmYwGKJO+Fz9xgQj
AifPJVildkUUsgKpDI2rtlCpQeEY5n47DYlK/iRzNP6DaseLcdyiJaliKiG3CXp5Cm0Pib6diLfY
unwSHxruk6y164gxIn718ROz5s++ufmK96fg6Nl5pcWS0+YvO5NrZ6QpdFlQDckPc+6hQNiIJD9W
iHuTnL5TJDHkuibHnnRVtg+ScqaiB6ZuQoPd/fKV/k03KIsj0mDl1/BSGlKfAY4Ski+HU2HlUTeJ
qt1MqgF8Q2V/TZbggnHl6L3ybknDkeX8vBJtLe+lELYuGd+yUIuhFNUiQ14aLJMFh7bi1EDgZq2B
VEwCewgUi7oGhEjThNvwDuEpjaEfp/lw2cESrpHtg87W+B8Na04Ejj21LcKOgldK2VPkzY6/hTcI
6h3CzM5I3IyJzhQQ4R+lK4CZ9X7G0kdnOjxj8ANAfzY1gB3WXIuOIXKiTgwro//GCd4eayw6ln8C
xjOiyrfwUsRN0m2H1s0ZWUZLO5MhfaafFWkfASKFbEdMJhxO8oAgR0IfiZlRYrvTasHGE5h723XP
QFDXKhHpRhW4w3y0Cdwrti1TezuWcTCx2wu0dKWAk0cR2gTm969W3emxgar8IsLR3w4AOuFCnLfD
Oj2VpLCz4Y2P3MldPp9F9Sn1n9jBy7mrrwnV5fR0TpOa/iM8ozctv/Qrmqc30h3zbxEeRynn4S0I
NbdR2sb6CGGKIgR9PGYMKg6tm1Trxp+LrjjJrIoIOCKblmvZBprlU3Vc5wDMHdxqGKoViWAkbuyk
V7/BATkAnSpMlWPFyi46fLy3PivqTNY3n6OTRPQ2TKxY9QzVUPyL/GJS9ut8t+09RX9h1ngWyFFr
kNV5BeqHJO5v47xHHUIY4yV7lOOOMxbRlh2zXCFrfDqoXqe5zCzgU8jU/POIQk5hxSF9kIsP082g
R04bVMFxd8mcJ01EqCdngbFJYtWIR8+2c/pSS1oGZ09u4nhu2xXFezM552qFJCZhBCj7llIsS0PX
2FSeMZtHuqivhx9kUYw5T6NFYoUnxkNj429JPr0PmOwdL6dGcs2NxieqyOFK6pEWhEZMB6Ubee0v
GlR8Le6jsRPsIV60BSgio3Pry8moaWY79KoePq8yTY4MA1LDbDO0zarE2FPn+IW310mCnuugYMZ7
pU8u6D7eUgebZEWDwGk1vL7YHBewgyDHCwtIkiLf0URo87gqJPcrkDvXo40z6zHrDb9OPvJ8qREL
IQCa4q55q25mbPHEepubKWQr8bMojD6p3mkW30H3kiJocKW6w6TR1uApG4O4ga8EX2MtxUG6UGqg
m1d4cNEOqxMafhr942OfvCq8TCkgjezt4yyjabhjnq9vKKFbJSUSbVWllCTyctHZJ5FQxrOhf//l
mzDfhwUmOpEgit+kZUNZ/Ia9IYRS46sec7Hu2ol+5/AVe+snQHMgN3Q+t7Xw80S/x3a7oHSzcPnQ
lvSbUYMVLQ/13SGiLgfzkRfyDnU29sGKmhYs11ZGeMxMV+KopFubT5tXd25sFKu/TZXaFmO1RBqE
iIcZ1TuJrfmekT9qEm7s529lqTaQyEdcPAkNWAoTVlFlXkw4sVniD2s+VZVV2B4xoqxYCMyxuDZt
O8o76Yufbdv0qwvLg36G4/nnBEWRVTp8eDy/eTvkcjELpxO0eTiO4lnXl34nJkqv520v3qVGSqzn
JDSROJVM/bfEP7CKCBHFKwr7E+CpAGrGmOrnCoy6fqQd4CmaXe3qt5zz4L1gf+lCcVgMaECglm5W
MB1gSvX9DxE8KorY/tmHjfgD3ReIFFNNPYw3WS15o4ba2K0cB8Ffsl3gy+52uNNu09K+LBJGfLMc
TcRIShHX2AeZ9Rp/HrwbpSwznB6J9gu0bIYx5x+2PHuGLFSeJ068WvrrKTWn4w44DJ5yBO/GJZLl
rPBFg/IXptcdigCK2mS2+9ffwFvy1H/uonvbd5ksUPMr+4OkhpwPm4LJryn0MwVKuV4oDJ5XzWf5
gEy/MHe05Lh5gWzEGGkYg9SRbDnrI9LYBgt4yGW0GAsTNNEa6igeT0bF834LPQ4yN+RG/c91W2K9
5NLXl1sQQ0MKKjsxG2Yf/pisU7ySWfZIBsZIYV42DYoZ+8KhcZvTzDZxz9Z5rcTp0fGcug8R7IlL
mBUnh4qxRxXp07DCposWJFnS5kUFV8ghDaLikAYnpI1cKNCK/p32ceI9x0l7aKZH3n+AN/oPQfTk
Pv1Oj01BByfN+/FBK8B/+DYHGgF3zEi0LvtG0CWkXc4CPqoAOO6HD1BZ4WXWeyZ15+izcx/HSkKZ
S7VWanPbSbxkt76/cP4vG0ehubbqy0m4vRIYvZ0EJ24TuYK3grBAyrF9C1wTnPVkisHS19dwLdMi
iAUaIm+me7K3lgslO2vAwPp4VNSY+TWhtp7QRy8FnvYmoecqwQ4pKKAVm0qD2a/m3CSixI96EKn0
6V9tc/vJ6FsdALRgX+yaD5flZoPMOB5KtbXaK54ELRM9zXSE3HKLyCcxrn7G9j+HPqCBIvHa6pIu
4+4WPR/J0JcpHOWXST9jxoDAG12GppvqfDR0UVfsotvrrAfnm32EJvmpRspWDKApQQR8BmtquLRE
paATJ7UpuZYbrbkLzLnw3hcPqztSqJlqY9F87SvcMHdc8a6hkAAczEM35P24iiqYh9cYjZ4RApXx
9Rvpjco53Doi+muuwAW1dhWBxNcK5LY5SxejbRxcbhMGKWH+URf/xsJG4UTnDCDhK3qbeOeCrm1R
0kNq18akzqZZz4T+lxmKhFY9kZT81AHfWDBSjNj2s7NPUShTaLK+/2yCGycPfW+m1Z/EUSVaLYLV
aQwGGbz6HzYfo32ZVco5/zmjbLoMGV9ph3MMNcz0jnVuL69lk+gjtlrTtd3N2AEFrPpjKHaPdlTD
fFHiiZWujtwOiMfsOei/BvTUokyKGuj5A6em9BNn6D/MB62tr16WP7dhKSR3Yit6DZ+g379i2OPs
+U6tBRRcra2tQze68zYpQxVIn4F8X0GpayXey7/P9oFeQNzxG8xq3gqNPb+OJmotIRK8ihvOjryE
YK+VduW/qSFkjlQHtWvsZwJKJsA7BS0O15Rlu2p1IAxEH935IMEfGXwB9cvTuZd/Iwg4ylNL35zT
vbRKIF+r5UmPSGtfVuh1HesZ5VnAjE4etSgD9Pb7LQXxjzKGznHVw2v0mJeiT1F3MJAPksN4rRDL
kRqeuCFNK4iANLdtlGX9EqVMK5dH+GbrP7xvvSnsg44guRbtd0w2j9y82VwHhPPk7fb4LtgfL7hH
xrT+3grwPpk7+DgjJXKJNKoEnS7axllHQDB286FmRAieWO9+Vxly9zmtzeue/KKWMaK6UQCX8jDp
3Yv6KDal+pVC33DfZKlbnp9tXa7SxLgVpZu1sdHGJhSbx+Od4hdLZIglpDXvgdD8yfe+XnesHyIN
MEUDI7AXfgHFCS2Igr5rVkvN5asGH5k4qo7P2Cw+XvgURM2t2C2laHbj+cPuGYtXz39AFKnR7CJ+
O/7rUID71oJkc2N4dV5HohDX1IFcoVFeA0Awq2l2q8OcsvCmQj0e7DdSQd0kbZ/0v5dTu+tcxuai
zL+pK888Q/0jsXUK0QuC5fiEhzyNmtTzdX0ws80I1pwKwO0H4At/uamUXjUgdhdSd5morzYTRTLB
rFL4eDjCDVBMONW+odIIDrW5Dgc2+POpXaGjiJ5hShk4ysu2Icxb6/BzrTWMWewV+XHGkbC+GLMH
Xq5pf6Zt73GKpGh70lpGGl+e9auyM/5xrZNC0bP8R1Bnr78pBelQi+F2++A2+lh5Syj9GDkXez50
nbDOjhTLG4K+NvNVUZVw45CdwblIz8HKdhfXFm2Vh1TZ+m9t9X/MhDzM6jW5hv+9nZ8Ln1lr8GlF
f9cmVQVMli//Ie+QyRD/ZD/AvJMOpdATVfBJjEU9jiSoqPlI8DhNij8B3ugAaR1sdgV55JYoHqYu
RzvrPfN7hKHUKwo+BilOB8v8Zv4hsVb5OYI20Pp0PzqgHzQuaNvS83mGK4VmnFRES6VviUtgGUlk
K7S+occIAuriqx00NFhXozDhatTJ3drPz5aFBpkaN7nWR4WIsW231JLH7793/w/pSjugyOqBV5yT
O0WpE516RhiCtmhqvODh79zMITD1x0zQs1d0TQSnTUe5ylkzp2lmW8RgWzRMnuuNwso5J2t6lg5C
KACVhuKgnjwFBet/zD4o0bZ9xNa7gWhCbqysmb3NMO9YimQzBfM/zNvp+mhH+piN8+bkaSOTefrY
y2zi2eWvTV0S6EIfeYVg8zXmoHz0AZ97t5f0aHZQm5F4sHhXOHn2WOmWAw2wqMjjcLXaHiaxchP+
oLHu354nXjNeYYQeIahjE1YKrjLAlUUCkWuPV27g+Jy5FRG8vSwxzuOQ3t+VBGwcFka6KxwUiOOl
ldT9sI28ys4SEZkODOHiLKLAZrFsTGo67d52YIUDJ9JzDcVd6Uvux9HY8j78Y+XveedfekAKV8wc
QwwPVK0lVL/U6PseCL26VJSxSdrV/qXE5suNHJSe+UtDZA7MLzi5qfpVAb4SLc10JBt+Jj5Mekv0
mIkoU55BwoXdB6rytjjA4tIvvZlmIQM3dzW/aUEuu1s4gaHkN76aPwn1QYx8ghuHkG7Q+fegffhW
z2UYyeVBrapKvW+Kft4HHDwh4knInlVcegro78ELRGLxx2ftOv3QBJLfBPX7Htvb4W7uP8pI6cf/
id7EYOt6jzef8oJXxohOd6RPM3aYxg2OwdLk5OyL4AlyoLwiNT3gBRZ4+0r8e15U39Ly7htHEyje
egtDN9YBLuZlzgZVh21i8QDL1EHFnEN5fMxyiD8fkg8j73mFjTr2ThSQ2rJl5SkgtLusXjOuR/Mk
lT+x7qV2B/Vlx0STp5SEyadO+pEcUpumWzsQ71+UfyaUCx/AUMAyRH4wkO+FmRIThGi/2JQ2mC5Q
NiXN3ab81pIg7PARUnJrCTr14RIhQ8C9U+hHTAwTUPb7s+S7v2RtHCAL8SlTr3kC1h8c7oiJ5+I+
1j6N1iCphZllCp0PrlQxXD7pvWjHZj7Wz0uM1xKVkwWVNDD17suwEZGSbDUm2E4kp3T2HMPFe6xE
/6s09GT8yorWEVfh0xRSHFrBeGHoy9GHMmy6umqRoY3+5IpbNwVwvg//1ileBY0zCr5V1/5HpXKu
mGgxuKyAzuv8Rx1yEDu8wy/LhSIJG9LyGw0wKHRBn9Kdu6nBmmbS+wV01GcKkGnSWoKGlbdo7g4R
k+KUZJdetIz9/uQmk9B2CWAeHLQ8C07cI/UB4vb6XE3YbY69H0u/jH3l8VEOqSdHnwhXb00q3nAc
2W9NhhQ/GfpQOQWpfxneFfxL6wMPs6yzqEJYaFFh1zL88491e96bCMMnCMs/ot0cFB6OGOnPusOb
5Bd483kPLuuEL/vJQhQ4Ep4jM35L7fyMFX0WF+hWRqyoh62d29ltzWURd+3zJoznNWl6mVqrOUk+
dTHg8L9PltjycB+ETnvsvYLg4S9WQTt2UrZaCayguMuClk02b/PR1GS3tQMMul2EUYz3vaPRH8A7
XoxkPnt+YHZ7v33vJ+nRifc1JijX1wjPwy3mFKNH86jg5K9nUmbQE3isDb6v+tKkum5Etpg7iCAJ
Pn63bW6YffZX55sbzzUH+oCjFnPwAN4foYCGtcd6YmlZcSt09IjQl9mNH3nAjjjZjP979q8Q5Q5G
yWognl1/KQayngoaJvlql/qMlmsyKhNsBlzGDhyDftowtkNHKHr3Zlvw9DHR35OVpyc1K6cNGjHv
OLsSw9ifycG3r+sPGDDUzsvyNAzkj0GGXhhp1gqg8y1UQsO8rMvTx/7zvFuBaNPbPgjQ13Gr9xAA
MeFWyoGVXfs6UUrd6ISB3P/dppP68oHu0ZVWMT21eI8tnjdIVsHCstGY8x2YfdZeD64mTs552BD+
7rvhtd6QJzzHszdoatqMks2D5JkIL/XwynItSFDaS4f7u9asnqYxNyPGGEYTIQoDxO8hztC4qMs3
sM8F5XthaaB0sRcrKtKmRSsXv5BsvjUyW5/vubWbVlj/yf2yrW0SZcZD2U51Fg8BUOCZxPELCe+d
XoEK2g9vl6a4uQAfdbYeGV/0vcJCjTZ8G8xzFpMmaos7gdmuUMjCRlP5TF3moTdiH110caZzDSGk
0d6i3LIOUAswvUTbXNKGRA3QL3a/21ZPQnhIVgB+mSvEIdfWLolXmBXp4yXf8sJG8dQranpMaTnG
T5a7qOCOlLVTA4o+gJdz2SHSaY+eX/UZB5XftcN3rHTACB0QbfkHOm1Uzk39U1IbD8V1myyicynO
6zoD9H1L8AHOpdZpCyvkqORODzOqDrycLSWTfhXj4DHSu8HXvp9C9IO0S2ipPDIcs/9wSAN25QNP
F5cYgIC4jCjg2OfaDZTMIlzFZeAOCgHtWjYTaYbfbs/bSEdiY5WbmSXgC5XPF2py38CGdXHdARCE
IW1Y+d3V14yXeP2nx9lem3IChRWJaQkwNhjxhYisduzetU68hc75ODWci7VFFj9cOS7P8wo51Ngp
sOb+chlAMSxUFaCE+Xaq9Srb71JSkffuokfiP420A4Q8G6BnEHHnAeynWjKFR27oLEuAPqoDC1jl
sU9Ae/QqgX6Ku1Aip5q87MJtvcUST4lgcSuwjUJlMN33n+nduAqkn36VNgeehRs5CmjhMF+FGULa
cZdiP4O6lF5SpV6b0LbmKAcg1m9g4H7UmBwC+rJ04Db97edM02bhy9ar3PFA8weksjBGcVGJOsso
l/nmvvZjjFoY5a3Fo/W0q4mAtQmWO5QBGrswgMuBUmw55XoQEBhDKVqvQMHQhg3H3I1rASdaBelC
d0FXQRM8pk928yXAXLQc8aAM7/JCDztawOIQaGqNrZnxL2Wxd84O3YzdFOQeIKvmkcgcyG4YHV4V
BxDP489MJq/zHwfNW/OHSU9cDkPjVjAOq/9LoMMnFwis4lkUPgozpeqc1N/kYY33dayXtMB13It1
OrFwaN2/7vQmTcIlVFOx8a7j9r2bqCtpb0/vAyAJGa34w1loRyRibhsn7oRAuPb4Sw3eL+TYB5jW
IuaNjkZ55sUhaRaMxr8q/AM+GhjSkQ5nfkEiXFkzTH+0EVj5zIwOeDzkQRGcExY3DJQ05riuNVg8
Pqq3ikSyLH8tSwHQT3Oufjj+HlaTGD6T7HrFesay4GTCNFAj+11abJybmKiaF1qfme8PbY0NxnT6
6N4JhQMnpJDIvuiQG0a72mpfl+kcm4kgxART+Gh1GywxlaCUudVDj7HOsilxMxWWFXfOFrhFGLeA
cDQdIqfGkKgt98JMxCSarcCfcYzYjmhRIA9z26HhisvAJ9yDHjLCH/t5U75y2aTM9zdgwCyo8fzi
YeTEdcAwLw0wd5EfZckycU2XxVPN2v6iZJDVyCLZLuTRakBOE14vY91hqEAsXEUKUSf5WXrhoxty
7pBCAvlFqiZDqqV6kOr7IsIdQ8mriBKsIwAezQJ5YOU3ORN06a8HdvoR2zpdV5iofVbbpiWVuLeS
SUeY80AdHEhrw7Ugy0bDdA9bYHkhGGBfrokUxxn0nFzIcl08Fmuacp5oaoad/VpTME1LIFGyYzoK
ZpyQtXrCDQ++nIwz4YTmDI6KlNIV/VNho1HowGI3LP5OwVH1URZHnan/4nLehJtzjWvNJno3/uxt
CPHw8L2EiXiR7SOCIlWWCQb6eYL0UnAo59/bLwtmtI+EUq1nUTtm9jItxY+fHvZdLEHIEu9tD9T2
mmXjWFiCAAAiHZoc7NW6uA5yInUeaXd2KnfBUE75362A4fl7bAtbQgKzUVAqzmdTuZWJxpN+kbgA
nkTlXXfjwR5e5qPbwt/DGlHcdPRIoCQFPXefwAdd5eipM3FYl+7/L1SFXJDAqVE8IPjOhbWsdlZ8
InAXXQXY5+QOrNymzEbKB/H6S+4udLcUkxZqN9OiQIp3ma2WppnizYFuU6T1qcqffNHjDgzTufjL
0iHOTcZ2nd3i0lZAms0N+MPGHN0bDHslypETn7cjJsrQIsNxZ+971RpkOQLSh2360Z2aI8Gjsxzw
loCNPItyaRntEg77aPPXzzT8SArpZa9GAXm2G62iDSPXyJiPInDsNrTOqjM8/rwuX6leK+OldM6q
3jb2K5OnIpQm0XGAh40tr9NjaRbMCMVWuKni1kDUprCzCw0NiPqzUPAs3dgOkHohD+ux8AecD35m
wcS8LOVe/rI87sMW+SH9+448BQqg7BimXFjtd8AiWpa80t9cXO++hUZhlVJHnDGqb5zVkJ9cuhLf
7aX68mluhyQUO0KoiRQQuec/OFqhR5/LljhaB5os+84zYDpxLyUjo+yVZulNKURdGmLYhArf58I8
URESuxeviYLuuUrcgmTwBxdf6Z+Qf4bvECfCXII7sB1LM8RsEBuvVzkJkC9z3+70rGtizMSOFQtJ
AJvnEczNc0FxlOKFmhEZFr2ck12xSXAZfFwg9DIV5SU/8ZL7HamUEFNd3BiNHzLK8p5uA8jtifYq
y/W4LW5BPpViHhYQ0P5XDQehqjyl9YrT3InHn7r+LeD9exUXiGL9x3Yz3tavNPNc5y2sXPGv+gpV
uIFAbJAtKXy6xxWsw9Snn9CMD+5EFFOtNsTV8gl2Pr2JzcgEmD4UNZhIAP8wcSA0k2IkNmoiuvKc
lvnwyn5BLS2poeRTEdJze1Hkz01lcJfeRkfGCaUKte/SkjY9CKrnNDc1T5PRjJ/R8M93hFTRoiiW
A6Xe87AHXqCo1fp9df+5DjHBLbPW8xWKPX4I3ieyaB1+NZAkXwOPXlgyeXWe76kFlMCg1OYQ+G3H
/D2SE9g3JTAm9nwBwWpInff9LVp7l/Qg+7i4kewOYOeiI24QhoKzhKX5CorYyZVQlJ8kSV89tcwg
frOgBOwpaD0zm6zqfEQe+YOCXqPFm2QsT02RHuGmiJE9Pdj1nlwPHpcyzXAWGt4klCzi081oDU6w
nF3FNnCpo09uwtm8oZ4RJQ7C4L/CEpJjchqz5ZbdF6F8EUKLO0UNFRa20ftJ7f634RSr1iUzB6Q1
yHumToe7IQl3qlukxthnzSGSs7M8Z0XdMJ17mfa2ZbmPEhU7MGClHVqKKjpIxAOD2cBPle7CjEze
O00+UGMK/O9DewFwddF2vUkxBlPH67XuUuE7iuQ5Ovjqr7QPaZolZ6h2hrBOWcxl2Hb1gG4EmDRj
t6PnmYvE8Ch1JMRjOdG6Rl6bG267aCFSvtMv2KZReW+mJ5XXutQVluZ01mdRBkxDgICVsIS0WTAD
p9ypbRPp1AiAG//QkKBjyC0xfBrXO4/HLK9UxE8AyeyOIjs8yh4Za3zHifAueUb/ozf6sTrAw9vd
12hx8DYpTRY+iy01KMWQA7hBw4CjCaFQiIKLvFVMsatMp5Z4IV0BXL7kUKnn7gC4CQLYePbdgYU/
+83+JXHDllmoHuKr4GeOckALEpL0OtknuKCQDwwF219jYACjdCo/U+FE4V6jbVWgZ76lVKjErZqB
DvRk/TRIl3jnY8rIyOySyW8eyGUvWxbdHp9dvIwMtxKGAlmWAY5WpwW0jMhFajHGeIPhZulqfQq5
r0cD4pDRyaWi7zg6MolmrHS3Eqn1NaKkBlyWfNm9H/d62pcSL+vCe3P0Fiw9dkPsIVwSH57Ra0Wt
CVcakvDB7hvnUHP0R6o8eu5zutvH64Ccrl4PW+rxpjPxOMuRWrdfqbxeQWN3R71eemeL49L4OGj0
kx9OKumdMj2WScPyRyDIC9gtTtfcyvwkZ+uBmdEmwmABHyI6LMp2FYRPk5TE1kkID5XSC63OUeRJ
2K8qMpLkUtxJrflmWLA/FjqvHbnR43PgtTRB0QRBfke87I09erAV2f5XP/31kmue5/urShDBXNOw
8Lg4yUpxxSfnkym33+t7wxvbpygnTGHmNeOVL0m6f1SLb68nW8RaETYRFKworIP3wgFsvtTDrm5C
kp3cDNInaz0FGY/IiXODdEKpFn6qbmbaO35zKhrsykQ2fBPoAj95lLSuZXELdcftZU/19+M9/EMo
3xrB85O25aW0sFqEUHcRRO9D4PgaFFEjEPs7r8rwAuBcVAMnhJVluzsW3JWteXzOInZNXPwkXuMG
CuXFceAU1IWAhwab5VbMRI+kCYvf+7uo5ICwGX5pZCzdIV0bdfAAzjJtRc1K8xS8GSjLvbfXPnPZ
XfS05M1r4HFtd37E74I2SNIGXQrjoOaiNIDAWMphTP7neqkzRCB5fwjVy8whZgyvPe/4SDSDPr9Y
BXoOb0HqEYNWEtYGX8lELATBZOR6GTtgcl80EkECQTDvFabSJvbKoaVslpOikIBszcJhtcU/Siee
wt8P8eH++BFevbYSwLaA9+B2Ob2u4fpuw8RaO+vvWRTnRD/rfQmYvtx5zXf12VBzNobTeRIZdSig
g1CYWncVeY9RdPJ2vNIlA1/lZykMyNivjtP3By+5dQdjC4tzm5pIWylsP1MTbVEenFOJZalNQ0uy
V94glFQ1UuIA1vVQIJ4UOH2e7S72phWsR8zkSrRdwoaaUrzknBdx4w6U8n65kMyvHqb5m7KXO+mb
HG27DHwPBN0XtbAOFbUc7pKbg57duwpG+HX64i4JCATq+EXOcbxDhl2CylAqS9Jr/JpPPGgKqNZn
M752jKwCly/dlOx0gszYMDLeyWTbWNnkaNVTQyUx7CDRjY9m7WTLFMAsfdSsiiBX7008oPzxt5c7
M5yG1F1FZBDtY0VxHcavKpjS5UDLxHP7zPjEc3OB2OJ2V4IM//+UHSf0w46/Jyq0hr+bwvSl56xm
3rNOAVRBJ6N/0E+EPH4q0/HqzeKIDm5Xc9ZGX+nyDiD4e5Fh/AgKRazdM2fQcAwWcL8G3jH6E1+x
Cwj6yAMrUu5Rq+JcbwpkR0DX5TLFQTNpOA2dX26K95aXex6GxyhZqxWewqQUNzG8IN3e23N8RXoi
HNpVtWN8Ke3oac0uMbtmsjnbBOj8sdyRYPWsQ8Ht+6ZUKBspnnoial3IglDuMER2f12lnHjsvzim
Znr3QcbEbgUd39wqQK4Z+2cLhMLapo4Sxto2+lzyeEhI804p/CUJUEgHtRFVEKYqSe4Y2tsC1r6D
P31ZjP7/Kjymq1i0vIAD1UsUUBShs6Qm8Q5PciXJB76T+Y19Uk4RIBX3dVNlfzznqjtLl+2vQjzb
YztVbBawkk6Aj0wFwXtdCFvn+UkjM89d5HF3T6Ha9U1Q2KPulmc/AEBw20kGm8q1eLK/IzKqyeAa
ova38YiwkZv8P2cDblAwSmyBeEZeG6ryIUtARgHRGp5zdL9zpzxeMiVMqdldmp91DVruZIE7lWTE
CgJ2DCunzjoQNclP4H0+O6J3J7Ihdi3Zv9itR6K6vCM1lFEL2ncOAw9UonXT1+woOXlTMpdj0lMy
D83ctf5GbT8voLcBJzNuVU8LNQkGHjX0mCOKX3V/qzRG4wjEWt50aN/NRNwDVAU2zEs+vEtoWpPm
P/iHHIDDuXexwYqWxVLZs2GujotZCrU2t1zQ18+ryzSN22C+4G4kjho4hKhRu19FOVQK70+pPSxa
sV6K4CIA/h+zk7ncBphrGzcVFo2Ng6yY5HqHRoAn+0M6zdxJSSh4m2pMxewZMjGQkZ2ZAc6j2vNP
0mR1vRkyV6+qgeTTLjJcFGLe4F1o+Dv9QCd5u5fjyVSvYaBGi/s/BfBvKCuYhP1uUYDhUOg6BUae
I/LVDDKFZDfhYK0TpY1X+54+fha/Tpu9g6JXPK5RtxNip/glbuNpsWh2hAnaeg3b9cYpGZ448C2j
DOTxKcTfd9T1XdQLtm9nU6iAW4jSU4V8eYcXkvMTW7cE50u0xytJS8/VoQTpJHjcV8WZH/0uzDAc
vZvEafZDAX0V6kEQtwZXzdBKeMNZcOCR7V+O8EAEG0VzhG5bcci0cLVjcRBvc855BwdGFsIz9B8i
cJGyEh46GOBRsXK1iEGNoUQGraxFAqkVjHwfXI77MG0ITiX5L2gtRMRJHrGFc/m6zzOJ8VQyPjsJ
gI8RYmYfQ90HcIIr/DGQvaQ/vku653mWjL30z0NBGBa8vAAOIoASCyUafuF3JrS4zk/CDjVvuNDV
uq3l2XoFwtWNElA88ME/U94OGrVGx1mon2FDRmR7SOwPFA/NlenrPHD8IQgvlbgL0ajYpEF+5EHb
gOuqDV4JMD3OWXkUpI+uNYP7ddujDVXOQcEs5WGDwg1wBw0ZzziQwu72YZ8azoVN+xUyrR+O6gpd
OU5dXswU/vyx+OOvLUU/xowp0aT+jpECwby/KxJihVX1iRA7MkOw1k9oS4KDf+cFdKLAr64l7mjd
bIDWb8RmLVpvlqMieSCB3CcnF+MLEZj2xtsZRPB43Vs4ZspqXbWoYJtDdhb0e0I7z4c9Lr+DUB1r
A6QGTPPv1kiQPWJt1SFcExQ5zhjTShI0rjm2qWiSUGUzqQBWCRedFoldGnDn7In2pp0ci/fy5bpr
CquVgB+hrflDkV0/iHWVGmK1Pwa82zBBf2u7lfYknZbSHvVOrrfnRLKzZgiqnki2txpvaZtkj23s
ClTikB/KZPj2dMW4JAK/i1xBlrJ8ONeDtX3xf7JlCyLDPFBe9Wujnhk3c/4bIbIatN3Fopepe7NR
dZ6/6oXUxD4LtWzmIILQSuKxYZ4cOAoUMHQj4f43zl9dpurY1s5Ei3uhRkO+Hmzaq+I2dHPSUVhr
MzHaNoi7GHehivJ583GUzdeErY0cyawzj4AfXUvJ5qHECT1PCvNKHxBj0TBoga5OpmTNDWcqmpXa
PHUX2+JskmU4moPhv5wE25fS7fSGzIT/0s9r2YD7TpKafNLPR7UKIfZiIoy7Oz5vT8iAbsXDtjOd
pB9HBELpRlKfMkksWEXT3dTIAoUowGB5M/spWgF2PEWVd017XaxBZzOOJCJdYx8IxdXQiYxoWiQd
baag6uCOz7dfwUn0dnlQg40aeVFbcaxE/dnOwZRk8PbFaoJ8MR/SxO0msIc4QVP0PYvKDWHqPs7w
E6CCvBHIxLR2Lc3AMsFGoe2BkdPG9xFNempJiHnsOVyKW53BUtY+ez9UcofeNsHp4eidAIySBktj
lX0BEovss7XfzDyTYBwo/zD0fZZCFx5GMILjZGbVxLncHxJqOpOCcENEkeSIKsMfqEJpOHq7SJ9x
Xrhnve69jnPN9gpqDhz79PW2aBlbQxo5WSVO2uV+JkdVYrkKyDXNbHai5WYRNDOlXXbTOJk7NjZV
uSibKJp0TQrE2zL/VzWzm6LjQx9eOnIGNUrK3Tn/GGIrNwzeIi4s7Vm1k7sm3X6ChpC3BZFfUwAv
FQm9xOYwCzL46eBz2dm0shlcrMsmlS8+8wCEd/9hZODI0MWtz0DsrWjMOGypDUVb6+6OhL09Io1M
vSxkShnk8DFUupER3BI++eOGmti1mpr7vsy3keGjkuE1i/fOmfwOFJWHhGTUgJ7Zf1cdEFz6ZvIc
9BhgWin1nhh7e9AgdvxF1g27rTFWgwRWwJTyRaAIRIRrHJlLJSS3xd+RHskZcCY3HjnUhkO75SR0
7X0587n8XvF7hnPffTrQ7qrYlVAE5qtLbnmWufX329ZVYSVUj2SVyH1l2BWYWVguZHeZRmFuWXlC
ZZaoygnQSjHZlAyWCljXJopTDSCakOl76FfNGp/ncX8YEJUTR6B2j/V5IFtMzO3MmbRZCSqFxm56
phdBjiCFiFv8WQfrhvwdB3EBZrQq1MB+GHti3Q6IFxp7OCQbiDw+CeeAHxJ0dOG90E/K/ZVXI6ms
k+NJxvSSMTM3ZcT8+/GWiMGxxRFEq0VxFhAwuoOv+Yux+wpcPNYg8j1E5zTEQ0cBzXzk0CLNwTKO
qzwa8ZmZDr57oF46oOokjG+87VlWvEQkpnVFG+UBuChRG/SIJQYcG7xQZ168Mvb9368s/6uApamb
6r99zQPW4zZYvpsM7eZoPbG0WNS+4ovozhHEYDrKFXkaY19WLwH85Wh0udI9h5ArtFeDl6XO3oNv
Lk7/y4ZdUGxK2QknqZwbvybIq6ZGREEoG3skjZZOlEIwAWoqI8JxHmgf/uTtxrNoruxXVz4mudjo
CQRnZ5bJ2K77bSIrr8nTUSTrRno66qHt+V4Lcr8OTrcXV2luPs97v7eFFbM0InTN5RNc8F6YTcQx
O2oe0rL+99lJxTvJgtHi62RQR2agGJsmjNrJEAp5bHGgGwT4cv3wEt17T+afGQ5aR71jMjLpPtn5
NN/1Q5KLfkzMYGHmvjdaImOpnI3WEKZM9W7QuKBKtL5snZaeF8ga0Rbvaw1A5qhBlyyR/temkuWi
X6KiHLNhEEn/TH8krO/JUQUH/RnY2hj38c7pwx70P2vBTk7LJuiNAlWOIJn652zxN3tyawsyUM51
qVewCrmpcz3yOyBd5XAt4uoma3eTKpIUgLtNm09xg4hac825IEwcOsLw29n4pgeLUH0vI1rawLvX
8p8xthTaR51ZlH3sVXuaMduojzL4U0KZgVlsdetIxmHklczEqOc26/gaXJBEx3M8YcHZlXkxcKbe
ZzywZp8GCeIzXdNGAvhN5T6ikVlAGmvEd+9zgDmGayY3BK+OJdwhBJmH+Gl19TD4YG8U/RhNx7N1
7gqmcpScqhqJGVhVBfC+A8tc17P0rmkdFXDc8GO18dgge7JI8cDwaWieU+kCQVuXMXELgKDEOCIq
RD7dNQNumQYH1YIUKh00JFW3bOawVh1L+m26pLc71NLWjs8DKxVe7cTgm1nvJxj0mRfmvPN0hChN
S2gA1QlYPv11nn2wEbOXS2gV/0zFDEIl55QOf33GwgnEPjdWNm1gKDg7aMXhdyTjFV3BH4akBha9
uGFQxLP/gvKyv1I0mwCN2lpNqA1vzqz/riIBaAKSUrKMdKprqABQHViCpdPw42IjrdStC0YEGB6z
PqYp3h5p4JvcFbg2VPqKf5WnwG+gXBzHhGgkrD3JBxEhiUZuURZ6k1qJLpGlzLVOGMlpsU2R2Svp
qmsPhe9MLzYbtZK2dLVGL/J28vyhL5gX4HxQuxz69pm+2oy7bbBJkpLR5X/AcEgASacEBvVQe22E
SbcERZV3RxZAxNDaooPWSKIjIY1in6sae3f+KNWenfnZgfVinje833LpgvFthhK0Io4nF3IbiAg2
0e3cViVb4IHPp5ea/f47VSH/3gsGRLqFa6xtU9EWiduM9qI915Tgv4+zQfxaE50LKYUwLF/g83sg
kN4tp90dSc5dq+Nz4zkLIIYlCG9bsLfm3UFuc7hx1bIBd1FSDVXGl3KLO5vSgYhIVl5H4BGwJXMh
mDvDwzFeSQ+N4Mv6V7xA/u5DgWnVEaPL4DqVwN9JUC2i2FYEABSeB1DQ7TTqbJhZBFHn92Gf0vAi
lesHKZRblX983A+tryD4aQ5oFsOlvi7+bL3aWS4RrjIA5cHQV0S5ACcP0CWVz7oEyMV4sSVpcSyk
QTDSk8WLa2wnj9LNyUwTBFfv2FfR0d+TkOnn2Ndl312AsZ0dM1a185foUPyoYVNL/3RHBWaq4Uor
yybGHGIAb1tgXNhfG1PzrgESRKMLfHTRW5BQA5/FRoCsitJlzituqIMGHSeL4O4ttHlL8h6z7lPp
+M4WAs7LQVGQUVMO2jYXXOHsjeckrnjNN5FSDE0a9uLhRGy/60XRbC0suD6qCsCWxHoKPZyjtlYV
NrIk/vprHh3eC/01A4lULpU+Vot7wWDVn1UezN9Pcxd9RPZnLzz24RZ30AVuHyW2rWFW6ue8mSDy
Nddx5g/UBWkaH+L5j5bgAilWuZddSdy+t28ihTF/ubRGsEVf10dzs5nAHn5CPDOlLlWZ9JTggno+
loR9G+RAqvXhC2w8fG4uroviFVMRYKUgJIilDFBfLAckQ5OC3cJLX305ECvRd5OhJojQ1RqZN3pT
XP0ndQldk+RSj7je/rP6qPB0uznHDNjlw/Exq8yBGhPyfAzef4pUUS+XMBQ5/k45w2j7GZHTCcZY
MqCj5QW/uGE+giVVGCQkVMzijLdjgVxNowOgXdQlMEI2XqQQ9CjDQMWJtd6Ml80KALPSWFl8f3/C
Zl5WhsCC+oS6WUEn7mz+m1O2C9JRNx6sn4umfwaGb3/gJvY2Rt+aGhC9U04/fvtaf9Yp2EMBSg3U
TXwtFAEESS+5Ksmi57hJEr6I3wRGYcNMAg5DaHW+rvE7uuaw8D3EpkWdk/+l/27HHeuTUPsO52OV
WjbILYo4OF/DZf/794PAB4kBHRe56W9ofDXYGkS9KlRPzDchTLT/TJyXuEAlqkjRyNgb/ltgUb+Q
veEmwLtsAOLGXueEEEBcP+1Sy71G8OM/itJrw/JJ0JD4BS9ws1rZ8AK0pOFTGRI8TiX3fCWcwMat
s2gm7Wf3axPiNu/1uYidltyj1T6BpMnXPEvCi7vTfWhP61JV+9rgMilM0RVyng4/a+5psjqCcpCn
XYYgKLR6UdYlWGPQU/Jh4BAroQTm/8VxT4pDvPPZnwfaPHawNdtx2g3ugJpFlI+Asmr9Eat6N82T
1EeZ2yiDyJR1SZ//9tbm2mtp2l0nhr2N1RfPF+6rE3DnI0CzSrHE51sHVslu84oe2/I3UX1SKIfl
rHaBskAENrP/OvQhNcJmLp1HYpNztqtg+3lZtI1N3pfWsfN7xoudGS0YyqNmeb5/gG0+RmyiTaZb
cS6FsAYLqLFYl1UFX/ZENgESFD6K1gxg+BfcaWjB//7XiKQfWUvTjFO0RPQnB2IgwWOZX42vp1tg
/+QEqqY0MumDKwcVnMPhBSNM94A9oQLHWxMC/jDZA1LwKBIZH6Dfu5h0eAblR4U51/iT8TySo1Mi
eU6K6C+Ow/C1PL6/P+pE07ocPde01GozxCLtEwMOAfGdXL2aSFAaymXNFzMVGWNEnEOu6GcIMg2Q
YP2O1YUuQt1LAQdIoBejwn3ck9jDEHgGAkejTz+4bXHY1Q3RlsMbaW6pLCRWCzvTprCTEZHLLfZt
IKr2qFhT7risoa84ecOspTzFomLuBLXk2I5046Jte5r8Kksb590vhGeMw4uU1KFbzpEbA8yAsDS4
Ej2qUngB6r9xE8nh2CcDP9hfN7CY0k0niHdQ2ABOGehjzsexTPrMMBRIHMiBty7hoSntROHC50Co
VsEGgJEm1v1W8FjxfNB5dJ/ZnMbKMHkb/n0Fqo+07J8ISk4L52AaKb/RLqcsLW79EO/Cnh6gpGlk
ywIGyprRKo/zGfZAgHYFPDDWJuOctn0+wKbv5BIK7M9oSUncbJJM+I5SKdcYT5KirlEirtXW0eCP
RQxAXXHLbXOidZ94MSYll8BRLm2Mp25U4uoNtL7de+F79ja+l3lI1rcOm2ocyL5iHk4KV4ZB3Sk3
3HTbjrX6/MtSA+vS1k9PNi6MVWeSdT4RF/BdwgYRdGG0S0oRNFlm+57GqBeTdoEmn1/B6UdEi0L7
qQk+jQZdLenf6QJVpxvLr4uK1AVBQYo3u1Sm8LJbUdtbU5mZX/itexwy4ivMbRrnLaB5tf3lJUXW
svaX21vkMUjJXVU/DNxRsIYotIOck/ZB1f5PxIU5wdTFWZgVWWUAYdqzQVoz26iznBKuqUPmjima
DP0MGOhfXkKluXhujbYPVE19HCNU0YXrIoLZzMGLH6MkQNyFWpuN6vv/lHc8nP1oszcDji7ZHXZN
BK8L+A323F+sx7W0S/gN5aAP74qEPK/0vVjvSEaz9fZUzWp5sreWMdG8yy+daUWp4PpUFrlRV4hq
Ux6OZ4ystdyEzsKUhl3mQuDn65SJbhiTUzdusy8TzG2vOPdVcys+09aUrNFOEJdLx+YrBAtoFI0B
gG1/1b0DF8HkLgVUS3MDFtrK7s5blbCk6Msfd+BI3rq5k2ZxGAaSffG4692lJ1mQd//qtJWoAADo
aqbe49e0Ey64zbmkp/qf64fV7dXfXHWQ/hhMQzy/EPJqlbAmVhob0DPosIPA0u8pQy8EQQmvD7xQ
+xp08vZh/2+OnwU9N+Gc84ML9sWiCC7spxNYGIguZi44JE+gZ7UN3BVczaDqdH+O+9QSDUx0IeVx
wM62PR7PV1p55spj4nvgHml2kXznUPEmtI53oD6ZKxFje48OcUxsO9BT5sL/3aykLVX6FukNPF9z
lXyBYgFXFYgFvwbDXl+cBFtyu+WQqvXCvLesBn+ZKFcGMDs3UAQlReaNm4NbnM4fKxviFeIbXut+
LgaW/J9tHSokNBioxw0Q1FyCWY0Pi84AuR1hdpQN1FZTmG/IdUkmgYTVa03kTAm/8F4QaFaZFGQz
ClagAn5v/rcPvqMgGbdWbk8uETiv9S1nfD+oKzUh969jjtzap3cZPt7lwHkMg3wEfeWXCIIrcpE8
Utd5/5c/TUArUBP184VclBSxizD3mTYGvBD2x3/mRTc7KGUyHEuKYgt+gnTC5XoIa8d2Id7lGUVH
mKSYOodrVDuPWUvR3OLluTf4Qn4sRh+ad5t+sIzSkuv0eIBusTvrImrs/jakRX7LDmp1QSlOgwZu
ZA9ErXrNOQte3e1BPFA6vJNQfNxrA+Z0B8xDwXzO8VtbbJQP45B2klby50FsMBcnUOlHLX+tz7tQ
u/n7H3jOyycj8Io3hKmEdpMTMNO2MeKTpmq0MZfgbadfuEeM0gyYhP0i3R3co1dE4yLdSNBQhxzZ
IXkRvJH3mKSkqTxeoCmnJF4wz3vhMGVXT4ZHbPocreXqoZqy4EMNbClC2z0HTV7xQrKRv1CMI44T
alSvSGsE8uelCOXrMew9mAQi0n9HcMQEeN6LaFlUV9W/m2Vwo7dZiwPjposYno2nDi4PinZv6C1J
lkH0ndM98O1tmrKGuM4BM46aWn02YRd4unhCo6KI8ujHETnLBIxmJuQGdtaKhkYrF1euIXFgtulh
9UkD5ADj0OWGTsW5lPyJpLVsfI6ufWTtR9aLCLS4HzLhK9fiCn5KjS5tJv0BenmPTUDHWF9e8ocY
dF0LAgE1nNxlPJRUICL6H7kTb+4NPmaFgjdvLuA3pSpTtfaxtVMJft8WjRtFeLlQnB7+KyvwXmih
cMZwBnQwBXV9Dt/KEByJutpVEZ4MDOmm1mXjazN3F7Yb/qkB5bNTibSxXwJcCMd9pTetYP+vEx8O
xsxVqkVYBTx2Iupvivz6pzlKw2GMeOPO1Q4HZoaqM9Ilsoe/NadF5UdFGlgM12Y/xFaTWsrfKOWj
r0aAN4vLYNP4wBf5/AYJBmXqrg/Vgb2+jNJPlxgYghLsyV23xWAaAJfUZK4iezyms9rsYUZFgJcF
SIZsq2l4n/QBD1e2Iq0Pw8jCRnfhWQ1+e4l2pqzI5xcPLdwA7yR+eFnS5luXEGSnNgX13XOCLWOd
HQ3RCOrk+tNP1d4clcbXjigcQF8VA6gGREmPLRMrVSy0IujA1ZomxlP06GDqTzqFM7/V35LLPOgt
4ccjpyagmKxl839MLtA7b8lRBJjrgCpOxvwJYwkt2Rj4yz5MUbi+WCIUXd0KV3qZ1KmxYMpMYT0a
yjFJJbQFA2qA8f9sOTquF7jFcNrrAoqTAmYt1SO/FFVEozaX0yOgY1y2cJedXzBwJ6QBNFtwXONu
3LvwEoBYKzwB7nY1paF4JsrJG00SHR61wXnXil37T2UEVzWjObjkvrNbTwQ59iKAfSYXE99L1eib
5L4wCzPyZaW7z0xi9mBD+NxeMy+TpN90G/a7bQ/bCRBo2q6Ke5PRX+WD12BhBwGLDLvasFq0818o
RnUUibvKCmCrRs35Mqv0L02PE8YNUJIgj4/4mRrqNgRpSJdULA0U3hsJvnd0M+c96pzHPkzMEQH8
qLvXU5FF5rrvNNVBg19RG9xlFSPTqJNH72ktLsu7lclffSFvb7EINz+0R1Itec6gEJEsNpXVvWYO
vlFG6H7BVZwmtHC5GluViuBWFXofieAus1QrYKk3v5sril+fbwLIXuHzsQMTLF4ab6i5k28RxdBl
37WbZsxBdXEpuAQvIgjJ2luYvAKbthwSvRjdl9V1C1Vy4wZg8JDnZ+GIHWgXnFzSw4ZKQykSj9Ng
je0DbUb/SkL2oTvre/c1nJxsY0eEiGqcjzcFKx+DPd9PlXbvooYG+3czs/h7JM17M1wBIq9nSz/c
GUQORGNH/imygGQQ5p2qr56R5x1sNh2jX+eYAiMmrbpEpuGDyqUxFtZYRC/RhbmixGcNyI++fl9h
PuXAbSY8Ckrd7DLSYVGhAmCIWb0Ouh8KIAaDTb/UaGumL5cxfY8+zrMHgV1NVL7ZX9WY4v8ulPBP
fK5xLNhs2rt1i1bTztYnkW59M8Fxhh3YKHxd6ydKrue5Xr1A/VUubZcnCzNDX+QItY7gMQFwu6II
RhloiO9hDcIb0oplAXJGVgN+Z2H1bjMs507TrEEFNuo40fdWjbMZFBOwWFPGBTFmKaUP0IkiPPba
h5KLX78lJddE/+2CZdoUfOyZ10nZgeAYg66R1in+QSLNOK+GOPqtpo2X+NNlY/04TFXe1cnSXQkW
7MnoVCg5LytE7+B/U5hmYBniRrKQTngRvmuGvivUZ1QjMEOO0IVyuGeJtNVha8cV3CIMMPyaK1uR
vpbIjivZcq08QFP6dvn2OLfi7ehtefSbfcGfxRDeZLWXOfY3mtbJ+IiL7O7i7ZNPEg+3ctganaY4
k9JM5LoFh53zj+IsbkyH7YqSNsq513uPlfOVhVhb+FKkP8dDyy/eisrAYmD1T8mRSSOzuFLtCQx8
MThG5TyMizNCFTow+Q7K7/xvxGlxUutNbQybxXriHLAlWYlfhXT7hyKcufjqnitnE88ftnDoDmS7
8NB7hJOnUyfgNBLOnUnOwthexM79NwT6sbD+RtkutRdIuF9zLkjGvITnODDzSefCTqIdahnVyDxS
eNQtG2MdYokqCyMPpKTi3L1jehQiPpjuXKPGQ3OR6GxxsOubFN6B8hDICdCZn5lf5mWNqZ8uqHOw
64WivFV19ClyuhQ6IT4JMdXWAw277DWcGNVFgrGY/dcZ3aRQ+AQxx/9wudAr03184OWT0YGXQsis
0LzcsEmCI/aaaTlH/ohTCV5nwR7VLwb2lHGJ1lPN2vSOv3/nLFDuaFUeFDmZQCEmkStcPQgM5UEG
9Tr4JgNmHrL9sHx2Nf+h64P/DfzpDkRJ4wrrm+7UTCspBBHE8RD1jKWSRfg4y+OCYD2luRCcsFFX
k+zMrQ9YKaPowTjYUtiDZq2uFqzTi8Etq55s4OU9/H9Ev6cOesk6DxMyxOkVjs9sr5At3Sj29r/4
+vc54WdJOCwvuhaUQRzh2DguDRn304NDNPRZc5o58+HR6tr4lop0Ddr9dWi+CRiYV46f/Jxf4OTP
Zvu1JlaAQKriYojGAq9EzpiS8xIe3JMCIcIgu5k2Smj/Jfx0PwdlfQvg3ikS/OSv3cY5DLZclDPZ
BlsEhuSROVHFpQlwEhQH7LZXTemvbaFr6u19ZvvFts5r2s2dPNN+bXfYUOXljVxeMJ7POK+lkpIg
WrR+r6GFxIyvD57s2MULD0iZgFOosOViKgSCfyC/p0N0HosKzIq+hVeN8m7esFg6LBeqVvkjELCb
vWpUCB6gcM0ZemDrft5DRanWpzTxAUpVhv15eKFhTyLZcicAkVg2TYvqgwBHMAnRJaE232QZcVUg
N1IPp5w3dAQMzEWBGZXukkx+Z36c/BjKfQbH1RR4Zrr6Ozr/UNl7sZ53hD9nSwYiatwsMbljTW8C
BoDQShSaQsm0HWf6MQTXMNVnDUw8c5pLjyOZXIdJ3pC9nEZOzWQ6TdocTEqsjUxAEiVJVyDbocPN
lSXsv0MR6C30TFgVj5vNwfx6OF6h6Zv4vv2jf6qIvZUgvcciY3lU5xSkW+RVVamLjTTGB/zVa9Cq
nblKzhIxeq1rNXO4Yw66tRVXAi1IplbMiSCzJqpNB02wehwaUBI7KleJf7MZLIAOYI98Qr9VQBa1
ulxWuiEVNfd7BULgRViZe8OqdM1u8MVYwukCjyeskXEsqijIFIF9rBhribFu4Uam3MPKkZGWDt/s
1HZB/GTibsIzdvE3WflRZxSpPr/yGLdV051IFIbZVE8r084VtJFrojMjnNHkjDs3A6pg/51RTCRf
hu5C5v8FxH5bDyWPI+IH4eyVMVKpso1tp1ButxE2Kit1lSaLUKGMtFdoglen4SEBSJG1LAn17GH9
qGlfi9of3E5W8WTF2AUQa1Dq+q8+aaRTX59+BNfG2DUcskg4MqSouQztL7e0l2S33Hh6gpyz5/tJ
+yyomAX6ELsXPkM/FnfOvoksEr9pq+Ml4/fzOPBgUay4r9W1oO007kYOoe4piXe0UznfQlTUPoT3
7QlCjqsG6uVfqlG+U7qjxOBxTjLErj7e/KxN7kIlfTajH90mBMepYhTLmcZ7z/A5KqhmzoWbvk53
GrVrnOrcXsMQo6M6LUvRXGVgfLy5gv/+MfeQhkBjmxZBFSzhxi3TPyY9i6u5OFFusAlAGZ/h+/ft
AcPRZcpcKewLKetra1PpajPza+Hc1VdGbHT9SJwNLIPpnizk8zt4Cuquy3iHl+zMwlhQoXbZwp1p
ZQrCV8XxbFDCxmeSsUcM0KucO9tFtZ9BjhKO/ctFSTM9jZsozeVwAu5UXou7w4F2+ZoCc5Miv5w4
RRVO3VZuXT6Bp1OsoMDPjaCs7FVFMWSMG/XEJ0pABBDSyH3Dw6OaLjjOBbK0/YlxA8fLjpu5VLh5
8rNNqBI2Kf45YXK8nUFZQDau1qWmyCROaAyeoAi0FcO/TP8iL7Q54mvBFn9TXvc0XmziHBIRvtHF
Yy7kqd7deha/4PZ2g5EBKRo0tksNVSPxoG4piKnQD7yqQrd1HmUkWsOsiOWTnfyFrrxr5jth6Esz
JOwN0SnBhzooNagzYZ+Pz/eQJ1PrQ2MJEdpdGvDfy7Ihs3HlBfaec4VY1LWazF/HN5n2rdub+RoC
Vr8N/yepys8FEx6y0ddPHAWp3+JD4eP8/xWjP2GMW1hlkE6pW+wKXhT7bxuqbAxHwJ6q6Y7JcI2t
eTrJVDatm3KejDQZd77TfewxT3cdZ7IYF7uKbf1fLge9diejR7n2FODjN6pQA7IP1pLZephnRVnQ
tZHe7XZlx03mrh2BrzOJu4uWoXkOt0H0AIehghkH8gTHd3ADwwr7C1JxNrwCK17XboaZRqdvQ72H
JnoILOaNIesLXLAbo/Ia2oDvNDNBK8Ohi/1yDTmka8HrTxYbLnTNit6frWbLSIosfC0RGQOvzgxs
ZEGs5KDZkzO2EWo7a+in1TwqKR3jjejAJsPr6d3+oDmDw4rOEA/3Coq/3plTbcnGtw9cNuAKj35s
e+rxyYYEJlMnwva4cUDUlKTxzIz101z8/6N55oxlxpqQXtzzE8lwBHqH1CzKZuk9H/6Hti/EiUhZ
rQsQKWFzC0LLWfGICELcGAu5Y/zjwkpZ7Y70J6JyHVuQTSePY97PDggYfkfMzA2r0mbZ2NwOdFQW
khmpJuq0vAMzDBF9gmA5SpeQQC77NNOuPtNZKP+BOSN8PoaOH0NPr5EwYy5Ro3XXE2P1A2yELjNF
LS9vwr50PfHflovhD6U+yQl6ERWDK7zf4EzSy1Y6q+jMDMbppFaKLL5XLSc/03vwp0cpkcoLjYSm
twpx2TNE4UyrN0P+UN7uM/j1fnyr1xbojflcWuhhg6ptBz+1X6tN0vhQy4x68bJAzLcxADuHlMmm
IrEm6eLKRNtNUJMDrrEzuJJ7KK9c1REEjTWyY5Ma74acLJpvpdwUsdPxSvXY2k5Z3ieguseXGt3e
la3kw0bLDQfKfjoM8eA2Xut+0t0K0r9w25/w3k0H7QXlNYls/eM6qjKBIFafxaSUmyyBxsokPVcO
puj40dKWBwe9kAJi6bZQU2jCDyL59vgid8NmO/9xNI/FRkximvfM4qJVx9Fkn2osGCEqBoC3eJ09
ksPUTj4HJphdcI+xXj8lyW4QuSBdkWK6TeItD55eQgyCOr3BLj+D4rQpNiwj/yRQe5ofsbTB6C6F
/5ID2YVHqtOAqEz5MFyWXQu4wzzj2+ffO1Fc0+g7MMvtvaPJt4twlvZIpGa5oC6r/3uBYF8KolQs
33OecKkB/SZgjbxaO24BPxSdXoTBRxqfTn1B+rvLG6Yx4QVWCDucuDpTBvmkFcDvEe7lTyFzK5VX
EUaef99hUGq3OgTqnWU7cdb6S1q66kE51lIae7enwt7WWdKlCkEfdoCljrTh/UBXRCL7iLkxVHth
3zkX7jA6I261da7NJ3OzyEJzxu+kNv8ls+M80gy8gKoJgyi8xWCSYOrGgeokWGY1VJzoxWfGpDOM
/R41e/1qtT87KRBLlqZkZfVCmw5re99bfAPLd8cp0UvQ4Kgtrawxzwxp/jHDCe0YF1KKFicxWr/B
uNUGJEcMUt/nBndESKvWTEWxKJteZsRbsTaA5EnYFfRnk4hsuhlFWTB3ZpFq9nW2MBCBA8L2ofUc
CcCEqr7YshIZxul0IUPNQHvWZD/dWvlbQ+qki+NrkeTWb1Wok191G+ZOBIvAAlCggFREOqjT158w
E/q8rZF/4l0e8aa9g7hhMOw2/Bf8OeCKnjnEbGynidQ8tHQXua0rLkGG6dtWjS+TkVj4/ocsC6zX
TGoV2n+JxH/OZkw1MrtmDr59va8G+krTJEgfu63Xgkhp65dv1vedUz8k1/0ukRds5ecaLdbklQ1H
3E4uikvDBDjkLdD0+lQklYDz+zIZNQBOoAnEM77cyhd1qOvWmYMNAO1yfXVXegiAMZl0UedQvnVz
DBbo1NHugMttZwcu8eVc5OXYJwZeteeb13/+jBNAK6CHhoX1R7Fuinr9IWC57eOyPjXp+Gz7Uk//
QErjHmqNhHNGTzTIUiAfsD9wnGhrNE6l24LdXC4odYihEU+v6iDv2/fLJ+BHaRIeC0dy+5gGz/8r
tiqW2vTtZLeQwDUIOXgPboJqz56higS6OSNKNFVc3aSLNfzPbnPJcsmF+lw4/O6ZGauUZuxfAyej
kAtECKi7WfnLQjZCMlKy+WV3pPqUYD2ahAHVuB4o6L5vDBIVYuONziJvuZzonem+sLk3rpasA/+c
bvHeSjDnlnWgtfLcfweYcdDvf+XdIZaIkr5DP1UL+o/DMgOr6uO+K2qLJC6WerMd/9hLcINSCvUI
N3IGFhkEE2AWqsaOqgb5/er8jveA6ti+kE4LAOI6fPU7EXkPW3sthS2NIzplR9EOvhFs7K4W17w0
vZXcQK+ecYUYwzHZayF09J63NPc9xL+1FDfh/PZgLrOThsMkbwYUypjUPGGS9iVeM+Ql+7NJa839
5d5kn3xszwMMCkw8TzfYkL7ZbNDtMGU1CGdG1c8hJrGZDqIo+aeDdlHxPYmXfsRagcISJyg9igBY
t34P46A3QVm4+tqkbSkpbgpanpyi4vspvcCEsRaKoY0byJ21hayaOy8ZVwU8eGbVahevGlG9EaC3
zHiTE/19JjSpmzZvRa04h0TZuraGpyUCiAOzPjsd4stvITf24/Q1JJQSKvdDgdDovSnS1V+qh3b7
+CFFMTuIwnCsFAsYPn2kie9JCDPevCUKa+7y15ZizW0wKcoPq70huKJOE9MfHs8l5uTkh/e1mHyE
du4MW8ZOSc0tN7pxhLq1sYU3O+r4BiGXG7pX+EyXxFWvWDpcz1XQNVSLU5SNGpwO2RhxCLRV2c5N
CqIGxnfUQQwI2hEuHLb/sw23nSGIPaQdUbscTp0jFPuYWqMdxGipDgzrjnFhQu/I95WSEyJf1bo5
j3zIdLl3w+I+H44+QgFtbikYF7V4iduyslDZ0nIIggiyY+Xsa7z27jCbR4gCAg6wGsSe0psqXOTE
GvtZ9EUAqGkviMj1/8zYY5pucJB8y+Q6TYoDdA3VzQeueL97YwQ+s3gFWFmzhGwtNGRsmAPYCZ+S
bZ76rc5IYzjsTIeS4lwZJ5CgeicnYIMSbw8yUC1BUGs8ojkpAW1gLTzOMWj32/kl7OKeMfiWx0x1
EENQ1N/sC9FLxMEOTYqloMflrEBATZcbTr37dhJIG/vS/rGiPHes4+iZOm1l4buGsTbwHKYJNejB
NhOsWEb6YmxbOmKeyAZAbux/IvDaUKgTEi9izCMZG0A5FswlmiZogUffo0UQ05xO95+K9/ix4yh2
6JeygDyMzOz8o5c2W+3s9R/I7rx4q2ExWctuLIk0mI5A89QJq1kdy1PdqDrc3nC/k7f0y8Wnaoal
u0DElfvqqy7gBxYTK4CZysmS0KGWSJG8UrzmwBpVuvJXqt0+haXtsfmskNU3nZd9EAqOelfRrFfe
Q9sfm3PqkIjDSHjsuk9hpza4SL1h1QX0a7xywiiPV7hE1gYoZw+ig5BNr1TIag/cLQ5uT9IwwTkj
fAk21ii+EcfPOMlPGOAqddJG9CoBwbLTFeNaAOlBKJ802JAosdgF3Frlip+jqlYfRcPmRgBYTjcA
YI8F6ZKQ7FIJGrbw1+1I7KuoSVRs1T5KcRV3q3OVaQKNnrGlpjN/NHEOzJr3qukEN+bC1MbTCt8H
gd0W3g7MonmH/ZJvs8X2NyaFJQJcFw9g859EITncpmdhnBIhPnpL4d88WC0YCPxpvAINXAlRnncb
l9+92XPBPOCCjmkQRqJD9HK4j/qQ6DBl1BwYzvJ8r+ajIte9VVCnraiu21/lRz4Mfod3m1ep90E4
TJLHvvHoT7k3ZZHRdY+jdHhSPukzAlWRg36ASjEN3ShsC+MxU03sEk3LucSfagkogBN/T5wA3Pmi
69KZjmROnk2oMd15CXuo6+MUGRDbri7aqUS1WX2o+M3CgsbNDRZV+R4A8T/oGG9bMwm7Z06qKgbs
ylhDzqcROm+7lyrjL6Qh6UugUzDe3A09ypdrn+VDlKWP6XmzbK6t/UzMPNvjabzQWUGyN9luTfhL
gm4x13vYMt42lAM+OF3r1iqOhxCGuhxvgSxR85ebJZEkALRGbaOdIoZ/YX7f+f8kgQgQYS8G6Jlv
Ni3ToVDsPJadldynKdsRoDZKT17DPAllNLsKDOkYziMIrIIWFpvc7DHR/u1pLcuQxW3eJXvxBY4k
cNDgWv17r7eLI6OYaRuDp9SV+VfPS4tJatcSwTtBGa86Cr+Hhszm2ToM30XEWPx/APSkkkkP4eCH
Ac+YlowdxK8yRvrnW3H4zalKkK1tRl2XW0hgjz0R1a3Hz/rynb4dPdQJb/CFRBR0aBdc1R1mPKka
2jLX4yMPnsgUc/BcWHsuBXzjXA6XcyN+NrvAKV6fCLNfTamn1BkK/V+CjJ/O/gSQ9KiavIMb5wxB
I4/tRsV6ix7VVKlx7P0dJz63nBf71cRxd6yQNHUzMXDDwhcgmEXjBn239d3RfubtQy2gcrLyUGka
vHqAmjH35pEQl1FgWfKUiWmUwJilhOKddWIs/GAn8rn3fmmROFVuVjt07hr4pDCz4zH8L5lnYVe+
AWpMV2gQC9wVXuFMGwdjm0JlzDjZCisqnMyo0lrWu+igVAWt9POgid0MS5hxHaL/uNC6VWbxW0Om
VL5Zt45JT0wNMKGR4W/v4htBqcfxysgBNpzuiZXnQm6heQG/G+weRsoaP+3AShb0+JwpkkbClvTo
/oRlClV8jZdMCnzXgtGmrZywXqw2TzRpcjgvvNg+dVLbPvlE32OIxCM5Qcq4z2cyQsRXN8aR0FBO
y+hytGEIj6QOzP8PRYc1BiCMs/t6O5sElufRokodmsLupV5NgUrAX7S3fW5z5XFqTbUQwhBtPtPH
7ZOyWggx71WxTTFWnsK8arkt0N2wQ74RaMsy1dpkW4w4r8RcGULUytR5cXhNDbuiu+uJ16syn7w8
txPHFVOdjLi6XdYcLAMNha1Mw97DuiR9tArGHM25Vivfgo4YguIV/pUp3QMH2+gpCga1JoAlHXpH
NNzAFsKAhuNLtfcIvb0kcQ2psZzPrW1x1e3E/Wz4Ux6UzniMsS/wl1xrg3yQTV3eVNRffG0lOYOo
ExnY+jaiYoM2927mgcsWQrPB+Wl6fbyXdA9DhlLQVjbV3Egi0sIn7Q7SJDCvnh040NP1kWTX7a7S
TZe+6V5FCbvP/VoNk+UTSSinzV2h/IhktLH3cgqp02Rsl0PWv9gZhU0Fb/ZEgHU4EsdLdKwXw4Zs
zrbnKILGQW1WciJJQQDg3SFXaGzj3TnX/69yavip2p5vVWgEgDABZLeoRXZ5HolBQoEZo/L/c61m
ICNK7NcK486+5DvuIDoULvtCpTE0IokrKuEzwO/3YCzi4gTfX1xmiNgwUjHqxIpVg9DPZnyZcDK8
WUw2ixkPq4WgGrGajt0QGE3f9bEL3tlKhQQd4wubczHE2EeCO7eb2sGkmR5Tt7He4SctHjRlvXKH
+4/8pAraaIdpfdXsYHM6E8VD4BeJXBJqylu7gM5DZNWDkOA0twf8g2YEYeIcn5pPCHbhsICdhUz9
46Zjb3DagLhKfvBAlkFYWUS7/oH6bKFjvxV73La46+9lhzcA0085P610NSgEsMh1RRmjt6IXMi4J
UP88miO+NZqLtbhD3d2hJiYwxugsoKZkG4bgblirFfa8wHvaoS+HRZ3/xKZI6R54p0Lt6B3KT2aA
7wK/sber0RAAqyMX3Apf4i81F6+SNeA4nYkD7ILBKo9LnCvzCxVlZaCbCkaZfwHmrmKEx72o7mKd
4C2bVGoHwWGSZ4OzcQcIMMnzVe9EKdNrPJCMu8sv+MEndjorIfQkPXwdTNWFFGs6qLsNbWTLyodG
VCpAimRQUI8cXSLmIs43/fTMWc2UR3yfFicqNgEpS58ScdHWP+i3v8s4+SGh3AKOmAnD5b5M4xaH
7it0q7CSIQ0RGFt73qlyh3zcIodv/N6PWOEklGdG3fE+WDJfUa8n6cyhhiahIrYC0nuio+m3Kk2Z
1/ARIO0bZXbFOKFdcErFhS00DcTRhSv2D55ugugGE5GKdNlJT8SstJ02+ScAkNDQ4/TmcRMQvCmv
y/ZbZooSA3p9ESoIGCp81BuR2lVgDJW2eElTTy8tlbjMH5c1Vqwe1zbi2suBf62FkXxh31p7045z
nAjEHKHiJMAqBLpHoq9ECYfBosh2jhsSs1SWg5bWZvHU4Av7UFW5eihe7c1WloiOLyrPB6UvO0Od
uEEwq9VgYUV3f8zBs1gc9kiYV6xPA+canXsImugzahNhwDYOAOSz3A/QUmHrW54NDPC3yWoESQzE
C/o+eJGDkmLQ2yVq2etcbIur/xChs9bxP7f5udyMJNbu7xE/0wIL/76XgpuMkIHNAqRRSTixCsMe
RqLgse8NQIRyLXOAtGUIZYv4juQnBINlnYBjh65D92A0Sk7i/r4gEZw2TQh5euNCd1C/I2reXB6w
EJUK693MN5QHf4Z0CEUOe51zYpxfGfErnaYQ5ty1oVLJZv6wj8by58m65yWbrB0S6KJyjwloCYds
nLJnNzy0kQMYQN0QEloYL9oyn1HjHlWXrB+8uUPBXJH71/9VT7QnkdrNlNEJbCsknRWDmsyzIumq
9nqBfsTvZ2DcQCXX3/IXlkLiO+IEtGzvBYdwj6rlkho9ZhwWCmuVSxRe0dBft7qzh+KZi1TnkvZ7
WQb0h0A3GuDJPeVnIT4KRLF8L3vpmoR6pO0LoYqK2IOPtshzQEawBYdGkkPOKZaUD8C8iMsFEVst
34PDBTJeWEkcB7GZIyoBQN27/BjbdB8wrUus3N2LxZSBQ7219xKcj+XSeUXDbgf2oS5yrw3RBvCi
eJdXhrrtbklQiWSJiZ6/cBdGwFK7NImzXghdwYiNWUN0+9E4k7CLQaCb0fYCZ9xTuQLRp1UmSQHi
mU2v4cR7tD89HBYPhWv1wW5fERczsL3ciBHAv34KC+lvKiF9xL5kscCzoBDitY8zlYsSPHGofgHS
UQvU9ewZDTHYUAYkc5FF+R/gujMUMT09O3N1Xw+uv9B1vZbRBEmMcjS+2y2QR1GLzpyZGU5ID8Mw
SgW0b8sLX/19t3esIET2M18ZoLbJZ13+XtDOvXcXJUsCgdLzKgBd93+gRPm+xiHrIFyED59RoTZm
+AH7cio8aCHDhPWjWVOo+s7G0eqKEX8QsxSsg6rFkPdY/Cfg78NCEA15jNxQCISvjtNKmSiAUrns
kzO0sYAIr1zHPQz6YuT84ZDyz2IWJt5kBY60hNrMcjNE7UHIB7e93UFsjieXFnwpq6jnisiu+aY9
4R1PsSjjIkIO6naZVgU69Vgjnxk71HyUZvk8gD53VAwb+kE20vOlMdh2tvgi9EOeUzBa7t6tOxPY
V3lJf+dLZc8+xsnLo/SNEB1RaNKKYkKp1QDlMKDNKHGstTuQdGUj8b7BnwutjHBxtAC08MMpwLyp
3KcxbSMHE+8umMTqqG8PlP0flbtP0oKtUpUJkFDw5JAjBNeHDanniLc8g+B01EqpFrxwzX5ZsAzL
iyWI6+7O7YKwJJgypuH9qUvolP2NduULdj5Piupd1Xo1PbSmMIgF9XW7xDSUQX6TBxjA6wX6/a/c
1EmnYAG9TV/K5M4JguX4DiGycfPkBMwKjjBEl39oVWgUBsAgna/5KjAkORu+4AS4Wj9d6GzCE4ew
otwd8MtxFQ9J+2At9V9AZuXqxkaZCEj7hcyTcMIc3fxGN5jCXR1KCiyMy1Busn1jTaEBOPnk4rtI
narmTOT79JluPZUa2UZzaa9mk1Ubc5zRH1q2YdD8SaLPOpIA/uKkoCoz5hBpxiU0itIeEO+q3RwP
Q0s9VNICV1SVvoLEZPjVLePXYGgxGgm1UHWVttu0ztBUKMgpIzFVXeh9iebkHrCwSQYo5YY46ILg
UMyVnx8bkZArM9xn2w7dqQWsBrHKdtdZ+CwgbyKUll6gf8IZqbLLN5wnazT4KLFKiptDcles7rAk
aCuQlSbJUObqFV6xD+MfHi4uOaueE4tfLeeBzWJdxCnrx/TVYpvGzuN7C9GQZf1ACMFUoj19o9uy
TgYbZk8mJ88L0E/MyN6YSmWQ7nYJB+8aqUY6DtSfJ0rjV5HB6MEN4et+WI56gpp/ZEvx68PCIWzN
RY4jFpo/Kn82dcJwhvazA1pLgXRJxhIVJPc3ZxGY6eNXz0N0i6OeZ21AC9vMd3tpfQxsk3P+dDAI
y+uAZsrKLmJYI4rBYajysHgV1CveQUas+VgbAkep8WaNnD97EMDl3a3r/uZWrajJ7QPtQpW80aZ3
YG09wUs+R2FRzZObcNmZnrKazfnOLCG+94xRt7INUicGkDs0D484kkdNyHLu8i3W/ij8b3/OnsvT
gEurU0z8/qGXL8jXQdPSegRThNuRFOo5sx7GDE/69oKKb/zkJZ036ucRd1oS25iXmp2gkQj6QT0M
1CvBAHbwgqCvS2BW2wyk2QvwaYklo3n4Ngldueesq8gHk93cmMxbf0L/O+QQTZH/GgAF1W8nEmZl
STxczVjHFh8Z59mtzyEDHI3lLelTumQuYIOjVVmSlrZz4YMaQU/sRfISlijaM+R69OtcdQnKuudF
DQMFjLLPsyAOb6zrYBuvoKOqazBpe8vhbC2BYwqai941j50rFooqvCQdi4rZwwZ/Ch0i/dtgKqZ+
M6d/5C4M8AkpLlEpvnKxC/vi42Btyxla+bKBI4ZHQwDdqrh5RbWXc1GFON/kVpQwhdMvz13BeWQr
NIV9V6PTlWnQat/VgewY1B0gkkwMcqSFyENs7VRnpnOf2AuUHi7OZn0ipoM1r7Qedet5RWRJON0K
zQQkM/TIsQ90IM5PVKE4qIcbttKnspbdwMNp8yCB7m6iZG5ldqDAxqR1hYFB3htwhE5vtwoS+J2f
lc8IUWA6C4a5+KE7InRS0GwfXCQzU1kCckDGvPnKUhLLarOCT2ZyQ8kcC7CILzKER3ZK9kALirJV
I+zX/jKOJpRxLZyrWdQCimuCplKgHrCtZW2MPxAdRXgz6/Zog0kJ30QQ3oGKU96j76MVQiG9mTlj
cgLtscwN8hFGoYjUUecZxn0GRggVBtLNLeV5K5ZGysfQsm7PcLFP4jKpsJv0hVw86WbmdnbkAbIp
v3+x7ibKibu5vY8TqZn1r99KKLXksCWAf1Mrc23Z1w4aYATLYPE09YhLo+XMNahvnBU+B7qlKnO1
XoINDN2gd85PibsNysiUBvWSNW29iAztazFOwSnJy3mBXLsXBnDJp5da/IkG6OytnIJdD/zMJcch
Dsskz+HxRbFyzFX5cMbpPaLFcTjjEauHbMHKuOksm616zh9Oc+MjTxGq0GsGPeh2tK1lC8mc14fC
1biC3oAgkHHwzbZE5Jn1B6It0KqSFcKHwI2a7V/3R0hZVrCAI6MgVlkIpO0BKfmBjDbwWA3byLXT
AlNJddbGLPyK0EYozSLuEXgOV0JzY+/4zs3YurwLq1+rThyX0K8bb6cIRdXgumu6CXF3z4vgj7id
o5cbHoPsnlxy8OV7R6h7+FNp+YRroLT0qJQjJsD/m/zRhDOT3UnxellP2Q/nO1LWoczLgMeShZWS
VJlBq0n0GB+8RC7+G2fRpCTL9bB7ZYxckBMpyDtdalflOrsc6nqP9fMGZeRskso8qSRTbdSIgFHA
KPDIQcznRxkcqsLzhG0EL680z8zyHlCYuZTaGTj26MuWD+ywxguTd51gEfQAVUyylI7mcqcjLMdN
ZoxD+vEz1jgudA0qM7UTbrdg9KQDsDrZLsP530P+L1lv4VSKN9w9JZ+YM1n7s6GIAFdqhOspFRVS
XtJHY1sFG67NmWALBNfo+B5lmaemWT+6h0vNrEpZqep6XBbdA6FRjBm2mJBbtexY+FuKVSFT6ajP
TPvGHl9E0kmlefyVcNE9Wj56P0tjFuAJ/V+Xavr3r/pSZgrszWc/V3Ok2brvyZd4WKAJJeUYY6pr
EiYzFVgZ8iqGRD3CLNodK2U1xKOOsCsceRBD6M8RZif2tzVYVmrglnuEg5Y/R75e0r0MblIEz2Dv
OFFQx/OmrBqcTa5Pv3AO3DXEYqVn0JGtRE4DMMSyF/1Ig/fe7tM/OCaUiyUZLKtPmUdXMrptB+wG
M7v6gxfqrEIvDOdaD+1ToYZoPipyGiFCIn9HeM/XKLQcQ+NoOKG0yWAbu6+0PWWzKPAkxI8NM5Ri
KdipbYavPpdveTLAf2FMp4WBtR0c4qi6loLkXH7acPuiFLban2nDqbA3XA82TlNmX5WWRmcHpyqe
8n64q0T1Ry0yMJqYTbJrWg9zenIJ5vpxPvl+r28bNaocPokqxd+KVabnHiLKDV6QC+vIacl82PL1
EeS9NxyndpjJ1oB9KlvZNS3G4yBSN+VdThrQI44KtSbSA+Pb9lAaFDAq36QeLXBbmn7p49w2Z5jP
C8hsL/7fcTvYiIslPP+Zv+/ITe+x+AiRUONdkzZItA4cPwt2SHDFId2ZSMX5ENei9tJWk6yGplw9
roRyWevhCkiXk7vidkqJlNogD+Fhg6ROqT5v33dJCV9QkB/8y14om38CMsVcMknlHLJ6Gd5A6vKL
9dvDOG0iuL/epMNbzdqtfgExjLe82S3VOlXwwIfHCTw+ZdGGKGj2WsxM94Wy6AHvnKIIsDFU+GRU
qceQzatDzSGe8kY2re4Lmqfzzm17erkaR5FYV1ee1BqaZDu27d2pTt6oGP/ZB2lJMd2qMPWzV3Ne
Eao5fNLXkonkInSHdTEtRhDm5WmhjpliYvHReIiSxvKHRsUcLXY4vsViSPUcHA7JzWmh7oG0S69p
zZ/XvBDduCLnqORg9OOl4NDD9pbeeB6jlvC3TVohJxdspf6HFCcLzcEezqz4Fm2/MoQX6SaNYLvo
YQxhS3Jly5+uzkbw/8gfsHPzpVq1J+8F88avh+dnL/OCVB6zOzL8CrqAnR2PYOVR3RN0l11xJqTb
Hag+59mIPa4PWsZxjTEB+oZvz0xcGHgnax8W5Bjrbw7mt+C4j1WVHqiqdkKf3XwFVKKrRySr9WzT
h5OMlLeiK4K84urbpwKam7n0ixa5cLmbPsuTqROC7075EqXSsOUJixT2lwTaT5MP3yzVhQSx/+SJ
CUH416EHXGqvt8nwPDb5KPAlYZELhuTYPjZzYDAPYiA04iC75bGzho5EJYWOYnQNPTsTax4jmE/L
CYhFPteFys/qW4SQb0mYnRGturd7mO6C0umCLO/uCR1K947OJ1WYjJ6AsjEeTZUa25JcUuf6BHuL
fivSDhy/U2BVhPi+cDiyGcH4omZ5Pv8i97bkvL5YhPdPNDuyVmGtqSJJEtNNFofqGO4coEPNHyJ4
yqBwgqiXptkdk45gfSh360+yg/nB+gMoSlBI1WweK1M8NlGuFyL8Xp3AALtNGWf3Qcl7cOWXI8Ft
jBeYTWRaLtp8C4YXseDJu97oL2B6F30NPGyeLeIZEc1OxiRJDR26ryTJOTqqJg65uAYKxaP9NSAu
ZHSmzy4ThZpWW1eVpIeJtvIeW+wgmGQRBkZWC5vuOnCDpP9wbKXwNkb+OxSXakkWHILA300Cf6bd
Jzx+cLW5kekcb+AWccHJObtGKGuyohonnC//USl6bxFhV1VEWmVuQ111wyjldPxp9WvgSqCKXpNM
E1ouKslYjB1+/KZxMv76KtgJ/rIE6lc/TSlNFMRwsCB3kLs5wjmyLAhPtmokNAOVpzSsMmEWPs98
Y85CBtuMd4GLL40nrBbGmc5BFSMFgOuXtQbrMydppDwQ6+chc+8PfynWnID4gYY0qW0PI+kFxvHJ
QL9TCUYsFeBScOTewdrEfxlAPCx6QNiJSEzv55D51IwDbKncut79MH8l+eIG7Ug94+w38Z6xo6kV
txZcP2DebcEjTS8S2R1U2aByX/hoPPV97DjbwwSvt3XxEeni3iPYl6LfvnvQb9AWVpsa7vXtDlIs
6HukguFDWt/XU5JiLavML4v48FeT7TORt/VzFTL3mhB4m/GPRl0l6iAVqUhrL+/H/CPfACfbH2QG
B0pNecyrTvnLWMYXdCP2TRlhaHHiQQz1PfHR7oROMUMek5ckZCfrGCyNAi46fPoJd6UvzBAFs7Io
0WIF4AOeDAtz8E9jXK0Ptjkb+obzP72pVH9Xp0yRgqcmZkkBIhFIoevFwtREu2xeyv3G+3oWcsU9
lWtZOqByR5chJnb2kuTkLiLbww2SWQ8XAZMCWx8+B/K9IHepQYwEI6wkB/fBKzk2WzxeLn2iGTul
ZxiZCjXVRxX3VfarlcpcqN6m/hEA+poCVTCReFXiEcZg80glzcjQT0shdguRu+BMZhxd/KbB9kAn
zPz1ZeyyZV+E2gN1n3p2tkDcL0gzOqZDOw2/JghfxYBlFZ5O3CTwosXv/s2ZpMrjDyo+XQbyCSXG
cZe4BxYDz+q5ClNsMqS/uNXSuxvqu7Q4Txi9YTRFEqzJOmnxsuOIYPXiLV7haGTU9S1wK55K2bR6
045+BkbgoCeyimhDj0W79qLcHywsVr901wXUr8IQcbNxmFGyNk8y4ReFXsS86HnNHicB0c7eGElN
a9ab9XGOTxTWFhNKrcW31cVUai5fjlkCGkRqJU1JOdSwAL+OLB6pJ5Ww0tiyPwc04vrHeAvDSx0E
zcAT62/blIYFTag8afFueXvWeeADXBNSYd/b1RaqPK4Edjeq3AK1tqLXzVmlUqElQeNkerke7+Z/
FU5dNAyjD0agKWKvjtBcO7RSe2TE7UqqWuPPpSvLc8Qa67R/wVyqEOoOzG92i7sXj5PHSCI458Uw
MJ2LYatRTrL2x04zs5uj/XFkVdJ9qweRdoYc7lfISpCu1iN5MT+ajZnZSvojcqHDx1twyxN+ILMA
KKPgtFqu5KVuKVfcSXRUWXy7dpOhVpJ4JlQ5BOZJqiv36df4hxNDPGBaX4pFK3OYgKjhh/CCHCC5
m+9+HSNBbBAl0axDZ+jAn8lS+iRhuYzVqHN2JogOPaP41kM0Rr/MzaRTR/Nbc2LFo8VqlfC090tJ
9Td2t7+AWkzW8BBC8H7QR5dn8FjisZjzdtgh7pP6wcs4d8A6gYqPxFiqyJxetgDq/PEQqC/N1HjT
qpczRftCkLfoXNB7NUQIHKAWKa/Eo0mPPFLr3v4Rld+l9pR1XFfp9xu2nzFcNOK8DP79EOWpwiqs
q7lWO2BHJMfo/KgIhRjvyfl5JbC2pRkZzLiLbe+ryRTyftRukjzK2wydl/tgIYjpOy2HPYpLO9W6
DhlJ3b+lJzEBvszt7uRZlW28R9HXhCfHDC+2iRg1XQVeWPZ0ZHktpPtSlw0VrqnrV2q9MTBgX/Ok
0Fp/y4N1/gDxq4aYopsZ8G8uMBzZWcUlXjmeou8fKDXifTUqCAmPc9AeWDBjyLkMPt2eESGhxh8A
uKhgzFts9cq/npZu+Mv9CDPs1/jOU+lsXr5msCkawUTlh1Z74fvYoXUZYJCP4N4dcCT08kaXC4Fs
NNsxwL3jeHlqK+3WVKghInSogl9Yei9kyHNk2YwLIMJYNeNjXWnCuq1sXF+3GNmvSiuqfOhdPxnI
47eUuSaVXJeVaQ2CVc8/7yh/AaTcZtZMt8sR6QsCeDbSeFb9p6Z/FOciaYEu8TbW3IgesvrVbp2T
NF/wG/HRGeTEMIMyDK61+YfKsytgK3WxpTYGlRvINMN12f61dGjonJ/BXHGbgilbuPvtW9FjCUri
+B9MXUJOEh85UNjORaosV7qO//ERr/w1JCPxXOnouekZiTJ1BOCYAo4sL5fOa+XVNHgoIiu+tMtv
ix7aJ+hsOnnR75r7l4dHWjTPi3QL68f4nwL7o5J8wQ0WJPYGbmva9LwUvikkbcHKiga/ss31fZL7
m3mFe/8ygk8oDV7yIS0K5h0O8cgvIUUOebfdDNVzF1SZVaiB56fNbGZCA9Mna1YEpLZbHHNhkQRB
KG7k/8n4UWayFBh1I1NbA0HeTCBRS6rUG08Qsc473MmuJ8d5qJ5dPQ0m3ap1FMgFWXCOZBznH71m
nPifK5tKbr4HBj9kd7kqNJyS4SXhVlwKxKSAqYmkLOeNpqHh5Y5Ku3X1RctlD8Yw2otqT7DdTSIp
QPpkfi+UoL//dzvLEHeCtfoQcs1vUEAKNBWy0cHP0fpUWp76ZaVaTIdeINuoD0mr0JI5/7A6x4FX
oLsXMJd5ikcLVX/V7qMXXaCHuXklIN9H+3QuSHrUzXvzBiUf2ab3DpkgAWqgTHyK20E1K2cq2tVK
wCpyL4wC5s8CnCSkHdVsjN5KPv2z5RgXASS797NjlSdnbOFoR6Kstg9E6WTm6PmGYpEaLsgUoeAF
lYSmq4Hsx7n8a3REHVZJQEZ8jv71CLBS6JU1KUMSvXdtZeFc/nvggmaRiRNt2LWdDf7rvpn1FOnx
iZ0f5WZmWYO7+HrTXuH5DhyuvSIea1tUaK6Zm4NxR1fFHT3vOLPx+HyfW18FhTBRassxiKvj8FXU
7soAt9XIgkaVsjEl2NKjZ2IrqKXLOr5x/CX6JU7NK+dkjlg/WUbpPDfe/oeBBuK2vnHiW/JlSlGa
XFBdthFav2NPstr/faUCda5VL3LnfA6J5tpP478q/OY5eta/AhApQWJjkNk6yCCzK/CpZ8cn3UTc
gWQ0kmOUH3z04hi4X6gBFKTryUinrFy7/4f66QKEMImikrqoeHZTaWecgZt42f85MbmOy8Y3QY15
L+nWHStYF6GEkJvAEriSqVXr3aCFkRXUO0M0ibVOWLj/E2EdaEk29nDBOIakU5z91c72HtyTvbNO
9bPNqYomjJKGMftXTiAGfaZGjaFQ4Za8kdOyVLOytUEvAsRypXaZ3XXJynE7R6VrEPXiQ3m2Mlmd
6JfkO+TdDctFKMEOOD5KAZ/Z4l4+BolqEDmKJ8xlwuLuLGfUdqeoM9dCpjaf+b/qUNvdgo4N5O8f
EKhkR2y8myoT7HUylvuO3pxJ+4fMSoPVkAGabfCINI6MpBABaMsJSLKG2bi0KaqJeiCUyuVy7aAH
yYwpXuRxFbkYlWcju4dtSvFxQE5kMx2UQOVDr9IqQSQFOAYSq1uhoPaKMDZ1SNVANqJA4XskRv4P
eO2d5o9IesyKZONe9qiF/XI9qnrZEa5H8xB7CM0wbKpH0d5jyLLeI+nnOewIkgv3NXMc2kFcTMnp
ShGWlzsLu16rIvbccOFEhEtEuslh/wo4d+tHZsbTMLwcJjV2r95kemveN1V17lUE42/9l0ZKZ2AQ
XEN9RDOw0iAz05eDbbeRK+IDi1kA8uWe0AQ07Sk8HUGukH0Vbmr59WPlmzWwCaHmSPIplXsgh8AP
xgENPdWO39M28vGvFE9iKHLfjJrJ5ha5eX6wKgV7NPsDSRrVvjEO76tOi0c9k1Zzuj7RLSsdGG3t
95kVF5i1RKJmBMFAqnu+HkqZKm+/z/ZaJ4smH8t2fUHnbj9eFlL7xgguv4f+CqH058n08oXgKBe1
w6p7hlW1sMbhTZaXaL+/juycEdhtUwwncC8GZuEwKcZPEBhaqo612xERv234mna+NzLhKJVlAYlf
QyUSDH65HR3X0VymigX+KRnFfa1mIEHWLJhGmyvlsc9754JoeZWomGhTSeKlNXezcArB7LI3OwYw
7sFaVn+Eh3mLzT+LIKKACfVw1aq+GItei/UXV7xGxEVQgqyUPKTZQy70M7ddUzyHA0lPhBghzG4u
YncxxhHR/PfJFvVmOdyIb5B7hhyXiuSu3JQYynxLt76bPa+Fr8+L6APLh/0x4md3YCilcSbUiLP+
7My/grGYipTQSstMGGN80P/uQKGAW6xeTj937rM4kmi5v479pljUTerY26n75KKdrCFuCjxgzFav
9jTwGC0BHciFC56YK4Iugwuqk6SLthqmaCQj0XNAUTBVGy6MApGY11Ee0p16Xf+C3aH34jgaNpcI
lOPty/ZL/meDoTATN/pmn4FJV9b1YoURHnpo2f/QBegi3ddGaUN5xjoTNQmt92zUciLkpR2iddOf
Ta8Mnr3/RrgWdJs+1mTxJM1ITuTsMrcSXLnuCZuiEBw/NlPaCOYEgviUFuJkoGsp2b+9LsshrFn9
hOkTPDEKn/N6qi8ZU2zSqXgLs4aWeaBOWqaCLM4FkZ5AaPHvOdb19Qu1TwhonkaYtxAiVeZO79go
agp41fpdvZP/99VgtkWXDIakCj1ZUMUiMl8K4AizDlFO+PlbMcRKd7znOJZXjQSyLDL8ExY3ASwe
TXQaFWdoQzrRVhJnIPlz4R8W0ORuM1E/Fy269Bb52nJZ9dPM94QIPXmZt6oH6lQLdVHrtRl7Z0lp
sMPBGjsvPpVuIGuT7u4GKYcNFOp9v1Jy4gQsiIv81swmxKQu8t1tnI8baZfkJ66f5l8KMlZGBO3W
C0A6khkTkimYFDBPpAP+Gqk/SrRZ3nx0kTKLxhjQZAnTE+C6vT0zgie/+cZQLAphzOqYmzjoEkRt
X4TzUfz4+TQz5wlATv/69icggS2flER7JgsMY1kBpnn3ATqRaiyJOoud3GOse8cbOIo+ZYa64rN6
xDHXEW50oWp8KHDOVcbZ0EU1UeunCnHbtteeBo7+5dhNDzUyhjEc/6gOEhNcC1GoqCSXrkqlVYW1
ye3JYyR2iZMS84hvYOFRtVIbA899D7NKo62nYGRsqV7nBalvfjA2NQal4FWwxYRIWibIWj6I9bc0
rxOo/T/1zJ8fJFV58z7plRdcjHZmiksRgvBSPO/LFgYjAkgIPnrBABZh8K6Rg00KHldnDCtLInHA
VtnP3v4elLRZj6uOJsXLZ9/9v/HvkpOusNVI3QsrKqKGoELiTyN4KBgYwzaX9Lu/dEOGUbnLOm+y
K74vTEyzjvcdWlvuBwtJUF97Fzj36PKCebuM4YCBfA6nvbwiDXb0LnIMAMuwr2usikqSM/60rbFi
gm4tPJ2AAUiUmGwYn12BMzSzJT8J0ygj866wM57Xum14JtQIpFyXCbY6k7ODOPZ/sfKzD27kQv3Y
Y20Ax9tY9jlaUwLy+dSn/7u+YktaMzN7kw9J5B1B9piOlK73oFxEZkBnM6mILD2bahbBr7CMqhRB
wFjq1zSQFKRAOC7xnt0g+RHqjio+Mttmc0FcrbHDlTIvCS1Zg+tp+wW/TIU618Fspqw9Uc3FyhXV
XPsMs/RxG4p7w1IThVF5Yh1HqEq1j07kiNg3RAKuwjQM4K7KfaVlmTDwPHN+Va6Yo8Z1lu0COj5R
ffCBpFtGwGCxOv8EYLujyg3gkdXYMtgqz2CwOvnIFILTVknpYD60Nq/FNnYl8+6itM+uRNsGEv5w
DCEanqoIGXUM64a7o/uWCSRsisd8F6aIy83/cbAJvybw/h8nx4heg45vZU3EY9p/IF0sXPPOERd0
cWj94Aa+3Y3e1gpQpZDSK4H7bHkN+BTnlVwTY6cuh9th5797dRGzJsUUTV/39E9/b1wMavwildNl
qhsyNxSrbUxpOQa7CqzGTdh/5HsVCaaj5TFnDcocADFPi9f78+1yOlHTBZbg1OOIETiulNXGcfC2
z4mCP4TLNnraNa0Q8INcqfgO6pOh/nFZGH9uz6NXbbN5rCwKz9G5J1IWYlHnnVKQD8VmZ/C5Rsu8
06zhDO4HMj5y5u7Z4K8D/975boRQKca1Gq4kkp97QtzB8mV/XPJ7PGiw1r30S+wch+o33Gtvs0dK
GMj+qCDktFNWMmE9Jvjefprh6dfHt7ZArSBH4XM1rl3xBRPB/f1pE5cEl5GJwaSL3Enit3IiP/o+
mSVtDEfhlT0XgRDfdFQkLPfl9yBcA4jWcgaPl+TVBbJcB9PuO4ngQqPJH5ZypaOIBHw/juPBgP8R
FsemvjyNgeXxL0zlXyvKWPHNvjwYXAhdB+erQlYCVwizKE0pIVgxJwKOly73whzL8HUt/aTFBIgF
urDYzQRD2DJiuZOFGSo7UooFClVFeUIMTpGwC/dyTto0L4OViWXvYqZ4Es1NP3H/2M2wRn5e8O3g
JYE5ZVqTPndIATQAK+eyIXsjCRgIVLSmQgAXFoDFe++V81vYrqDxfLOqayjagZjg5sLBfPNFSN+g
SZNc6s+cl9zZ1km0Ai2DrF/rSa+H3loI3GJSZjjjdFeb9e7wpUb+cfF8U7IOLC6pHDhHU5pkpOnj
59MQRGn7ZhkvOrhG2BUPHo805zLAfz2bHkcDugyPbGpclfAGCg7uHkpe2bq6M2kEEpAV7/xPTFU2
1OsoeQGFPi79O+9BmEddfnCiXRc7jN3Z1Ofwkn/AVUlahO1UW3Tuat02uV/yG25+VYWIuAzXbDJe
rcfJyz7HTxkpUY7M3eci6yEQQoKBTUMx/VVqu45CEH6XTgy0SA6vb7xVLrgkLDgAWciIh/UEUHEg
rsm2IEMsTEKoAe9Cg/lJ9ypCOpczQO7eu8nWIzlOizr9tWBqwfE1kpY19UborxdFYBgO45NUetrc
P3t9Cah3w0rlVtAF3yelkux89kLRuQ+PL8SQSnQW9YdB9nzEjzsgQXWcuNPtI/4fA2VGxkzeRVxO
StifotivAh+Vt4rPH5KaqDVGA+D58CpDVyjv8n8prsbeH9RA1C131psWpwZy0y/alQcTksYd14s6
Vg2S3iechm9hewSLIAP/HtY5W1Cl5+i+3dul8SbjYfLdze70jEhPEzsXjS1Uo7zcejXREJ4oIuqL
dAtX8U5zGmhO+6KeTQ3Wfnfas5EvuQFuoeoFuCpePwOL8i7BdfXxuIJ+B5bmrfyz1pweTbvdD+84
2KZeE/tN8hAcWlBFHI6E//QYNDM6E/rCaHjbEIb/0qTav7gsdmo7tDg7g6K9xgQ7j2B3Mp8vB2bt
BaaxVQBQjLe6TGyMIuRAf9Hli5VLjNAat0t1o90nPKbqY8ftviCCYP0nUtz0fy0D2GbZwkuMJTAp
9zdYugYMMFchNVUajseTY0LpZtRVVGg68b73ZrenBXmZvIs0M+C7xzRDc45rW9D9etKK98m0eKH+
Qbe1EnJK64Gl3/o2rSYHLpmxkoBjL6Beuk+qIRGp3P5EHra0TmVV1/vXTR9kdTOGIwvrQ8F6exw5
cEI74qggfkfiZowsZA0zAZxxI0N96Up6ttI4AAUFasU4I6Ma/xpixl3peUAvokbBFJLkCLbbpGGu
QjcxJmTLJsk6SU8q8DxDrBs3Z39VwiW4zvdw+8uTFR4nBEx1DnuKmNStA1G9T4IXHa9oUmXsksnb
+Zp8d4LCB6bgGUQT8LF21x5bZYPcSJingtiDCtbuAjAg3pVjaFOW+rdj67m5moJDncI1UbpwZ2bo
rnq9/37CSHGpXZeE1O8E2NOgDxOA4EmPzfRA64FGeiekYxwNcXjZ0ud+TxiX8luSsCrUzguHg2gM
KY2x3SQ5N1ZpdOYd1o1s2zi1TNChg7P0VIUcp1oqSnVYggSOQpK/2fcJfhyqU6+KYR0UXRhFl2ue
gD4zjOXYdnNJUCz+q/1LChOyqs5t41KyInA5dYoKCXKHfP3eeq++jcm8cjP5rKti1Lru+Ts+H9dO
w7T8IsZuubCbNHDeo+Fq1tumyT0HzRY5dz2YIXAHRpfmui+hhtudL0kAVuCZWcMUD0ASIh44uM2E
rJ9swoT1/BEXwYYouYs56Y1BP0Pt8yler5/NNYQ/kRxwv5LJeFu65JJm+0tNG03j73ysXkg8fEvq
iqy6EkSf+Hu2dlcY/AbSUazcek8muB+Li/ZsJSGkFPWd1CAVV1TjKxZQn2mwIuQ9jAWArgrSY/iu
z7HyjldBMGxY3beEJGO+TUDf1JOA8FTvIKhDjR2bcD5AGOkQv0LhtmtMq2tXsDKfSx7c5JIoxjKh
+uQkU1bgGiDve4P1JYAfU01dj9HZDvf3O1HRBNvMYGGtQ8ujlBgDn4SXwp/5f/v0uQzkr0f9OfJS
ztCwzJ7WdAx1XngplFv1iGWmt7OunzVN6EH7/98g2s7f2HPv/AK9yK0OrbEQyG6oXAQudA5Requc
Mu0tI3Ymp/RvAkj0U245Dc6ZwtPhnHJU1AITBaOg02TkiNdJnN58YRmEymkkJgO7xjAfph4pLXy1
IWfl2vDNeR9sFEqPlvs3PT0C6RCxsXeJQ5AYxYgw70WmihlF+K4X9159AJjOAAvZCqVuJWRo746/
7ee4bIZxvHsm3A1SgQLSpBreB3boO9KHitbA5rfFoXJdAQZ1yjlezH3jxch1xThLOI3PCY7RPOvf
M88cJZBlyR7UBnoy9SV47i1ij2mMVjnw+8rO2JRZMQdZTnJggJjTu1xWuIhMrXg+vfoZBz4NU88F
O1VEbbbc2Z4Gu/Cx9XKoEl7MijnK8bl4y6XFejExjTbeuY/xoBmy4jtTITDXWnaHZiQ7MBmMyNRs
lX+ByIVBTylyE21HzQ5w+rQxDtZJtNbIzzEd6EeUg5d+821mTSVDihslT/5z1dhzLLadavfDkumW
YpVL+8Mj+NjKsHBTMh4qulWk8iL0Ui+nJY07FwmLpEfzlY+MrpRbZdMgXzQD1ygvNvPlzgI97Bpo
hrvCFGOFZo10lfwaPuPkijOv4Sv/x6ZXq0y3VGHelidEUWqHYq0LxHI3yelD53DLn9XY0fByG6je
nJL9zbtnD0m6jR8AV+k77a4g59bnHh3IqD55Eppgk8p+Ob1zhLPC+Hdp9rIm6HCKJvDDbVcEusry
CHLHixdEQ7Ihz1tgD/1kc3ollSFPT2FuzlyTGHdm4nztluTtLHR3ajaApvQ0BGZy9Oojq4LH4hSf
9BPfYXbNTZYd4apNbm1JOpTbrYzissGZquSjKdVghcfzD8YjEPOjgQpitmT4IOx7f4gUhDIVJuh7
Ki7mtVf4KJcBnLwk0CW5y8BXqzv8yJYOJQdQfrUzfAbwzpMimgStQQafEeroJOpk8DRPqFnps0EX
IARZ2Y1/96rKzUvlTMKBSS88qbxNr3nNCimBEUDAUNrksZlN50EviqzAcSFLacDwEBDfkbHqwxZu
SMzXSN/FoB5p14g2bq+nWX9tFN0sb8pokWxLKbw6+MCNX9Kj1eaptQl8rIfkVsPA+lk5qqHYNwcn
blvwKtZ900+UMqFl+rwRO/EB7vnCQwzNmLfQso5bfe18D8YDKfSUe+JbtBR3feZYVc1LaVhocSXj
1MjJyOsoz2L23iLPCkqbZ10xgS/xCl8Y5o3MYROli5Cug1pPhXkYtdkXDyrV8smx4gopMx2o9mHZ
my1Lf+wSzeXugIGZ+AMvPmpxgSa6MGR8FBWXGWaMJiyUF+c+V7vKAfonmqfrB0/zzq1Bfkq5j4D5
dtw+l9KhnbJ0+bk20wHDiM8Ghwao8cHKf8rklF1S1B/z7qn5zHv3dvKLrmF9h46lQyFQtis4llPK
xMlpRbk0kff+aOTP3XXHqc6R4SZy1Sf4SxgcDKJ+Yz0yOGXNfpnLceljbLm+6/8T9hM05ACZD2ii
ETk/3ZqSx4RT5Ox+uUNBHY5POekdAC99hRhXtgVM4Vtpv3h2ph2gGxungDJzpdWtdFNXU1d7NAy8
QtkngGi+g+wiUOEQZtJIOBnC41tiEWdTI5W5xcz8A7bqvHHEtDmxDK23EBMcoQhUM+AqKJpS2M3N
ODF+8euLwt4W3zjZtzJB+OH69xn9DsJi7jJl3Vg5RNmlvJ/j+FA3uuuPgLWmlhCwISl95HYhZURO
Eyvo1RboTzX+GpHMRin+lnrKSQYs6EC5le5RWZ8kPpcDLLkM5/Wa/0AoaFVJJlpKtdCq3THjD73C
R2s7MRkQueckiPB3YuMVXw/UcFhUjE5JnXii9EPgOkqSyYJqHOn2scWbyiWenMIfqD32XQ/qd/Te
3/32/GwCiMHpjGLGeHQmq010/2/mhfViymltZ4NKAYX6ioS5qWxfg+bpW1z2nIyNJhOVfOMHM5ov
zQjkQPyuDEN2qBKlxW3svXhI9ndgBkrzown+EItI2KiCyM06db02Ljb8aQ1/YLgR/lQXwonR/IAw
uF1J7aWmTKJW4W0Py6CCLQtddHAPDMKddA0VoZ4UevmFfnt3QnArKsKv8RCXhmzdbs1T9Fcsxttt
jMUb3GIa3cLZu23CR3yIKMy1/n1IlqainpPHevBYSJaiaSFuKYCcfhAKPVdFFvXMIzjMblbspB8T
qXdPuGdnyL/FlKhnan6lxaTbHxVoOU5Zi0Jkf0esYiyULBmDmzmiFjfKLmkaZLks8II2slTF8S55
ANK/hsOJ2MTTRLkv3HjGWTuuBBzv+CsHtJdClq+JIHW4F+UL+yPkENdkMITGveoDLOWTkLYbK8wj
ISB6ShYINM9pQWXtA7NYvI1wSJZPgDK+B8xC5PG4mcI9RpVUyELxeTiIrHjdByiYyAbFpiKdsZpj
f7xCr9Z4RV7EWhGnn2iXqYJjOBroWP7pc8F6UvSWf42e27a+/sYMDfpkvSuJ67at6JlgSe+owNin
P3ho44PBJ2N4aDWX5wMc1BCej1RPia3Q2satD/0bgmC4k1QksiYf2jH4OwEcb719NFoTUB6NXmj6
AagbHJj3KOhRlpoaSjR00fijUO9xgJBaqQf5vSDvCIJuBiA8rd5vWc6X/EHhQytpuTP/ht6Naitq
bmIGzBfm+ZdX20hgXwKL2ysgSzgasRtL1fDF5AYvUiwLWZDqjBNuJlJ7xy1VH0mDg4HHB7etuKMC
yjg9+mEc34yjWxE+SA9IUTAl1pxPpaoqThmENdZ7c9/5NnnYK9Y5izyWuHHuDqOL0tGXQJF4SJBI
mK0Fa3XT22qisPZ+yp9Ey0VzxigBHnR64pr4ZuMuzBq7eKtJsMYSw/kstWfiHcsqnCd98bdVMKdT
930V0xoBsmlkXDkhDnGuKgy6NA24QrIi8zvLzKH9ANFjKEoouNSEh1RmyOIJ6yKgcdT9ed9mWYSE
5TBlM63XPSLc2ZPuj4sbOD8gGZzMmvAOWTHhJsgtWH3fFSvz8MSZgbp0Jglk6fH96dLzPaUJcxVV
frSB4zp25lVKt+b+f7dEQ2c0TIjidpZcXYSXGNLtyICDN+Auw3rY7Qo4c3y+Vib7uF0Fju6fVXxE
3XsBJKTEM15HIcUr1NapsOEoM8a8b8ckB7GMTJF+C8wVafyNhfgq/jOsqBTl4Vcdk3XQxecuYAvq
9c/TK/bXPM2KzCed+KEVTPfOWc12J2i7deBAC99QEsDTtRcT5d2skHBEjGV1UHa2HkSQcYywl1dC
mlpD0UWc39igxetNK07uKx1eFzIaCtWJDYMT/uIcVXCI1kF2S2YN2gUVN3h+diTcNJ0TK0+lGaJB
uugz1i3FQyLcaJyONcQF//BprWvm0dsmRUyrOQcQpM+m7vWPjkAJvE105DbJvLPHVpjK+swWlHAf
tLHdxRf8quEUA+LaftBl49QU6ALmp8pkHQ0A7B0gd3d8EnQlW4icMRTLbcmrkApG1wrCqvoEzpca
Q7znrHl0/ZXoX/NGiwCVhLUS3EW+Xck98zcqiWdSy6x4HYEjXKy2x+tbj1bUqtmddu28cHsbt7HU
5787A0GzVaK8WAo4uHEzIL5v6fbGnEVSTPe2vw7MndkEiPXMk449mJGYkxOMGxSBbgXJnJhsk5eL
n+T+T4b47Y7fzjBGGArGTwTIdpCcFx+htf2GMVGyyu2itbFX92BO42HkqezMu8+L1v5Rw4IoDBwC
DgkMEQ4bMRc1yEWap3gMFeO4dWC1isjkSlWx+I0JuuGdF1jSxbyU2v8qajcuNlDheHy6u0IArHT9
snMSfoTStKARfQ3pdAraUakEV34jYOy9DG2kQPV0XqugMXpiL73qu+IFXtIfC+GfK6Uo17DXEzTX
D5mBIK/20zS7rk9tg0zklGyukJb7wegfKSwwioqGUm5jWOvuhMdUqXQEjfaToLegvV7JpmQINYod
Yp8sRwd+Hua4PMrRlPCZh0uppwlu/wqf9EHa791cL2hIeC/tXTsGb8PWdOKPJ/Pn7QuNjAwnMe9p
aYA+7DLl89ta7h1z4lTLLgWFHxGHqNP+82OZe6oJH/Gmu1o1WoAlPsuNXjt0NMx0K8v02t1JurrO
H/MFUeqBsRzgxOExrI1EXh0CW2jMrDEi0/R3Q1ViE0At0JezM13at8KGxNjy8cN42qJDI+bqMY9n
4Th85ra8r6hjWo/VcgAXPz62gUysHqrHtWmrPcFYKpLbF2l1zJvo2H3qc3t2UvInHqStPtHzovhI
wdHxUdTVnwKBixoDqaz1y94xXcg4xWpCcREse4Dpj7rZOdk+OFa3xhA5dMh9ci7NvZgviawcMluE
ztYpJusG42vSPj2Kv+IujBp2Cki81jKhY62wIaX6TPYyLzN+SPhTtGWQ81Mk91aVEVqYvUgDU1Wk
wHPpkg70RPvwSJv59e92UpPRSvXNWwmw7ExdnAfT8pBzazMftJ6umqPQusNrkTf9V3DFj2faRmOA
+lX+HFKS/4oRY0UGPfRpry/QgVj2EmyV4wwnoHJYXqrv3ISnux6Jd2H77qz8fQN9oRtjJmeMA0gx
hEu/d5uTPQqEXN0W2/8qQmDtSLlCVT2HxRpD4WWs0wjwuRNn7OGdP2yj18Y2KtlvXph7jiYpGT4S
msQB9sr6Da2rs3sHmz103raAiCjY+TU7sx0ImOWzJGoFcy1MGIwSPBt4hFYb8u9WaW2ivYCnti81
6ZEIcFTrWOu/eDHC0ac7fenvVepmsVMFR+2ar9nUEHjMtdhdBjltbaEcv/9RnOLGqabL/P8TALun
drStdaX3HwyFErFYoV8Z/vzHTVYPzsSH5FxNS04/MX3LOkwFZruigtqa0o0GEs9bKbSAzwCDfgz7
0BXwDue02LKenD3mcUOlsSE6agv3vrAW4q2LnS5V5QHGZ/XSymH5kZonuwMPCNcKrV9QAIrMSJxe
5YVl7ovQYbVy5Hpa7dt7DkGqKppt7SzxN6Wi2dpcT1kZXkp+rYth85kdkT7VfwGiJmCbHx0hkXj4
GvhTiNxdcZcDUtBpeBddTnp5XFeb7tr0ZLshY4/G0RZTzRaO02PG5t3OVrkx99ewhWPA7eQ0qxaq
KAshLPBZWMjRoMIaE6poaiWLAd8TwKVRQJY/ol8uKZeLeGRi9YGiV78oY/hjsnuz6b/bUWbVdJjq
quwPeL7W9K5U5dHSKNd9u8YtfOohrIWv+LGb6Z/xG1tLP7E5WDwp8d8ofgP0D14FsFFpfGmBfMPB
EVKfxCfnmsSATDRiizSJfAl7cie1l7KfYZwWEtBOv5RTvdEKU7cKGEu0+dEhmbbKA+yXvEKH06aA
O8jfvDqTKcvsDTjZksBh75FBMW8hTvYK3iy4YvOWpWWNBVYQmAy5KGXWMA63tb8wQIMohCoOtQzb
AJR271N8NczK5Ghdq6/sy/Jn2Z2SHMymEZVv+udfun9sOKudmU8948LQfMvv3gppvDDsk3gZrN32
2BlXdk8+RMRbqW7gJwj8Xqn7GOlekPnvfLG1Cy6y+3mZlKRo0q38TjQVX1qOvkhiDaPIJBrR/JcT
41pz0QWCMjSmCbz19pY03bLyrJbkhMMn6MnrU3n/DB7zMKQFANXErI/yKTAKtJyCZ/A1pb56CikQ
9jmrDk/Y81YWCjRygrvz3BmrOC4NkYEzPTUkZB8hBRMMD0UyKu31IzaCaecqUb5HPLrs4EXOY/az
cOLWzNGL8MwezhXxKEI40FuHdIdL8u/mLFrHo5/Zc7pyPQakznfl0D8Ket80OduP3MLlfVc2D7yA
mFv+zNu/Sd3n3XfrrdQ5JX6FuzqJDGqdTgaCO5GALbGiWpXwKhzKpT8MyzzmYAs/zHoGefRCD+r1
Nuy9H6Qc6IVDHY7WpZpRYgpXGamRD3VvnMjALj3Bc/xCj3FVmgDIVDJ4akbptEj1cUwzvFyXZ0vQ
Th2uuLFXBaXk8dzFz0xdAVQgsjL2aP7en4lvlOJZUiY39Bdv2Ksyyzl1nIFRq10lubog/0vrVHgb
y1PxQAi520ibpL7SRDxNEBE672ofYK8/VvtyUIYW+E5s3Fkk5akmIL8NYI26RemnHcmwhKFvb+WU
XlWAzGTkB8xGiRM0en4k55yqta8Q5b/nbtDXgDh2iJjT9fefhyNRTOQifVuIs5nheJ7j61bcXzpT
PkqNRMwEcNtkdtrBjQ1LOegMSvkNPUpbyybfrdTeEZmz9rxn4zHWbtLIL4+1s8ya2SSt754xYZx/
IzgbFjTph263pcIkWaYg51i4rSYprnBj6HK7v7FDJK1TVmvg8ZzCFLKSVf3sGS41zZD2fid4TIoh
G9eyQ6Y2951VX+DyHc/IuRrJAQEJs6IX0Tgu7hNU8h2jr5g8cufGneGAjCHuZswEmIrJhA2U6xjs
vjTcyVQRPDVfk9CiYrHx7plRcOeJ9EAYPCOJDIxw+DZPEC6HXXJmnEdGOloRP7Wf0/ksOz04VqtW
R449h/MilmvoGNLlc2VOTdNcxPXl7I4D65AXloF2ogr9tOqrg5LsWkODBDl6QgACVqlVNgwfNLvR
9EBT00+VyQFBctyvX4r36W7bgpbv3pCXsyhCE/OA0lot4EVV6598UAvFjRofUnbSjBwtPnu8dcmG
3FxZaRaDucxr+nKIN9M9s8zTRfSkQMeJI+0PtBu48wsyWnVPFFtC5Q2BES8W8/tx3A+jb62cBrsl
QPy4x8JeCOFT3VJMbAVRrJgdpgEE1gPi7LOU/TUnGmnAJiong/kjXn3y5oeuxy9uHDeHC+ZirKpp
ylHk+mP177VCpP5IABsNaRIdL+abwXxdAQ3nyWhK0yCSBJFZu419ZBpm1/y3/4CEfmEtvrO4v/l6
7XE3JScCscB8A9squrB8ow3Fdyv3tQGFrsc9rm/wA5iybw+dUNXeShQiAOdp7YOUYtZPVf2SJTjl
odr71EfSBUa66VwRq8vav36VVwhGfggZS+WAJfZBf41MF1dx/2xxdWEtmKvg7p0z10BKCjirX46M
gPlmEA4AqSxLgvYUIt8QMRlv5MqxX7epi9YIAtAHm2gQiCIneIj9OuZ88vWEyTgxn0QS/jOhSRMK
h+kxJwzR8CtPRoyU80oFREV7K5TL327WWdfVv6IiF+L37zwu89EI13l6BtrbOgSdv5RnBE46hbeG
iuHGVBxcv7GiE1JY5TwLEWJmgTy37PLtqaaValYvHv/MrNT92Jahet6YjO4iVvQpkfsDN7rc29rE
nZk0VC7GOpKWielVY4H8IMpzfG0mourMyPjRAFMsGwdMOD7ntZtTmSWJvpZAu4Ypaui8jLylOnqR
yHaANN7xGsdFlfkZxFtxL7gxHWosoR/ZQJVPkQxAvYYnhhgl51vnoEOrhyfsjbP4yCjXzPjuzPaa
iW4Gpkelcrz/5OX+P0KC1xDB3z9Z52lHH+wdbsLI5vz9r1eXZdKi0N/yd846RHxcYIKQ/NPwMuZq
r1UzRr1zLurUjNZLROmcjeDYWEz2HE4PZqKleYdkI5f8061XmNtmAqWVNuCmwygQfXTAi0x6Z5HC
Jnn20Ef7wxdVBXppNh/CP8cxmL3b//gY9sEQctu9BZllvBtpe+opunjjAiEodiOK+v3xiDQwAjNF
nrt6ORy2IIDMW00VIulSIH3aNGTxz3slC+/gDIYSExu7JdsxtCJfpu9U8el91vKUUQoQZSmPMvX8
lPI8cTRhF3xuyhGOKLy0RkyaPAnGduBPnfI0l5AcEu9ssmMQ8vOWEe2sGc9cetdPcJRgOpHPfQRh
GOdRXYGDNeOZLlL/hqf8N2nypMeZJohcBLrHNBRQONOrgyae66VVmgDfEFtkPdtmTfAvzXLJm7hV
YogIz+5q7rgozp0hyzOfhjoQot92Q9AdYxVKKNBy8MiRFkyzlujrUPP7KhMmluwJjOqG3JW8FDt3
boKE7ANPQMTk7Rkt3qbyqemghmdXxh/MRNXMxMTfXiRGx0/ZB2imrC2NG8cCvf9kMvFvAxGBZNkL
PD+UbFZ/IsWTAKIi21dLirasQSTM3MUKBw1Hr4gm4GDa8593noifbCumUZpEkGC9OpkIf6kV2RFa
xfvpmfVfuYor2a8oQj+zbdUvVPu6gFdI5WfquYTJAaZ3IEY45/TMweGV33//tmY0Z5EsbFwaAcoW
jTB87JWN0xcZO6jEKBrvEZhck8jme7/8PSAbVyezIyyvMEhI+h0ffJcTIy/EdruWeS31r2LDpwNf
cnpjq3VjYt+VHKMg0XtChHhYcGJyxWbXuWPV2MCmbu53lw96HikXbrn5H+B7305bdaGbJ4YWbFAv
tZ0xEZb5KnfVSXPxSCQFY5uNG9SoK70L7eyRBe0QpM8XskqZ4rKWNxSyXeHcpSOZsaD1BF08b25E
xym/2kGGwvcYiQZm/hRPHfyP2jZqKJyrR/3lAmAEJFknpUiYqkArm+CWLzNSWJQgMYsi5RSgtiVY
MALgAdIR1NC/s4jIUePRkhpBqo3psqGmBM/tf2tR7qpL5CQdS8XtzLZ6v/VNOcNm/8QzYbpk9MJa
YnanLlxq2FO+PZqok5Od9yyhCmeRekOk6a4fAbSZUx/R8LFEmhcfQkweFOZeZdv+DHENBN5E0hFp
mR8CZnN63rFqjhHbKnLJp6w0uoOCUO6zlRNExadHkHgGZ7pJuw9VWlBFf4uqAAfIySeAcd1vJVMJ
venqNL7Zqtubw3kLpptkRYsN6shZu5YhkCHGqCJRrpxFUqfI+Ksahw0QmWSoJ2xj093GGDZCUMTW
YnVjCxHTks3X317LOuT3LVCMhMQrTijAJ+mJ30tw8SEy1UPWbktYUQyeQekHIhIlZiZCIQCvI4YH
2WpeOD+YArGqkBIeH3WRmhVt8naL/pXUfDhERvuWA5VvnAReTt6LyUozug4usws0x4+4WsGPnZmr
5iQH7pxDjdV/FnsCNVYbMCq3FfL2YieWWs5g3VZYrU9BMB7LsTJa5hLEPTQOmIQ6vVU1hfmk4/Gn
9dKoTPE2UsV8Jjx0gI+jyVS9brxwdVnFkK26IICHu3WhqK+3LP+yvjq1D6UI/nvPLQY1EORrEdlB
ql0tfucNOxfDIfTY/NV3WmiOHa4BcTJ6kncVquHJAKZV6bdu38Zf5UhWoyQrKgT/1YFdS55pU/BH
icciZkkxKLaF41LDMEpsP8iKeIETHHhzCTs0uLFbT5YL+He+ueMs9gdmz/j04cf3xE5CYisV98BU
S8MsU3mxxGDg6KLXXqfBTZh2GF4qDzP7tuGXbI91Rf3/I3seImAjG7LWz+WMQ0Rsq6/XCN3T+G7f
M0jgnixCFLWAEziKqzc3jwlq5GmDwPfJP9E1SNqrjSPwJdy0pkm+j+z9paB84jMq/HAOPxGLXewn
NPhQbJ4EdA7I3iVNol6XwAkV7tUUb1P+UoNigO5dVKCSXYi6Rmj+MEbS021hy8dJdpRyaeulclJz
COjUG0jbsn6ATHnpDjDImaouNtvlRG4sWvFWFO4su2IYJAo8A0DleDNJitEWh7cs+61pitMJ8WqD
cHv1I8oLNxYbMhpybHTt1JWN3o0X/H5axm/46mSUk+4PRAc+/XpwAR3kpcP+m9F88uo/tZq4fcHt
3B+u6C84jZSLpJFhRHQC/92/aaUhFlUebevpMpS1STE1z93LCNgg9bRrwCk5JcY4gzpPh+9gIm7M
eoM9HfW5sYpcau/9Z5YsbILph1lqBjyHPjf+eYy/16EIVskGfzy+OR1Nc/7oHOdQnH+cEMjYYHrA
c6nzS+zeN3OrS0Vb98PxUgB9+21o52nyQofz9olmo3amGta0aag6kMJg51yN6iX5zzVmTfJdzbIt
Wn3C6bMBVlyQ8YuYwRem2sGsY6bG6Y57g1lhXkS3AtAFUj8msq2Due6sA0+CEsDhIxHu1U9lVePo
g6I0iuDlyf2y2Gij22xnV8p1bIrYMr35AWc+UkpRL3/e4fVz+v3GDIsTOzkLaH+aP5pgdUb0UIvY
rfyvJ5rHvD1AJLM4vfXU4PBxeq6sOzSjwweGNF3ryAzRWy40okkqQR/laKVk7AqaRIq1UfTjG66G
e8WclxMzZel6nJ1j6c6lMFEWt2RHDJRindbA9XDrEUWk6C5RjwHLgfvvASEQ4AHnV3Jo/A/ij+YE
8LoBOSslB6aDz7caageCQbxRYRCK/Hp1q4TzCRSWDTo7YDqTQPOPSUKwY14nCH8/5HNC+FI+9rM/
wL/JOUTJ2rLWSjKMmO542Qmkakh7bWVLBtCt+KN8KqmYbaohyXitPg5APvOYStAPBVoLTlEGdc32
5FKpxJ4+yPhdwrul6uXsEuIWoIZy2t+EaWz5Cz8CR61Be9dbAxqqzOT7th0sgIJs6S3jGdfPgiM0
6qYyPl+3Zd+vPQHpK3R27xiSuykmz1gcZZaFE8Nge7qXxPUSAI520gMG04Yk3dOIDrmeLh0xHbqC
B7W/AjAYJDaV8OD6ZT6l6VvB8cWqVX/e2S9/IZfOn9gm9ctjEnN4c7RTn2w8ClDmpJdSNhOP/pnT
Hcyw51gcM32p3N6V7tG/XlFh7KD2qmprwrwRljZHpaKYvAcRn1ifohCLhesBfFCNXlvZqJc2qEfB
amrzggMzjJ7Dz9kb7RzlICiE7tE9ON0d7WgejGdx0FNCH3AIkI9ObSYLKcLlQixCyfDgqBhiaTwp
/59AYlyZWDW9mZmLX7O6YmcTucCYB72M2dwXQqvjDn5OFIwVs8SRrVFOaAOLeBjKK6E9doKhDteo
NKiWlkm57tfU4e78wVQ1TL4Lk7SgKM46JpVFJdOpYr53IaoI+xeO6JaYQbJW2YK0lzO4qZHTwP+9
zkiCnBlFrzs6Yqrcj7aPsWmC1legjQ08LDisKFdNqGemCW87DXRNeXoq6P5nGnXN+rs0dkZTzo0b
Pj+dq1pqZ0Xi0t5B24f0Jdu0mVdIQlOcByjd3plma2vLtjYzXjE/rhfk6O8c+IFMcUE2B+P65ACQ
Hxas2Xiye2edGH6tSh13+retq9/va97KfVcYUkoMETkxnMQALf7BBeAibmSaI9lgCuXzloeeEttg
LRMJsReVjiRH8HSakC5tQkhyOMhSXNwihVOs3O2rh2rDP6A1v7tm9Yf70sdnC9s6L1g8dWarWvkv
AsJC9tOZysuZPiuEPm1BHc63kNZMzSxChjrvWOC5V4eIRjfo08+IozOsWPFCcTU666WaGXr5E2uj
tkRuhjea4A0J3Nox4MctvzrrF5QqobXGz/M2fGOxclzS3X2KiW5nvmGXP2cn9qxUvQO5lkvAtdoN
EEnDWFK++kHC9MjwcgPyNGJ69roPBmfNil4Zhg7bUEobCY60aUYgNyke1RRvKXeyxYE/by6j7h99
e9/otMYPQgX63tyqjPLp+tFYPrB1MycBOtd8Fgc+hMPoXgTwC2TQuGbKC7GxuHDu+PuXCoubZfM4
L7eailDfLxpUv8uN2GKcj34zsB1SlSluVxR3Kn+4VhEjUIzwz2AC4y5Ts+NsIweE8kmaeQCKfgs8
dJSlSdFwyZxqzkWBm72c9cPWuJmfeFr6MS4s97zneoPVNPsH5zc/HH4yiLJLBWaAkU7fUjHWeJyJ
MiMB0GlClxCzGP0xH9piXq1ybHu3xbu/WvHOd1RpCakaUqd+VjXBgCTATAKaONQIGx61B/51FMOw
6d7H3+W013L1Y0l/L7CT4S6O91QMzHgRuvmqYBby8UHppHKa4hdvylHoc0l+Kx3Kz2N56N4r6qqJ
dZwB/5A+YK4bDAd1lxD31j9+VqTBJL0UGPOCiRgnzUFV/S2cma50g9CYBzU1S4kq1HQO5jBTmx+5
sbds5exUPEZlaLlYGXqMR5ltPk1obfbvkrFsFPoTueXMAD8panN8a9rHHc1PV+DjBwWQ6q4dL+z4
gwTCmo4gfoWndpZOwImjSXmQA60r/TebgbjeiSJcEBpvJ0VQi2Mqf0iUnjrSJft11wwJqCUGU39/
mE1Ct2vMSnPNh1SmtuAtvUOAroCgRH4xwH1tyFRwNqJBUCaotur1Uua0bS4NyeVmuETNZ17O9uGm
6c0nx9yXg0oj5knI4qiaLoQx1Cym89hEBXryJFvrqS7pMX8gmqzyklvg/dan9IpxOnUtaLsnPTuQ
DJnY8g2wnFEdog+Kp53GRfiwBfZ1pkK5YNg+sN8wPwngS004dofNnIoei5t7w8kAMjUvCSMwtkhE
MP1gtiP+HJb4hijb+yiYPVK3+ArsyFSjC6EmKD2ejztuOTVEbLxvkSojtqiN0621I3sD8CTeDK3z
aMl1go8J8w9TQ+hWF4MFePoYCKHJ7fOOdYp17iakhUSZDqwYgvX3Yxl5/ucwyWVVKScJLoj1UfDQ
H7ZhieXpHkBge1TFObGppzXxIfo/2GTNuHpUpTxHMGI5MALF3UA96uPjiuSEMCreFB4z6cGbDv4/
1+nlTAA64NSBxocVZeoUCqX9BBj1BCcUYuR++ubFoPgRWDa3CEsEtQzl1EVdqRtjEmVe/sXNbq6e
JmDUPXACGuCw/q6f5O1XGNn0okuCBJvwxN8tZvpgqQnNb/2kdj2pSaQg5siWy0e9DEUtq3fI0qDk
MgT9C99TFtfBL9DWbzVjoIQUCt+8NNcZeHiE/EK1VLNl0g3JoMU10i8JMKllntO01qaUnfKoJoen
rcG59HOs/b1jyTXg6z3OshxpdXM9bKKZgcXVGn72ugVmLQL37xK36kJ17sRccy5x7izi7309Pcci
2tq/Q3aBcDwscUgH/vgeYr783cbRQue8+hSKZ9cmAEjbZkQ35pbanljaLpM+hrACYrwIXfHF+OQb
VzTuuygUy+wfbnrGIo93QtftaWDuHJa5WswD5JtUxpJI2gviJIIfw4EpyGpDloiJgr4/jbyLboTc
yYNBm3ixUoX4EgX3xQucvlcnIO5/jGZR4dZOwxgpI0zRM8OVC+5l45HIKAz8Fm79OA1YYbqKDDS4
XdbnmZVtUtPx8UjqNrNP4W0hT0vWNweYOoU+j3VdAfuh06H9fHVdUswR+3qWegrinEglOHg4wgwL
0npAYRbrushgH+3agxFPhdxo+vBvCjt2qOVqHWWI7WLXNw3N9sp9eT9EviTP6zy+zXCeX5C6nM4y
I5hQ4mKKtB+I0HTWHUoUG7/iJMG0L6jCaYvu+eA2+IylrIiKrEWmgVd00BWgLf+kqc18BGG9vG+U
TKp5Q9d11p/uPWT7vV2uTfEtxRPBwLdmqiqDZGb6pFisAi9pTsGF83Yq7I+8OUrA3a8PKD2tw692
P/kzh9bNS0YVi31O/Sw3qCflncTiteQNlAKOhy5syqMzpzA7hewPQeYfZXbbWmwsPDjYEsgnD1J2
WDJPST5KfzIItwLdANW1lOoR/uPJzFrrv7ZbnywSEUMDwBuKEIFsNiP/GtGBWUK6nTQRPb8gJN14
5xQZsJCCSg50TgKxG3Rxv5J7umgvzScrZfNZIliw0QlwysluncZcsdoDHpglj4LnYdI8DSfei7xB
Q5zyH+DU7NYWQNVjAtwwYuUrByxyVkCoxR+Ihc0gy2Jj/4Z5TPFPrv1Z1J8O2s8rwkWwEFjYN6l7
O2mncgpvbAgckalssoRW7txW2JP+vzuuFbP3sbjb3txLQbnUPT45QsM0xJEDTyxjP+50WzhqcJ0c
xVUSdun1RONFzCRObrehWfLER8w/BrTrufh8g0rxkuI1wUnA/+zVx+re4zUpWSDSMBv2/sQgKst1
4KEt4QsYlz2irOQw8aRDcdIjmlTm1Y9PcM6n2fOP5ZBKgpq7rSzVrB+kHrgJ9qqB7GwtbeD05ShG
g8/fTC1vxX7AmUDBPIutr8m4/DCoVMOqkDHnyKy/rfUKQ/m7HwMpenEiiH1q15DsxpNvCt5O+lCu
bBKT7WBC/org3BuEc/xXA9zCCTCHRXItWyIspEujthkcd8OuQ8cNIw3p5nuHqUHT9ravoMKBLqI9
Gj+TO2LqGRN2+uraBcz0vlV2wLy/i+axsAlOQXbYiMj4rZeBy2XziSg3udRE3unekOlAmnllLCDt
6k+x+kV5AFczE4Y8IENtA+90RvSdl0Q5c2wVroA7tZatsRG31xyZdf+gaxS2J8hFA5CuFTjfYBpX
ftegwRPkvrFD45O8trHKGL//W9H02RcwaefWDtWy51M7n6CMEjRH6p17FnU7yrBkPmxg51XYU4Wr
mE8heo1XH3mtYzB05dkKsjcnrpMzeq9N69TXNQvm3UQL1hHXPwBYso8U1AWh6ArB7E0R7YwP1uOt
d7LvjFBW7o9WZkIzKcrbYrTVbnagFULuWCkJQO2v8Kxp4UxdqkJBBu1DRbk/zC8fdK13Jd9C2oDG
TBAayhLgFgnts7leQxP+0wr8Jiz/GW8ATv+25uALPhZ1XYicUsfUsoRkfAlRvlXxJdKbiUsHiZM6
z6Bn2tak0UrdmN8bx5CoKEP7lRExMvXrtov1Gm7PzYU5yiZWQarZhj6FD0naCnYdDM9NJLjfOBpF
QHF6BfFWtXtSnNTi0ReRyaxC7QeUIBWkaTEQKNMe+/JVhVaiLKxYBlYz8SsxzJVq9+//bmYET14T
QfJwA9h5kpGW/Byc+3KuJudiKiBWZB3u5IwPTAzi7Jc1yjmadRvUGiIKtYRH631zhJByhm7QYf1p
O0D0QqKiJA93Sy5FK/gOra+X1fXG0ymLkg6qMjmpFsECOvoVkWd1BjVJXC3xLnHmk/9lWDIbl7Bf
2ho/RCA0q7At9l3CeKFTLxkpfbsu226LCWDKbRSs5b7V7FUOoDpkrfr+e1mG2jG8pC+BV9PZOi23
qFi6cmbBgO1PAO5oi5DChMmduHk1e2c+XBRL41z52Tr9PPf3gPKr3xWXYQpVxMte39RH6eDy6Z24
4yKR2yhQ3smoewzOoBMAxJrgrsjjTixyF47TzL6kJ/FQm7mGDE9NcOQYJ0YQ3kVttapPgZ9D843B
kJwcbNoYPUpr5UNYeoYXwIH6EkD9qaptTzcHBmqRRZA0QR8NlZ6RJGcw4rQ9Vj36wO11IXPZAkjT
zoeMvo9KVoIyaE2IK0YC6PprKU6kr8Ki0Ycs6xgUkCKZHiM5ch9eEV54Dxph8nMLMCQy8z39VZ1m
gUkWVbWDxwgZCOeecTIZGDQEKYIFgR66Zaha3JDfhCLGVgqyeNdEX/jfoB4Hr8XcLsJsdzHiS7Ia
hLAh1LtSXJxz5kN2ylxUsfRHPNEJ6USKB8LH5pGAFK/ySQC//jZgLjoPDdtM9Hy4XkT3E5P95PAC
lUxtIvC2tM64VruvunKKJSwe4BHUb7l6KRc0JySFatgXdyQhVq3cGdXRws0vRk0Abe6d9bG4PjHN
7FkNaxFpGAKsB2BosimYUsB4QAUugRhX76oh7MTjdmIjhxixYVHABV8wAYHffUz1srGBfQ2XLNb0
bV+kN8eO6f2mzyUEJZqFgoBpp+Zb//lY4nqBtq/VxtTHxbu97OQz6nf2sTo0rhJSg2zlOI2pVQ1w
6eAWsgksTL/z3R8W9pIECxmgIM4jbgjZ2xVrVJKVIgd87kJAJTxeVBaFC1n8qhEARDGSS37on8fW
HGxJyR2ivSZSt5c7mv6VaCGtu9G5ntAXvq1kWv+0xnbDCeo2R4+LmsxSGH5ehQOMA1EJybUIhB89
6joFsxVkA+cNEksmy+Moy+nkSCdjRBwvjtZy9/9wBQhn2FcUaiQNT4MwenC8NnMYTnZvX3bpm95O
s3dkXNPyxQ//2SIeeFu+6X2vjNLTQ35wlLjKR/e1xqN5B5Bwhd9yxh6nMMSx0doQrftVzm0TqhmM
1kS0G60kESx3MdQUatVUTKU1h5wltqkL+5j4ogcPvZ+Io6YoV6y1rUZiduwKIrkD+lrZ+kZcwm/E
nPsjj3i35iTqJoPLpva6+uxiI9MNvx7lSrpG9/HAA6vVkN/rwzt2UwUP/24jIxi/jXn7vT6ae/9+
436uHmbvIpZPceOiGLfL/5yROyGd/A6gK0684lkW9QHKsqPsnmXySrRJ3kUBOb6MdkbU/MpmpOsk
Y/WYJGwD9OHwlNNc2ISjktkMpRn3gN8f4FYkBI7juSRwojjimZL447jGAnYSWdijoZ6L3CA48je3
0p9saraBLjmBwdxF35sipsSvK1ixS3wxoAdUcilG5Jrou3RMzlqRrlEp3bUocKhQQHU0hEiHiXoG
ipU0ZUXZzYq2uZbAGKvAgDOCOzftX/WVM+IPejL2IVgTbXQYV0j7uNWzd78WNByB3b6jQCQVxHHV
IvAkiOGD/BtgRtM0i8FwirQfVHvwBokygy0PuAkBg9JjtaA+hxS7nDxSQeRQJEKwkBk/OrEy8Vog
9qS66VhzNiCU+l3Nns3C9c2qZ9xoE39n7qFi9dFYHdYjjpogFIVGvwxtssaQSF91Hv1TmWP+RSkq
L4v18McKpDbe7rGw20EpbR2YMETcvTFWZPbpYzyqjnI9+aDs+/dch6HJJ+hu1MwlGZ+7ETSVvPvt
LZ1J2NLYn8ftXqUR9bjXNSmlh1dyqunh83SyTuzarZEPMglXE7RlN5WSHouHb2Ff8GnL/S3rKIHD
DLB9HhEN9Vfr9HpMKtShnDapb2lsfWofzNMOd6xDjjgMCA1S75gzp/5GxexkwauEoI0d5VBkEADH
Ue9NQ5c1iw1q7QFjUptwIjBhtBC6RlaSh8gwxf57gHoiecQkbtluMJYIOJdAXwZ/IJ42aa0YVtdn
3QwoGZDRJli2TogN64tsMsmEsenTTe/80LI2aA2cyuZEg9stPtvbrGqWFimU+FyKaeyAxabQ8v7f
iFZnhzyMceKBAl9brRd5q61tlk1N/3JFJcfr7Js46iAXkSHYhRnstQjt/Zo0LvnNu5wXBEG9lI4n
KZHRlXVa7xbLEj8/571GJsEtcofyzWhA95jQvEfBocGPbVrh64gmGepsHDCcI8FvV3zc/U+YRAm3
7egpz+vFZrLiovxjlxIrUAFnJyl9Rhj1L6x8hp3FMhpKg3j4xf3qz3lTCWfD6ywNuO8PZgGb0ll5
RVBSN171XsXBCnPB6Bx4XrHt5xp68RZZwTtohKQLpNbTm3aA2VA4PWg/8dE2OdZttJS6uAekcna4
6ji42JbwgQ4upJ4LpNPfqjoyH48wEHLEg//pa6Sl+eVrJELDt43gF97L+0kSC6tiqHrJvEYufPgg
DDtgFSibOWKwGrN6iYjPsmAjTPvPKS/7UaxWYDBCvwVUL7gIEZp3QMileb8BD5f2zq+MRRBCty6r
9qk5R6e6sPVPHVhbUgsBqlCJP0aXPN5y9eeAfQS9cF2FYg25ZHYOqgDUrJGD7MDDXJxCmb7HDKeA
fUqG10hD/hO58NI/9ByZ2brzu8DkI2PuTq7kNQaRDq9/rWwWhhqYsKTdnqM3WuVOPxYbOM4691UP
XdvLSqQxT+6062PNhteaJbFdXpoNEgoOO2hT/XVQGnmX8ZMdWhL7B/mZ0HxiAMw1cFsQQh9uJJQP
ZECXHoT4oyevH8H3CONZC0ALNWgFPnjzYjsSGDoQeiR+iRqaKXeUyHNDyPRA587FhDAaR9zbm7ce
IppU7a3qaiqR99vGoy1tuJ+VwlPvtP/NfL34gJus9t9PZedNBa1QMjEXMo7plRhfRfOu1FqmaoSh
GiAltEWW8Gaur8Byv/86CpFPfafo6nWlngRYbzPKfHuOfH1AQ6rqzMlsdmXOmDxDuF5jm8bZro3k
VkF+lwdGuw3Ay72nMOVtSF5gI08Q/1MiMCdWxgBizrBhRkwRZ2yNZW80vGX8j6S8dGzA4U76gIX5
WeCgQ+1PsutyF/rx4VKHoni7p38e7ZbvOl8RGrRG1iRBJx9QVRksFMjO5ZwHEevas5jd8Vq7tdAM
JumZBKazmJo+qyDubXioqxaXWp2CLqDI1C9pvCVHmyZuevUGSsVlwsq9PJITsZCTy3daH0g01zhH
ickIkWu9J61IPS4nNXORv6d6h7+Uyar8xtfn9b9E8+H0zYcnftUhlc4ZNATikfrpG0dSzrA2s3GA
mVdmgj0P5rT8EW6eyGrLXoBN9V9YqE9/HehXM8s5B6Se0MqQira7L0JFkIjbIbolhCwWuNc7sMY+
AIHlSHwqFMKlrPfP7Bu35KPj3pDiEsU1ybDZi1+0S5wu7aLgjb8hkV6vorBfki0G8b0orHas5UQf
8K5OExnbts3fJeZJ162wZOB21nx3VKhY2Vem2pF/P2KFAJ2wBouYHU2U47JWc0DvaCF1OgB0Lm/2
x8S5rk+hrgebi3Ffc1QM3Kv1I9TKvUWL/A8KDaU+FWVSFXL4nxcYi+6pJoVUpgoU1XQKYrmdMd98
gwnzrVehCS+2MyRCMIeUpfhvE7eot/btxdmq9tqwKNckrTfl9lP9WSGjf2vmxaw94wWeD2qzpxfC
K9pwsKBbTCGdIm7m+sC7kar/Mib6rtCzQ5EdDkBuh02ygTtxUzpPAsz2wv4hBPI0Ih8MBBOtvNbc
7twRscmnYiYPn5eTc7g+J1P+wwovOzatQIx9FMqQ5zJuAy1MLvyr53Z5qAkpcpl3FovszhfZRGwo
ASdQCnm94zbaueKG0w9koQytJUbAUsBxVKCRsJi0Uipx56sxE4zpFG8DjPVEX0AwfPyeEv4n+GUi
pO/aWWawOl2ngBrxxis0VUjTQZI9AaJkjpZtSxbCWMCtoXD+TOtj8n7SMTe/GlKmij//apWci3cx
VTMDBXxZSxFQ1ms+5dVgsq5X0SR4C2AZ7Oh+0KIT5E9d0TrmOa9wTj6Cqx8f4W8PUCtXUSHC8deK
ksgoVLa//fU27cUK3xeoIFDQ7M2DybFr5jlJKY/LEbcrJrPFg72/79W4PREacq6O0n+cfgFCyWZS
7ma4vlLXnU2SPrYFokrj98ykwZtDNeFRXBxGclD6g5inT8p1QnvBDAjaehrHHFo5ZfsoJyqveFz2
c48Buyfv09rmYI1MNlXfpOnrRuDXHklC9XEiiM6gGicd2jrLfoYw3LCvUTHPAaLn01x+Ife5zBhA
LELkJuD6LXG2GaB9oIy+Vik3CLJIKrFOSmqFR4Kb45Z+KLFSh3Qzl6ezULIUrz6dUixGRWdBJvaP
FOhgFKIUi0HIeUXYTHCfHauHqutF+S1bFtQjjUkxbE02xSW3ildjh0pp7ggHGrNG5OrtzD/vED22
RyB/bRp3mkRacpy4nXJO9UGZFVu0uWEUJurdwa0R3BKP1E13QIvthqXyQNm0hfWqBbo5xImZGBJc
ZqJwVu4TUmpmRaqu2WusL9KlX6CgDhw12G3jiwK+1+hYBADQ/2DdsT8/4omtljdndgEBFTFoCiPd
iNxX+1kLxKrle9rT2BSnlxK2yCBKxnAY+Tl4yWRCgiZsG3tpW/6iKpuTiP3vmfitUOpZa0uvLxV5
3d2zNU+OXabQ9pRSSWV6lCF9NcVhVSwlzvVej0hpIbtq85NwTj92FWh+I+exU95NLF2OHAfo1/WF
r4XLOeSFotQA3ZJCBN81cmRGo+ryqQA0tT8TIckaienhbe6HEIf9MKMSAkQesRrk6lefb4i78ASV
dAj5tnXNRN5Zn3Zs/TNf8xpY/Fxn0Cn1/vx1FOJTldFSiG2iQw8GJNmwp1Ob2KPkXJyQ/KR8lR/y
p8LcWedIJi41jPEvOCwClJJxsrxzGzCgIbFxQTtFeXPpUc+nFBpGLOjhC2b2cFABi+eL0eJhQuEt
ilIzmyzHQW9oJL7++KzxY42ONGzO1CLQ/VpBD4PK5ARNbNw5Y3QGSkwELkRTGA+Dtc7mXevXKGtN
MG7yNRW8UAJmoadBj5qGdV7Ym8AtL2VTbhVKPV0T6Daowlc363etEl2cq9vv67GFx5fGqnpygR72
HtLJUswuzTaMhmkrg4rbQrP5g52NRiPDN3JWOibXOP7Juk1JtzpXTyFGbc9ZhvUTVnOtrjA29ciT
3A97X1h1hOi5jAPXVl/R7H46yUkbQxO2X/PfzK0AgUobWthX5qPlAqpMOv2oOim1wTXzDS6pg+5d
R83GvMS9Jp3Wqd5283BS7BFMeilt/7AC5q6a5ioa3XSEDZf2XTPsVvvXD9wfj2D2BTP/7qzlLoss
Dh94dcC7kVa2q31sIAH0IjO5drAJuNuzKZck+mOIPSgLeZrKo2m8/NDpeEMOgGHyMHaDTHUN66fd
1MF/VbZilI90hpftWwNU+mvSyiDddM7Ht/GjZSzJRETEp0ZbIQr0+/Vtil6UZTO2cBCFd9QNZBgL
NE6A4lB0icpfV3R/LhypkLQ8+zuyHFTbYvxKwyllhwD9MKzw7pY0yttrMkW1rl0G206KeSIM9j25
d21cwlTzVQPLFDWXmSJnb6Q3KUGfRhXmlrLgxIcLwvIHpZuTRxyA3uCd6DbigzI4YVrSZDQKpvVt
/yPVUUHs66EkcoSGyRvKmavea1+uWfxP6Q7L/WiImmqowjl/7AgJS21pUETKhnqDe2ws5bV1a4c6
JdqS2BxMUu11A5S1HI3Y1TrDXB2n5IbadiNOqwneU517jvR80PsZ6ChUl/y2FmHlAckjDsvPszAL
DJvXHUKUxl4Ilplw2zqB/Dkt5IuC2EesdMWnzxF36CVSm1fypkqGsXwrpoB7m8XYrpTU5f18kc2d
siFwKm9Efk2E7Jkd9FpwUZAl6CZgr4Zmx0bMkFn1Is5WiIm8LUl9ztufafrY0Qfo5a4c/a9hmxxM
KIJZ3Srxae7S1+2Efhzzp+yqqOPdH3Bo7K2ZF7v2ncTza6+H0Q1WU+S69wgq4GUBizFgkRNA2LZQ
OGH5/fD8+KQpsEGAkUWnOLDfh8ns6RB14xM9Eh1sC0c8Wd/kk3cQPQby14Cghzz/qWadwYkXnMN1
i+s2KW3NrQzyfU/KX7z6ufX2+qx397qvWHXZlGjies/afjXi9uRRK6BC2vRWUpPT50b2GzDvoBcK
+pUkmkOyf6sd6fLVGWAfmFfua0UqSTja7xrBpEzSEAwrlNTolTMPBa2m4l8mATGurc43IN3Lc8Vt
85/wGHqsskhXXbruM1L9FmqqVMlNYdXlpIk6+IKXJn0oMtAFin0+RYFEOnpSbt619MlXrbeckePv
MbADK1/jA4qfXGmY6sZv0RCx6fYR2qX/2KcuDWIA8VfhPbxYbqMgieDTMUxn+c01+2HVR2xIiGgO
V25jGVtcleUnI8ufqqoYn3vAiNKsXKLGsYqV1lYtJEBSf2O7gueBofI0ABcz4vF/ptOUp3Iy24ly
x6ETa93W8K11ds+c9HmmAFrPJYey69/D6neza6jYM0ThSRoTpOD6CuJu6sUeVUuSoFcwX1XzQG8x
eEckBLd5vaGqAe9InvmsBFXh4dK46brw2HaTyfT7Ft13i52qVh5ZHHPfjUkzgeq6MF4vXbKL9hTl
EmWFCHVlDjxHnKPHujh+EBD/xNqlavrc2HasrVgrQcGSSAP+pl3/VOakAnKLlUU3VvbgZpcGSKGO
u2aoRGpETdBjcPkLIj5eVkzwtGbLxzCosjf2z7Dp60URophqPuKbcLb7hgHSz8w3j8ipEChir0Hu
h0vZ1POdRqn9tipUHiWe7L64D6EnZX/X3+RFw7yZTWTo0hIynfAuhvpOyjxV/uQ4dU1yeN6ycwbb
OqeyZc14aJN4/3cWt2gJISJk9JQ9zXNWD2RBTmnNX+7S1eEDc8/FveiXR/s4BIk2Ay+tdyoTF97v
+OGN6jjPZrTmzHiJu+/QNn/k+5BIkcjduYQj+pnRXY9+lwRdLn5XJKjDl76ZUIWhh5yR163QvFkG
8N3XQi0H4ntnUVED8V89cAVHO88RTyjj/o/wR0ZrkbJE58AE4jkTsdOVxaZ4tvROc99CjMrFWGmw
2TFX+XII+j/ydqK684j+Gw3wae1/RAuduVyeaYGfT2tPgcJ66Gkay81jqsQU2MOO42z7dwtPBZOo
v8Om5LK77fO/YEaoFhDEBt0Ew/t1CHBOBqk/woXgRfhl6brPM+7c4tIAIeCdMtHCNQbFTc908rV8
pWsdOkI1Z114Ai3tn92aiMWU4i5vngq6Gzsf/srEld6U8CQfgScOjsdiqQ1vNRWAZN41r7Vkr3w5
IIF5NnzgEV4E7Mb4tsaZ5K25wehExjdNpscSJ4iSprlt43ZWLChXYsSWxZy9cPlqJyVXSISoDjZ5
O5buZR7NjkGhunEJAHJ2pn1CMYW52Mz0vW5aUmhJ8d2p9POTfDga4nj6ikcgjACfz4DRROf/MpeM
/4/UK7XWyFBUV0+ndQm0UVCfVu/9LcfozP5BWKgYZuhnjtcEV3fm/J+DQBSO4Z4hcgZcdByGuOxE
hg5rAPMMEWIZ2q+8FYUn63/nS8iwEF1JwF8ApvjxIsjBUWFiM3lJqQY7gTAfEEcADS0RUQ5GD5gh
bBMvH+8spZcvRAfnciruKxna8rEUzCeh6nlBxbKpbTdxIEwq6fhACeA+OfyUOaVT5UDpj3p3x/lY
End1J16wK+GuMKJW/jSKaq6mEwiRJsc/KTuXvIY/+Q+tOC+UebJaGWwbBNnFLYUvZPlMlHMAuU45
UMe/IQKjtmn7YpzZYiAYUVdWONp2bIMy5r6gGOTa+mPMBVA+eTJT7UdvYNR6DGDZuxjE+eh+gcb6
gRZbrk43Y/T+ccNmcwBeRiFnf8rKg1rec9KqDA+4POcf+4rJBu9Xle97MwLervLoCF0mjZMC2g29
FQ5JIJ9v89g2/1qpzu4tU2zPDrZKI7OhvHMwnNS5vHcwxlpfF/BiZbBQxDyfKZn8pEdwMMJb9C5w
De8bNDEoSyy8SjF3OOa24GITvkO8DwoG4zjUqHxAPcsOrJOzFGdVSMfPs3rOlnuLCwgVYa0ce06B
Zu5hEHjg9I7B4DQbBOsip7IXN72SMgD2A4iqbSAurHQs7mTIMmahtkRkybUT3gAQYuknsK+2eKRU
pB486ZC8xauMoFjQUXi3ItJn2k6QXvnTIh9F9NJFRs+yz+pLVTh5HIZfRTu4a8RSoWy6PuTSb8xk
N6g919h92O9FtGswJ5WTqlzspPdBU/lnq+qnH5aJb6gnJigHdtZ2MP2hQ5OBsyFZOP5pw3hUzBNN
xr217M7eNYxsL/gzB7sefNU6NVHYCTE5zqrfoLuXKb3SdWadO6U6ZoYY0e9HOl+QCqKsq+dIfEo6
yXw9Ud3MPffNo/79yz5qPGZmTFMEjmQIbC1ccMa3/vrR++Qz1xjdR46Es5DsGxsDQuMNyRYaWZYo
N8C++YmTQx7uJ8LyU6NW80vYRiWtn5o+ki6wk8CAlbxH8kpOZwDGXJSLiCqO4NeXLiDLtVtFYx/+
xLtRUJMy7XvoE8DzlMlQvF+/zM8piEuKj8n2sTFF0/BewZ6b7xCFW2t+aEX1IF0tKf2LOcOqdd/l
R7PKDIVznRPWKi2NQm/vNHA+U3GF9Cfnn/KOchViFc42LK9eul3TuRF3Imj42cF8TcHuWO0sQ1tX
GxEtIuDlspgvr5YHLROJDTw4tU98jQvYOKng8TCa/A5tP+7c2wYVu5VYqnThFhIW4bsgKBNQtAW1
cMqom0IjbdEtw93nSBlBiL6PdfFeYT61+dW/MAJMdLioy//cgCjvLjT1zQWdiWOOxVGlHjb82qUz
WrQU8qz/rc0owNYvnjEMpNcQtDyvZubnxv4z1ZJkEx0TIQu3dIoPEPimgG9lKztlDwtC7HgJZagZ
WKPCNvLK7wgtjUZ9vqqVi6AM3weW4zMB0V1g2q0Rsnn5e6cLJyOg6ma8uxaLLvg1yO8u72q89ef+
c4cINCsUaqNPG8hNgzvUqI27Gzl0cshKHOtANgBc+3AdWCbxjKZYxS60mowMX5SlmbWbLLLRa2bw
5lMKSTRymqdZCl5585bmZ1h9AMt2TP+QwrsZZaCT4FlgG6vMuZdMr3/GeCVrB1J1wSWStKVDdZfW
oaN5ezEJg/vPuUv2eMtIc7o2JfPUybISBFUqEH7yJcXOheEmkO4feqWibrmYowBLhbZC/kqD2v9C
PaTqcBtEihVZ+3XchrOHTJyJo2OorP120ccz3XFCnAz+c76wW3dG6Gkpn7BYpsMJbTViAyOlje3G
28xZxl4dsVixkEqA2Ri50rbhTST90z9Ha8+JT+PhLrVm6mCZzdzhDf0iIGq7oTUwAKTWvi9jUHUS
OXW+MmHc1VUJSxG5Mm9rcJrQhgwuzm9QKUxl5o/znkjySlDTsO2U0stNQ9PMqKuTm3eeqWRpXsRp
TrEF7vxMT+5oa7O66+ND8FfganD3rGTca4SnEekXC71OnuLitvWxfO6J8CkFfz/spAbW8+Rp0GW+
o+z3ww1guFAWan9yNHrtrBwebg8VIIsuH6/M0xSLGnJA8jkQ0fd2UCysI2NDukbtqUtcqQ+GwcTc
RapnGA3kRb27K+IFypw4J+DJHwGJ/sF+c8j2EjLcewh5YQOXupWcwQ8r8728MnypuLikFk+6lCfF
KVHXf+z86G0CPHFiY4n5/m+FBth8EYM1tA/bNavCiwTxauNueGDPjGOzteikc70oEEIAP7rO+ieq
iS7mfQOHuk7CIhdxpMjnX08XSdjdlXio35locm1Mz8PzJfYcdE5H4cswg6fjgZRxpOWTU1idr1aC
5nMlBjhNcUFPUJZFpZ1RiR68dIeIQbl60d3uwg4bzAJPZ22Oul4RwVVKfXn5q8WwaDoSd3ZD/BLn
2cjKrHlE0+M7Gfg5jGmQLhMwiVXAUHHLa/qMHfRlVHM8Q960MJ8S6tmLgJ+WUeygvbGeX1ThKIF8
+fMerGPQQBu0K+RgQc7/nb14LrvRVYqPmwBiEgUAJAvrI7FD0FsaFBExlrQkrdbALxeRgtWP5uEn
RJSE00QII3eB+d/aJkto1CK+x9Sx816SQxCHmlYHZ6mVO7TBwE6+BnflAjgLCh79GjKAynx5k2Pt
9NM+5xQM56hzv6U0OCyxz2IU1TD0Eq0CSIkGbmyn4R3GpqgmxtJap7ITaPmVuQE1/pTmhRs08PK5
mZrVPjwY0MFg0KYLoRtZAyUryNPlQYTdwzLAvb/TVb6Zae9TbBoVTBbLA8gzUuO7LSVJhxC590Sn
L/qNvm5AxGRSqU+nDhlaM/+L2AV7Ev3dmgccdip5A2OAMYH0zaypDy/L9NUCjgrLzHiqkZumFx3R
4vCQ6TTEMsfYsrktI1HKn3sh0+w5R/f2IRySieKHYBbHAEG8I1oaUxa5jwcISw0ZxrkzbCg0VdWG
VGhZ7YmRHm0jl71hzULWauAbf7v+eftAkAIrRxuJ7U5njxiuPo0HpZBIg9a2J+uc8676bfBGqn1w
cHoQ+gRJTvhtv6vLpF2Ba0ckA3aH7+XVqlWPMeK/pWsoIy11WyAFRBorPtw9zTHlWOtkPf/H1o8x
NXV6LalPxQuE/MqBvX6ThnW87JYh69Yl/2bQtsyhzy9b1ifrBEROsogyEFncpTwrD0PoNCpVdJbu
4hV28bLwcZpjUSzv2xpCTTstzWKzfy0cUq95xask4/dhQOVBsTyWqlxXxUaCI2kpjMxRajiGxISS
VX66fm0CzQFzhJaNfze0oBLmIwV3QPPzjy3r1s1lv9rmrIVL8nGtcl/sjBIHutnQ9ZE3t4rcQuKm
R6PLSTrz7rPWe7R967ZxC+Tuy0snz+g83M6M68ZdsAKHSkDpo0n1FVTNoILyMsk5wd/wpsBq7OOn
Hbc2+HtbccRejCiY8yYbxsFXSzvCV98GElLJkSDsD2EaYO+DZMZVu/YpvHR756kVKvbyANeI3aFB
FCcXT1VTYpfNx5S9l5UlLsMtmBtOGpujFWmvvKzihg7LsEjOw/eQWKEwYoG9JB6GmenYp+ZmzG2V
34E2DtaeNUqegBzlrM4ZfqnryNLxTbSKpW/GZ5y8dymYoPx2B5D9cGDVLLe7N4dBGYDWDYu3aI72
8fsrWlJBP5+312DmFBGGeG3oB3Cq+y2k/XYWKFEnEl0EbNLw2mkRNI1MBoXm/ls8z3WfrlCighQV
VPVgh1IstP4fGn6DbPMmc1BQkeCYNVMcsmOM5QP/Ya93NbgE78tzoEbsm8m3gGTgvkV58LXbwxos
eWuFECo9j3p+QMeWQE/8ACtfAv9Rcfoh4+xfm14zjqOCjrDkNwOCj49iSpYIL5RcBDh8ZC1X0xer
4KClxQBgS0pWooONXcCSVkvfHlcGMSEX//8eu9tXtYHaz9AHXWL4DYDHwdCwgQapzhWo6pqlSPF7
NXTc837uLzZI0JcCmUxv3NCW8z43zMlBWQNjGAHanmCzPV19NNghkiLjDF2aR7b6SLFcGv9ggYsW
7VUZpOInFsfQpIncwMGoRAAhwZw/hwtrW3IHhSmxKg8lkzn71VRB8ILdHdPiRura6QtOCExUCmke
7RjJJUK+mgqxfbqSJXqsEbOCKye36o3XrsCHVioPe6S7L64eWNVgSLw0fbTnbwuj0/LyNxsJqM0f
fnm0JrPfa/BiTG6u6GmuNvq94B9FyYy/o9Dzp/lgKB1gFlknZY+RhY+yb7emxnKmaKvqUPQpNXP6
No5orjI5UuXotvtvJLcB6G1rkW4+ejHob4N45aj5eV9c2Lq39aPB3IJaA2Jx1mIiyPw7yTawDKW0
Eb/QaloZPBYZEl49J7sl3kRvgkbl8K+UDBx+66c3dSccbzjojePqzsVQRBUdT+cMA8xJ8qJyeu/W
u/+YZr4JBlJAmeMm/kLeeFZo1hoRTUgXMuiqDDh8BRaeOShHfNh84L11Ce8V53LLDKiN6kqJ8ell
M3lgAUh57vqQBouY+GilkAFnWGyvoajBDcz5iKw7GrS2Txq+spDe/yvgfdWl/xIVNsyxAT903s44
ZfZSoF1+qVu4zTZD6lEvW2FT2i3tyxi+NnTjhw/YQipnrLcAw0snYz2+xM4HQTTi5nt3EC9Pycax
tqXI0kAH5pC17urYZfi0MhP1p2LobXhzi/KKNUyYShej1PcXVC8BTX/g6Tf/XA9imxyVxN0wpefX
VwDft6+weBOLwhMfqY8skCzsVByaiRQ+SffFYR9YKeIqzJV7J7x2SvzK/u/x6fL+7QkJZNcyELj+
6xp0z+SHZnrQJtgMtpsfXYfbCdg/0JTT1FQGgpduCo5NR/naytzAmsi0hy9nH5w92nWg+X8NjBN0
SjWNKo8nL/rchk7E/vzNudhXW9hupypKnq2GfJ1gn2K0xJwxIHOnqK8CvHIA5c87nETgjCwREGHQ
l5wn8DrCkauYee93OCBm/8SRp7ZXKIDoHtMqc2hPyG6zqTv5bSFY5geupsPDwxWqxJqI7oceqBwg
BcwHOGJlfJSWG1Oxtpu1BksJQX03JV2FioblxfsFoYiEd/Jj4RuOuZTwG9PC1nWUwpWjU5SYii0P
VZIEH3UbmCQnJJgDx56C3vAYjEEPjmKBBhp348eoNuP06JA0+y6meFdv1bgGYfkPAB1FjGPe6L7S
SA26PyAEwhqQstnyIfUdynEGm2J6ps6t9C4En4ljgFbyCTe1B/Gm2LpiMykxq6E1a32IXIdogXdi
zXJFe8YV1C6bM+kzfyTmfmhxTPLcX0hkUZ7bKjB2ZPQzR+mOHVIwYecMgPb7Z0MHDTiLPtxeme2o
uOKAAviod8+nQh++PMRrK6jtrTe5FaSCb954pF0474aOzBUyLuI9lqBkejSDJ3j/BlkTm/RU66aN
GFAMk85l5swsGapS7FqBK6T9u5BsKKOMAbny0fgS7WrGbm1LIOFH1JFCXSAb10v/Vfy+Vr+/k4OQ
FOlo4ATh1ERTprr8tfiyGq77EArr1UUItE/es2d16Ydl7j80ZNJBlzxEoPTgCO8H5wDIPeO64yCx
2rAYVsM5D02GyiE04Rky/LeSq65gfzHPK5kiCQWLQXAh6/A7zUuMKsjQ4hhvDWvLjKwKqUVdbobt
F6eXgN66tVNQwm3s21iURY5syX3f2Bx8L+lQBFfX79tDbiY5GmUtpJ2NB9frrRp2HVJSqxIGDBg0
RjvgBdqsuFznWSo4Q18ryKSmto8xCLXLNRsyezvofZVa1OzRJ64cC3cGnltHBlWtaQ9UPu4LIL81
4G83SuIJ/FqaPQ7LzGreg2SrZFhst1tRE5gxIJ+fN1fks17+/h4kl6S2zFth0E12ILjnsuxhKYyX
xS1koWNmvRI9TyiT9XXY4q6/gvkjOt6uzcNTSy8toMuSXVSZ7u9q3MRkUZs16qPmFFm/iXCp6NeQ
ju2NDF191gFThhR3c1s9IxyNUkDc6SWjDNcPDzxNSCERN02hxWOlilpqZigKfjNjtMf5yPQ6SW7e
FeiaJ60x2rsRkse2np6EQPu7ExqxDipEfKEUc2z4D+uQpGkIfS+D6McOmThcpuSujYqW0Gu7jH6z
Lg03iU7xD8KnlSe2REBJXuPuR3iutRpsoT56lHPmLceXMhgmFrlchrqp1YSMZRTt1xUSEodvK9Mi
7uD5XEU6E4Vf4og8K/hLwkHgzdY9Z97rWom62q52uBAUcVPD62uxx3TS5QG2+Qk+xBfUsKMJGJaq
DAOnmvcy9b38YPntbM3Iu2z9o8dsjhWDYED2ZpL04DMUNVL84pPeGxz03x7Q1ZDQbFIrMC5acQn7
L7IH4ZIMhKT5vgzGrD4oekEmDPkVyjy+rDlh7HsBun7U90oJGQjgQhjdLdXEahzTwYvQ5tYiSU44
9HyFTRiL4F4dFgD3NJtXuVSCHsYG+5i/ymLYKu6BBTEV9Zu6l2A9iPnBBrOxlahfBpxjJPbCGtLi
IABVStPPRP0juhs5uImqwdGh21t8utsNMn3eMO/geJbaIoltWBLZUWP4w0YV0UDJtbo3W2vMsBF1
dDqfA6l2xg096QuT+dV8+cMCP5hIsviXYXZkAN9dj/TFxD6K5UVDdanthBoYWmui+jQM9DJxQTJh
GVYorsO5FE2gg2XDH5Sw9F1V1kvfELugejj/dmBzOi+jtHvLxKMSBOymy97klZNFTh/WqUR9cEAP
euYlc8xgqKH3PamegfzetMyNrqsXeVsJTgAfbjVG9DKxtqUT0hX0vb2UIfW79aOjvDnInvHWiSIv
QUIrdpAoLSywTUkR5crvlRqX0mpB7JkvTPF3bWd3HFtOApcsZlBxkvFpygmQHLFwChjEptVLLJkw
j83r2pxUiC+uM3UmsgS+39bmO2IPrg59aJrHeIsSbgwasSNvcZOv4XiEgrHQGydqZyBV7I+exSmh
v8Yqr8MLjaCxjXx4GtTY23MgKez2o6/iR3WlQ8AO0uRGCnXua/bXwnkGrCcpAozscsz4bUL5XtTz
rtxgCntMgc18ypJuXglYQDPig9uN296RCS0DI3IeuBMU7xpsilNuxxqXbVP/H3u6pMXnkrlQKMx2
Yt8eiXp4ym1Av6LiJgcC+XZA/0vFGJvTgV6Q12zPA+EUYVyQy7aTqGH4m9S9ygehoNvkEMIun8iC
iO+xGrtZX4Szy0N7XdxOGSoyXtGNvTkyEDdRqpOWDUD4xMXsbFAoRv5QFCqHFVusEFze/GzmBHUC
nfS0UsY/QVn7ekFbhyK92I+fmPbQxZ/k/A0S/WxZdKrGjMnkAnjDKUUK79F98B3HOTgp0QfW3k+M
cjmszwQywQParNI15SjRJEwS4OfZR3d5LPF8QPfT14U0ZX41Sss25spoZ3vmXFeRCUbCeOAqgpb6
oICAjRVoNvVJUTre8V4xcEu00XT2Bsa7kOt3syjI7JPOPxC2eZ8VxK8U9l/rXarfuUVhpBEEWToE
OY2+uQOm9++ZcEAffMLKLWIz8+4p8EYOhwU+JpWMTXmhYhpSo8nbwaLZywfAvRYFIObOhge4fNA4
ycY/GhtnJL8w70yw6E56pQu0N8lUJmFrrI3/356jc3h8pBCZAnCcBlPIg8XkAaW/F76AAjEUnT/D
0+hWOESml2sjb67uY1Q8LrjQJqx8TBZYEw+hyukPFPdpJn+IhZm5jrtjV+Lr8vzI/H3C6f7AdSzO
emwfnzr8oPc2rfWvwqU0g4m2aDDvhdRB1Aywdctgu9AjCem861Pt2fl838kDADJEgktup3EBRWkA
fRy0ANKgXZ4rTjVpX5xU+TrLHavMPK9pj/P9VRprCqi5OOpdyqkyW3ymcRon46yjxH5gd1siS3Gv
Eqvf++/fZh3BkuKjmW/Xzf1UqPoqZmtovR6pSc3WXUKms/si0yhL/+yPnyFZs3TspyC4tCeKorOn
peFRwXKtc2fPa1hddQhl+CvFZWGtZYsmTNzikPi40WFPoMTwVnmvFspQJ0H2sNrE7pYJv9Xrarlc
cTBS+mwnX9IGxvfV4ApeAR4bapJz5Xy29TJUuHXSMy5zbluf6YGf+gr/eO7VRPXGgVOiL+/SFF8t
UtByx5yV+y8BZ2cfi5iy18nfDnQkE6K4Y2zFWhf/YTmC3gheYfcN83IMg9PfLhEKoa00Yxm7rUxI
tInIhFq7YrTlVX3pE3vAqZG9hWlp46mhYdpGr1BTIZ7OHMavoyGguCzFYSrUapn7PrKGYQfOLRRv
ONs78BGZyT0XHgntLzGiTjueWp5zjEjaJ/es3E5J+DQKWiNvCBk+rrHEynMsNmwvMqdHnBqdhwZD
45WNWlu1qbR0LJ8swxAWd39BISR0VYFUA1Sc5s08LL00RGvtC9FqEgB9gWlmLRu8dU0w97wbsoEO
SIyvfChd9WdgK5VyZX+P/wAg81YDyKgtIDZFasTfw1MrWeI/tOIKSwYtdyS6/FDycwlg7WHopHR1
UuOybxii2XHyOq8wFtKFxLteubFAz+db1OekbwVGjD09Q9o1673STQVMiGOjsjRos9BrkQrkYtCJ
vUeYzJ5auOQkyGaFbkufaf7AD4gxaTlA1h7EdElQ4272Ip4rTOoIVlf9Lon9JoX3krOn3CqzcK6N
ujbpIQsU8PcTXZdKDht7RYKLihK+viGlrZV9ymUBfG3qaXZHtND52TwCQuPD2K6964/8jcT5uy8N
y98LTFKduGjocevG2azvXnKybhXdbwpkS3a96tQr+qNf6ujNKu5iToJhQ3qKY1UjwAAyI7+l39ma
KU1bU794BMPX29LrbsMZARnaDZZMk36iXjjAMjReLB3mrCa99pASllNAKBjNyi+J31YcDizm9HBW
XVQjwDoui7d2CnCPGL5S+QYEuHNYBwEaCcvPycHe4TnQmRCo19hLLhncMzAtH4lZD2hsA5Vc8eOY
0ZLzDw9jBx7rNL1CF3uz4wjDrZC8l42HQK+ViOqFFilsszw8bJpLzlLjStByXNKZZgslgfxWmnxI
4Y3MyR9CXsL3E4kb7Y8pZa4kziM481xakDR104oTQsZ0yyAHtfmbDWsiX3aaTF7G8ijBGycnE9Wn
mHmubaEDCIXVyCbs7zpQZnKovBAl14BRmvjqm1PC1pl9/hJQ4pLfenjTwxjF9C6KZQ3dOlcqvhv9
AAFQAUuJnCjcz4fLZiH7g+A59zMjDxMeGhQzM8i6XLJPq8c4G+gE5i4sQdV3MUjK1L0wivslG+FD
uQzQqgaUiMa+uwpkzI6kIPwGJrCF0qUOvQF8DG9erfiqrm+em6duXp3nacPb5rBK9lrzzzNtXGAs
DIKHi4k0e4BtiAxxDa/ZJx9oKL6geh2GhhrQWP7/wtRMaFmBNRtpWEExrRVCYmq2maUtHfRU9eOC
5bNYs1Mv1XR26wT+k7kcW7L6DrQrWT+N/JoYv4tCRKm7+4zfCU9AAuSKR+XoRdNzcGaGKv51g7WW
ISlCft8DbbU1+W2LkiERcNsfJaVA82fnQK1/hKiVvrUQJjNYqsTmmGFYH1HPX+wb1SolNVa6OREL
TBeQRVxlJhEFrLqAC8CVB2peteQ1uBa9OJKLPNCXLfri+XAhKyfcAIdsImyzFe9xLnHZS/JCVLFs
o1yhIBwzoUuIOyyDOKx+r3fe44YZmXsxQOh9B1PeXWVrskQFuOD1dizDCyhKwlEbV9qeF/ClaRq3
2mjp8UKG8gvzuFHTzlacBeTuqh34+xVFtu8VuSnsCnawXKPkq8ldRP8PVNSF9RHpUxu6RTZ0rycS
Loougey9J7cO7/MLDeH3T21Adr774vY5dbkottwTRFhRa2F2xCYswavye9OD1DvuHn0DJ7nRzCDK
jzAZK5NpCZmquTO59fSyuQEhuW5Zgim8uanDf9hhwPndcg0VFnWOeEjDvzmmnJdLcQBebZlPlz77
GIKS59nOYNAMxUv/Ns6AjyMZDDpA41FoV13X/7/SFfrzVqElTuYTJ8mpX88MDm6zaFUdj46PfD0b
e3dxvYXLvFcd2GK4rJ2xj1DZEhYt3MWfpFxPWqQ9odXuptzbkm5cW1u++qbQUb5S6aA75JhiJx5p
kbNMW2Pe/b5bXBwEunqivosuSM1SEW4of0Od3UwUNt81/UGRKEN/7JjiIzxV8cfpNYcMqzSCsIHb
Q2yAumRBPXPQGeJA4fuZz3jwgm5qxQZ0QcAP99gdE0hqy2wAYOOTE7InNxBDqfVF8ONDcLpYZPnH
nIhDkvzPZS1xvnhgFVQ1jjEJX964MG3cWoUK+V0Tb7u23/FoAPahoz2gT305fVq1VWtQ/ciHB5fe
O4+BLqXNanfMl4jfFMZXmttae3nJbGX/mcZgBG7xZSR24DEh9s6KzRV2dhuopR1WRMTYkqGHyiSe
0heWjL9/WQ0vScIojbSfxOPikVcDJq2xuxTHTmaYg53/BK3UGXjETcZt8x4865pYTWYGUXTO9gxO
Vmvrcy8+SxbD3HRpq11P32rmrYdyspVGn9DeN7t5gVlIU5nWZfqGtM+PnHi6SGuU+W6RRs0WnPX/
tqiQIhdQkzG7nxVti4rVYW8Gkv3J6WlPkz7xHdQZAHzzS15kUfC7k5E663DvXCcNZOMbB285Mdb1
pvrm8gK4OiExZXGZDX4p6YViA94ht9nr8ueZhOE9aXiTDrtLNyN6RtkBINmxUB64gddLBlK7hPd3
CZBt1NmjQEViQ8BD9dAM5btkzUgbwMAap0bh6PYllXS2jWPVCLkAIUvyst/wRrcRAeMNGyoz8Ch/
at9DavRwiA/d/cdFiuedL6RATpOEZQYr7on6Mvq+UB2FrWv21jv/88WaeYt8qXP0pXXA/DqTFcCW
8cnYpnkbFDO2XNKYUIlexnSq9Gh8dNAuPaeb3iNs6iYU6s0hGgpmvbbjty5Cz2J0OKfppYaerHKa
tJA9fOd15N2ThgRNU6gmuxVx+u/29cKXcWEhQ3kJPCxsW/mzQvgptPedIyOsD3UAcWyO91TsnXea
345aGCqn6ZM2YY/RRhS+Lo9RPOExWBT9PUIqjOSMpszsEzGRblAnqz4ea4rH22GAnW4f1IfbkXab
VkNF1vRVPb5/tjbyBM3ZQHvSCctUE2poADc5v45789p9eKcKImCpQrMwLgmEH8quEEQdscPQqJhM
+PDFrqIHpiV8TIgmyxLvjbZIfGt4+KIdmozsybYW4q7+C0cTHiM+Sn4846AMo1x+eNeP1EKv+iG7
YATJ1c9X6RNVaM1FgOg60EMJezKkmNUr8MQ70O9PfS8r6tFttD7quVJ9ro+3qlTfF2S8L4C98Ng8
dCKEOi3toNVjKS9IJXE6b3TrAMLZX+eCYGFHLvD6A13cMsX1pzTkhGBe0YPF8te0D6432JVL3d9r
W7P+3dcV+eRgwHjCENRbLzmFZGJ+H1Wgsww23o8fzQeGflxrCt7dfUdQTtFYEVK72GZVkGYfdvjm
D/cDRrWdEUrJlX+pusCo2uUSJfqHUuqjb+SiqSqfTkgzF5u6f0YvR5dswBgphDo800HdaCpOFY95
F8blk2lcWAmrm84r9HH0mY460mrD1z8fFDYf4+JSx1tlEJ+/O3uiUpL2NUtOxxTMJenKtasoZMHQ
orST0ecRsV4lyLywJgnYuDIOQpbbFi0hJDdSPMEHVdMkv8YocgUiuqnWQ9KIq2Xtc369lH94HuKR
rSIDCk7gwnjv4tTvnIUsquUcnRJqDaxtZHGHvitxjq8NVsIzxy8dkccadiScClWLGvRLK0Fq4w/Y
Qga1MwT1pFK6ZcZkRTkB8yb6mOenPvBLcAIrqVSmqoyFiQoSVf/QERXdINHi72J3jFdMOUFdxXJ9
nm6cpNYU4SWU9q0uKz1xW7dVEoJvrIiymG8zNWFBePuWrbmBD6wbDftWV845FHfACXPpVgxv7dg4
lJ5VmxI932sjsPjEI7KvpdQHrWWSGbdrg9+Kmus2yyjp13axzlFMUhxruwxNwpaJyYcRmCSMVGXZ
T4X3aPVBrTI0aD4TxjYnNVmhSk2ad1+1Y6Ql4Q2HvVswxOtoDo+hr1zh8Vk9t0yBALpDEPJz2ADU
FNeaQFTQ65QLwzc5gdCDDpA4AGVieMaRChc8iP4w7qIbtti3EXg7T+kA+u/MQVvCZkrddcgYhYdB
J+ooKE0WIDikHVnGwv1uIna48XGiE8iJM5O8o4cu90SHfYIMSTaqWM7X57OgMnmJeI7WmBm7C0HF
GX8QhE+9qutnN1XADtiCruAWx/jQGxz7hZZEPgEYocERQCvabQRon9BCx3WxVX9iyIxrK6RV8D0x
PF+ueUk7bSCkt1Fostgg5QtPtEB1IsO6v2g6UTbvqK+8lkb80yVJfXmysbE8vrGBt4HaIfZCkmDm
Q76lE6CqP0l+JyX5L8G0+H5U8NHXrgwhKHc2meL3BZQeWvckl8csiu1TTYeHMaBRVEi1xcyKR1Ht
2xxXY+Bje4TE4E8gspjJyQrukTEFTIuVlypadTE1r4fm1s/ui/zSIodVkGaKUudhU2yVT4uqxaXT
IF/LR710vBM/HillOeuK7FkbmZYgggKIQV3p6+H4inCj6TeDScaOdc3BS2GqKTUGZ1r6QuEd5yM9
hKL0/btIq+TWKGdPxeB8BIakAUPxHIWiqC86JYibtKNzifvdmv0J7YmMzzJyHGP6pJAX3/1luMZ2
+O3P9vbITe5EfUZ8MWeJTPjEcsm0iR+FuCFGYXUBCtj/BEe6hjskL6jjQ7Xk/o54DxjT1OHJMsJ0
Tia0np4ueq59fd2jdbefNEtH4b8qrEO3wNnI+MeKm8eGSkRZXVbiIrR74/YWvweYezQsqdqslpLJ
Q0IlTWEGjkAeCx7QfR6lRHv0i49DtuP4XUHN75hsDTTsYhTAfV2+mzM7S7WjpeF2AXwWKAElk1i/
RcIY0rzTue3SZKkyS8NDZ71oca99MI29b9PwdH95k3NQFlhCaNWNeHgFRMYBYjusDk2M2seRSuVZ
QxkkwOMOITQ92+Z6qAPZZBTlxX5bQphiSvq/RFJttFvPxpcBUTV7/qDgB2B/RDUS9RS5LZI4y0p1
Xwp4MOjsoBQ4M7OOgCVQxtde14FjU0yz8m2COQjegMOhoEzAig+4E84R3nrkWgJQbvdaOK1pk133
iVKV/sOCqdPPeHd5rWDX62NlOpP7DYRFHgDn52YzhMMxXaGRrZUXGuTjyBfANm1tsdNbr03X8fU0
eKHegvPTZipFa6vdFkLgn/T0zE4gZyyZCg5cgF8b26ssVDOW37cFxaZa20tx13l1Nwm2yF+6uWrt
gtUJfriN1HqQrtUIpPuQBEjHzPk++uO5RNmvb8KXgJZRLcRvsYVt6VxexEePMpwm4EyWd29fbC1O
3UbqWOfBM6rRg8gKq7Urt/m3kvawABPnH/puH/X8wAemXk7NXfFrXopMsnqY7dYYAeUhS+ASXFm3
3siFBiQIT2djpAJDAnlzXH5QbuQxdenH8mwTE9Pk9Kby8UbP+tavhpwMCFU0B47E1lTmJi5X3syh
Jy/SXenrQNvQgwBuT63/gFkeT2dLkNbLfpiZzHZD6yhOl0SJ2FK7qG6keBRzr5JsQMJxKOtl2SO+
Yt2iI49H9PAgxNeUwKQQm1Qnl8C+LeLr3wM2tfv6gPHS3yvhgQA/OVxU9i8fNyJsVWpEWs09JjRW
WyINFJfgTTHX7gIpcMZdefxBiC7q/rTYd9Q+tijtfuHR62c4LoPns0yghQU6NF5UXYscudiDatm/
oepmpEngt4dMverg8X8THvcjiFoyRzLwqySbYcpF5U5V6OyU8x2RqAApBhTRb7e4cJF9k3bCeGfv
qvevQwHFEppP1W12T6NkshQCHZGrHmqgDIzM5c7z+iiS6ouWgb5Uzmpg3B1yt0HZ9lfwHxD+gzmd
R73DF0vN5R2iL9mpcDnqnfJ1eKMDet5I2XSz1iK9tHzuBCtdl/tC0z/4cwcz/EzJJ5354clxGRCj
z52Hex0UEzCwW6jlebj/CPJCHQ49jqlJWWjY9QirFnGggTmE3pMqtWxupvzptISNuMr+eVgxEqhE
LzsYgIfBenH4qmcFRhhEZhqpoeIZn30v1Db5VvXRvGwW17AqyOB4YzJfSL27BwOJNwj90rFVtYnr
bdN9hXyLwovitUEy91mPTzcDV0Pj43onGq//dHI2G1hGk8CaMdo5TJJ9237vZEATHyWmW+f0Ehcy
QeAFcoNxwtV1dDl8a1eyqsTftk2W1x3HR/ZqgL59sH/7kG+d+/6wq4KX9BBpcTAaCGLQ9DEMlbul
pTQafK1OWB6zb/W6L41C2+3bguot0QoSwx4c+iRjY/cKzmpuVTiPzj5ETt8J62WXIqdZ6MlPKQ5L
jbtzzEbDA8raKpGfA5mhwyMtGwVYWqwSUj/XZOqQ85HcQqCeHwjTW+mojcm6bYIMlUikfaseWy37
itMyai1GzPlFh+VxHvZVysodHw4xGoaKAJzn3Z0Z46ZrTQwj0eLLgWvwl10NKbdGvuPmf1v5LBFp
+9WnxGIQ9EkGsfn0OAu/4ycs1qxeCsj5nodEY2QfrodtDDXJY8otop7m78fk2hn9CbyIqNPVtGd2
6JpBWfkX9vLXeHUluhb/jMmACagEX28FtW493NWvhLUTn9jnE9kxMQQXKAioDIFPu6XThPFyQIlQ
RrqOFazmr8M18ggS3dDcVMkXAfYvbthGKb8Wvo0CeFx4OtlX7V0iKG0QdCg7uprOSaOGKU/Hviku
4Qi02Zk3q+Skvrbdl2b79STRzcuW3GEDL9HZv1MTZTnFpdjriOb5M6IwqDCIsAJeb5UXot/G2BDG
Cm/v+vvTUyuaidIGvHI+t5GxhjpS9Fqcow1J9NCqKly5PDAfZmt/ZWBKR4/WzF2g441S1qmNztVc
wLXdF7NpaCi2YeKKKqxuIedt2OIbK0usspJCDUYeeGiFxDPa9ojSAabbfOQvyrVQuaKwl0KKbZ9c
9JyZIvmGBf0ja9sCUe7WYjN1f9BhS35lCz920hOTSloNhXAdEgnhfj0X2kZNaKjxwmEY3coDgxF2
q4pkVBsBXpUUbvB5djx7If6ToLLpHDnjxaj4WhWty0+SYYwOgodo6mtB0Ufv9q7g08GHN632VzPx
KHL9N/kza+vO6d/yOpBVPcokqhS/ZVkg9vT3U2BCbknSyvi61BMSerdSoaMQtVblkDZq7gaAUqws
tP8jIPScTMZ0nhlPSsgBkazpbjSPNY86RSENfdUagSVxFolm+O3nvGvbdOJpaFVJNH7NbHQv2luW
7FMm0oT09g+FSIBXTpO7M5x8XCtmm8q3r9U8j+j7kLk5ArgunfKDWFaqSm+B0LEAHyOaKdf3LHK7
dIpi1s0lXiOWZB+ASUarHGDi9jJTa+w2qmTYwQCez6r4vzD6G0bZNYN5lOfFaE4Mpm5pKPnR+umi
BFjyJNNdHh/B4RrKERjUR/AHLdWUeWYXOpQuEcNWoq/T9KeCJewWyfeBBiCI3mcTr2UsMs64nmbf
bJWZEuljyJzJzH3LDaGMAlywerCzpN88Omq95VHX7xcEgiR4hA2fOPVCqBxZCIyIqMYUpbWy4VIb
+Nx25WM5gDSFUHmq6hUm77CxX22hob2kbfUVd1dMq2+BBovpruIhfqlCR4JARqUaQYV2Zmeqx1C1
tSN0gM+f77aDssTHRXqtmesjIyQKh7ZAJZpJ2/6KDdCpL9FZbJhy9HBJRx0OpTTeMN3TQE/hXprK
wbFWYxpPVKFxXs76ALirwzAWhOm9KY9HpP8G3jTuLVa0rVIDh2NOvYV8RKYUYFtqcbwtoNKC8shd
Wxy5vsgzi4xmsZxN51+Mz8t13ABkNUDjKRrjyATqfx6fbjcqiHhV7TG2MAXBcaZDPEL25HM1+LGm
TNPCoYbibo2H7+xft1Iq9QqyiPQKYLeurmRL8Lp/GGhfYr9gttAS0J+fGUJsTDgpmN4SqBq5hKlr
l9ydYcI4klfCHssLXC3rqxJo8zucxR3B3in9aReoCNqt9xsw+uJDkhlNhKAZKnI+nmDrSgYFTwYI
VFMka/z46NUPqABOG7P16ODwsvQ0Kj7xXtZuyS3WbmhPBW41tDDQWcTmPfP7b85HWMEM5GcYvYI1
DibB0cKhfvRXsUdJx/cuy1dZldnYJXI3sc1W7WycpNhiYfjmwpJtL37B+5AYytRZTwQJV6PYb44j
CYlQselhIP18lnYMhq+wp08tEw3sJCIDkUt+J67JWI1ZZVv0kV8Sd8ymBqzo4nnWOs6ge2V9O3YQ
B82JVXee7k/7+3ZaS+DnyT0dPI89sHR5TXvS4fQ7sH/TWe745X6T/EJnWRIRJDusP9QrLVyV0+Z9
dX3XN9qPO4t6SWvYDosVcidfamZPY+MkwczeBC6pRs6L+YbGKwfLTkirJ2zwJ0sRODeOJ44ahZ7j
dElKJDr0KQMMQD72jixMLIfPF48uEYcVQOJaYx2dCN32Bi73oZaQFQEUJVv1wsdLvy5atNM1urzt
7UL87DofPAJrv2E2wg0pheiDzetuBair+qMO2I0Q2ifHwJo35QD/+TWcDoBPc3gMo2s1zJjPWFbO
ao2HUUH4JhYF/bdSwb92ozgtLxiq7u+KPpdoFY+w/p3BRMvRq8+UZSa9hzC3WjZ0AdwQxbSsTMJB
62klsa2ULBMa3ZYM0xtqqy3oDFCnJyjZzmBfWroNz48LuFBj2F8ZfkYaZSfEp9kUGcdF/+I9ar7k
Ysek7IHO+Qe3R/bInya/D6HO7xPU67z2VyVV70A0nXKF3bWISDNI/XmKO8y2TYqYP8GBgMStJZO0
9d1CPw4jso0fomv1jjKERB6aWuX36BNRqPvMJQKysl0v/c7ZpnG9XN2zTSkaylQSO3ZUQixyPytA
wP3M7a0UrWjmEmpPkAK116WqrHeuzdQ50+gky0MFZXsdtbAJJ8ks4842NBQoknQiK8QtJr7yQwqh
hpbvoeJSpWW9GDkfjsoY/iff4ZYqGOWq1Fcwzh7XKuSVWNNe4hqu5C6N3tfutKdgufYpFFtRrvpa
M5wij9ltjy2Vm+Fxr8UUX4rhoMugVlfvIdsWbS0b095gkDsQkNM51aiJEE1dacqPoYwA6p9I3n/i
4hWPDCdo4VUstii4D9vxrhdDjPiBpujN5Z32Sy7sa5H31Z7zLVC/OwZERU+pGM83KtyhGz+VCPGF
tLwkT0I1hk8sPUYpHEkrsed3Evd+1U1DQyIyanpa0x71OhEU8Y+hVYAXN+yBdVjGZJeeJpQXXEhS
hA6v4SUKXY7sa0A4caDj3b+QXA546rczRxr2XySIzfxqzpQ1j/9PS4SKPeV/9UdiCMZr7VoIpUzG
nLpvYghal/6cJ2gC8ezMdk8lmPctuu454OAs17e+YTNhwUhYtO4kuRX1aaeO4tYSkhfEkPGP1Tg5
cdLUcDYdEtQ/io9C+bQ4JL8BjCdv15xb0dl4iG7ydxgdJFrBQSZS2vHpmZDFKWyjKytyO3dkUSmB
Dsk73o1g1E7FcVBsRRBXd+5D9UbY79l2wAZat7ig83iA3HuEPBhR20y33LyxbsotJutGg/3hER/7
Uew0w2EJSUpM6FpsKDJK6ypOKuZWQSqLYA2hISxhYADX/SGVltdRYehioe2QBCwCMmJjaUh+oRhe
TEjqr3NlnTPZl0zB/QppIWbFatOFCVURURFeHV9hxlbl+dX+fwov1PGC1JX9PYIFpmnducKL43+k
pnNceoR3skvUuC+wxIiAvgLfW3AqrtuahGz/H10ehMPy+gtyFVZ5PBcwKkZoET/+QRGb0Kr7cCZw
b09iYoJspvhGnCUGMuhZ6O3N66mvhCJoU3VUBcx5kNHCmOV6qFKDBfL7RPRkaYzgDMPTGwABMmW0
X8VrUrCRaKBWkmi4PDNjIF/v7t7uuMIp6kQ9PV+8UPoGJnjtZz7MXDsVuqjpsbax09bNUAfvRUnE
YlUmt63nhXH/lJEdS9psg5elvchwYuVvqxYVgYD9Rl9IlhJ3Ow+AR188EYEa8nLcMeg9PfLa4HMI
n2sCEAsC/Rb11/QPf2hazuXuIzEamPsd/XlFV+2StMMnkb2iFsFvz1FQZX+r8FZYG1xQuP9G8Gz3
p1gGa14r9ad1hz8ltLY8K4rYh2jGEEzjxCbA0WNwrmM/0BJ0QsEgq7wyaL3+vre0YQmu+IuTIkuT
9TyOdwMxqWTAH5pebdTffvThyZPHv0EF0TcTWmyMG1bK61Bs36RqUYmNiawNIxn+2bXHXgukBWd9
gkquJ8IK/0WU9/HOcpBTvEwaxSFajJcm1bhZjWsuIm7rm7musy7q3ho3dcncKj7wRDuVDvxv8ze/
4FzzzfN9XI9lSDwGRM8sFk50XD0uSMvAwzFsht32NaPaereuhc4myWLiXT2ce2BomWQ5/oz0OEAP
C/spX6ugtdVE6/WrmWhoBjS7XvAHSCf30QmQicuQSFNQgV9gx1Diwsim4Bbef2YaRaxEhOIwanYl
u2n9DgesMlDrHbeaAfimsYwhwAHKXIvLXb1wmFBaP2NjK3Vcq+lQnIBx8kBPbdzBr0LRJ5+7GeG5
ZWKrBK3Vg11UE0Cc3qIUhtqFNEvQqx7KOk7dmMjBmwytzImernXzAh/OxYgeGm3EL/QSo1vh5Q7U
n29ZsKjAq769RPRfSkDJKfzDFm8/u5rHjtnwz6hnAxMIshaU3lFrcZWfZPfdqgLzrJN3WTT/7WDP
sPScl00/Rfp6yNMhoJm+wVqCcTIfmDRwRWdCkM/57zjXjIRBIC/BRd6NzJJ+T6BWjhYL5nVTWvHk
uZpMgoI4WEINP7DuyXijZF7Hj3a4oKJFjSc4BYHQrnI5hzBFGXasUrT0O+Y9GdtN3QCFFkDrf7hw
+tZV2NA60Zhg45N6cxmW0Abx1rNVYq8RTwY0WVyPnuGVnflEURDWimPli9mRMzg6emSdzCHlIqpf
R/QBYtfzs/y+835zT6Yyjh3NQ4l8ljAk527UNA698yes4wCX2LCwgopZZYvDA4VWED1MStyveyld
NTISTAqG+VtmoIo1fDsqYUrod/AQFr9oBJDC3bW4o7zIM+RsQkg5HCI1lQnWzqyoFIh5lu90vQCb
dDuR+yO7XTIACy6e3Sov2/Tgn2qXzAwyjjYVufD8IqaCBLo6OYCMGNiEaPtl9w5LqZluohTB5oO5
7FrwnQiNQD4fJRqivcGDkNCkdICDziOSiNAUUOhbY/pjJMtHlGbBm6717oC0KZFrE76NrR6NwbRR
pfIAsQpgMQYTnQwvzVfDNgFafZGmvpq4Zt/G7ma8+3QkRF3pNVxRp61M7id4XmzPRLS8zC1Kalrk
QJ+4HI4v1Yj3Ww8OpdzV89fZUegOvjOckCmZXwLMzSp8J7noxDKWSoLUbSEjJvMdctOZp/YkMPJ0
tJ0b2ZnwtTPBL6eBTAyhjFy7e9oqO164X7BQzxeZnx6mveH06Baqa2LC//mrum0af06uJomUSe/t
a6gV+oe6Dk22x/rw4edga9oEQ7hSsnO51MT/36LXpAqUvn1Whnv8fSeFUNGbmFmDuYvqGWDFSDb5
F6t69ltExYbP+fGPTOysrCUXBvKXiAiY7HgKLPZvNWOpuotbJjOp0pn6CJMuJwW64bWy5FgVmvfM
SDxnlJQ+yxi0/LCs4cBTjfxU10IZtfVX1t4Divr/B/U1C/rzGUPaUlKi5uDaACziZ4L3BXKPyEjS
aoxawQj/t/j4NxCJ24ZOraQNPBKrrIlAJE+QP8fkNESvdl1huxBmqq3mr1Sz6rJFEiudM3zAGN4G
vGuGDmfEZphZX9UtcdGKolugXIbQmbkBcExIc1hPN+xgIIelMKB4ercWH7hjE+Tw1DH4osh9hgeO
qjX/i4aP4ogHn7ALPgCMkAcnQsMD7ryfSKF8CiJE1rwYdH9wgRvSj2ss4oHpTy/1Zz5jNbv1vy/s
BC7DKDXsNjER91qDxKAViRPcttHHWOzy9pYmax9/tK7PxQ4HA0eqPqXwPQXT1imc73pEZpdDgMsM
yntnArEy9xXLW3nLllrxcVR5LmWcQ4uWVVhjIgCOcuTKMfdmbcJQDKAGIniw6na/oxvav3lrER/A
/n05CpcMIKVDMoBY6UfJrXzFGOdpy0Y2y1h+EL2mXemysOqAiKm8L2eyjTRjZGoRioYvK1ZsuYPa
Fbb7Mwx0fdIF+sYuexv+goo5HC6shymfs8Sbk/nWAI8jeJqsDk8xMFSkrSvWMDVGjCvXO1XxD/Qq
ZRcBJOtH2UtSXZhF0lf8WtMuMTJMBj80FH3PWeU9fGWpKuXWtygRYOSOklw2JHRB8gUgKzl5H5LJ
JgPodtkPwd7dWH9VluixrZKFg/VXSyWC3w+ebqWBJyKwghDaKz3OLR6b96pgkXWr6afYcN7dLnGO
RAodJATcWaY0FdLxkxf4xWZGJTZiijTjnuwjLtYi1bWemhL4BwTs+HkYpNC0oxrCyWs3Y9VqW11F
ToXnxq8t5+lmAiL8mWK6p1HyLt4V3/vaUp749T0uow9b5eV3EVDXhnA7ZBcJwfJVLubg10fbmGwj
j3n6NrsgM952ijNcsXLJHCXclgdVYxkqIjNUUUZfIXAejrJ2BsIIY4ez+m5UU0ORZUPXIcvm4AEg
AOCXxh9LSeUzWLZgA0TnLxDObQKjZ9fVkplu1vxXDuz68wuTaJYlXK0HU1RYKkrxbLZbG1Gpi0W9
NJELPWbNZ0AEpKvA+v+BXbCil9quWN8BZ93+GoUgGUOWs87CLwJQl/8VtSqKbN+B6LSTCM0s1TUJ
KglheSXao1D68iI/T/i6Rdg1eJ+zMvz/tpK8q9P7kPOB37sZJioSio5LTW9/GVRH9zqHIY320J5v
HvU4yOfoeklQy5OYVLJeljjycLuvErkDNZRLeOCfyEae8hjrmhv4E6NJciZHV3LuIC3tJTWXBs4S
kVPvn6zgaPUFfhsF+CwdcIln/UsGhEIlDAPTnLbdVM78bNs8BHEMMTBi9vL2B5gHLfWE6w77t3+c
2qWJEBNKWCdcnwRQHC8Cg5NKc5nCZRjHGM23yfUvj4mk4TryLDScrhCr6oscdH9Qofa6ZMuVAYNP
a2consLDqvOZc4fpgrlnb42HBFJj/EJw2POkzIGrA15t1m/ZmWCFD515JV+ibM/SMbAV2fC6pQx9
XaTPuBbYcKIhwRx8kIyg+WwQoNR85RIAJ3R7++WxzlYArcOkAG0GGJcCtPDpc0TCUk5YOkTtniM1
K6Q8Cu/dWAQAZ11lK7ZKqjr4eiOZU+9LaS0fiTQMrL6tHrzoj9/9AwnYSpFBIX9Irgp4M3USCmPw
osN6fNfMwn8ge4V+6glLLQLFJGQVbPiNvgxxs5g3k9gzPphbF6Ib55Op5FRvtFBVrvI5OMB2SC1y
4R2NYnt5FaES8KGXlOQ50wb2XdpHgwltk2wFVAoSX51dKXhyHpifub6hjBzuNkVESZCb9L+cu9Jr
KF/vQb1fBJtsW9nTJ6T1scODWGqu2gW8th4HfLs3RUNMsRbPaqxIxls617/fgRkJvpDt2KODiVh8
YIsM7KEFWQn6nYZIbmIIbw/WyXkBX7ncTa8x2mAy4QGkDxf4nmnDtSFAOAJYpoNalrgQX0sJtHH7
EnV7cAjyVLSJxJA/WgwIAn9y6y8RpL5rMIvDWUTa8QsUNPdkpG2vy7lssU4FXdZP2uWQlfGVRGjZ
bHe1boWU7aFiV6fIGs/uPGWsLuCZp3GZ79lQCcZdAFPXWd+K4IRSYM4sKXk/cjInqlfLQPOe7uEZ
Q6lkdMcGtrXaoApT3UNHoP21Ih4n7ICq6SVmffJR4YcIFDyZ2UiQl4XnphpGrSNvAHonhn7HwDHC
/HQ2ytm55tYRD+Hzm6q9AnQktQnbANoiDtX9KjMB7S8fN9DkUKTaqRKfredtLrDrTuaIRUsAw2va
Y7aVtPdlE2UVVWtdo5HhR87hdkMJNCM6nITNa5y+hGfeqXJ1u2StAkxoBoN5KcCwU6mKfpSpflLk
an4etEKsVSP6StY56JpgyvsqjVTUtPnJ4lQ8RVhHHD9OiHvG+tmlvNAeh8k5OqZ9GsCZBQmqklQ9
K4hRUSt7wHbwLF+Oi7YLLnkc4Zzdc5kpA35KYYf4MuVdRlRvhWS0vO7dH3l/EkrzdVP/lrVRhgiK
QaABRGanwlgwow/5QhsL8jlQYsfGfDd1JOF2DvqVlWAJMePYm0Bu9rd978wv2jPx9NnyKC1XpkmU
gCa6PnkrLdc/Ghl8TU+nTnJq2CLskdcrIfXiG2tLbeh7U4Yql3ADG1zpc25RCt/lHqKCl2WRphdt
ABxtEDdfXrxvG/bchtfn+/aGQ5OcL1uA/bxr0XGwWBRMITIL0YZApHGIOhDcsMOVlMlwcLCG4t+3
oCJkmMirkz6TUkqpdkDPTzGzTuukuwlhDkHk4tAr64q+KB7a4s7xEAamRbpJViVGR4EtAytGC/C2
HMveJy8o4m7HWHQymlTjHbq2nM+khC5r9EHULLJPuXEoXYnhaWKU0qqPN+ISGg/pNqju1P3h8E7m
nNRVvyC3Fi5lTqFNge3LGNPCJossjIvO0h+pFXbuKm1xmOy0oervb8wLYgCfLehNuF/p4Tqma3N+
0hx0XUrLoEgimoVu47IbTh8mvA6Cq4YLgQuLSRv+aC3d27C4EmJFgjvysIo5tW83VDAuUrlyk/De
rrKgL8BuQLarD5Ge6rrD3TjfQZh+7NDT9eQi93geIHsadHgNjTelr5xenyI8N8i7BQ/8uPDNADq3
J+B/o8piPGtx5Rly2nD62TI9o5LF8ONEvd08z8BVAwD6mb2d6rq6UCiRrsc+i+7QiZDzxXRJDv6X
RmKSILHquHRGguiWzeAPGwu0SMO4GsSjwiAlbBG+kozvYJP1aDkx2B2SUifKQ8lA0DLI+yH8DWd3
lWPEOYVNuF2fiaKR8iDEgskx6CBXl3WTbhMEM38oC+0nSxa7uLMK0vxOtHz+r9SavU4VL7Rns+Xl
aWGxZL13Ymew3XB+GmOP8L6aGO8bMelc1N8ASO4FlYHDHB5sTUWgApcXBUvO3sc2UNLZqVxl4vPo
GPQl+7DIzha2hPOUfKJFu6Ci2TKwafVib2h8ZegPkGUZ1LKAHrcvgNurZWt7svra/M+qBI+xpMRq
Sor1BH7i1FPq5VmRZyDvQ39sLWryHueTPwp0h/DTV0k17Y1b1ExBK7ISWQLGJrgtKbhjJYT/kiKb
pfJR2XEsN0nTmbYk3U1EseN7me6wiMvgkvnDUgV7v1Zsk3TBcY2zapmk7mVRIil1gimiDLKAeRgo
Zs6FdcqDTEkO3um69IKk1klahcjKzTWIfPAknntLRnWts9xoh/V60obznq7WObWuVAKLLZQ17FSS
JHSSUgJ4H5bAo+n9/Dv2gW/7BVklb9s44WBADJeUg/gNhpDHkgBeHArF0GbPg3CjQIMy64xWIz4Y
XxJswQsbmljSiIA552K017LvcKYBAVGoW8+D5GrRHiY8z8fHDEpB8IwYjxx+KTNXpmaIOFVg4xto
0Eduh2ysL35QCuI7rYJYO3q93vRib98K9FxxK+ZPciyhwQ+THFHFCdgFS1Qzc5wEIrRqvfbYSypP
VwNfBaD+7aE4fQzag3DrpKlgnSHj0kgWJumRdN5kUlVsg4vi+SrXOIy8aRHC9NPLzEWUqHhPIclu
nsm438rRZA1ZL6m6Ya0tHtJMyUTkLx+kWZJGaxTqwSW5is4sB/OuUlXv5BI7PQ3chZ6T/m+V0ndf
PM5fsun7Xbus6R610rZ3pgXnn+XPKKe24/h2mq7ovhQpRdAYD7KFREoYstJKXw9qxCNSR3M5y+Qq
7dgU5dY48e+73605u2Pl3dsT/MwCOCIc36SN2ctC218xIU/ZmiQz/J8/0Qw1R9b7OAwOxbu4rz2D
8IonDDSHMK3KwTmkF8AQXZwJlJ16ewBy/vYQl0jhk6gkIcqJJzTnZ/35eRfUng2+F0u9ZWgmV3jv
+p5HIUEvpHNksa1kce7oLub0/SH+Ge36J1lGUVdivXTc4rlW/FqgQffXrTEEGE7PZyKBex4kXQQU
9DY23Dpxyo6EkLiAVV2JUoajkyQz93N1LAf+8TLPD4WkQqOLBdu7tMXgZ5doy8ruAbH2kaA+gzNb
6rYdJGo+mXfngh44ow5kj+7GJvPQqfUoIqFuYk6XGTtQQhuvBjTnePXj7t8TtJChyWK6JpTyig+4
ihbTpGrJiSWOhi+AdSMzge6y/AZf29Bes+7bYrYo7lBzUC5aAWvkv4mebdmrJ11DsqQ6dJQQtmhU
3i/N9AzMkLPoa7vvdqq2MsRkpIl6eu46EBy/N9trs9O2KkoHINudFRrA05uVdJ9wRng2yIALexnv
WHC2+qfGr5q7XSKvhBP8LToWIcZhMBpRTklX8mEZLeBV8AXg8ckj97cFTi6C4Mimbho6f5j3xv5/
TvtsxSWNgOh/AlLfBlHrCA+TBmSVOhmR/W3/q3TPRajzJu1XqPgrtzgs9km3iAVFtpkFpZOE41lI
qav/4myfkUA0ybrLZ/JFmsmlpiCnSMjofZMNzeXFVYdM3Rg8zRPmc9sF4j9HXMcWL0cFfqbQclme
2vy6aJcpsZFr8IfjNxi5S+sqfOqd20bk5n8sk/HJ8WIGVO+Xip1ZAC7+CH0Z3iw2/P4GbrCePwwv
yd6cdK56Q5/Muz544vEei823ILVh9wmG/QltQwVBHxjlem/GrHeo+AGD0uuhmxfLKg0c/uYwWBN9
RblHMMWPJjtks5T1CYSNXC6dCO036dzxGa7/hNl/YyZX/po2hiPHE3oKCGbyVRU/yzzYbdcHWP3t
Cp/Fezk8YaBVOIdP7C61D4pWshWBlyFZ3XvCxLZpu1QQykiXjjHobjkv7D7bTFdgLX0YluukSACC
so/pWzbHmQSLONfaFR0ZEN5zsYv9cDnCLenf+LNVI7nzopI7rS5sygOwAGsdF+oUB1HTPAO1ZGUb
DKmickPfuix/IyaXH5eThD8jzjd9bsYHqWCpqGrQDAVzvs9Ooetx8Rw9L4U6i0h41pzhEZN3I5//
LFnV6KIdGSGUe84uZ81I7YmdqoEFMzB8nYpbkeQlZQUWIABEtMA7msqTpRmN74Ip42XN+1P4fGyT
ZhHeC5TgeSnR6lys/MCHuOhWI9JfVcKKYXqrtTGUOBikWzRF3ZZh/CYAfJ/hFNx1Q3P/FBXrNRxR
rsUaElbK+QYTVjGByiMq3zHL85dzvc+ifK2Z+BksFwqdzu4ASURnBaju2Ppb8w7B51tBMOvIu5+W
OJA8FCtFRKPxsf8Qa3fg1f18yTZT+AG9W2l4H30Pai5OucecwapjqI901SR71HzfyPW6crwdMK/B
rCiMB6SZvlLzyblpzx34jq6qbitXDbAWRIKb6fS4WqY6EUB/8wYi/w23pFreKuGogS7OvMfMbQh+
8/f2yY6ZphxzZgMiCESkZGi1w3xd7BUP1Uu8t8nj/zOlorpF2YXvaF6lEd3H6IjK1mhioQfXpD2P
qrNmpHCiCEYoKvdj/bwuhGHrZz1LLVMbPmeK0oxiq/13Ro0eV3dk+PnuPpBDt61CUOSf1cL6am1i
q1+9y0fKsS0og+zA4U59WAKUe8qpg5ZvHedLSLSCrDTb+ceibjkXVc4AznSpUU2W0PsXBE+m8XSp
/ZMXFk+0MzuIAGidBKZ11NY2pNGU/CoRcNfVr3Xiuz2Y2CraCnzWl/vte9IVlA8A4D6MpxOo0HZe
lswQED4qA6tiFlIPYMo2ewkOBcEbO6CUVL+0FEVRDWFt4Yf9E/UJ6QLVtiPdeXBI3CXK6BwP0v5o
ZrHwqHjbp6TQ4ERYJYcgdTUdMKtsSNBOpD7Jr2w409sWcPdngZp0qnRUg8br0ufT0zEYxpt0skxD
1SIv7T2EeaEaMs5HDTem95fIILDsySSXRQv//4TwH483JHsC3t9DGPSBCABFpn3ugCU6VU7AR0Dn
XudBHNAxoQftChKhUf4cCmxrzcfKkk5xNpuqMa0WShacUjYvwcneCxGd61a/eY2mVdMjMDdOGKDl
tvfTwpgE0BEWtV7tWmY/4d8cTcXp6eit3osyzq6F3uI0wVvrUgfgrUEWPAlV9BbecxtPscxgu3ZD
kmOoS4YBLxtJLcVXPwE5DpNFkUcJPG9DGSiGjIYew4EUHyqxRHFCIIBgw8wi0rgkzcHJxYo2QQZt
CJm0nXiUHuXIEuPjL8qTAAyfzrb6dzKIIlDaGE165nqz4o9+1obkfoTp4uRRu5PyoiYXZhQc04Dq
7bysiOrgwdI65YfEL6KixcWSt2ds01IFvGuxRFsHIhDcKyq1Zt7XyC/jHP6tFrYFrNBTSRWK/Vlj
1bQGaic5jCkmBsTEs9TmfViAdjobr70r9UbDse4r3hJSUl1TEoFgQAyBGi5XcHSn5lEH0xyoHO0x
EwsErPn9v7uAPWAT67Nky2wmkUwFGnzkp3pBluiwqWVjVxD4jX4WhHPZOUwG5uolMd5Gk70mTFvQ
QEvioKja3nCV3BN3GcQ7+WxwoHX1zbyvRE7sJzY73IE1KmREEnipiYSkiHj2fcb94zF9dCeCTMai
6w2vKdORDEjCfL6jGxz6SWVmTQMrtRHCfbFOvSqljKZf25MQ8s7G8XRV8gAc5C1Mg5DAs4z1aFpo
AKsi4T+Dgu40IzXa3KNrwY7nDJUB8RF3Uv8Yp2b/RyZw36MTv0/OBH6is/x+1n+oY5XNvMQ9pzo7
31YkYTIjBUub7RjRydw9mlPTm9EpyZAcQ4gZMjgGvofZhCoUNlm5zICPvmVUUlvBkmPrql0WcfPH
FDhhtx5X9V26Vj7tB+JS9j0uWswz34Kbi5EgV8TkuQ/jfhWkpcWNs1GdhMjVXgt187Tl2CH4bPAw
TDhQznAnWY43dt0a6LROXoaM441ly+t/zV/yJ26OhEaV9eEmk/Y1KgH5BM333LWlydD82/t0Qrwu
szt9LJ9MTrVbsM/Y9XN3IA30EVIlQj7BmJWnPcZsuguzz4d/mpefUYpgitOAgLxLY1bEE3aBgXYn
W/fXKbHDNyRHYdDwyYtKNXwRjZANhf3q2CRkerlDg/zR0F0tAukuoRecx3kB+AiDGilbtgSfQ0tt
eE0jYHizz9V0G41Ei+JSRunN7Ou+EBhNjEiywW6DECZjsDVsep78eRYbKo/bE7p5B+mWUmw9+4Ht
5HDq1C2NXU1SsaJ7tlSloTov44EBmguTaSs9oOnvWF5AL13Zt9UTReQWQX1s87ycj2IxUGeZYovV
j1UGwMMBTZ1XAsJfaEYvR0F45GTzX6PQvVaRZvvLVtS7xwVyh5sBONJXyXC8o2YCjoH7oreNDxHV
zplTttPlbcdlnqT166paV473+voIABuDfL2KZAMNkd+JfDoQWyUmSynLIrAwWZeLhPK5dZvzkf4y
E0v7hT3dD5XFO2MFTmhFAG7IEa13B22LJbHVYe4tZf7xDpVo/fr7EZ+sJJLJvyowzi9nTZ6LwHtY
mU8wA1DXvH2wgmSOG4vy4zsBRwGtJMybJvoKfZXwxp7yGF28DId4BOzeUucd41XRilOkE8hoYcuV
MPJzjU67fpF1IowSgN02Yza6vcfG/qmQ53s6rx+tx3epy/WmJ2qkpQouhuLMB0bZ/x2uICsD/yBw
Ykd6I96YPN/Sf2Nu418Dd2bsYjkJdgGg0H7HiKOwFhTvGtkoj/vALtmVDetQhlSqYCgGdLrd25YL
MsXuXwkEUamcnfJkSbm/2p3bGm6O16ilbPB+vE4sZjJSZOzWtMHFsBRSvIW7yAq1fpwrJC8o3gWk
2gKWJZosBB2qeYWTv7oT5VXVMqpp8+ac4SYL3r2tAK+dSxUeEwJHgScWGJJaAFtu4fMEm0wV0CiA
l4ztUIyc8CqsF5lT2FrFd2ntSbIj1Im0jK1e+ZU/lehyjFxXlujrtOn5zjz1vQjKFBoNpB5kX6EG
HzJE00qUmuBWR143+9HVCMXdewOn5xI40gPrpayIba++zh6yP82BHr+LE+AnpLMyfUKxGbucVToA
fqgTufmfQAUXmjU0NpVbeSGr+/t7WyGsWWuvcf7mMhKdjuPjqAawCGwNMeVmJJ29s9iFtSZfYJ1r
E3vlA+IQFUq++OO9+bQfQ4YhN+51dkYziTc1mPAYucUsy7JNSVKdYdJZ8lSjv6OLue7I4qNqKsXj
VctbmZbrlJ2wtbzu3GRXiEAX711rPu88x4/MIfxlTGjV1JlPlNxSmIaQc0Fsalk8tmQjIoJTDDDw
7G9bbR3SAc2wpCxiRcIU+F8U1qXOYj9MtGQz1PpR2Ga+ueVqIv9HgN/6YxUV3tsYbTJK1R5HyWG5
fkxVC3R9xia/5hdHNtM1/HEz4PGhqKZ/f4CHS3eJiZVQ1hQwF95v9nnH8rrrOZEAfzHV2r+kWiQi
3L44K519drt/mWCKpN0jpPP+cgxtXq6OBN4iVnbXi5cRhbzfqTWhxUfPvVTIyhwGrjciVSFR8eDk
uaOVdOQPbDMKlMLXB9uPAKq/d6lt/Fn0g5ToVoXNnmN5SVkja994gSJzX3m19SplslD1OOFTsnql
ZzK5ZPZbLKaz+Ttu/6jg6eyI0izRRTxzKxyNfaGNEgcjXcP3YJJtTmbcg18rb+n5geb7syrmyj4r
qAEjBqNvd1xX5cpTrtQMoV0mOHt48rmmaeQKkWlBQrmMRX1seVGUMS3u1zm5OPA9tGc+kfQaUPUX
Fkw5EHzjCRf1HMcQpbe4S5hBcLNEHlkhGxE1K7R3Irms7QBYpZbQYl/kjb6529JhhuCu5nfw4QKB
uLrA1g7YPCW+mO7o8uP/yxXW4cqycODiEphjdBxwS/E6B3nGs7tydKOHeEzyxAwRHwW2Uq7Ogl8V
Eo2Kjtadhse8xmWJrkdlaCcT2w2drHccs672H1aScm2AVCzCa6xb3bQ3G4oe6G87YLQXKDm+XmjI
2H/3Okig7zRd0LAcEqSp4IUXdmbvay/KRGFC2hPWaWhkCyMRhL6QcznvOlu6Ou78k8gJEjkw1PTs
qL8owM1WmYvVzg8wt4NOvkXzQmWyL5UR2nRX+Bj4akvYN8vRBLUfeEc9yWah483T55AQ7qua8cUW
a7J80lToO6/CXqeZHEIlKlhhpIqhqjvig1GRWByUHVq9utdVUHZGZmRKY+Pabl5xY7z/LDeO+uti
MVgmgYL9to79sKKYgmIdk65cpomRrJiaZ8AKc1P7dzAreCA3APEyc1ngw2cmG4+21aT+jVcHvFxV
5XDtm8ZX7GmdSlcmZKFF2G7upg3vDlpiQ0FuQtX0RTe1XIU3Q4CcSw2RzDqKlN61t/k+3NHIokMI
2pyPOGMKAuAQ2afTCfU+Dd6WlX2d+Mtry/iiyl3d1WowHUWkN4iy55rn36CdJuuUs0jdkPm3frml
vgwWcSq0rEBxa0qiFiBVlO4Q5qe7rdtategNLgDoTDw/I16bNQwGXZasMW9WnJp757mT8WzBe2qf
DGoNqt2Mzpj7iWjNlGr9tZABXJISYLqPZXc3oq2ytZGIsdy3/rPLkxYHg3Qmt6j2YjdgHAo/3B4q
VfU4y8eUW7eQLOni4nfAV6w9ybeDzmiE0dSo5FTphz4XxpxOJbNaCE8WMKqgXtDl8Py9pAbYCjLc
7uRzJHNgu8Ke15GfZHr2XRkH8YYr0jbYqlOQX1UPrpEmZe33ItE+T+/juo8B20aGKLc2qkzf5nrD
5RU1aJ5/pplYDWKLA73MB75VOBlWZTCCn0UsM3av+OBbmamPH7JUJO5i62D/AV93oYj+aiKrH5hp
5FWkTzjFsxr2idbW6IUq2TMfHnLelkF6Pices1VycRYhmMyliKGZObRBy1rvElnpB+rH0ajVidvW
1dtIJaHPIhnCHVHL3VlgwoB1+E0FR+r9H4EjRty5OD4xFnV32eNJrFVwIaT/9L7aW9E/0fDfojgI
RuoRPDpBeDr1bEv93HktyM5Sa/LS51KPo9rwiJjCJ5dF7FZm/vxBkn9tiYQzU/030nKGv23KcWzQ
a3wythBh9ZW1zYV+nZzwan5zc+llRJMO8CCD9JhyqJxyHZBR7tyQUdR14rDMAzSxWygk41bQH/bt
3692K3nYJ+s3tEYd0HZvdtN07gjtrCHe7cAvn76uDPSrP9sep9szHpNpHCRTn9wx4igNFna76tdT
EavC8Nr6vKB7F3aN8v/1jNJljtSF0/mpkT3iGaxw9LCccVSh+t+VuI70VhmH+GhwUchi13eLeIeR
RaZbhhQ/2yeH0AsQus5BcnqmVTMf9Luml3RgyWWtvjLsYUupORsHVtyZ8VXTbKv6UXcOFO9Pjk76
lPM9CK7AhKvVGQP4YB/HQniC2cBTMmUFNS/NP2xhCW9DmE+nEcqnFvMjtMWLdse19AYx49XRUiIn
U6qlf/1Ja98WEvdtYEfO2WpTMHbTaEgm03RW2vBl3zu2+9+og3kNgrD458xLmFq3q+qyQmsJMstf
RqN9spcf6Do8ky7aX20wPoTbhP1Qsq8K6ayeoXNP9sf1o9EuV0VTpmPbchz9QvCSDpX9MXE6VvIN
H71puSzhD3YLEzpUsNFb1zwY2Tn50BgaszI71CANg014E1ZqzZ24fxOYxaIjnBUJA0aU+sUuGj/T
7iuXPaoJ+KTnlKWl+ccqPWbftzDKH2NChLMJ7t2eTBk2xaHpS6kObuAQV++K0ZuSl52nCEoDT5uE
Bm0Nw5l6GSe3IVioqK6URUU0kI+ZipUHMP6Od/E/OGU+JCv2/ciy7RWvHLZe0v37JFn/Zr3KIn9e
9tg5IfCqXvqg9U0VZQuGLgikydu9JkhPzlJF3fIbNfT9p+iwtng7I89afcISjH8d1vmLXUKaF7xb
w5C0zoBG4RXZs2C/XUp0D0jQ8Uf5IemFj009cxNeC+30kPGrC5KpIHTlHj5RONWqYc7cVHD9pm4d
Tge3cz2Wy8/4OKb6l8PknMBCvg0tAoftq6U80FspdJcBDrPBSPOmozxos9K8PhEma8wrJrcfYjsh
H6RiBTn2qHy9I2AZQRT2IIJiKSO7IPD1gZZBlO0YVGnGtJSyL0jleMPLi0qEJxN/Frdh2NCHFON+
lzGDeVTQHN8WZXrV+5n00y9jN7+oRFBnh8NK0kLxdArdLCZCEDwpkr81Utm+mvvHCBE5f7mx5INR
YmtVK+mOYz67DgoY4J0lwVRlgjfxNLxippVZ6GB0ncWPoY4NcJLksQgIlvVVHWYK2QdfcRYlgkWO
ItdXObN3qqLPQhyNa7Lq2XGRR/ZN89QI3H3vO1mgF/l7uuhbFtFmCbwKxKkiouZ3nLy27LvVDgFZ
RsSvtiffOJjSy8HEI0lXrPzpWWh4pxkEgZ/Qg9TKXmIYI9+aYzI+kYD0+KlVocE87MkooAFVdfny
zEFVn4f0aPL9YYiWrbht6OdN58TPleCmIsBsbtJEZ600YSTQd+DmGYa8/phihW9oKNiV5Jm+Y+b7
2VaxytuX5ugP2jhlcSa6be7ijNp6IPI2rHy6nkH6O8SWmeESk4xls1lXRJ6fO11YweaYHxmvVNLx
m7pQw7v8ZiOt6Z1M5VVe6oZUspQJq5Ops70gtrHlcYFxinoB90zjKaT75JXOpAU3t+T2DLYIl9/d
Xyx9Wu+cPMBjfFMzWV9yn/i+u7+jAps5cOjOclWaKVLDPFy7Vd4p44HENJL1CHworlSnnSZMpINj
VVAaFknh260C6cVE2Kts7f1NDM5I0LctA6bAQNjEQqPJzgjzshGaNt3VNGWKG1aEGKH1EKBp+ges
rfDie8Rovgfyy1zYiVVbuG8eoKey/I2wI0S4QNQsUL28YTWEJ3IIsSVLS8Bs3XJjdnspmXoRwPyd
m4OtsqnVbQ8Jcyrqgl2VxYIiU94NjqBe01JVGDsmvn30nw6WXUaMiQiat7I+G0pisIz2WwKKnt0U
4eI0KpP4oLPtfwhdi08WXv/9w4XWM+nQy9GQTQC6MJ74LBgeCzPPDN5uVyH5EqLenCyOEA3tGEfL
enxnCTjx9MPBoI7qVdl2RM6JNQ3+wEyxxWLm6vLAkHGhWMsbKDCYjqpOp09+psyy5SjYELwNGFRG
4mZuEDgUKJka9De8aEdk3D2jFCtcvDP9WzRjep37X1sTeiNFe+0WNS7OQINQ3LvCo2KhHbgCmYWW
rOZNWLoxpSxjj9fjkrRYMZU9kimrdm0lyAnl46yAD/Kqnk8a36p7qj+TQrZHGWClS68mx37y8t6z
Ww+dglBpoo56zsM7i6Fw3rWDhbbj2wQfvi7QCBHP4vgjQx0dxUQrJ2rbrxqEDBx3qaPxA/dR5j+G
TnwmD8by1AXDRzGRWStWAkf/jUqbZWwsWpC4QCi5d7bihMCfecEXH/tSPH8NJPsTk4ttpfAAkB3u
wSxD4h0svCCLcAlNkpS0Z7B6tc0gkfTeErnld9mALyRiZST03OZK8DOmLWa+ivBKWVhoLdnTaFHr
1wP+ZCrinp9beeU6A/0A+LBOuhj56rcFqezVM8CGDAY24Q57A/CB8ZiS7li1G214/WgVQIHguiZr
wGmO9+FTGA3HhQYF8jWbH2cAxSy6No3rkOulKeB1FGrV8Wd0l1AG+6R4RPtc5nXR+mAALcgsNgQy
hf2BwOnKgPTbw43X6/0SpHPzcKHqe+uUTP4HhZaBV+KsHJpePKLI/KpQaVezcPf0nX2jEku6ivC+
IZrw0CgX8JdM8voHJr3DucaWgOjJHB/T7GniPa8gpVIaxDJPLyYb9FbZsNi4hu6EDtplm1quMhTP
fPbfE1CRfWorjT40B8L74ukilZ20TR8JvWC9LUYyHqEj1TL1NcDmYGPIYLee3dCU3qVTGJKPOIvg
MmwGaV6dStnUsffpsvj2aNW7Jk5q09/PM2O7jYdSgHGtGozeTaPSuJ8kcuTXnu58pllEUtO8fgMd
pg94oMm9+vxbqw3jP21WiGKhtKTSScWEk6j9cl5CKX0SYV0vIZj0JRC84n1SKe0avmvXyAr0dLV5
4O5RWFctLzCNpZtQFMrIIhlTRTYUlUFdV93dRFLPedIadAk06BsMVWsRruoJzzjHr38RuX66vuR+
EUZZTH9jVq3dQFW4bysZVR3J6aHnEdt5HnJzRZlq0xDv7JwVNykRDXN7JNssgk05C23Teeifcvdn
hHih9i+pU5zxe5FaYQJ5kAPoBl36cUiKewUvh1FUJJGCUcFKm+NoE7qdNfllJIfDVbp92t1d1+un
a9UUBLIzwSf663pTfU+1CEQ2gh0MRWTQBWW1inV1tdFsHzMXmc8hSJ1+DYfPuYVeNJOQsc84gJYY
HBp0QLJXyD/5CqIP04Y/AsUi9ue9LTdl65UHBvaIbHlpqIOawYMYpSC8VfEB0769UXv5rVmZL03Q
ZZ3uhSJRrtar1gSAmJpBPMZLSkUzOXhFOy6OOBYRkm54FBfpTnrGKrJzasmqSMIa80b7lERNJ4Nh
YL6BfXEhk+wFBRuoU/NhPOWcUGDungfTrB0ainawy3jhjovjh2zpYyw9XsxlG9s/50N833zVtRB7
OBFw5vPXQo9FLJTq0ZyFjDDjsAkWPs/P/6HpQWNwY3zV89fNFJl1Dp0iO5ACjdjkOyIyYTEvwdfn
aJtYUnxPVtV698Uw6q1ZqSQrddyJtO5UekSsMLExDqdBubX7S9+pacc8blkUbXIJ+tKFPQYdcJmX
aUdExBmO25DoiyUCduvaGo3+H6Ic3/m8++gdtPfQNXaX95BSI/DUYECzchilnf96noEz3i8UqbOT
HE0Vn7aeYM1prQbYWc6tVe/LZjtx6DRjo6i0DKT1LNLaFXZqm6E2A+0jv/Cebk/KRKjf0E50/AVQ
7ZiHFNJWHKoo7mTUZxQmxwA7VlUMhOp0pazUSPZ1R2uYjC6q/Ezz/W+7FA5FBR/bubt1B8YULpAZ
gGhVGU1gS+nQNRqhck9Uy//7+vgVvKVhBcXmoAkg9TbqAfWocZL6MeNb+VAAtY/hdxxC/dgqm6zJ
KTtgWluLxCXIFt16VcJRm9+8kH5+tX1mLxzgsLL+aZMocsDDw+nady8XUTyqzp5F24Lep/3WYNls
mzA85FOOQTvguypi79mkVlfMT8lx3nFHBclUmnHPMglYFV0cRbvR84KGHi0ZUKacXtDHB0XnbF+y
EDhSO3S5u2nJktkAg6VmbusCypwJyATpzk6fje1jq/lCi1eC/KJpecWKOGKQoISJUhQvkgQkVc+V
8nQTbZ02vfMBuv92RCQC4+/qaWmij5wLVQQFzhz5FZejHhj8ElJVsPFUPLwWxIa/r+BSZsz8rNEw
4UGB+VZg1g3u/FxOoGCSmsTLi0Y7WUwUZR7K1hPd2Fijn17aA30P30LHP4YFhJv3gysADwSaPMK6
00V6TZ1b8yaFXpMJc1eV9JaTOZBU/HlW0jDAhN7Of3nbgr1u6TexB3HpJJRnDPXPvoJbF5qlhMKf
SIDu9qp7Q2T7N9ocZihRAgCuPQmUZyqizlToy7v1+S9fhGkkPh0dSBkNojTg7MN5+sQJ5p5CQums
IePzCaz1npB1In8z7PIhsGTnlCszru+gj41+H/7oFj8TnsdDpU2krpRB5lckEfVwlwyHc4/P6DYu
LYWhg4vdXm4VGkboEwirJ+rygbrEKLok+QEj0hALxkLlPOplthx/dXctq3NSryJ0HgXYJHq237Or
SISSWcfMa7hvKDGio0tHv1u6xOl7KqAvn9KoQxikToqW+qL1o3QlHJ7Ztl2C4UGzVqIZuq3xVz3o
l1gqMl7GabTh1MHj44IF9sezsZCbhNc/j/eX+Tr2luhhn0olhI7di7bBRn91mv0EJ3p5yFPDkiTW
nCMH9iS85J2r+VrAwcafUPpy7cPWRCDBBzVMpXDM5UlDSmeiHNRMkBUn1Kywyv0gKQBKx9DXNHw3
9k/+NwofBqq15XjTFQahspfQk7V3o8TXwjLdMDuh1i0yv/VQj4Ncq/hnd3XiWwmI4bHqo7rGmgLa
ebaImC2+3wEYkHE8WDydT/NU3nf3BFP1U+wGZRpaSKJUCcxDqeJ1kgyUKEqD1rypqASstNK6Pbel
kn3OJ6jVFfgB10LybEnrpxukBlp2kiP1ayPDBUcFArsE2oQjRk61P2i99CG3gef9UcD8RJp4L2QZ
jvInTdr8cAvMuQoXCRBi3kWuYSmRX44J8PPVt2uE9AP8Ny7XwtxOEEReokh7/eoFZymvtw2EgXzd
g8Qz7JNCnRZg7co2L1lCHOpV8NUmddQxJsNQrXXBZ/uNLwCeHSynqo3+yKyeqN6U6Z1NYqWlmmAC
Ki9JJ+dYKogKlzrGU8eRdVYdqxnxoHOfqM39C4raUGt3dfvVswBhrjI+aBBJb509n4V7WYY4aGxU
HygkKSXCRVdmhPSJcxdnPnhWW2YonsOkuhUhDX0Rd3i8fVxAZtXc5Rd5OKipoCGErDbgOJhlCD8R
9cJb+5m/TOimIxzcCeBMzTK/Y5gQNseC5OUxOohGgCANXYe0+J5BVWT9gQSk+4NNuXIRngmY4nK4
a+wFtbE8CYh56Dp4z7yOX4laJbIVwpMRD5D/Fiylo9SK4UBWJ+516FHlV9xy0ilTExv7qQ6mqJs2
z029CZWnM3cdZ+TIWgK7uvHooTEv5Z9HQFfpNqWX7irv/kdlriv2TOAnxd43MIdK6+2VHns1WRJI
gYvE6SgZA3vNN9bluwg+6Yay+qnq1oSyW/C4fWCp/hdOfxkKGQUkcY3XJsGN09GEIDMv6MkjBddz
frziCW5hw0gdjIEvYmqp3fBJj717HAtb8oYRIWNXe3rOEpuDJ4cXTvShadM3ZK7C5T21y+mtxz+r
8YFk+xKEJDYo1EmHFM/cy3Clk1t8FoyMiYpXONemfufPwGjJvRrmGinO32hr23nx6wrYY2dXrvXb
0LC/KxdrAEhe13qVn6Jc8ftOFU6fXPheZh9SytAheaIV1r99bM9bMNaLhwUVjj40AgnPRBQnYMoV
T8wX9a73DRorT3CuAJ8z2wcqkHVH+C6yuRF9tJJYiH3xahgU6f4X0a1/4eD+lvfcg/TPfq6WL8kO
mSVtFrw45zVDMEb+DYKammThtwKGp3NmJKgoK+wvQ+xJCJ7UTGMMO8cMzzCuPae/Y1ZqDZ3gao8W
CUjw6aycdiKJH7SY6wJUjG4nz3jOEgR41eY4kRmvN2O2W4eyMQj50IPYaX6kuNX+JQJvJTO/Sl9y
PQm200ODMwCus41vee0w7OZZ52fqPLlRgQLiHBsukmrTRlihNUWUf3H1Yd+4+z3AsKABhDiE3Whn
lFDkSUOIhrfNYknDPZ8LkLad6IlnN75fCEr/RqXhtbFShNmZ2s3spLI2i/dwVA9B0aojVeMpN1Yf
biE9oMNJYTY3PBh+4S90FUzK4lUY1RPUKoaKwRekhJJ1j1/SZb10fRR/KSsM2CLYVVtxPPndLm8u
Clg9IR02EeFyKcjMRBXyFwaGmsSS/9L2RwWHkUF7AFguXqCSOKC4lNZ5zrOPSPJLj8f3V3VTnGDc
gan8Jqf6rQJ04e6gkMNOYik9j6PqAQPSJ8XDbMcTu/loETIlPThPtNBOceL7lP+OtvAFXRwX3feL
IJSFuANFMzPHZEDdvzSD3coyUCqUm/jNcIoRjMUu7Qy9FCmApAafoV3gNSeZ1qPwLhXXlXng+XVV
aekv8N9XLfRyYDKTokH0DVohS0coSoB+vnRSkG54URKuGwZetkD9Vzomc7ZL8CsEJ/DCgfxaDtXG
EGlf5O1zfjiJl/AlLLUEGiTPlb4WYnoCeKIhWXICPy6+2Uv4ZLx3oNur6M7xyTux66M85H31FIm+
fG8Bv5c+H6N46f1sahrK2phFZrPm9ZiXt4uClrugGIX5VMvMSuWWL0BueokhxJNZzAJHotbXSuy9
I4ex7wTk3FInMDz0umM0EOb1j9lzEVcoXoforbSvdTHERQvNxK76FmzLO7ymEbC7IYlEXOLXAf3A
gpDAxnsoeahoALI+zaP8zuiE/NjLNrtLJikta2P4NCBwQi4rYRd4Gn31Hat5fROUme++FDTZ2hYc
aHJVDft6NkdOPob08IjKruJpnFr59Bw093yRd1YTw6FNHEaYdOa6dnzulYJ2h+oZ/AyPd2IB4g++
tg3fUD2SVuCCnS6pMostX6+JbzNMOUSKczF8qV8V8DPvDYtj+XtxVb3FqJobCUm8KtBuG4dHQEM/
rLJYcg+Vz8BxqGSrqXVN5FYSLza9VYDE3lBsNDjkGEkV+6fs9RD1kOVI5mBhfwKYTz9PGUIv9jX+
gLzcNlQ/9Pgo7lsS7opx4R6rm/ZvD5XFLxE7FligDenirpfuzBKbbfXjxXhoPQ9Ix5xzQPkysLJ8
ADUoOmNnJIuB+woWdiVuwLk7EYycvRMCt8+4P7/ICMQ5KBwAP543mbrADU7b4ASG4uGH76NdATez
8ezPQbFSQgvitpi2IqTKoMDYJt81ltbSAHF/tRy0wBwxWKIi9iyoXgwzodjqEl/4EI8cIlvxi19p
AI4zl5D3AhxU22to+H5gRtOG5yevOPqg+I/txOOhGgvm1TP/vwZkIscLiox+ASrr+SsubFJpk5R8
7qnuHVCx1K8mpqtqe8iOvHYtkTtLfh/HVmlyad3Xxhgx9DKzoEnm6mA4qPHJKZXAEoJ88u1UNoL7
XDOWfGKrQgAvn9H27t0qDCDfGDr7GExu0fWiT9xuLyBDWQp3E8laROT12p8ZdxNPP5TBJblZSXvO
+3pglerG+/48iZkUsvyGcNb8BRRNVoKKwbVUyBpxJXczn9QDcSKK1nuPbIHr22CjNQOi8PplgDB9
uv4qWEt07Bo7t7OXqmIjcha9w6FWd18/fsRyu62RebPPfcj7+EemhPtorXPnbT/Hh4FTb9qxWGsy
tiAnaAqHFlGeRkEFFz4Wow4Y5AVO5jVi6KdkaTZf3gcgpRVZNuuhDVbH4DjQixyw00kZJC3kmiHk
EONaukP8Yzaiyt8ANnXAux5L+3D7uk7s3hIFYAROHBX/fj0U74dkcU0/vdYUvjlrdwJq1alu5j+A
QVJaL/hTdmGaQOAZDHxamttQzOcQTV6vM137BVL10E7NVC5oz2V7tVLzBZeQRyUAOfmGP1JdeEtX
Vqebex+JxAtLt/yVwWS/YrUEsLKUM8cjC3Q88aOqEsbxMzOnXslBYVajHagK8VUF+SONNoR+q8XI
K3e2X/9hfk1huxutbsam0CNoVRdbK1ccrti7NcXuwv3VK22v3QiMIwmD5L+h1WyCnJod86ebgZ7U
Bd/ZUV+fuFvYHNEx7BTnZSSNcM6/ElVvZxP4uiMbJJcC3QvR+JjbCRZPBvCNrJZ53CU4hYoYRPRS
+cvkmyXm3CjyCoWTlWqee51CYnR7cSOiL/cOG3KizRi9TQ4l0YG/TS15q+MXd/5HFK8/5wkWyaDo
8APJcqzf+yCA+AgtI7vhqDbf8xD/S0WzcDXMgMp5ZpIvzkwo9I+XmlRVUFnDXXf7JZS1TyKWc482
N1VjiyJJzmGIx3slQwsaScdTeLRbcMIJyL6swPCnPMnBifuLkYH1ZgUpbA4NCdd8wMmTxduLTEcp
lSoBd/X4RRWQA9xX+9ICUwKdSFi7HMBedggiaNiQwota/J4+Kw5d1hjMlL18RtOasTLK2h7e82UF
zDT0LzxtFHjyWOpJO4s8DsdDkU+OuXAg1de25fqe9afkTTdde3cnwi7f0HKKqmKKuIzq9hQwxgfV
oF8KKewZN//P3qS2Bl9QXkaBunp3R5N1y4e6nDaDQK1dbVTKD0o93k+9beYl8B3Dbrt4q5wO1hjR
5BOD+IVkorDrAtIBT/D/mZQ6t+dyy7PVg5t7sT9tZnaoAOPhTfaUJrD90sSGSGMMb/zmSEzz+pxl
7IilUH54G/6ITr1wrem+LsJJHwVsgf3EEWFwisBjYd4W+adHpe7/2ASUrONrZnwM6NM7cibqPUd0
mFBiiq3PnnfPpaQbKidDvJb/JRqHoZr4SxYSolGD0Zx3NGaOcpj5BUdDe0eRu48/chDnBE04fxFb
d+ZfBp+5CLSUM0xtxj+Ly1Hrt9deZjvJoONk111veBMG8xkxcKRcTjde7atFFxDbazEiwvuKoVe+
CPIoJvZgXAopFu/4QaRFRZ6ZnUOf/Dlb+Qh3K/6BDTteqANN90/YrCHWGs/yzVs2hyPKPCRiiwS5
7RIgxmnRjxsB2rxhROrJx4VM+dvpxeTkI/exKteg6RwQYRDO/4E+rPQTJhA5rA1xhCqHkNBUHvPf
T2NxM+BMATncSgAJM5vOw/VwOoKPfLh8qUeV3QV+ZaFVSclHXF98NG4lVbCozh41r4ErwPfN+j7D
uqJHM73jPUsGnf2fIaISRyKOo+MR10wDu6HhdL7rEIXCRyspQyltcXEvILmTHpNJqOkENl8At3I7
iyLwVD9DL1rEpG85qEmgF1xF8PSY0gf+wFnwDfBRu0WT7cwjUDY9n8sjfMRL6VRq8o/fEp/nVtqW
D4mdcRCr939iL92D1y2RZ+ErFvWqwdTm/0gtzoaMogtarAjOFwOEqZ5e+kRkqmh9N+6t6cRfOV5r
jF+uJGq4sfYCujY7hnoqXO/x9yIMmOfxR3xej7SnTKrQjwthnomYspK/gZ/CPs94jm0oiQpGc3y4
SHurMp/IuzA5Dx2eLvIZmLI19NssWztNiDUxq5XwW/JRGzJT434VmLRQs+UMpepC8YRH1vwFmEWX
jjq9Mc3MMcUc1Oy9yk6fopDDTToNT1N3pmhFQj51qmY47nTpupQS3aqI/NiE7T0IBeWQYvq2TlDs
fqs++Raiysb+cz6JFdkqsn5TTw3iqMV+EfbB/pz5DAtRartUFEGRLOVAF1WVUSdiqdkxPINT6UWA
qs8H+bMd1DdmqbcDs8kr5oRIpZkHaW06cmXsxJ7BaOhLL1fEr4aIGLVkOkMItlk0Drz3PL4ncl42
edWhBqftUA3DWN+tKcZX94UeRmthf3TKWu4afLQcxkmvoYeI2SqKpxeFognYXXdLQdToI4OTWRuz
EJEIube7iOp3hkNbK7m9WDVixg/ghIMZQVL/xIduLCTfQHFMJ5LsWkNBxpfccPu/LRRTqQQwb7m2
R9TGk5J5LnoTNxzDmROAD+SN7cthnbBUFumjk48EpqnEL5qSVDx73Sjmg345V2B2dQeM+u0Yu4E4
WPoQs45BKFastFclLWUywm0Al6tk7EYs8qFYCn8SfhMhZa+oRiCIfEtmpEUKXiHbUw2Q92y2NCN4
wRU57VbuuojdL3qtloNP5ThzDQOeKNGNnU1Wxrl+McweICHIn0M0MhJY/3CcTOxkst+HYGefqis2
KC+RDaKys2FI2+YTFiFj5eyAAAWhZR07zWkbHbF7W48xwqwwxy0UK2qiLXCA6L2wNzomr5KocSrY
ZMm0KO/Dm8ohzSj8oA7cMVZeH5CLrFC7+dBF+V/KU3/Ih0Im6usxZd+e/rjpS+BjTalv8LYb7ubN
7aHt6+MFp88YIyE9cp9F7g+mcsIT9AxcT2ip5P+zYBQpMB88/t4mtHZ/xz3pMX0mtDCXGE1P6ZB7
rxfc6BXuBeHRCUKl8khfT/6Q5cg9A+LCurcb47ufRbJmJkBmstc6iCoTDuhqrvRhc9k8Cky/X6nb
XSndc+2LjCkDpZfWBHE3CUg7Zh4i889c6niRUsX773YnMkU5rSmnmFSwu4fHqOjVgY49IvlJziS7
iQI3i5nn6tPTJeIWjydD9YXEKZ0JsE7mVIB3EmRKzlqIi+xnHWwh5KejJ8nCCdQh/zkH29hdiPka
KvalaT0nzdACcuxZA3lvKoHoL46MiwPbCHMvy+eqQW5+zHaftYzBJEmDzeUdaYsDDYHPpjL2qr8v
++MONL0Hi9uBzTxTKniqKhpvNORlt2hdnyoNkdqbztkqUBfBAa/rGY4Cn5yn/XH64DBkhSEQXVK9
VZU8Bp7eNqG1WR1LusfmEg5X6gzHVQVND2WL6aHYj7//b8ebAT47PNCNps/hjj7xBiVhRxqEHn1U
aa1EHjglBNgDEpcZvaVW8+3I5RS/oRdVTzRmYMvb9wZLsm+jMhmkZOPmCmJ2NAuMqNWGcZScBG0q
NRk+WIBOvMd1F0enM4p5Gj41vDZstwrCwLN5wz3pxThGtEnAV2j+/w/x2h3My9xOp4Adrm6wML+p
eTO01sFXzQ1cnfaIskjCQqnqMcSd5/+G3dC5eBNW3Bv5KygKH406lrnJinIlNElFYWfZg7Zgr6uy
n/iVx0zaDG2pGMtbXeCLqEVpa0ftWEZfRajSgAlcHNtpcutqZmFPmIZqrUK4Bd159N6G0vO1UHxv
7spDSjR6VqVkAR785sZ498daw+7Qx8tdyEJx3XlSURh2710D2AlhdWEGBvarhgvk/iq9g6S9X5dD
rLuWEZkRtQexW51KwbdsjNEoYB7STBkndM2djeKpxdhiYEzoBbz7wv4CKWjf5J55dCtiuxMXucXX
Yx24+5O9EF3FLBqG8o+C3pG1L0/hQ/NX6buUN4xEgq6qmcaIiY7Di3ofG6JsHQhQkCxO8KSsPSvU
QQ5tO8IaYs0sX8ZJ/Z6wklaDSAQP0L1M89yaGNJ+d7kdG9Dq78LvMZaLQHV+ir/+8wL4wOZwJMC7
FTKOYRsgk865CoHcxdYiCZ0fpqUGU5WloJWTcfpwapqIE19JhKTQgZqt2mtBsjgtcMNtjFnbzQ5r
0fPuTHPI/wuJsArlMManKZE+bP4OR5za3i3FrmggBR4ODZw6ri/tqZuZ6KvtM2nWhHSoUXBUQ6Uk
IHxFEbYSZEf+I0Eclt3FNLLlCCRiYRM9BYGAPF2SvFWFe09tQDDP4bJD48+eFrVjUJPbQdWCNBvJ
10i2JB+vuv/cCI5S1kVjZ1G1fZt7vKLwMBH3DqHxBpXudMLnzyT6Af50Ejgh8BABF/uKKlDH0w5B
BdQDD95DPwDJL0cfURzkYEQcTl++YidUqTyMqZe+wAjlOFGapomD2agfX43O8tXDGLyDsFVYyEwy
dXPM825MqGu/SUk4h/Lw4ATE5XmuOUJD+kMF9eOPVdsbD7Yzpc8CWM4uUyOjADe+JdjxbxWjECBl
DXs51pUcDRwFvg82y2Bbj13r/DjrQM21/7qzJOW/BH0o5HaNlPExFIL/3KwzN0k1CAqECmUfJL7w
qlXOzKgVq8PXZkqHfkXZICA71VzBV/nnkiCW8hEIWN/KmFHPNOMiWVJXK0l4knYWEn51ptDa6khZ
sL5yF+jK1jVqipYY9hwwKzVPgtekiRk/mGddpy7SkBZgQ8nSa5yJQQr3lMUoro9CjFTEgq95Me0u
JU69iI7+X/PxXJ0+HH8S71RfGdN3L5MGxm/vMQ9ORhGTHlMatKB7a0L8bpIZtf/lFxruelHjIFM7
3keaaPkhO0CYGbuMyTVcKB1UafdbvSRag31/t/QQW0stoFk4wHNlmTthA0OEMEOixZTzzNwmti7R
LemUcbwzgofoxc3iZXhuUMBUEoQoB8Xyruw/X62QRbUgooyxD0n8esJOKYv1oaTc7dAPQbqZbzzo
BwqSb7dNlDjjC7+1RvRdtd65U6YmJ0WJMIzKIzSWXPeNktr4F95bsPxbjdG3M/xZH83KOj5cr8wZ
iHPmZeEV2dGlxnhyVBO3Z9gv+yz/RTcsUtcZI7aTC+zXqIGWftLq6LR8WWe1yucoRd/BUPDiKS3T
W1uoJOYfZ6f1a9+X6q1oL2mVIR8wpSFaCb76d4S4mdiSDw0CDtjU6OpeJ5ZkJ+mnurok/XCVbEki
cY1c63OboIj5QDM50PmyfN8epkngNHMkGA2AEVy/peLcW+5mgKMWlzR0vCTHoMrAeSn7x+Wzamxg
zGTlNZo9/6HwEU1EJFZSnqQ0/qlt0dMmotRqXRTTSSSw+cUPs1Ehse2fG49EdJTsW2WmH2lIVKXR
O/5wrVXW5NalJlYpDyzHgpaLIlUGmQYdJX7tCp9R5R8YaDz/JNBwDTT90grKrqFI+FUTf8N9ojyo
IGAjs8yBWXAVODy1bABf6pfmNy993GQuGfzc/VGSHA7oNoGiTnhloO74YEY8dA6pxvvhn4nXgVMs
s9cu5INK1Bjv/3LF2g9+QOA596TpiJzIjhaKMSWHpi+F6eiscGf2Lp5rr11BOyDB32nWpv6y4tIP
5yc2i5Z6CsSRCnn8l0d5adDqs81+NIbO8NCmDjsJs3DIsoTOofjnEENtSwUFhrCFcCmFVQly7tKU
v3edqpQOdkofB9q/oLEjPV9teQ5fS2g/inxqCorIUTgfUb2tIe18Nfkd3GGj1fBprXxGgx7OeyN8
V9GgPzYyZrSr2yKE3t1hB7+ec6oSfFV+hfeVI/iB2T3CJGfkXrqVmntqhtXdgkkdetOGcguCElEk
H7w3lfgKzcx77o4qCCDbIwujf+F2kR7niEbwS7fH96YqHwejzNmwA3ZVfD74OmVEbL5xY9hjswGl
sFfCMR4/zRihwinFMA0kZKjjzVYf52F+r3U6672+bXPr1tPBB7R1Xtp9MI8nEjuwHYZl8Etb2vgC
QlQHJ87MePztz2e+ObKVGKnxTO0iwO70QWeORBN8damLdM5NleAVoL+P70TwvUiYOOqUX5lC6K7+
T+66kOvaAwCRz5vsujjkxiVQ2pVBCQKXLsHiaC1Xzs0s5G8zKasRODTiWIzeucPEX9UPPTw0ItkM
2HJOAYko6iyv+p0JhSMFhv+SyJeTnTo9CRYiMsIupSo2VdtmNpiO7/VciTe/XLnkhiAY+K7HekTo
K2YL4peeVanlLXQX/UuDkAaF8G1NBcBwYi1uzf8cQh2pLbKRWpFrRWPoajPcJ+aro/mHmf6Tp++l
ZVTwnsdx2LRpZ7bGX6ZKmPr6lhZEtaPVXRmixNUEmLSazT8auf/+9vV9r3hw/AqY2qQQjoNeChq8
2dxldEwp0lFfTl5E7b0npTszru7lJ4GH9Wla0ltFoAcFImXTwv/BLybpNeBMr0Fi/zw8WO7q1RAV
GJXdMwS7NdTLzbMGFNwvKp1IMfYcNltSXq36fNlGPu8YlCJehMQHJbyoMg/oG4dNmwB+bnOdSiqR
n7bNxiV1bpYLy12U5Zti9DDAWCsK4OdpMNPKwUBOPd19xgIYffnmGUYaFb/uIBQvON2furN7BdFS
meXovWxPqYe0lEJAE8on7BfOX1d3vSlLjx/NmCkbvQ3B1/jpgfQwQsm43LW94NhNh2lV7R/tHp2I
KMrb5Wht+Z9l/xFqJMCaoZ5dEYGKWBBeQ9u+aPWECgZBboTcB40q1drX83UF8VLxB6XHhOrhciUD
yPiXppHuSQuEfG7/40T/v3VStjlo3855LwKyXSl00mqFWC58PyV/YWVA6HQ7hzmuVAS5XmlqGicI
VQSKpqGD/+BaFsr1a4QcI1mzfFqOLi5qVzQQEhpzq8aOGb5BascQeKv8WeXGOqUQ/euHoJqsBPtz
2lTjB/XJGXa/BViGtjuxeJrpCqTXouYR199zte8lzx/4R+0gxcDK8GcasczwHN4inqJH7a8uVGfL
yVbMWBV9SZ4ZTIfuvpNwc1VIz6rGHmd0io/+F+B97B77QkdrY6biMEZRlT2j+8uF+W3KQxKYnCSE
WedaKF3X4aTXAIegBbgQIsyRP6maldMJWhp1XRqQBHS1vIAaQL1k7STmKhtX7rl4pKFT/gWIOQUm
uV9qry5OP5xO7n+1Y14ySHgiCssp8IUCgdfB7Kyr2SOE8WZeaBCQP73RPpfBsWEwbLLCCv65fbWk
SrLIUONtF4X6OOhDy9Ul6adZrdhr42G4L95P/ElYCmNuNflNT9LIz/4F07Igk8rn3kySbWqovQ61
bIHxjtlKnuLrnjMd7WKdPEwZpWToPw2EwkZ2YcijZAn6E2UYUpMLC3xBK+sfIUC75SNIdGWEnggF
Ya90N8ZhykLOJ0e2U7GtEErQoOAaCdcL+0n1imaN0KM3OW7UIN76D5mh1moUBARqopQI6bW/MAiT
RKgFkdZGhH4PAvXzkTP1IKVUZm8Ftye7USYNeccrNCxU52Nz7VaGMDHHdEBlf9OE/kWL3aItWitx
nWfPvPAxtvGYIXLk4qGV0tftikmm8xh8wiVDz1NZ1lnSec4MVneDNXLir6ilROPv2MiFF+IpJGV9
eGB6wR1GiUeCHhCk5uvc3rfzenmmEqpaox4IAibOjVUGXVbWSCu8wjRM5QMo9TPIOc6+zi6NDNUz
oVxUfASV9dG1WOrrbSmZYHCSvYguTaG/cfQYUjXk4KUcBSNsnhKpAVoXGBeInP+bpON7dJuZJRD6
LktgydTOi+73qfFxS3AJrQipVT2Uby65Hhs+OHe2NlEYSO3qTGb9AqVoJmAMaoeKgsUrIsvbGjqz
f+yR2UTY8ROInSHaDlvx+ONgGIqlCSktr77LlulTpOwrXzoJ4GFblCcbX4TDo7IB8FzpKINCnLP9
6dzo82rmiw2bFkq3Nh7LIsKkhSrhgvSyXQKZt7z6tHAWuNv3M5rrPsha1FhUn2bA0xdv8NCG1jL5
yyEnD9cubDpoMBpJ0tOGRgfgPNyQ89tCD4dCLrHl+p6GeTyJXfQTNu69JrP0ISizGfb+AQrO9ZrG
gvtmv7Fh33Dc2AFxxUA2dVoQE9HftKzIljNQI5ZR/VnywvFhHN7Fo/rBLXiQ07NXvZpnd4GQ4fCv
UHO8A8I2AA/uc8VjsihzsuomIokW3K5Qrf5JRuwZIuDkie3YnO01zHI3HWbL8LaKBOKTx5RHMifQ
Wr3lU6TwA1WJhLXHT2FN7Qol53QH0Scm7SkMADpJ6GtmVFa5kBFeB++C6d4/1mHJJ4doyGzAv2EB
grQKBXESJslyLdtJ75EPN9qnM2BxkfkizzlkiZqivLzpxAfgC4uO/Kx2QiZVo8/hLCrajB+g2RLV
HE2gzv6y0e2ijZTvJua/dmrXDXrCkUTgSQggtDx4sCSC31Lft0ed7LeZ7RQTExXTbDKplcYs9PUh
Dox1WaC1rzbCK1uZnFom9RC+RrL84zVud9yU9Wl1/xHAmzD6tZ+kx8ux2x0xhh9bKvQfEzN1xq74
3pTR6k/6nmWSijZhDeHaVSjqEaXh0opSBZDFA0JRb/rHMaH3v1Ks6k+Jz3/DWKCxrO/+TNWAO7xY
MdO+4K3AjgkCgraM8qksMJcX0Gy/yPE5bIGH8v47+Tu+orYwji8hNeFlBGa9WIbBG2J67bEhd3JZ
u2zU6ZIU8YM94In91M/Yk/TI6EAL6zUFZTzV85TFVf7Vx6Lws7VS3t2wkM/YIyicmCFrtli24mM3
xORrSDksBb2pTe/txvGiguBh1WKpwIi/2fsjqMHYAdyBYK5VJvanO7d8DZnEWOD6NYNHEuXX2nhQ
7bQoglPtGc8zr9uHUGca17ZQq3e+5VfLE+0kyTZBP/gyHXMtR2eqXNepKkR6Lji6DoAnhGL6xZYE
tsfpSHsTQ/CpuciMUglDAGv6XudOpaD3kwxJOI6FdcPDZnJaIHkp/zkZe/GFg9IJejvUa0yhIAi3
SazRyE49BPoIIs9kyQeR59d+vzQjynE/6johuLbNv3tAaDWfbGGcZRVEK809RNcCrDAiez0isaJd
xcufucZsVOQ0XUbAJfkQmVbA3fMaH4uhw2d8IdHS0mBb/mDZr2bvgBOmoOQ6gNUnUvy6pfR3SMh6
AzvYPsYgsggThA/kcvjKH4k63mYu+kZnl4XpYUoOFU7gpvAW+cRhs1m3lZjkmh4C0CznHCz1XfVV
+J8Q2/SXqA3/4nCMxIbwTCcE5BhV0g9Q7XsvQOWY2qdqI/XvlSABH8erxphVR2yYi4bANJ1dv00R
ypzaeN+/6LxU+zKSZX/Zfvpo8vG+wNMPy7P5Rt1um9Hvv5zUvnL/XWF2zasY4Yy2twbGEvBTUrgE
bqaNra4UuQLRsv894zOWEvKdI+4OVLpM247iMaHkvMPH2cS0Kx943UkJ1h//guKch3cu2mWFpjdy
01FaT0zeg03raKIYHj/s0flK2j9o48ulethdHvmKK4U8Non4LaGmd2xfqRFvCI733I1uNXRurwdh
38j6OblC+LvoeU8KrnFnR1jHpcnbaR0YqGZIb7JruQ6xoL3G4HbPqfwsqrvws/+i//yl8mWCLtZ4
SEG8fMXmDnkaYxRBEwN6mwmLV/1oK9WTurp+PpBzmxzjloiLmAsj6MNp2WtbeANCM46/3tSFxKd6
l7b0NqBgah7vfysIFflzK0vXp1Ml7dB/m5S+s6azjSyC7oEIktAUCgIfn0C43FHYqQxVekNeO8r9
6ATB/GS0ZtuHDEylPulAgYTgIXAQfAuvIr/1HtYs3Y9p3Y8AQvjvmQgBq0PanzBOF1V4puH/yNp4
WGMxO1YNrRyHkL2QvRJVuWDu9zQO/M1JwSQ98ZnnQxiQsk4fnkU7YuZMWykuf5xXPwBLFGy48s63
Lqnihz4UkQT+aUvDlLMxxsa+Anfa+DbHQq7CDbp4WiZzKTWiDEce5rro+Z87NqX0XS3TZILaevqz
1QReMRZN56OfVrVUTfim1Owsh56UvBJFZ2xAoQ50x1m+80g7wAHyIWvsrDy7k+x33PU1tCgfw7E2
qTGjx3j6PnhIHdQ2DPyXHG9/BgU3CZZ+/BeB9pfG9mSPnpoIPcBsUOQ7Stnet++yGSxp1oGUnQB6
gAA/38/hsQoz3AJs828IuS8jwDJpA5zMmPQAQy/TCP4EtVw7Dd1eRNX3WjHJ6KglKsDFlCbZq5sS
ig+2WuEzDAJYlqSM+oK+iVJiuHGMFPztbM5jn3fILqAJ7rbQKftodn9rSdcDhJogL3O0FuBSozmd
MVoPkeSyG1mA/7j6fP/TQMxKKBHUCgKUDfiQc2/Yh4IQw4Jljzj5IuWoydlE3agGOixfMcm7ycDO
w2j11WOi9aIAsUOvwMt6tdbUWoGUBuok5RX4M6wg3rolFkmRHrpRfwdMoABkL+U5D6k7KC7/qqXL
P79SQld9Dy2Qaih/J19WISwvwnjytJSA4JiHGdZN+y7tiw3MvhoFdc36vpgwJdmTvDuFLxahVj0j
UzFWpOU9fA5e4hsVN6lYHU9bpSXlxB0dcm3P4uMMtCJ6ECgmkG9sGjEyDLUVEc0KJqA51KF38Whg
Q4oRFw++wG5vGwi1JN6DM4UFz3h7AjalnEtRYiDUQQ/eVgm5/g5ZShuYygCMibQHC8KHD9WY/cOs
ublsPQxOWBZ5AOo5xh5SCPHZV4QMFbnRK1kh+sVt0sJoUhJ4dZfrRzpJM+adE0U8QAPm/+9FjIZK
WehvwukxbU+9XwFuTuapedP54ljI/WA9hpoS3WmdqpadJxpQuyO3+DaSm0adtkpI6lxv4DT+/kc/
MiuhHoemkjGsZQj0S38+v/fj0cJqmhpocP/twyE5u4nNi1rVgs8VWm+Yr5X3HCYkEl6nWOsCXbiN
zVyfncZLEKWXWidAjBXRWtA18KWi17Ilyr4taCua46GCIG3JDY2FXWG49NWBMb7tCyHN0kTZU6cw
l3FrUwgxyfnYWmi79QuIopazyYhCUKhbo3VJt4uHROE5Cvaq85ZrJd50S9m/+zlisvR8/vehc/j1
M2xlE3shaQUJ89DlrdAYNTdPjKoJAd7L4xYBa+aYW7muDlx6RqHeiRwXTq/23IoCjHvYcStkMgHF
UoJ80gRrsvTUhFBdDkAmUv76qKra8ToKawqO7Jn656KKmnYBTZWfM/fEo12Y/4gBmC+kJfwYNJ7b
ziE1QOPucIRfqT/CLk2iA50iFUe/WQboA16F9uWCAmE2LZMoK0maSRQL62OdNjCqlOMd8wFKKYZD
nGtzt54EB6KJSzsKTrQ9jb63/39ztAs9F5nUG4tBv2VWy8Fyw9x/sTpsbo59/r/mop/Ya3a1eVxX
QPowvl2J4ThIjfMMvAyEw1DIii97FlbKJPAVHPOmbS0jMEYyBrDsEDVeezMxdksTMw0Ru7iplGzO
ZDm5J0RW3DUucscvsXc0NlthjhHpjsJv9tCGtX8YfF0PWg50MtTa4ooonKHmjLH792snLObbOlhs
CAnFD/Ufg9RDxcZd7BEydzjy4p6OsAEF1l0PcDf8e76+QPR1drz+elIPh/Afka+DGrTpdUAVZH1J
hx5kbV96E3lS0Z8J6LfhudMzHPS98vcK3ObJtHmPwA1JbBXToAkBbtmaTil2z2Mim6DFmLCvoRW9
IsACAfQelGug7W1Hdr9mf6DL4x9v9tMQrptK0J8ks96R56NeKwg2fr6CANDBFjW9tal35TT/mh+L
p/LiFw8+cL7twRxZXHLeJBeDe215ousCO7QaOkW9nomKgxCPcBG79fYQeh8jwHCQXqbcdggowJG3
O7vCGzrW/qj7Cu+GjwgAEjKe4W+QDzarXMLIydD4q2Qt1q6DSpecan19sLnt61a+Ak71nNrpHoV6
KkNmvHj0X7YOIuIijR7sGxUg1F6yNSUXQdqVwptwBhlv97jmuxHPgCfufmTRzmJlCEcdqCF5FeuF
q1cWC2KKaq4WnAqiEGui1n3ufkS/q7F622y7uQnipaea1W/IP8BJO4fxwFjmJBgMtBP6emxH9C5F
FcDt/lBbxz3HfXbxUFxALQ39tvdCGKsf5IH3JJVV7DQFE+tLmjTBop3QMPwIr+BkH6aYOubbnmgN
0Wb0b59Sxu+xhfpKABYFIT+B8KjA1jJugg0vbPwTfGeobJzgAm/2bweqVSOpIxh8XH8Lnqplmp9R
fvM6aOjoQpdVXcB2lubbWjHRML8TybTw/ijFoF3TAhYMb+Ob1Xpj/sEI+DPsrnmPmh0B4uu+te+s
Pmlol4reriedgcX0pC6NVFc8quEyfotYezNSUeQbcHWbumyb9IynMJG4RM2Q04J1BW1OHeKTev0q
SA2BWPQ5TBRFJwxpPIeGlNGY/Km0we6O7+H6rUW7ThFO8yILPKiYXpmxYUylb/IcF6CifbYSYgBL
hp7NlzQBQOQvthzkcU5gHQnHQRR2zE2jId3Q7lOLLHP82COY2bbti+PNQpVm1xFJBpgMENyyKei3
Tc92XuSmHSlK8uadl+Ho8fO1ye7w/G2GrSC698+AZzco4CdYYMZGdrU8F4gAfdYC3FnjX4HZ+Ngf
HmGygeD8dpNwvayh0Qg0FmKCNA5TKOLcIC9lIExg7wQk8JE/+VeSwbYop3FhDeyhEZiPQJK0oyPs
Yha4Z1MOhHRPyHIB00ve65k39L7vo2T2sN6J+WBPayrBjLxC10pJtXlb5yMGWStDQ9Z7vZZpcHCx
SuouLhPlztC4Q/4izx30r0hEj7oVvRgmVd37WojVnRXR6uU7iwl5pTME9aqMfE6UW7/aPchuDNpS
kM1os4ohZau5BtCIxBl42brfoFJ/TGAW/tnla5Sfo83tZP9In6JNScza/V//8JtCLNy7OAgxPZMi
yibJ6AqREqsnmiRnqVuHUfgKm4KwsKlhfxGGIGDW7wYuMHsR6KB7Ghq+/Bz9f7h0Q/mDQ8qXuiZT
pAolr5VIMK7hCwHGGv10I2JIQYmZXDCFfL3ERqhau8JFIQDQ75TbkCr8xvidb1TjDL4oQmgtlUv3
m3vaVEpBTKXspFfLqOZRKFNdSL4eH/f1B2zHsyTrCFZNzlMla/EyllC8QUdq2L6IyXwIpoeDcmNC
erlsQ+8XHikW9Rd29siSsJyQTAAHZ8SJSiyqAIBV1LPvQtQAaMlgMix9bNyM7wjuwK5BMtvAKRS3
9U8YbOsD1AgOk8aCF1+Mbk+ylXHJvKhS6KX1Sq0kjt4DJDQ+s8eToRfaJrHZzvMkwJTqB/OEopMM
E2SLxHZQG5+RM7XsD4zWCqohMN/EbkwwOXhnO+OxgllCoGYR5Y+1vm7dY30LPxUzh9f00S4xpxoz
W7b5CIbq7PDuirw3Idl7Yo/H0AuTVKEq+LKyOprjgH3CHbbXIjAixkUOXI9fbOv6CmodYKoFBwsE
VJBjFvlgMhuN+Twtv5xp7g+ZeJ8IPcdi06nanwPlCYZjFazzJVOg8MgVyNZb0id9hQyDPaHpflrB
77pqh/o+7vAZfs8ffzXApkTZitjgT7k3daSlxVd+ehzfy76a9xR81WEI0UicnizKbTjlPkCTuJmP
4xrI3yXOqgrzv9yLi4rTXxZtTIc5MwaRPGaYvNblEWLZbpi3+HD7rQCOnQZkbW1FLxdYpq8vPy6c
aCL1oZQQzoHezBOnVRKAvvwVzU3wXUx9dcaiMHVfM+dl6ETZhkvqg8d3Zyo+CI6wS4Yaihw4fwdu
UR6J6GNDWPgR4tdUgYRG38ys82Bthuy16lYq5/HT9RlLIaBi5qJOJ8dnvsG4Un72lvsW4eMzjYPt
QUdZBI3ejaBQba9pYSq5Mef8bSMfVzvmt8N7qzOhjghI2e3s3CBOyqqmZGGpTEnogd+wPEbtGyNl
OyGbocaupTQcz+J40/RbaAWtYKDQp31Z6UBSEGk7jnHfAiXyLrPSlBs9fwdGnLjgATtOCpXexDEn
fRCHOgwDRM+QMoxMVbAs2dgvm0ssYMNBHlZaUW5HEQROoR3INiVBBADaMnbWjzuD4XTwwN5SZGZG
3N0jQthOgDrJUH4tmDRzmwOoTW5UykivQbq9KiQFLaTJhjJ7ic35tpF5qYmU6x3e6SQlrwpRIhf+
hBhqcHc+ZLjmBMt4/ZYJz4BGXYsIytpRAFAS6kjWSh9qknuBhTzHux+snAwuQbunQ+y7n04VFkxM
isLt69T6UPR90NESK7+IWunFnKWzSOlzs1qNoI+lICoi7tUxq/JwUOwANqdYyIxnLAbQuWaYahuX
75A5/tCIJIMt7XxlnUKSe1LMcAelSaZByw8sWDK+CVpRs455gdl+4LgF4GY7NoqKmd+QuOPugR0l
edkaa77OtcIPmP1stN3F3BH4IjL89XaUf5PjkvuuRYnOs/lb5hFQNXAK+AiKqvTI2i8Y6JXP1l7I
Lo28uXhqn5DwsVyKmSKjrNsi0ZEs7Ts75vFQXetSP8YFLDKVCSYTg+u9e38PZkKFkrqlD1Y64h1a
BE/PZjwWqw3G7ewRA8G8C9x2AsDih+euivjBbQJadTjDNTl102c0lqD5xAdjja+f7uA8tR8qknca
jCEet2R+aQqRolW649qSeISLkS4vavC7s8miB0ZQrHRomFGpHckGA2/BDVUL2ggeEJB/r5EWDA18
aHCA4hPwvxlYeAswRiZvFZm42xg97KpYTIauC2Yj3Lr+DIoD+MpH3ciAmkaPRWdLj5lxxN16nDqt
DdayeFaVVShqG9POpuUfrDsHcaLA1IXd44S46NjMMNp7gAbj4xYaeYxyAB9HVP0+EEaaIaAi0Dtg
OPSLtXFvwvNi28TUW7zWbkqIBwBJcX0L0Dt4n64UzqGjqSQQOoZ6K1L48J1EyX6lnn576FZZKjhe
w1h6x2aIR4Xo57WxHg8FwGzDdhdzlHMlw7bJX4J0tLoPpO/XLWs7XWDxdfaHLooVCZHZlY/VKHwv
bVsmf3d2TFHKZGrXf2T6vGT1v2rX2YI172cw/GOQPpnq5CiUm2B0PO0P2uerXbyRDUsw0RF6Eys5
uTpWpfNhn5AJROJwDfgnLTZJTs7A4S5+S1zOkt7TSvd5u+ZellNE0R8wPbC4qDROESqcxGb9ewN3
bvVuKUPOqBaJ18PzklFH4ys4h2fUhjn4REaYeLUqKo3pR9I6rBT0R9H8nEjhaWWnpwqI318XWyHz
0VHtn73rOsq6gdJai1WWuwx5wpKsM5jFxVVmCJnQyNcgzRolYByw1wexqIapLOtlMwmB8e8XF30v
mFzV8EZyW57uWvy4+AR9ToafbG32wGuRQw07LcnkKGPoYMc2dzthy0a6i5ZUb2iawMoY8RJ0O5+a
2b3iE2ASuDvJEmO5I6NJNXWTdoSb0eB41v6zQ+9Q12iqJw/gOqlbRbAR5tmXFbxNGDYQZ+/LGJbr
ff1FFimdbR0KJNuz1J0YLu1rxt1Ec/B8xYafLfMACXa6Wxd6JYFGVGRgcgX/DuMeBPX2R6joHcQf
7pl5H09rAICPUWNJEjdCu89cgZDfqI+/euZaO43D9/hzQA1Ea8dDnxHlQY1Vm/fc/CuXggRRXUZp
lfAs/Os93ZYGT6cKDbb9pBeDXt+n3AQHPjHWiG+Ilu2J5u3OYQDsawc2MiIMRiJe5zA+gGtKFihK
VSYvnpGa5ofWANdyLGOxxQ18S1xFbS5au3f02HljaTuhUGPoSpu4a37W9TRbgHA1k4DqjxCLWMDv
2WCo6q+nvx1oujGVYIQm+8HUnyBLsLkTMr9ucdjZ+7PoKpr+MBYtrph7b0saBGPiD5q5zKP7Eth1
iqajFdRYNAIi12nqP6jhHt4GhmU6X5BASLWBZM5tnFEYRYMv1ry332w53oX1JDpqiSOOY/D1+yxQ
FcNVbTxatExkYsxkiFQ703Pp2T9SF4IMX3cA8Ea5uwev+D890QK1yPh95Fu1i9GjoasKQRmxU1in
Zq93LOwNMSMY4LdcxgPEsWzIFP148TTVVOQS/4rfAzSK4flq/yvjCn0DqXClb2Id+C1Tb2wmDRGs
VqFsKjIyCPSV/hc5pKiHxdLfzTckZcM1Y3KTBVmRLXJhbRCifAZXMqjXMF0eMXF0TGh5z6+IMS7j
WUGkmAaeZebWoJWgg9xncjhAmfPwstAkCQCwhMRDhYRjmGPPSWtJ8fTMMq6kgkQcNS/+sN/PsKr0
DVJ+9MlR7eXDwkRX7yi2I1pjT8c/gme5ioEpbcbNrxFPinHq9FWMt59hMuKIZR5fIk8VxYRlO4bn
TVZ+fGAfFebJYdipS3o+y/8U2TEuyBEyOlU5kRB9YhyDDrpKzKuxjzaGT6LniaalJ2r7FUI9JJMm
KiCPWXpvSkibnHq/mQUO8/wQftDg3hPKOMIZlXDRLORiXBVfnq3eARDQWPHsB2GlM0ub3gvuDDzh
U+Drv5OdiJ74J/ulZORziMmBacJPqvaN5DOA6+DnxWl8RvO8cZO3URctzN7WV3CxzH023Gy4+OJE
askSj1LhVwqNWDGhs1yu7FOAuQXHm8fr9TWwYCL/yrJZd90y9SHTo6xsQVB7NR8iZqAuGBRyJuXN
6oxCohYFf5B3IGdQYkYPyX1b/h8OuK/wHQo4ZuDc95CWuEw1W6QwEQEVJahPD6PAerLSUB0NAPkf
jym5t6FF+LTb9tK0askjxJjanIaeDCUPk91ac6jWZdERsER1aOCRlfSzbA7I+yvM579z4jrRHlVP
MDF+7f9f3p/3yHaYVWNgpAXeOwVUKzxGgwPX1IsUVVdutt4OwsHMaC2FC5GO1uhGyyS4/OjjG12k
GgktBULm+mtVdpLxfO8WDvUPI2jTZtML6sJiOZUQtfgl337A4noM/frpBSwCo5motEXNEnltVoLr
QOgfeXrcIDuWmuZyhejjpzc+zYnzudfiKyGnquHUetmaQ9z5uW04/YFhsnk1NNbkecn5KZRJRIty
6YCQNF4tbq1igwll3h30Cv7RILReFwLEm7QasAyjtAzcsGobLDl3AFrYJVECgRZffWlGIrcF/qwv
6BeOUtIjDVJIMteWOsaVIKzrjY7/zlyU5gystzHRw4OxTViEur1vGGpGN2EweCsHBDF40cEm2xkD
C8vv+cdnbQKktAZ6OinuvCgRwz6K4hWO5QRQjvXqNz5xV1dFxgLfj1iiCLLAz6+wy7Tp3Hn3aCvA
XnWUulVEL5S4HGuTwkLP+to6O8SYmr4da+cZd2Oo7qzGn8PoPutgne/xaIfZ25cPpogAZ3fYJJi2
xpoM64h6Cf9gzKKnkSvqJOlZIsxPMMbJdI9Zq0tsdruQQLrJlFQgYHlSsg/iwq3b+pncQNNa8I7+
cYlHQf2kD+U8qwOC/k8uf/diRKn1aDednIEsZrPfqFURNfnGb4CGgN7fFp+D0dU+O3wtPxgyqUzw
K4MuyolshbPbGj+z9C3JATEfo/8RcxNeTBvPMehZKPkedVhzVB13fwjC3pKPoYhSZMsZ0iUPiEb9
/Q8UIms84Y7bnW6WGF8YQM2oGqUC6xeHgs1QIRYhKFLocO1NWk0g0YSd0Mf06vlnE0qi60QTiHLQ
uC/Gnu4h0biHWLFMER5VXXBH0jfbbrQxm3vSzDLkxyELi9a1dDeU7BS9LMCy+Og04JRh4LZkgAW5
eYBxQuBB7wq/FE60LtphINIzczyQjoJTjVGKnXdgR7OVWcqZrG34Pxu5YLqtyot5QBw/djw3be6X
Wvv2BIgiDesJrVFnQb4nW35ZxpY2QhxbUSi0t2QHfb5iAvzB2SGOKxII/0/sT8IVavHWxJg6tSOS
P2MDdi8BxnWhfNar5Dg2xRepxtIuxRKPjwTErNyVZBoS6pkL0HuHSTkBRlaeCQmKxXEf+mBksXhx
rdRC+VFmXk0/vgoXTc1yO4rVZZuOs4pQv5IxoAyhNrS+RLMa/aQYl+x2bKPp7FnewVA4XoGbMZOy
HOGPsCg0LVCRBO6VPhQtn9Hayd8cTa74lsq0yKZ8Lb0En09U0w0QlqKBJVfefinMspB5AYUMhhJZ
AB+kq8H0k0t4NiOMVVBnqABnuZbqoN1a22MeMk4zSmSOrCFnu6juSgJ0HOc0EqSW3rv9IT3+ZjjG
2QUw2SV6TXMTfamwiXpvJnbtHOtRoaYJEhK6Qb27FgfjP/ni6Kfsq+xAdB56qJj0qNVmY/fsaiD7
ylRw6EJNeffYeg55OcPDB9nwuoZdC8c+HiJo+UYHQcUaBRGxv4lv4odFiMwxZlPbHi7SYrwzC7K7
rrC2oUKaiJZ3dkXkY4stpOquB+RBot656jWbPdQjC7516eLnwiL0sLabL2Y3H+nQtYHe/R+oAGZY
PXJyvc9f5uSx8jpiCGFm4VDDlqp7YBr1TisajuZdW3CLID5zlrPZE8+0Gg+xAwIXlC3BegYTxoo1
Auk/DEj2P9DUqjnvWRL6HfjdymHvNM7E0JXcKfa+N+roj0Yv3n8/JtX/mqTJMDUxy2LiuU5tMDKI
Ae1WqJpMmnCHZzAEhGi4E2SBVbXJVqoZEF0i5TCBqFly3OJZ/A1s/PtSkfTtgvMzlxfpBbPeyeNS
245FncOJdJWBs/Eneoh46pLW12WuUTJYGIK/ZRL2bfV3BHIdAycp94pBEPLeHP24aUblq5VyD19R
Nf+jUU8xB1PpKjtHXWuLeMvT6XnTXOneQvTwB1t3JjQWI/OYh03AFwQebOew8V3Go2GyuJCtW0ED
SObX7MlR9G6cwE7vYupqnMickuWJu5NTNnHg3iHzyb/Q0usorZzFZt3u8wRt0I0z+ycZxp2PKScZ
S/XHxy3lzcajOpiKQMj31ohjA3moI4GVnzZ0LVTAeyqYl8OAmI4uB6lDxyEhXmjkGNoiC0UL+krX
f4idQQkJFPbUAxL3ZYxPs/n1aaJl7VmzimjA3zqRhtDTdYnOP0konr5GCBsVbeTjuZ0wZeQhLk4V
UAEf7Q5P3Umh6UPfIgDByjjNRgWgpmIc7VzdTAe4piyNYyv5Dsl/eP+xw+YGoE/FgxVscla0JVLx
+O4TwqfkIiGO0sb8S+TJYzNsXkjLyuhkDcyn0quYTYJJD0weiuY/e/vYzOH6d0OHl7jIyYLsp9cz
9I78padpwkZEYLbWjU5J/uWDL1XC3vb55NO7LjjcZrG0mo+eMIjEdupE8rOXXyPlGAvmUFDEhTlQ
EokA24WilfnxiQRQCrenbmJBnmUnAV67m6oNWovI4T4Gr5zhA5rHBBIrTchwb1XHYppw/ZhDRxXV
viZP49utckRpxPeN0TGmxMs/DMmTGOhDbOOEJxVhGdwW9z4QrClaj4ufauAeDfknX95zVpk2Oo7y
aRNnZKj2aHDenmFI0MRp8chghaOFVwUcLxzckRzJZvHRMl6k0Ntjjpgtp9BMIs3SB3luIjPLWlGE
owFLHdzK8y/uaRXvkiX3bAeDh4/3ab8AmaFe/d4t0o2hkdC8lKy9NvG9xkeELhew35czdMASYy6B
V2aBoXnuXmov7YuYpt9XH9ZVrz6KFhfAsGFdqbfixmW5jC2FkT6D+OuYHOZg+r3E9ORj8f19njMb
e3VaOvkP1fwahW1sWBhRKkJ7GgOPRxdCTixC5P513Mz9h/sCpoVzNLpLCt2g1JT7SPU/xgJ/J96R
tF6liFAPFmzz+4TFAw8+IlM8cVTNToheJdIzzTHppCqLGCaF4cRPsJgUVo9SD7oypr3mDwNmRWas
1cwKH2Me3e7E8lh/qp/fFIpaQ2CVUiz8ipid7i+LYQQ0tk5IN0f9YA2G8yFmk7iMgMha9z0sFu1T
ylQ0rvs3zspVV7nUzQ5swYd2pA84MF22oqDInXG8Z76zFs0K6JfoDUc8NvXlx0tXOJA7dcJUMkEc
vBU+8ZO+E/Thg/QItegh7HPjSFMdkrsNK6Qr4faH8QTwBe39r+3dz9beFOlOHd2dcQd+xQgAI2Yu
JX7elnWWe3DQCYw7hbWpLT938b8oPaTfAAy37rDJ8FeOGiBM6aVSDgXuihsfNGzNF/PlKoexEN20
cqduT5MnU/SO2zhIPdhpzluZAkJLpLMFC3qbphqsg5jBfpKDkb/Y9Q3K8HF0K839yztDmjWZPxMD
dj5PI3o5/3LS4+l7Yve3WoQotV32eRfnWnfOmHnJvTpfgF65n81InNk3iiZ3hFSL1hdReU6pBkvd
aKpfFyhIE/DEoFotWrKTjIFOSb6HjC+6dx0fobXr1u/tMrpmy4zPlDG0+k493tGZXkhgM2shBdsf
y06Ejvhkl8HGNK8WRsNW4n343dPTs3R+Oh7DDttwoM/xRxv7rGT50/JanNVp9bOrk8kgY+uerb65
7JLaHLKbbZZfBb7gcFiCqoprnevAAcZZ3nAJw4Rnprccgsk4oI1rGqewCHDEVI7qAT4uIU/tZrrp
wUF2K7MVGttXAQOe9MooEVRiEsrrUxSKjAcMTTZzUAF2PIPqYmBCOxpWnYgqVIYAvTzWXrzLfRPb
zfEDdwxHxNdlCRCF3JfASbKu3n4NLiGEPrCT8qO3VCBeo97zRtnkR/4hLV0z18sinZSz3a4J8Op3
WSxmd1oO8sJ37aTADBFmxwaCA9NnNXPsM6LCHyHZpnzv1qFoh+9ntiZh7dtNWq/zwmUnv+gLVjXZ
awsB4Fd9aeFVUXTPwz9aq2mtqDVoraq0sZzOCdQDSk4MusBOSWLG0BCFiyHr0Vasr5CaEqICs91L
mBddU9WOUhYjk2cLS8JntaaZv+hr0QRdTWa21A75tbzVN+0M3rVAt0711llnrxkOKDbjTHpPthS8
niXLYK8aOqGVkXVzlskYfv0KzAlYLwfDDmFUVHi/AcUayuBjPDMOFbZxlpAwXmfY10b6WyC5JxvD
XcYgoBr1ZJgorU0kbWfcnK6BnXOpXFH30VwSqz0E2XfVV0z7VkJPVIpHgemBQ6mATE/Cku2aXdfD
+pYeaKkZDjQI1P+FbGTuIinkAKszvAV3JLHmi+m/wrLaDfHlYhBmBCvxJqRjNOxwKs3RpF8jprqc
X5WbIO+J4Y9VIPjAsfcLk51eA7LL4W1sK75mKeksBg+qctpzrNAxEtCv4V3zn+7bc5GJXiOA9RKW
s2Izl6f2TS6MZLneKn2dJZy7Ja7pQFGY7VJUTVsNfhG/gd1kY9qkc/jfyD43JPbbLQcwdkjOOz5A
tbLEK2/U6Qw9uyoiNQ6DEESf9+KQt0Rp7LAhr/G8Cghs/cd15fqSSZS4ihdUpQFoGTJo2TwVvCFw
rRwzPsQPMiqWccWt/2rIkwXhZeOOdYKZjn4z+wH6j1baFcBH+lwsYAGMrc4Rl1X5fH0FfTWCNxoX
wP+TrXgaY1+wcMfQvko2e0CjN8GYu0pK1rfEjEvB/zO9CCjFmBQlUFmbWmsn2kjKa9O7TEtMsmzE
yhZQrMubffEFF0rQi/Oq+8u/PnWVRfKrQMFhBN1h12NV0Gk5MzAKZailRxvfD+BgBNRiiQBECzhd
8IuVp+ps5lOaEwILKWu3y+jMJCqeYwd+or2lCgNh5uvXFckDBNNiEHB717tyzsUpsUoV3ZSPxCMJ
XQv5Q5aWSPy5gfWx81Cu4QZ6D8ujDf4iGIhq/x5WuQi+KVaiatfQj9XpcOF+T9HVhrVhcRJHT2HV
qrmRE7tqCmbaMj30m57rBm0R2hY7ICupeStDqqIAgV4hzF+LhISuSmbb+6GLSqqmSCYREVpO1gvA
Sx3pqfumMhTY66w7ZpXffaqLevlWRcYgw5l6Kqm6Tgj9BGy4fH7Lz85BnahEhbmav8mLFgo6CPkT
7NiFp8WZFYcoTb2XgqPNeeXCK1D6en0IvYbZ+uRkYv3MVlAX81XcRHxqjm3iR7/GEl+niVIqDejm
VTWVQZxFC7K1R4gugwaKCgo7g0Ups/bOlgLZAc4B8BYZvymPKbiaPBbscQmjkiCs1mikgo27wC2/
UgxdXclUsxVJcYMXb1acHnbExaTpoEQxlmo15S5aFzseK7324PpJd2M85OnlMLDti2Je9CKesiwp
nfHQ2DYte7mAgiR0N0Tb5XQq39SixXcz7Vlwuma5d7M9rTr7hl/7L9KmmT/XkkRdeLBMfx6c8z/A
Z5o+yt711iv9YV+5LRz0rATtFJabIA7B+XUmCuSriV/a25BQ2Hv1CIQxoOau2dIcsdDA+wVevRD1
hyo169q5WjR/zkZLsDL1n7ITOV9Fao1pBa8w75XZ0LbXKWCED+Xhx4LltWx+aSvwHYqq1UIIOz68
eMBZUcnstLnaCYyPdMsikbRvsgp8XYy9vtukqIFeXKRF2eeyLLRvvf0ZJRRLpgH2O1Jb1ncHYEiK
6EmPl9MYTP+k6lfgHMZiOtrpknosZwkaXZ8jKZJnpgXp9b9ngKnbGB2o/+UrDGgzPx8z92yK7iNw
WfRfSfO2hGDZ5DOuNG3+epXdRJzQRwNze0vmQ1KQXfyjid18xvGaLJfXLBuda4SYfLNwqDqUYFA5
qn+iJz7Sn4x75z+LE27Vq21jaBV08G+15NNGS4y+wS3ZmAC4BCyP409uKJkOF+mF/aXJmrP3JKx/
3YqaTBGffEpufNbJl0nf6M5/h5JxEDxSeVDhVrwmmrBYEGAsuZmC8xuAfBEiVE2oHhkG0Bgh+GZl
aZon1mvq3PxTHuiTwHXBrVx/jgYw4rGhARWlTi8umrxI7jJKzNKAKqByxfF5aRR3PtyzyKiCzdmm
5wqWA47y7lblQkDA6uRL1lXTz54DqhFqzTVNKKYs+iSnZrO5Za5hpyR8q7MCHcdQDZcIj+BzGmTg
QjeV8qmyD0JWQbKLmH9FQgHuE86EC6mUO+t0LA27esgFIsIzmMGENOuQYRJ8/wNaKFRZESIi9X21
ESxL87Z856EBQsRKdJbcu/IMbnYAoRN6nFnLZjmWIRzLtmzbaNHPmU36JCeiH8vYtBPmQxR4nUuH
fUzHNTHKyBQXlgkek87YunkAA4bSLkEcyYBKWPL+D+jfm2pH7bI2so7hBOXXOaYsaRrjDuOf3ku/
IHaOZrfU9hbiMfI0ZKhg7y8x+8DcLr/0oWyiynruDyv/JILvhX4ttUgDbiLTtS0hGXUguWqg0tWP
AXFh7yjjonROfOLDGWOWZ5WWCWUzCjkgeLziKuTlNFWfQPxjDTX0Oqhk3FN65254t5rVFBeEsRiS
a8CPugfymRjqmVA/XPm/b99Z/sR6NX8oQwPMCc59Ob5S0jcy/xloLTZ7z23B0jPe4/VeCCDAPOEq
9tygfZMaZsADXyWTAwBdezG8Nj5qfJaapTknzf03ceSaS8JWybhLhWrsstnOgoNTBAmtnu7sD1EH
Bxj/zZu63AqENMofQidmLDoRxvBuJn/wArKWmR6nAgmPfxig1TeNDgsXfN6fXaV5tdEUe8hVHoQT
ZKBQUl2p/JaCxCZg6GuTEDGfTL1XVKfM3VRiWMoGrW55oe/FFmfJBjAwm/kBizkPG4pubJaIKCPv
UbRpZXwKtK7PsJmXW3xkYzgWkXuBvG017MdBvfzKZuKLKx3pXh1xEI8J8Urlx7byhZ0RGEb75msE
ZkU+JngGYMdu4dKqbZEteUcINC/YTlXaXVGHrOykvBKf5MX0MBQq3qLVDpv+dRjRjvXsy+RdL70j
iY7YJ9qf08jXd8ETv9Qfw1aFJzQAcSVIx5OnBxosMxJa7Z2wTmiVHm2iAhsIJRJi+fLRFFgEy94O
N6bA7R20hyDoSUyF2lJYGvwApAqwyaoWWvW0RMwe7tMTo8kCAdywYp9LanY/wyT8ZexseonXSxaN
AlwN6s7YkcnFQg6nHimwS3lAf4vkN1E1l/7S8MVN65SRuq5oTEeKZarScUZQZEUUs8tuqUsAG+Cu
2zW0w/94GR9xRqTL12EaBG6hsib99yTlpdH5FNAvIKsOR/Fhi8CukwCxJiiY+W5pQDNqN1OgsENA
Wd+5qmd7Vw6P8qct/UZtacjWXBEaXGk8xlzHJSeFqgsR9XscnEBBFs11n/SOjUXGHLDclRTEykmA
4EzLPzuNgVQsxZV5CjoqlvF5WiCrBkFW+ZNzT4OQBcMt+cV45Ki1r4wevtPjcWcFvod9jlf4dCdF
ubL2DI1dNfiIbLN+VlUyCbqClWkuRJIJ75dUvQjATE/bAM8n8DuKxRaBDflsM0mv6/6RqpnjHYlE
A8ebEnlhzr6DoVQ0sQnzdjVqTAnEQDwbCTgyUGeFWmReeBn0LAMMLuI8h57TtACXb5XPvMJnw56y
KEv0qUDvkEr5Fw/ASEneHjMBk6BKLeD1YWVafhYXgjXYb87mjDZdAr+lszK8+NAAk/K5WL/WsOc9
Y0oSmNn32QQTCUbXf52X/H/HrQ1tIGgR89I6w8DY3p4dKbCq2LI1Bow+eQhaGU+onfQ+PBI73vlf
QMEf+CHm6ctYRdrIXjeOzpl3DwCVc8rmi7jpZ1PUldLiNw2hxlAIMoTNlX8+k1aGySrmpHcV3XBj
dv4m4wyVlzQof1LZpaX2QN6Oh2/MvJd9FW/OoHRyO1CxBGhEedQOx+xcOYOMLBwUxjD0LHTCHU3X
H0/FqKocM4xmVBP/LqwiaevpoRkeadp0k3GXhQrk5hvku1+4FI+vQqfe7Gct7zI4a1n1DbT3nh7g
MctghrZ/vFttK6P+DNCAAiWIptjdjtmcG5n4g10u0wwC8fUzIpTlnBF2dAyebMXMrYB5EJW26J8u
upJLIMmSFJLcrkHhXapFBhFMQFz//9bgQe2UHtKqS4vjeQ3wLJr7vADLOviNA55oR9d65PuddALh
RmpMer4ruGUZcWu3eYuR5fyAUsHzWDWU3IbORXgm7p+JBQmQEJgNdV+sQzn+xQhl/arqEtSuhaS8
ceWBOEDhoLt/j+pBlPymBnuJapZS8nsMzemkyf70CGwzJ3Xv1NUbgMpEDHzmdbskw7JBj2XKHslL
x/AdlWpYYre5c3Balrk0ZBTkEeaMV1BQHUzHHmK6uMWGmZZ5c1gt6NMt+MQ2TPuQcw6gPGbQc9hy
SAg4ShLfJYqpM2HBWDSEEsKsfdVrF5+mtcV7bFI322lcyArNTtTVI5jeLMRLnGD2OSwI4m149kiI
jKwm5nTfhrJCBHNyrOZeMdkFuNckeSpTUTDNbz7dLcM0RxCqQRpoyBS4mIIMb+0Zcd+txt1Qj/Lx
QJ5Zv7lMywjh5JIXIyMYj5QbTXk8OxiEjXQb2PvUXWJ1u0RUDgbjhnnEZsmyJ8gBu5auVcL+HGVl
9HGsnQZW44MTGIX4IixVbaasH/VV2cNS56kuDiEn9VZlwluSrUXC56Ee9yDGhjHzoHN7CXLPRMrf
npydWkBR6SLtW0WVhwxYGQbCeVm/TtZW8P7/NljyWJOIYhC1R3nb28JxZwyULBP//f5uyNj+eDU7
PuSXq2080oH1JBx3fYKHH8Eb4GTKmAEzeMVvVtj24m516UV0qaIJ+5+txiFZ6yL839c3JooI5+Pf
w4VTfKutR4AzjcpNUuZl8CFwLEYe4HewQJ0Asyrz+XeFrSYiGQntXb76dhowuwdrHGtvZuN6DhAe
5Rl7CCsZVLuIbMKzsMP+d4eCNso6ffqd16GNCLaSP+jfMPJWz5ghJ4BQ7hRYycTE4zpCQnYvAe17
BjhA7dBihmiWgBNyAR+0n3T107+OBNa8s9HzYAI3urG9R6o5c+KKfAkBhuFPFMLUdjj6CSv4Evta
nfmZq88CuZ1g6V5XfdlctWw+Opu3pfS1NGvf6ROL274rrbM9PtbMHq/sTMptjCuE4nqMjH4kM7tY
4eauELfgi+/d3MNW3zsKgocFNfbOQUj3MPV6gTjvbdclOcYASGCqLhGVb6UDpRmxeMNOgwBN/nkX
eqQV26vhqFeg4ipBByTNqYz4BU19s57+Pi88dvHsSt+bcn+dxjEhquhXt0L4VXD4yOKpBcyFx+CQ
AezVk1GfZHtYpHNHa1/AOdLH0/4crHyOoODTP3kIunWXdjGIoYBLv3+6Yg5Qfpwijj5RAYQiyPMy
qn0nZJ9fKVPnat9E5z7OSXf4QtuRecIgaQ6/vPlBJ3mq8tWiax1n5ICkWHqawHx52Jp/rt8YInYM
qos60mrn32D6roBOgKqB7s/sAg3louNJFdfbzSW65rL+rp2EsJ7AF6M9LwKx6zHqz6k8wYOh4OeZ
znzNH2oGHYa19kLa+eFPAHN0FOVOMlSRDaoxsjH/rfNB6oJ+1fkDBAk+OWeg/6TfXKunq+hNwgnx
iGG8I5UUqGXPPVCzR/hwuslDOSloThZ+BPwGFK4iC+ZREWALkxfxqMiMKvy/0WBS5qfosfJIj2zM
jr/8rktxazYKBd3QEctmlgFNDpmmnHb5gRPAYXqk6CamSuZWcCthhYZktMfkX0Svc4XQcc00WuVf
Wp6ZKRkaV2lA6XeH8zkKcKXrY8FqmQ2/H2XHVQbP/s4L7CW6xZxcchYOj82nZTZY4e2sIO7BRWps
OdpIjPhg3WSccCy7eAzbJs4VIAlf86dTB66I6Fienkkm27Gf0fS6e467OuHR2INP4gdaim1jqTkX
8Cdejxj5yPw/1THoown834eZshVS5YNMxzSEHs0oa3wwXUy/s0+A8fPzKKrPZP4Wo6XYTHlg8kwh
AnYm5hxEXnLC3ZC/s7KnXIFjElcIxal98/wTw5eMebIAZGgTdSmta3IlaFvfy8T5ZyOFYi6fqpIn
gd/BA+FEoqZ73x4DjBwtFLiAKP4GmIgB4Q58FK+n4zn2ftNVKiMQfKaStbCIsfI7R71z7xIBdhLK
nTSvXTD8Thbqb3+UNpQBmzzYmU4L/4pODrh7RLxytJ1IhPkMGEZpSC27Qyvw9wdIc8UZlT51swlB
xWiML+/Breal+Vw7vixROW8AfRhU7tXyEVo6QQcLJsn72jLayvnhHtCRzxBczSU4mnIyPoW/q1wH
Wk6KmEhNKGsCt77VzD36vCt15ti40SzioD4ynwfC6ecbxIMU8M9HGCysStzDDh0x4Yzy+fyNr9eW
ct9BQUAZK1tAnZE6/aQTWskhDNINH8Sl0qlwulsBKNdufoTHkKvmURcKlmVm3gZQ9G6ybxOxe4nx
sFCAKRabscrPKdVvzMH6CiP/kxnnVIwEITkdxaR3ofgCHZY4p/XDjjoisB7nnsjIBMhW1LK5yBbL
mw6rK8/xMJ3HWMNr5G3ekpjkC8PTT6AxDLJjgLNQoRfZf6L3sUwLwHjKPWuA6w9bnpg4s4dDyCMS
6g8nAx/3+MPRJDh//I58VsQ5cbi/5YnFhN7GnzhZiR/mjoy0k41kMJ8gqtQxzQbBA6ZIlaavY3iD
tS7RdgSPBTzMDVftOfAIAZ/OgtbFO2CKTNzo4fqTb9i8AYmU4RzmMWPyi3VflMvBiRQxImc/3BtC
M6IiIpZgPz+IHOI3S0bkcgVEIWRHSm++ZekzyGs7GqDBNPkmdPUZZIOSTpkOzcgt61Lv0glX21JW
N2JSlN7E21xP1aEPtZWnfU1iSoq7aDASQu9tpZujtd3c/hyr1I9zolPmXRZGHMz162QHx0JzNOSv
n6i/G0Vld8MvudTnqWD+yN7Sm1HR2sQu5uqKLRTNLHFno3QrBjI2KMl+FjkW+b2qS3VWXDS4LVaE
SX6HqmGvkjErU4s2May1Jf7yldl0R7sJNMQYrot+K5f8On/ilQEH+3ZPeQuy5RGh1K7vGkkECEmk
C46hcWlWXrQC9Uyl+Yj/uGT4ZRERLujpzms23VoaRJUsjt5kNqi3z2+ZrBx54FtedhGubctneS9v
98he+yhQXMBL4JV8zFGaRCqLAgUFaQEiTyY+Ut93f6p5k5vKeEO5qDwMmuMgb23UfnIaar6GI2q3
JJul6eYOh0m1nkQUXlO5ZDR+FER9bTH81uaaVGdhfUYIDvH3dl4LqCggOWvCzyDxwLIl06OJ7tRD
GI4HTt4zAUVW/rKjbSspgec3fxTWAzYJ0lhjC/phYZJNBROGsS0cOS72pSPunyZRF3TsKxXKJjyY
rUct1D02zA+qMMOZ/3olCa/zEQyPLvdWa6OI1fzMaNOZRbeGIE/qvVihxK7HlusJ015wVaUXG119
1wAoJn/goGcKjdLRrkjZpHm55ikdtMXT4QjoNp82llU8j6fxPuUA16VL5kVCsg98tQUWiHkppT96
mTaHQIjjHgGlV//BYuf/rQLNZtjrjjaD48pfBt1ucqxyZQX9cw0bWwgnzuUWuQuoMGO3DXVOHDnz
/obhqTBBvKzfFV9BSIyOovvKOf5GidKeCRq2vPv5p99u4BuHwaNzro0NtnZoyZtWwiIIH72rsK1W
qPz1gKwc6D2grbrCV6+S4Fqp1k+Ceuv3ykzRMWORzLro8wMRih/yA7qfWQ/zFreYyjjGRseZKozG
HCIE7lM3Qsm7VTWo6yi1SEBw13CGlyGI5awdgAYspZLW/KX/DuhPjJm/gNL55TdhUtQEReVuMw/e
9wGIZV86GX5NMqauY+WSLTmeSz5/wdS5IOlBswzjCH/Trh62vQHNsbV9SuLe0bXyw5NYkuVlgDKo
CEwLKyZSg2ioB1RiUXNWT6Lb2xs2/MwKWsq12/YtzGLRWi33zdOvKGPmVrzspNcSHE9ZNYE+xpJi
XteydQ8pO6SpLgu/YkAr9Q+nvzCpN1ngI0C4/7R0+vewmt4YM04ApjnkZS9aRDrNEsQ1Ao7fXdmI
NC2aJ0Zk+BftsE4ljLq3uLV3Tw0sd8MArMkjrYCSEtlKgPhj4s9qMe5L2u2TEN1Fk03YxHCGLRNo
VVOh3erEA5FvatCMYXcoh4GnUcNcjazoP4wWwOvOoLFIX5f2yBe5LnGyIsXXldU9tcsUZyDUt0RA
GelbNELwvkFB4Lv5CJb0JD26M76LRNurQ508DkEbsadKZFJjOlLaXDfPvgXGiLlr0Q4Ce17WmJZB
dFRC/nT/vyWvLxAEXJAKD+78FMt/eAtmv42kYSZHLBEPtKxmVFry//SXI8TjoXrsJdRcmC+BBUB0
8bQ3aytjCY9YKesYcetUToocq5yPw8JxYhH0ojzEy6yiPHFki1SBL2DWbMziGsyaeGowx/78+9z9
k1Qn71T42v66lRUAn32uoySYPeCgiem130hGf0IiVweBBDD0hOtqYv1CD77/GYKyTj+Go92pX9j4
RCQtF3RLn+C8DyaehQRlBKDmpxnpCtlJgQmdcSkkcRXYOOrDA/agF2wrlFEmtNM0aQ7ZalNlsdWY
Cbq1sunOE1ZWOOUM6u23yrziCgtK8ZP3OttLg6sWhG31/8D2zrRY9Z86OhTv0VarmiMyqK7wf+9f
r8jphJOH0hDgNAbqVnrirS3cCzfQZ6wE1MXe0+DiSBnvitIVseM2KMVjVXOSLYH+9pfU43h/ac4v
o+tA7Jx5CSP5qJ3FrfwAliH6BkI+i/ENxamFMHJvuwua2hM6GIRRasTkfgSmtx1LGdLPLYrBqY4F
Het5kw6f4yEI197ZlJgdH7XPqJ0OPsl9FlGS+ZiRgcbEAxYBPlTtLVXnBZbFjXxVXjeJaS4TXWOl
qQCZ4Yx4MOx2UMlEGp9j2A+cv7s+sXCxR4trPREqo5boyKjp46ES4D/yEqd3recy37kFKaSVaa/z
WtHF6lKRBEJ6YS2KByvlJEn9M3wdLo/DhxnA/MES/zCw5pm2y6GYLYcUsUMMdxtWJQ6nnswMnOdc
oUNSA0cNAFq9otIEPy02JeOryWY7rNGfFE6ESN++Y5TfNjXWi0XFbPFfLaPzFujVFx4MBwYwOb3I
9uOB4MSD18Jm1d5gAYQJS1ZtbQoLsSj1ufLCxlsPkq7ANvKTkZjcYjGolykwQ1/azMV/Sw/M6bbq
0BjAaPrDsFHActw6VdSPEYPeX3x/5Qddyublqccfhkkpp+pgp2rg7Sbwb6DYxUJ49YB3r3gjVJY8
40AIEoW6agowMtXOe+3ofkhsV21OBgwu3Jv2Kvsj/GKUdcvEG710ovqys3f5LwAxKcSJA03qqdCf
9oODXHPR/+3pYgrm7yrympxAiGKTnIuk7lTh3CipREuPrcU5Z1jcMvYT8yS29pQhJmuBXa6pEF+a
VVyk14qx7Ankm5Qy3w+HHvD1Y9c/5SwU8ca1wm4gB46Xc6bUR9dUa3/W4vMWo9kpq0sIFoBoaFMo
/rxFLt62qhihkbUE6Pjuze+YvuLCYA4Z5DPgt/weEltk2nCQL76oeG4bp/qz9dqYRtsn310RDavt
3TORP76jzdjQmNA6/Fb6NNONhQvwGE6S6CyLaet6WIdBaRvYJk2lg900lL9dd5a4I4n/VruZLWnN
DGspjjKdipwvopP35KZqmKdOAMnGXvyd97CzRA42Mq6OvazsZhFn8+LzUtZfQIXcZs0rDN2FCgv5
W5E125s8WSXGe+yfK9ne+hOCKDf1lg5rec3JmafpwwnxNF51cVueyGXovtrC1v+KAhOLC7on/gnt
XW7wJhuKLnHv0xJNrvsbjw81mN4cbkFyBJRASAxGSfVkBbDX9cD+8fG3VDsBY9DELrrkLbRZ3GsD
lGbnHx1cYuPSE9QWi/Lwr1dCs+hjfu+lqaVLKaYAtFPwQb0VyB5esrwdXOA5c/yjkIJbpqhacmgP
LH2Pf7fVobt4AHSM7PKmXQ3wCVoSiMdofl9c9oCWkTyULs1O0kAO31Xy5DJ08UN5bryKE3wG56aT
WxReVCAQXbRxNo941/YSWYgTKUqv8qH2QpVkXomOQc2Up7SCckkttJADjoF06DeSDUOONVO0M+DN
BQwXI93UAhUFZtQmkyVCiSVWn4facaYhJuTRntFglEFPOMCcMT+vtyD7I9zH5Q+k7XSbnJ0ae2qs
bNvgYvIMM2+WG+xb0s6y70onUa2Rq3OtJ05RUKcRX0RkIrrR2xB4cjxsXuPQZyzUsIVMhETd6w+K
oJSOuwBefpgTO7/n78YucQpLA4x6wNVsjJYYtxry/FJ9pJTKyKySzm6Vkv37aRt441WnXxm5hdyE
zFC/Prs5me094KNN8mM9/PvTJkNtR9guq2YwgX6YecdSnDIWfQY9SeE21exGX6pPGpvMPJi89c5g
pvC7VL8yktojr0F8BIkbU20oIwfu1whQ0/TGiNphmHbpL0j3OFkHjhLppHGZf7awSO9ty/OhlNsH
Xh58+Sz+HagaHs/lbguuBoLKP6rYTVPltJ7AzxEUaLKXMo6SEZWQOSpl5Sumciz6xj43HeJuYDKb
77WxV710lcThFtWy7qSDdpJo4pv07zdlcLf0qX+XmIjm4fB+xlNFRqZhsWvEeNO/KSejtjFcvJX0
yU2foIQ+tHJ7XpdROyKRO8HPF12ahPznRrBLIU82iec2k3rxzClrn0e4G/+LM4aZnE7LWQLPyToP
m0SJDjVAoNZ4ZVJ0v+Rh8rH+FFsF10aI4EuF/kmcUDdaflUXe/BEkuisLUQjQ3+0OqYu44vBjOwu
XtpnV4yUEefZaRqryRSUYi40zWXYie9ZXw6G8PF1nYGe3ccNb/yua469qiYKjWgsfqXkD7ovwCpi
Fb83lSic0Qg400jyii2JlPTyGrceLc4p9d/0aLpV328LALYpwgIb6o/qvvl1TxCQIZ59N6c4stRO
o+NPBsCt8Fsb6lqa8knOdu9auOrg6vh4NhuUfbvOk8gaTqDHdhMABv/cIUcrzld6cf7zIOLPtoNV
/JkWZJr9+QwQNu4vi2lUhfBm4yRrOD3honhWG7sJEHtJ59BtjdWNuRdE014HkjnkjQQeHZSEjGYy
a3P9QhUE791aWYrttDCf1P4isvpUAHRVlgRwtJviDsAHijSjAZwIVcUcH4DNiZLsQMlkKYU/2wvN
//ux3CPqNnhFRgl3J3Q0bhmcm7oYL0Nkt5F8r4JSHyzBjRlD0+vdRfDQ7ryBsVbCxhrbNDFKoyro
0KZHLtgcYhlVqY4pad+p6jxASF7FEFzrYAI8llPpSbckVcg4vA5x89Hcnjm1KHXAEelatxo3ABQ6
SAYYne+G+k2ITBLCKtd37g0sm+xy2ETred+gv4R0a7/KmR86KczMBsojTHOq+Zp5kMaXhVLxgJO8
pjxamnhQIvgwuj3aSVrG0VW8L685OEUpcL6bJgIp2ucMDJu4J3sEMzlLEaieNY/PIxSWG2zuemJ0
pXqGDhBbL5wc1zUe45tbUh56Kx8LQDkNJk/aFWmffGIlbFreN8Q3yBL3ewH6KyM1siQLP8gouHPy
6YJUA+TwyDsxeq5LhSo/3zng8F8FSCLM7jaxNjW1UMTycKZAA586FnGpQEeT/JR4kckeGvcv2VJY
yh/LpT7gs6rsOPpx3gdWYihdCryk6KvH/QSPS0Du6WK4lboyxLHYvTA73GqqI02XnL0V5btrkP4H
rZrNQZh/dKVH7tM7q5OvCBxpXzcRZx8nr+ncbw5oiqxRln29fARcw8VShgGxsbGNKW59b38Q4Gb9
yzABqoVKPLGz8/53oKqYmXwFZQYWoPnwTdezIl15TwDi4QwuOqpkQtK5HOftHzoBvrE5bWuipi5R
AQh5+v+Iqn0/Ea/tDSNsfLMKt2oB8q9iSQFbwzQ0aH4UbwnPhyGptSDF8H6OF3Hb+TOODQBsj8Id
Z9cuArlgPUp7RqNtyLpbDdzpyi+Qy4hfJe8hBAF+2CY78Ylz2yVJaZOXYdkK5QbqMmsfiHM033mf
sBSd7yz3iVLHm7G5uwER9g1qLxQvIIgW0l1IDnjLWnZuKijxtSpNMEoil0WuqwwMMcRQwlWIgFCX
N64YrVENbQgfgZfHxt4VYjrPb67yp27sjslOUSbxAzcjbzogtqSVEYfWAMP4mtxMbO8qeMJ3Dza7
Y8t2pzbEXi3yDC6RTpgZpsx3SZGhpy2B7kmPLVHdcKP1TLMzulezB2Y/7b6dqyR/ndXh6WQYwzUE
XhivNxkBL4pqiu1VeM66o/8nDjrTY8+OGKluy28ffY/o46vxnjan/E3MOGPus/Dy0P6gDTeYF7F9
zCfkubbrATuX7s/keM96ihk6X/R4dph+zfGzCpGvNYrYxr3RMMHO/t8ExsDth3LGx9u6u/xsaOJq
EjawyR7UJ23I1uJOHTZYhrgIElD2Xo/vQHSBjVIaiddbFlESAYgD+KUi8lrvwWDhyHQFdYLSg/aL
nmFa/kMvQ+jkUyxeSGy5Hb17VGu/ps1Px6NqR8pYrNQyaQ8BVgf+9UB6sdi9zBFRmeur311WXcWs
sDY/qL/Nvy00zj4kCPtigyI8s0zu0qDiwXUBi+ts9CaOVnkoLyR5xmXDDwmBqRFI0DtYJMEpF4em
pxIOIONxXyj0mAJIp1mVpkb4zDpgwHM1FGD884FpnuIlF3GJoqdntsul15NjKGXu00y62PWN4piz
otP8e3rpMUcfk9nH/veyz7qH4+UEUs3ZVsiGjE/MC3neZ5pyW6ejwzRiRl8qm5SB10GgMyRNF+UT
QnDOHExeyAfpPsB8h6BP97wmded3P3N8mUdsPiIRHeXh9+VwR6GJEKhN4M0CSc+UHjLSADhaVpha
Jo0aNzYYbf2V9ZLvoAJ+DOslR2L4VbqdVy/gytoHWPFrUoG7fyV6ypMdwtGJgntm7wf30heXLYsS
FgN1CxxvP0D+QXH/Bfh/7YmNUxi8Gzb0c6G+vztuot9s2DWv4QlJtU4F7IJhRR3EcKupO0MW42aW
fqLwCgYBuGNKqiEYf9VtqH3ccGWH/5e5T4nZuVygWFIg1eIC3BTQSdN/eKBzdUzwtdxm4s9XunvB
avuH4Ie+YaaverYx7GjBsJ7loVXgFeIuRoSf+sMKJfEhQF81krBoJvlZnAPwvvfyrxPIQY+xWnoZ
32dE2rwDR35r1nkhxAem0xNyHLQCcQHDoPfCkDgQHlwvQfvsvnaXaHBx7Xo5eNgQHeTc+zXc4jQ5
hN0qToxfj60KxX/eVcNR6swdASnUKyRF0t84hNlqGu0wfD4GexIhLEvNB7enCyBxiEYcgaLpUtZV
yv8K9hcDXfQdYQ68JuHlIeNxDEACxaCUIOohOhW3EOlKV3CG9QkLT2fkSqGCHYx4cCEY22x2s7Ux
y9MVCWMHsCOT3CXjuaNaIrkktZiUi/A/ynbdFoRUfuolPFE0e8EKFVrENoEwxLLCOrTmm7yOeaZt
3DQbyJGF92D976tyRvA9cVtQLEVhLy0cpy0kPS+boTv4hFL+poKa1NNAEQe16XEjUL0cKuuERTPW
C3cMsRGt37oiLZMV0OrkOow/1dDIEwZTdqo4FcXReJaIa13NZPNzCnobUVyfwki4jdEptOw/+Nee
duj4XBSlfAeRL6yetgl631YcGh0p/qvtjXcwK4Rj0TNGlkufeD1KVL6e64NKOaT1Me5shqjBFfBN
TDzAe1WxBg7+XJ6+w2kB9G/ULCa5jVakHzgUizsfohg6ChFus5lmRHzRuqp+jadgb21DTf2LlJxY
XxBnAc+WRJO6aEuX4mZy+ZwZN5EQeriHgY8EODsA77JzOXj4SXrcoH4Ixo+3AUcVdAADNkmI5q/t
7OtOz4A8q8VyG48aHHg5qSJ2s9awx26ZoTyP9+Le23KA0k1hYzVaNcxVIDDXw3x623cPgULJl8/K
+KnQ7EsFeEbEqyXU77+fEWG2V7TSeVXA6QYKLVZeoHJlNuJJ7iZLSU/i66c+ECGW7EDQwdVq/wcP
lZSBKAHxary3KuCaO+5ifV01HWz5DOBMTK6SMALJ8L1332G4lnM/DL797ddiY+D5BxvfzxBvofrr
YMATLQIQ7YCf/GP4SGlwAIy/Ct3RQNKCyn7SIg+1B3oBYT9/dpUE1EZHNkTzf1622oQ1oZ6vCiMM
oa/uxy951QjgqATVM/HrO7bnKrJPnGtdwyumVDfYBX7dYSsMVJMOME2dwibMnJ+X56WB74xBReQs
WB8QZbSPQJLoGos+lH/SJ8leuL/ycK9OiLKxzvy277A9gHD0DIFnxP3cXqugTvL5ZPQ9wXEDYg7R
nDUeIMRxnkeQKSO+hD5+NyXAlOkJTuniOApqkYJf0RnDj2WbkFzlgUCKMW1BQvF4F7YwjmWn9coZ
Z7yLKwlTaSzhAmIHRArfRy8Ul1YSdgkjff1pZCKmtmEXj80BLjy0H5QPtZofyT022fT+efNHkzpw
51dgkzMn4NrriWQLmB6wRrjyQWXZhX4LFMkjAXoCjuFWaKRAgKRzTwby5nYFwbZriwP6zj2Poc96
9Jlvi+rzA9pxNVcW/mj5l4tbyLvI+XyJxN/ufnpwnr9aS2eoDZyuj3AnXGKG8VKXEhuDenwy2htF
sgbFP3gbAnGFeOJYe5SIFR3CGPeK358pP4N+JHmVKxUPdmOMzW27XStfYKmwD10Mm6EMTbH8V6RY
k4/+882DcmB1R3CegkSTcbw/ZgsEIFCInBpk09pI9hKM9V3OSklE+nNi7zxOOLvo5NN67rFRdiI4
H3DzAPdKczbbS4LUomNlUXZvhr/2jCjBXI1x8tEv9atR2PaeDIRetzgDpoZyHLFPLZk4QfA85URA
/0JT8NvmdokkN8SA/ERYcwHmooSu9FNbfV8e2IEH7AzqXDNGRVa/tWh288WxaNoBRAll9NTkwxnO
C5UZ27Xv44j2df/Az08rh3ANpqA/r2sLHQYSB8gHHNacbnVw6Z4yPkHxDzmxzGEZfWtyacfT7Ib5
u3CKtKSTIcsFV3XjJf4U9D6OK2+gzulm38GCOYTUOZLTELv/FLlyHl5x82ViOKfQgnj3qOyRFwRt
7lH5GsLRcrPljpcdxWU1VBrt3Y19qORoadRx3Yx8AQGfV4ag91J14lPHw8yWLZm0itDeSV/dWFrv
7yBjw2Be+G+vA2ziYB5Ok6alFmzQ7wmOz8DZakYMis4c0PtaCQzyrpB6x9Nmq/lQfWHMMtyihx6Z
BKU46z7/hhTMd7PkO+CByr4oIPgH99URGraeCV+rsPkMUpZpsEOizWKiIkZ2LBN5s8i904SyTPQF
NkL6T9EOVo0kw+jpBsiOVaRZywF6QWgBRpM2nbCvUnBzwBogT5oN/U9Q7fAtupPGRmCw8JVfi069
N/7NYZYcnWxjxqbn/nBYcbsC84wLJhvL2b05hRHXfDTAVMsfUlJkconZNp8JWsiuJEDugNSQoERa
l/poCsOrQkWzB4+wHK21GQxxKSzaYcn4jLK7e2QpqwwEJWAh3EcebCHg2KckzKn+soJcWHQE0T4S
cqMeXc+DyM9164ZJNHAUZmA6VXC5F8tTOY26G+GGyJuW20BpAcODLY5CkcxIgOene8AKCaPSovvI
yI+dG9jNlPewltrSBFJozEbd+modRzCt6U6Yg+QBR1itrnX95dDgbMuO1XmOI1JffDu4n4Cxi59a
hzfn67swkjRydajsRiFooavgH4yj93BIz4UiPNbqkVW8x2noDPxSgjEv7w3kHMg0ZknAOXjY26Oj
7ejxLNRBERb4dKx19wsKQOazlucs3nijgEdZQGnTDi8k3i3x3F5LsVLnf/T7lbtDJSpPowuCCwxR
VNeoNLwZ2NSlW55/ng1INWiGzAZXHTU8dBX6yX9wvbSKnEIdZtE/F4PFpF1luOsLOoyIX6/S5ujD
CtAR5eunt3IuiJnxf9JAkgQAokv+Eq4WTukzdXtZo4hOO7+NAKqPsLk/I6KTTFjL05bk3UHQY9zJ
zzMgwmwf/xiMeb04q1VcU/7t0Wg8PZnlAU2/wLbfM/+iFcnGJLBqBFmodVZhC17BBblt2gw0Maic
rRl/CY35ImRbViIhqFiPhrCnXFAYhTCEoEWkr2iE+w0zJBMWgSrpk0a5b44/BwkMt7EJrCymLCe9
HeogcWItqATp0adpgGrco7jvgfokxZZtoA5m8ecWPNgbhik++c06u4dHExrW2VNxiv7FlehyFg+O
XVhs8XYi/N4REQI3w8UPkVh3jtykQLrMlTkgKI48mg0txxYEN3ZYxs9EzEdw2VyBcK0fZTms8/80
1PnzvzPrGl3y0R5QEl2J9/aQxvPyRaB7wwnGjgC0x6yKol4dO3paoQv+3/Yzn5WEA/RkJk9a5kA7
BxUnGQH7auO6SKA8pD4DHXrNFtUA4MFFJ+P1g5NvDA6jbSFM3lQjb3kVWcmw/0eecUzerlKuZt6m
6bvEpdgn0M/x3AX1ORQYN1iAzOXp/40u6NxCQoeBa5b45VmTwsuTGdvC5LwhGynzNQ8aFIL3Dlzu
orCdFZ1+yeB+8P/78YHmq4cGGnNs9ZOPEEeTnPNdeI/hKWBKXMPq1eiwGPonUCWVtRTmgjHrDVNA
NskF/PLjUV0XPkh/0ZXxWsAiKiBCx2Rr8Pe8lRs23WlceaTKNYCxSXSf69+6fRlu1/ze0ZK0SLPH
CVN5OYBbCIeDnJjZndZx9MXtcNX32b7l5rMsv3FOk3H08QlxEarcSnbZR+4YeuEDwoMmfarWxiy0
UkJ5HLELhacoSds/0hrcXml234ppddJ8etxb7YoAFKzqWz+OpsltqOpZfFhdtcFQW8+zsYUtBjUl
zZtQrBCmPmtMO6S0OuQtwPFj9TNlcDqxO69eW069JHNrWuzxIMV+IVp5OBER1Xjh9HqJAZm5dJwG
8UzatCRgPo+2byCLQ8IptU5qI0UlmOliDYIgydFRfBjISzSxRh5cM1jg4JqiLTRz48A2t+e5MGxb
Ce8vjlja9DTVstHsO29AN0/P0+2tvfKhRVELGozPuz0AcQrZIp3Y9TQrGurJ1bFx8z5v21SyRL1l
QT/55htIx95u+wXYxpyzySge6w8F97kJFSucHMXRyNnKysr8FlHNZUUj7LhiVI2EFH954yJR7VYK
ogGISLRTPCXU++97yFLrxVrvaZieJusbBfvP/sBrp5rVtkem14Gu288Nkzvdl30z3gee/GTh21YN
SSOPG5VdtvvpzIjdNUK0AYkzxhPINwlZUfbFwQQvMeB9tpetRSQ/+sq3hwTtew9iWzaNizbEwrwq
oKGZKAJtTTfLEWnpPr/lEFjdIgvKzAty/W74TV+kMQVwCNF7gXrf6Yy4nb/VJWT2bhnJVStHkTLH
LKVhUG7jGEzEdlJcNNHa6kVLDUnnrs6LT22M1ccfTe34FmADhSZbR16A5kBW/mUaX5hiU/tSwdPg
zkWc1+zSwOjym3BzPLLFs22un1oPzpHW2YqN2HZlgDVJDmEmfypN0Jhpk1po28eOVFeaD0NTfSaj
zBkcCtjwu2I1VzQlfdEqfY6g6wdkYiMI/g9fSco56KswKpw/4UMtmg9twiPJ8cKmaXjmDcV2MMqC
tNKtKYxNQxYovfRh+qJw6CQ/BnPUR0imdvPqg1YoGJ0zQ+XjhWeA4qj+w8CyV9LTKSDTyWNb+ehQ
w5UC7KZgNyy67avsmr0GG/0zdTMbCgjRg3dXDXEYnSZ9KVv1CvoTWn8BynO+NZytCHTHLh6AbUq/
h56zi64p/fytKI8xv57XozM+XYq+JoMSaP2vL1TnMiuE6VQh88VKF7FOvYK7Zvn+kwHprm86rgn/
xHRfFKsFLq1nncYrAOqtwmFctWfTW7L/1vGsF6goj+KlSVnJ+HJbUwVtEEAomLdYNJPKUBUYr1BW
RR+aTfnWxvz9Ai3Y0ZBliLbKrgkVH32OpCdt06XGeThr6lXIQk0AMk1tQ0zAyudOWNDJvVXdPNoF
YvFd2ZAR2DGvCVKvAf4DlQrc1EfvzqCSCfVuukGNIa23A/YTc5+zRsZfaVJemyUTARegzMl9dhHa
2WACgEzhaiEGVbl54r7L7t49YmgiXrVtc4fO7sd+NOyYmdXMzlUg05mV3HkXtFE/6nU2fR2/CDgP
OWVgD3FbP94iqhEc38nKkZ9gafpU7mgV8Kk3lk5b8RoqcY8I0Frp2k0TTk9+2lnbXWKHCDbbplJb
mh9PQjv17M/xofh/IWUm1041y5S4RJs2Kp8xgav4JZC9agWycHgAwXmwOg5LhrE4YuldzaPXXt4Z
BGJ+DQROiqHX0IIcaSdCvQV659UJW7aQz38vQz5oI0Lk9XAF6/Yz/huwlS43JZi6cpaJXp041CV1
XXaRj/oRARQJTlb7B9Akjg9yJpxWJxe6K2rcVflXqHspof7OO+IOHsaCP/Uks0TyuhRgQHInXAlz
yGl4bfc+5TOZ+/jFiids8irjs6F+mn0Ua1jDL9arQTmTFSWF5Yl1DeBFKeLnOWuenAeWSD4l3uM9
Ycq03SAaHMhtHn8Z16OclVswrShFSlX7BDccrCJziUEt7a8TzH7MXr0yqbrnuh8g9r7hP3TEozxm
QU/Noszzh22D4km5VjzhcOEBLugVvwd3OroZKDWARsrXXsoQ2Z7FkyJ6mLJSWaWNe/hm5I4mdtLH
Ix8co5Z8z9ke2Dotzj4xNiZqu7QpbQOneWLYqgXQhqx/XcUVQ4QcxCH9pV7MK5zUHNeJ/lxQoQbc
AKAM18D0b5IwY9sKtio8ivjj1XtsHJ1Y0TyeofYWioQzYAOUWXe1IBAF94qiDi9gv2r3IQ0GKv4g
7yqGJYJa7YuPhgsbgiyQsbxW6rh6AE8HmP9eF9Xo/EKrM/CPp0u3upWiB8LQuUsJHvYCXxbvvdb/
3M7MFKOumfM45A7BpFwMxAJioAF+trFTxXoKO59sRnDm+jjHsdr9OYXNVOldVlpGnZeT50MY+vkG
KuP3DDfMYZ2P9W1gdYHSCiFCFL5Y662mxbssXFtUq8GQc9yyO/Zf0E39lshXZ8mthkmZ4lhNEjUL
u1R9yIW7fRk7bTfmXd/INcMuSdCkZG2IhHbUPi0G1HmMn5hL1MtqUutGVi732fhP05zRDXRCUTnb
tjdDAUsNuknLj2a1wzzsRhuLD7O3zcFMP4N3ZgmCVG78aakloD8bAj/mxTIHuM5/42O31dMKrMKh
4vPDogawq5R2VLgW/vF9QT3DKgKywvKRUeLJIyjyaXmZpiSF4JPsps87ZzdMCsumjUJkQ0KmRDqd
mplWZbnazERVu2JFi5oQ5h+lFyLJUAQqSeRp5zsm10aGyl2rPTcvAB6udRsbx+kYTlvvKvBiYuXS
mT0foU83tGfpBVAuUkV2IteFWxNyQlwiKwEanKkFQ0B8vHyxVA9xA34y0SfRqWtJ5lY3sRvGoLCW
XvDK2YqBTebqxAkdb2IaJgywmZUPqmT4Z9l3SUN/wm+H4iqp/U+by5FobV/sRRvSQoatJX9OfhC6
FsJes4cSxN674rkditz87oOKC7w8Tw2ex/AG8ylG0nV5nzusuLk5qaVYKmrQLxGgbmyU4HoC1u/w
7QTBphtqitTaeXdKoh+1y3JtIN4g+QY9PlGXFDSdGVdPeFzzFufnI1JnmK0Qm6LW1wP3ddh9us11
qygMviU0CEr9tYM7aCrtBB8y0UgKKfiNlb8STq2eYjQQDOT6I461LZXn7X6XmX2PhMV3xBvT+4HM
t0aBArtSUTEHiACiX6jHhn1Ap5lpef9ZsU8Q1MjPs/HE8E9qUgeR8CqAKQMx6NT1avFRNBuRV4SG
bFPYjjZeRvfrszfXgUyv1qmk0HBdFC+2QEUtF1xH69vCY2BLszl12hvp+6JcckYY8B5Nif0F4wxy
stSehl51LXA8qDa9dFi+J+EZ5Gl3GQcLBSGqzoVp8O6O0CD1x9EpzXJqUO1V4kgBkbQwAvKNU50z
1lbFRv4gg7TGedDbE10yLNtZqmnaknbxWOmPjki5DM7DVJG8MiEJuILCfoFv13Otm9P7R7YGI4we
30ViIhDE0pHXzEX8EF1uYEp78Gq+OIJNpGJ8QqqKvdHfbFHfB1e4X+gYdivj48QpbC4mgGOohbm5
TrVXx2fn+Y1wFNcyzeD51soRk34WQ1F+ktacMaQx1YePH9Ep/pmhB9Lwcpi9HoaFjXjAamtqSOZY
lCVeUecJkEANPkaHtB3Yc3nPJxm2g/IBGzvWG6KtSzqgbyYKZwhGlAoJbXmPOFV5Z/cqz9R97xiK
qWgHGJp50pseZetWvJJQKeMeRSpcrmYxikBna14+mXTCelgqgI3AaWimEJf3sUuPtmWHztN3UBpp
7spKkCwH2qbZt7IVB9TY4EJKs8D/liNKWOzWY2ymScobWTCRFrxFjV2Pp6BUjfxvb1a/wZAm0W+m
kHT1JQ6mhxC8m2Tk9NgoSeTG27/sIHkIkkNCZK/IS7oasyRDP0GadACuvWE9gpDmzDJEJvRGGUV7
6jyd1gxvj0pyRusP+lcB4hgz1xzesu5xdfB36rVpypGYBHuLFy2B5rYVUQ5X7BTa5kAqz+C3XgQB
YguNeiTl5Kl5euMnQUt/T3jNmUAAPzNLIm8X/zTsrwo2grkxkyPo1XslJmBtoOUaTo1Ux+XQkNeg
lFJLAKae9jvmV8YVC0mMYPXUyZMXepga6EjfavQ329YnB1Q+EdmNfp05UkiSswRknXfgGo7T2np0
XwNn2RwV9LfI2Narez2swLqiMOWn8qif+L0DR30PLU/smZYGR3iES17M4d62SNqNlNqh+44b5LR9
q4pezIT+/mSyYLCO0L6Py7pYqiJy8t2FFHVAYbD880RByCeS+cvoBQITgRjAAk9KDB+Fi9MgiLIX
iC+hRZLfNWMt5u2AmCPzk16K8WXgrfylrSZWcNSlnFLNnky4wAaZLotMejbaKyYulRx1adYqyRFu
HfMkcvB2JQDISJV52XuYp1BSmWXeDET1eHNaqUl8NPSKjPGa+LF8l5RL6Ze65wqJINyXxgzanTBJ
aIsaKY+PARExVnTBlzXsq+MbNCvaJi9fcquBSmIRtGOaKLDqZvBIuQDLZTnTLRb78k+AQyy/6HlZ
UIj3VACLo8tmiZDXRKgaNzF6g9vEM7dFQAl4UUBZmFrT6usn2hsce8uvZkkP4Jz7g4iFUkksARny
8sqMvvF0e5hScxtKhGYBkd9Qumo+jlZrWFStre1y4Zyfz0/sGy43nAXHinkxlw6ZBmrFHWMT+lJH
DOUuzc3lJbDg6qK2Q6mgx6WZaO9ZS0KcEEYDDaVgSfNtZsC2i3h3YJaJ6nojEwW5eE0Z0lAVjwRd
HEGO+z51tAMg8xzDi1L5Q2iB4pwWJq82dK0ESeMOsYCAISoVy3EA29SvZrWLl77UOLjwK4e0Htn4
R9WbOSQRhn1XS94dfBUA7fuMmyo+hMAT3BtN7Px24jBXPmVm4mwAwgmjpJ5QAKMDylRzxSpnt6lu
nRzh6LlpX+qoNYgpmq0F/DtDepWuYR0nULO4E23J5Djc9VD2gmievksJHmKDk/SMrCQgOKG7XrAk
4bDURr/OCEAgu4n/BoA2LHLM2hnDhcxXBnF/o/5OC+AyR0P+8feCJ8hYO/FnxdW73ywOnDEDYg27
6vgZ0URGJe0QIugY96zKat2uzIf8rEjCQ7M4PbHRWhHdCNjGD/mGflCofBxLMUAeZ6qHmpq8fBC/
ntHk9N5O1UvDfkgpZlzANxpvFg5r5g/2a5b+MLD+vFmhv68p456GbYOjtc4fXqMA3HqtymNtXGhJ
JrQobrUJhD2ZVHHkARqdAvZhEy8MMlSScNXgElhSh8knCvbRTqrX8BumilyLroH/G+z/QJX/Zwlj
T5k4oICGA8UkXe8t7+E/u39QroBAWHypM4/2eKfR+iO0gZICdkznuI03VJK8zFgGEOU31Rcqc+zh
okNHbYWCr1V/EEFnhOjCn2Ba9+TniByUkqGvSSRsIgwiPcuYF6hetPcPdaC337P7jQ8VqccgQfgm
W6DFiqnGNgisNkfDZdOKjazwpJz+N6AqY7Z07+Nx9JPEXKzmslO6BqJMAKpvc9A0eblA+CHZLZU4
ZmYkBdzad2tRIliY9yxiwFxrYoG5DQr3AANWgegoKJrEw/ri4K4NxGyj6wsju+f3uLbSJBHJAgBJ
CFvoOTmI95cNk2MsmkijDRujiHZzc677qOnmJlQ54v2cZKnJidqo0nP+XmGXB44wEoAQ7WEuxfld
Fn+R77wRFHG2QErQPULhCpzvXkhizk45Zm2co1OM577KZDhUovTH8hNKr6HiF+I12pZBdU82ugdu
V/TXcdcfytDHFmMfCPfCZwycI470GbxqpJBv7PaCkaCCN2870HI5qAPvtzSzPSj8/xLfuguZCYZQ
pSNqfxYMgbjLGVes3QQuhzkLsr93OtcPEq///tOuLUF8bBUv4gVshnkQ6qwrSV3F8vQ/srY4bPQR
s5kE9AHgiA8scErGSJsZzywEwHlCZY7Vc8Ma0pP6aHXICmw9muNijNPXt4pO9N1nMdbOFGjRDjrj
RjLsBkVyHPGINYlkP1F6FSOKQJz6+KDa7hNarcZapxec2BzsBhG9vv715TeJVgnyIusWrCIX1Xnn
toCdPg02PASmW3Y0j65Gh2V1UFQ/HrsVOcf3qPG5Qp6ighnA2Vh70U6yHC78Rq9dfT6PRNCVkc17
zS9AwvE9v1q9ICbyM9x7LCNHGe/22Vmkxlvc+6p+NBQw8R4UnaMjvviOgY9A7IZbmzt1v1rPVplN
Gm8W7FqV+cFrpGdtmmmw+276l4/9zHWjRUpyGVkjaIUDAPxRFyNSNLKXja/x2XcsTzFCkuFw/kii
1Vsq1LUbTvMVX4bbF6oLCCFfkxhmqlwxXDzzraDGqXb8GJHSAHzEkPybgsJgXfIwAAUlS7mjnglM
NzytCZMuTzoXNrVk3KCQPPySrAnQByuNZkY/Z9/2kRcoYsajPp4kiQKkbfYtiw9hFiKD8EYrqLHZ
NwjqN7eJWCHQccuIHzejqI+QZtZoeOgcUs8SFQBkD8Zym65YgoMyfPpNLmFqc6fGFY0JGJHVoyKQ
LU3C2+/EDqCfKumwbHWYXg/HWaRubVdDokALSyCy0WXNWM4U2f+1qtCy6izE521VKINshOJYnAzk
TNebdY3UmNaHx3eTTpumL6cJd14X1zH8VZNUyi8HsJJvnwKLjWqiyEg8pFeGYsIkWLQQq7z8iazO
KaWYsC2GoQjyE7iabdOWSTK6mo6qFpMPV6C8XXOCzACpmkX1G2xcIgJfiyAy6fJ4gZ19mDVQALUD
d69IQSuJARuM7nWuJw/K21PY9muKYMbQU7hi+Q+3SrI4Stv/bu7eq+SUfHHcoK+00SFjeAHQZ+vF
eFqd3TGkaxDueqCVo+uL4+8vnrG3Prv2KAB9d+mr69aiEKhJVHDuv+DGOzNz6idjglSqqcHP5Jkj
ZrSqOGwJ7uUQQiy9+q/9KqiLR2aUnV+2uKrVjmBNgZ0zR7wmmRdkHkLL3yoEX/XvX7umKki+m88M
RRVX6MI5Sf2Oy0OJSbBDCCApaJ2JD7ip5EjOmXfEYuCz/g7e+JMpmAyUfnyG7YSf05Catu6FaCbA
VIe3OyNZZ0NuASqXnnGfnSHtdipd/AD6zzk7hO/hXg7ov33op9Nd27pszw6Oix31nhZTfZwKT2hR
4nxh9cMeLDrxSoMtVJCGoxaU9kOtgkPSJJX+A+c9ADNDhGdykqbhTkeEs5+RjsJN8rV8kEjbUhN7
xj4E1HgvRTQbDZ9hnzMPF+9Uf24Af4SrXxYl9QRUHAfEBivmG/h2yqC4xhmCnqZstq6uxHDIG5nD
9zklHQbN51MlCCYmjhgwF08WfejWmkGvv8+EqSOlH+ufervZQAu6rEd7yZmqK3h6P9CEGeEoqB5F
W8bGGejFmjI9fZPG0eHBO8VwvOhXFrdFwu0pfAno0cJWcgleDMMeHbV5xPDhWDWwg9TwapdpAVAD
vGIbcSqJNDLL1ex19lUpv7gY3R6clkBRFLpg72Z2t89hc6AY0BHCA481CAQDomgFu0QGRupRaU7q
/n1sPcmO+oKrVeG46G/OGex0O7/2ZqJLf5GqWvOhEAgZcZm58aVhXz1gzWqklrOLSBLb4wPxSrLW
cZPVJ3CKZLCVnS+16KcgKj8FFeXWVtwDQoI9TotYm7nT6JQp43uCezVSPBH1vPZqzYozOkDkeY1M
YbOgUtjRHbhdF9TSDNQWeS8tTfLqTID9SnoemgAhjYGkRouYNw+KJ0uC6EK/s+Ir/TG3UFjP7b1k
kiqL9zShYO3lkwrGB3k2/Bya67YDqQMfU8poU2yP+pSMgHgj8YoTVgUEZq58D6kke5a2oei4/zDE
0CDxdNfy26jFpaT9TpfJkwM3WmrAnfk6ElBPeYLU7Om6IH1K/hXL6BYfWeHaB93SB0xS0k4vc/hP
Fq+o6zdPyQpEEsrdUtEW4qaq5UKLse7DZ01JK0Nd930uEXZjIJybAOZM7YloXrVuIFiFjDo9gCMw
QUX5elRie3+bOR8W+CC3AYQcJcHyi0smYj6xIoLEXWD044pXVNM4qE23KOerNx0MbOk/8JzRawIg
dn41jEjacGAxWYLkZYbLVc6a7McEV2FAImcGpG0apwZZy8RR8nzQ92Q8EY//XNMYiR2u7+hl9IVS
zwu2ii8ojEH8bfXPS4XDdKuXNat1ZWwr7k1lK+e/WPd1nj47gQ7EbSV9/Z2Rq4XL+k6BIbEsrlo7
Ki4b23zk/OvFX7lauK/VM3IQhAsRhl6469FGlOGNIfgypNoW5wFMbSz5DZol8Yzvk6SYPLoCGGYB
CeVrRHV4ug1T+u51rcOdsoXfBtGCLL+I1ymmRD6q42L7o2VrKj0+0v3pVmgwcCnL2dvQgc7YsCND
K2RZmyyqBiG+qAEYc99YRXTgufuf718tWipN7KqMH4n1MYSWFzthVRMXxEVCvTjW9xdpQISz/YAD
3O0E0Zy3UzZbZMtIlmejsGHjE0/uqT9c5RZMyM+BGiGolJqBjmnjMOUXidHXde8WP7IBhDovwwrm
AycgsAyFJG3utlEmgDWaF/q0XZ0RQeXuvgFWiClU5+wfgDhJmzrbwPCbv8YLMppXfnbFPoiy2UkC
2rTw59ZMYT41boWuRFcGcYg19+IIXLZR1Deh9ARI9dSkpaUqJmrbEYwXvC8LmY9+w9k+vBSw14W9
EEbSdbD00pnMQrTNbBb1/DMBvwXZCt8uwxiYqSg8I5AhvVTpMPluRS34mkaMhT8wnZwgFe90SJZ1
LVbGYdMUF6lLf3tszRj50AcqUImG2uld/X/wIMQpKLVohn6j5Z0825+lUOoUaKhR4rVFuiy9FvTJ
NkjoFej9IB4WdgwO6N6atfkOcEipKdrI05wBe+wQrl4MZjSMurf6Vf1kUwn8/ti/qZtFHdPM63Fm
Wku7tKZDm4uUOaDSxZ+w/YsYbMTitBG5dmqgzRFEOBoZs05IeHcpKeqDYVPRzYiedbxFcPtuaKuA
Ckl0AjCIpEDwbq8D9jW4Y0vDO75VBut+TBiiQa9XdHWEZHdypOVT4BEK9hBayq+AJCphHZJMKtns
sZUh8pB/DAY8B9IpArbB+lzqJCs/nN+MDdexUFjM5fxDY7aPDh7/GEbgEv/kvL0kgTUlV6+eWbKs
oQQwhuXiGeD3SMYzgyEXqb7TAiXlPFqSB5Y+zGK1jCkuss50RcBi74lJxrJuq45ThhRkKK95NrPa
9gqMoXQT+iwHV2gJ9ebZetkZmBKFepcsU9Tq/S12bR8qc7NHCCTijmBEt6rOjQOQDx76bQDRXKc+
e4NkePEuiJw1AQnyr/Y9lRQYl5PXRTj5WvVVEUoL0x9gVAx5dDcmxMfq8ayaURmAH7rYpZo9ZvWv
972ZqVqSKxy4j2hv66+X07BoVfiRvOeNpVlNOecDFYCFKrF97iJY6Ydi5kfZZXnVbeUVlfIPL82M
WVADGT+0oCLk1rQrgey0owe2omeFhQ/YWeMe0GPc2vYTemVXB6wjXJLrBHPMOMKS4T5/CDenff2E
i+5S13RyAEpgDd6JjyPaZd9ez1iWwiNcuAEWuWx9qLxC89E/skvuWUll0M5ccJ2SzqWtaDitjf1T
l16er66bZ58+Tt6zU5XjU5BIjAzKstGr6q1c/RaETlr1s+DvMlLoENR+4/dvghJbKnxWYhclswcd
uC2X/1boYf+2RFL2fSYe1w4WWPHVJ197aUK2GpO9Wj9qXelNLZ6Ia96G1Di/0jNtPJFhtTx8RV0C
Hmf7bGMZpT55aVXlez2xfvhQp27JzJngoosInRZGqBVecE2kE6ox7/RhMPiIw8YGAqgXxMJh/6HP
UnVHnqbEJES2PHl4VqcgEtcc9UeeGR5J2ROHXxdTQNtLGMrtHAhI8fXNYnmXKw5ukSRdAYvBZwZC
p/yNgTggoIPDIeJuddA3bIepeGn+pHPZ1yoKA+3NPPkGgQ9LU4XjmRQ4pTS6aAJal/FBG0BQYJet
cwsrQmtm0tjY26nCNr3Tig8MIQ0PBVoMJBJ5TAyCDcaQqK8xcC5tPXX9BBZvFfD5UGITJKMxUwfq
yXfvwm64Uu+r1fmfzJPuyTPCnOrgaGbbXI+GZ3/zB7KbaMYQLjHP0f2a9Mxk12GK6dRFjQZjddL5
zYHzpYfUAZ382IOU9mI668iGG8tWMPmnplzllZvI58d7ilUo1iU8a467/9hcQSMSEIqSc6DNY+Qo
o2uiG1qZuJlltpJYnajQfZe/ZOIybwtjVvtgoHOpHJK74W8oxZKVDJctl7G7DJ1qPTA1QireVw4M
cRoKDGDwJLnH8id29VTcQJYfFKqhL2fdawdhJycVIOcbz5rayvDv7J23oXrRZGiPGcWysGlrU1aE
x412iqB7v5yNllf/LPura/V4KHeTx+AYGsfCnNq7ohPTlpJAj+rB8VL5vzvbRmAa5SEX8lDjaoX6
hobo4Oe9k0pXwbU3zF4EKfs9ihr4GhPXzvjUYC8pcsu9X6jghXFWzb+DHKY+6nnrK0pB0rH10Khb
ps6Rl6+t+QftWD5KfZqf7lmBLAHeviZ6g6wbDdCsOqhT28ghjls7KzVGWea3pNzi1RWvJtCv70Ts
Q0dZNv2uo79iF5+QAZzx2ptt0rI/HVr6kcwjcDFvgZWa5eI3tJ3Zc3sSFmQuPndkO6HYh2G3INjp
qNjQgy602xQR0fRB/1fku4+V9K5+VBUPqNZOW8zTk0kEYxMqoU6fQSmkdx8Wms9Sdy2G9EOzfFkU
h+kxIw/JqK7xcEwiqZEFuh/bVU4fd31xELgVZKDBGY9mpV2j4KeInRRd9dkKpNggb6hAWsNSkA6d
akQC8cBAHQhLCXYYJSphfiMm4fPL6YV1BgqihQdZK6dI01vOvdOCXZoZn/77qUqPzebc17oa94Nw
t0Z43n0/FjoYBqfDrUnTVZbTBZxxq4htV4JGtwNsxu+XcbXdKKf2dRtVUbnDUatgbgPpieSNhT7K
cz4vMD3VjFFI1ClT+mHQvdJ9cBF1UPLCPN2AOxK9nLJn7k9dHSBxFVwEhKC7vOj/CIctZLLuG11P
p761CoRQnuSWmlFsTGfsqoIZQaI3y3Nam82dkEWvS+5NsTZadQv8PCtuE/G/+N4dDk7ZrCGggRss
UttN71bADQH96XCtV+1N8FCNqiprFMAYzogJ1NOr71YxFzwpn3l5mVpD084Gsa+miUsfEkK0erS+
gNWpp+biYyRAteAk3KunDGNMpjnBDZHFBlI0eMt50y7WP+1FLdzJJ0gj5GYmP+MPi9xWXx98Xbrg
28IUqCK9M/fOHZ1kX7lJx+v4dANvH1JC3ob48tOjwemK5l/RioxznsvyUvHOd1cd4b+S4QuCDPtS
Yvif7pQ1Or/ZCn8Zgn/IVXfHGYV4/KJjiI1pDejZiEPJwx7efPA+W8UG8GWrQRHN/vdg2K9cd39M
rPYtf69hVIeo9s0OjBlI4n0//C1rSxipngYFaGvfubthv9wgzlxCLAAitkshDRYPG/J9sIqnMbuZ
PcK7WRHSmdaQ9Nnl8hLzkXdnBCpQUaa+Vd83Dc9/58kXsG+pe35j22c576+6QrN9g+qSTGpfhZah
RGHi9gS4zBlbqL5b0K+4SojDCqG5lER4zZgqESnucmCkHfqff4KeDCFIVEGQCPgFSFvipzw2OKmZ
dfKMrJ3YcC0gLpuK5FLkwjSITAz/AQ+GhZX3sykbMdH6CC7dKS/gzjnxsHaRuaFynTFMI2dsJrZj
M3MIj3f9+ASJbeLi3GYz7euYW9pz6nj3vD64X3NQpi88jrwZV3uWcmVEWQm/gRtEPKxEGRFYdteG
KycPkk6NGJQmIXoxu9LwnYFywp5HkgiqbbCGL0Toche6HBItUkgLRhWOAK+/HmPALif2cAB+372N
sk7OT8oNLKr9eJEsYgJEEFTdaXmWbvYETQM54kpK5uxNy5HiDd/+XCNPhE+NhJjA3F9kTDQU15g8
JK7upoAZCWLsdyw4/IwbvnVsCENSipq64zYXyypz/ySggaZl5r29uvR/hPD+BTnuWuaQWIcm0U9a
m/nwk2QZ1IFk863lv04acnykcKAIy/+W7QJwH5yE9duKbXoH5+bdDmmhjSGBXra1Fd7+f5UL3qAJ
0hzA3Iv6+N66E5jzYdw01hujucAgMvYI5PFoXt3TMMcfMC2Z5Z81sJHKb5FtcgCAk/ko4g32nMO4
xrto9ljOuo4btprmtI0oom9QoS8af+s0DNRu3Rx0tWHHzpa1DbrrN1afVsJEGTApTRscyFan22lo
bffr9wZNKmNw9PqbG8elFiqC2Bgq9KAQErSqyOWgO6OTRqD12nMuaDV7WXlLSIuqkhGlKFHluagz
gSyGqO+KNbATRvSrTGts+3zOljyX4mR3F3RoUBVst/G2YqDpRzcY6MdoVkMn+hBLc2EuiO1fHSBj
b5pB6qPSNYtdE/V+DyCx7WiYQzwZ6e28+a1dcWbH0gZgXrCqnkpWSSbsc/0Tpics0yNEjszxrF4i
bQvtJa7k1J0mubG1u3mNipRXZdEl3unOGunAzwYRPzsFnUdE8qpdH1cr3QRwEWkgnydolfCJm5Pa
ByHBz01NCQJAp2KH/EQQOZ2FYz2ifChoILRA8ksBJcGnaEDWgASFEh9AbxglW5fUbbeT0qZu9CzW
K7VnG9CFV71F4chlyz6S8KYW+0RLcwUJ0ACQ3z3qqvf2r8Me0Yhyst0tCptH1Y2Lb1B2wu/JJOLH
Trx1ptrSh6JoLiYTP9zng0mLO1pxRskFW6LemBU+BYdJwUZqr5I81DawyGCwb/rg+svpYFzxe6eX
W9AtMfpsCMSY4iFWiJy+DqAopFxZNw+31ayxncATOCZf2bfcouIHzWlz8WTjktrPZxaG74NZ+mJG
J/KM2BmaxnvGV3Lbwg6ayKCN7cWkeEO5oU6Rn1AuB6aNgLUo2J2fYU6Ag7sNbVqMhdeuuF36Xovo
IOERtER4wBr5IzmRIj9tAjJqjcxeR9X+ZM1GsLZYylYbq25cpRMhRslh33uKkfk1IsaYmv7lOqKp
DJeURWqkjfdPa4+t1JFenT/Te2bR3F7fNy8aRm4buZqhVYOQM+7OglSgEvGt0ef0eSRLHrKOEBeJ
RAJNWn/rXI8gkkWQWEDQEO8TCojIeIppl3mj9F3ShS95JgLvQsfMbZzet5p7rZfxk8ddXtdricy6
PdmW6jSXOkT8YGIRR8lKUeOvt/FuOY4WzI6Glh8hm+ZJfqgNtTOqEytyn0sUA8QenNHDXhKC4aFn
3g+e8GYLf42J2mh9NiJw1SuatptOKh1/rkzgBBMR3FHHE1mnUCYrnCaCe2l5vAzHbHcwLoVYbzzd
JnndjBxyfzy+VF/PGP0GgjSDAQD83SCjERL7o6oIH7iuRLtEi0tbN/ruPvWQmSaCdHbmmX/A9cR+
iunHFtAYotS+tIg8XZtlV5h3YTv7uIQU4CwpUWOyEXS0eUgK1+otN9XjE/2AfiZ06SJnDaY+McMd
B45JyTYRzvG5lK/zB/1pGHqYnASiYfwZCfMT3bovrTlLbxQfmIL0DkcL+xm3KKBtU/LHErsBKrOs
d8eNEJPmQu3A0Gi5bk7cJut/Hjrc7z+g/D1jY/28ustfTvDlcPfGCKMI2LTC6iphSjmKIhWJpm1b
URrTTZpryTGPNaA6LymMXbHbnGnJAOTK0d/9PkJaJywNm/phQLF2/Ep9oLxNjpvKV2fP4uhLNl5R
uk5thd8D/LA5vWyk7EMmhayPLOLAqyigecdoIN17J+wDXic9P/RQA+tVNqgf545d6QcuHEGxswMt
X5Nk+6v/5TyIGJcJEOWP5rw0LEl8KM3LHevjCfvO2CR4OHkWPBb2ULd4t8raxRTFUn6KXPCuO931
87P3rOAoINdvXyd/T8v0a2TdQpkuyyc2b2DJRfo6ckw/WXBn3s+sddyGrtH56RmJAJH9uJNyTN6r
Zm+eeOLB3KoP2X8HCIK22JjMdwovc3dgrNQFJ06nlUNzSQpA32PtOoBMYjuQMLvB+fjAIs9Zz2NK
OjBQI0kdvIYUFfdY0olZlILhAGuVnzwAE4ZUjCud6zsyePodCqD/L4gdaBmr56elFRRnPT8ay4V5
pkZNXuKu2oFd3e0AXgAF5wC8UCD4CmvFzBeZ0W02vsaxLygUgdQI/cXHIOzh199eBSxoNHueOnGT
Q1+nGjrmW84XVTj8yDYvwuNr0qKzU4nhHJ+SDGwNa+AIaIoZaLYeCZSd7N1lj9EVs7Xjrp15tgWd
iopdA+aJOJb39XBovp5MdBapxui50z7XEP13BmLu76ucwOiu6iqJ5xjiKbruc1KFd2Whj9NbuoM4
sLA43zQamb3ze4vPuTKKptgLrecehLpdyxWZaxNBG+r2hmaguCrY1vt3TYss68nvB0qEgIhY2Tvk
WTXQqc5BONCdJdgkz3OJlOAJZVNc5TF098EEe452NNhJrKl6gOmuFOwM7tyebDr00bZXhyISmBbD
Wk8JanGYUVVheBma2Q7oLBV//N4nPe+O2y+87NuSe6xIWZkkTNJsDzNOkU0PAKkAKv2EWr3A3GtY
7+3scfO2Ck8IzqsQDLgd5OCv+8o6weEAc3DfMUE4wsNitY1a0d3R6k+/0L9ilaGqe6go7w86euHe
bxyU41GSU7FBF8LMCvhfqbk1tlnexDaWVgQIyzXUa97k3qoFhpp8FzFDCNKn4lyHnCj2l99vGoBB
SfscUEPqQ2hfdlPb2QefOAe3cJynr2wxTvb12ncALoyQ7qNHiadq2Q5J8NelcZrqjM6EBUakhhjx
+9FakFG2cVYa37sqUns5ECgnnZf8bPdkg2YcvQcf0UkWTcD++enHNGKqLOrgmSxlGvIBbsdamJOu
VeWH+Ik1JtvL81p63C00hwPIWySbEF9/V/4l8umPgYmzqjBmZu5b2yfRJWYnfkJ4+cdTv/6QcM2r
SxSXyeHIgLAfygOVUDO/IU7yu0yp91KFM81Bou7UNZSUp4pLsEqV4QaFbkYh3SMOisgdMAf3UQ56
a8CY5kwRWyFYbQcdJE7RF8gzHd2n7FDRNkr1hQru95zudW+F3/bMavyItZIiGScF7zibxIkOIJ7z
+Qqn41h6Pn8nw1blFL+zy4wRGQCZaxhVKxV/rnE25MWpcoShLQZqSC278fWJt/HXiCzdkA/nVTXO
7EQcj5OQeYS61KB4yDLN3h1hpMfesZuoc8I8wzjrH+OUjV9LuW6z50RVSpcbn2/stHzlpC80BO2i
3isBJIGmthFOYmFClcyQcotH55iUNrELTZZQe4GBG8DagBK6e1+MIi+KHuNlHAf4w2dA5vZhVMZI
IZFiuT3X3R7Sh2YbMOYN4M/nzlS9eyMQMI+0BC+W2X+CrD/OBRSYsTfTiVtJzgHZ3BEJ12rBFdwm
i6h90x4iRkoHfzTTWuzrG0n43ZW3buROkYZHGKOFQMncq3bD69Wi9r09R3qqFLd3xuf0yKEoNIu0
rlTDGH1euETRvDe3cG9pi7LgzJ0pbFPQ4QuRR7aRyiqTjY4vlxSgiCpfeGEcql96TXZAqH1f2WQD
px1HTa6CM+MvGFSSV+gmCMgOdWE7+Tn/qXUU6MTROeEaQcA9arrW4N28oO7+vxn/J0iCwD0pcQ0/
3RwqaLWI6OGr8rw60O74myWmBXzWVzRDYJMq7ZIWysizo28t18Z9U+7ZkcklGoQpziD4zKyqRJTa
VwIU+fE8bOXUbAhn7G128GFzpYPh3mFgv4UHW5jSav8owoP5/ykGpb+YCauy7n4FflnpblB3eEBa
LDWTMX66otVoNnYA4fhhe7ut4e+kz+ZlYDDG9r8nPJR7fymuXHk0pdUwY9G+TnAa0Y6z/BOzClRz
NsIJksdzzJYATiusYIvMWCvKr71IxMGda4zXBOnRniCFFP+UpHUXrZ8yT6AuPXXgY61EJvpJ+FZI
mpjsEFBnrA+hYfAEuDfceVvm2mGu7JQUKEuWexGxiePQ5x95xRx/vOoYbpGaAPg9tDCveDFyrHkY
BJKXiag6AdpMLAD3LWOzlANbauijuDISiTtxyBmOvuenrb5NMOertrgN+s2hDc/0gYmWC/JYUfbx
3Z/fvWcurW4GEC8R6zizDZ5c2AP+zwnstNFUhIueYdeaTlzhokmGphWCavilDqV1gOsZEfFfxPKj
0e6gjGb9VTBrLKwMtQK4pIS59PUCnaG6g6Dcc/CSOGCpow9q5Hgmj0UyoQKhBSLmmFdn7sOvMZ+N
hlfW34/cQkML77QgzjNC0VgFubSkkNVEsZBEkWVbxXamgHG39JExzYntAdwvy9wS8zoO3HO4ep41
IVuOIEWYMmOi8wo3SE3ePtbHBykwulT5avwKd97slDCcbQf7BpSYjF3hUXUtKEGxVfLKbunh6mF8
Zq1m+Z2F7iM4fGHUqFddAcMBVRvo5F+7JYkjUzUjs3LO3Baj4b/EAz0eF+w67ubAFuI01hZwXAim
frFgwAiJwda34RnTLnhcpEj7lf31XsMUsnqzvmoorrnjRYVA//zm621CTA+++Enjudzlknu6uec7
u1sGRNe5NrRf/j3pygTfT4pOQ0AEhnr1sB1Rz3R8VC29qItHfk7ElP06ZF38wpAKNPnK38QoTGee
kBhHPvImpHqYoyxbwBIVD0WA2r+APhu1hvYlxhY8lPWhHR5dEZTk1JVKph/8Owj6LsYpup+7PLH8
iOvV2EpIlNVVT+2vUTbT9GOXa6i4sbNhRYjbeu7LHLAMw9lNWnGSmBuifuPSQFViBiw+clg7RhZJ
rNJL+TB5oCkAnZPYtwGVtXz5OPhhBOCEZCX39tGWBJY27A+iCjhnXH96ONpuqruieNnTIQPlFmz3
+4odNRsk7DPCx+AyYBA72RHDKXTaurYM6geCl4h36UQniThyGgKGg09cXjaoQqo80pVo5T2lGrk0
wXkBM/8vhu94++2OAXtPenmp/mZYQscQ0H5YtbLoiCZqEu3PR+9yUUDlPNqfmY1U7crhIuJqPScR
5XATcFUaYiiif4xt9Iu3AK7HzQWtVZT3sTGDn5L/I+UCTm1hGHEFCTxFdSon+ocvAjwwTx5n/uV4
yDEONuPr0KyQwLWe75jCyw7O18I9Iseh2W7BM9pdEeZaLJbxpKjB18RiqJk0rZrA2iTcZSysxIs3
jhqm1cZ57Sy/y2CckBmF9U+yQq4W2QfsTMZzKKHxmFqjQ5b2aNJdsc44D0jGHQo6iRAYZwUOebEm
tB8+gqC1dh/uoVvx0iX5OCpTdVS9VQuDkXqFIEeINgh2uWe9VdDxXbgMBaWPqzerBbDojuF+HPIR
82AsSpwYMbszbIUank5YGVlbZtivVZrvjJKKoZMHuBVMHxV7026FHd73UCgcWv6u30KOc2tppO9K
w9dnoo5pcnim2HCo5keBt05Cn6VS+QXwDl1X3xEWr7SRAEPnxWrym+Gfv4AV2cYdH2wSmQ4bJ6V/
sI0K0FKGf7FQPe4vdl3fgvTTxzrGExKej9PB03gMLCZlFzzPNfY4zTQMtBNI7UPO5nFvcPE2owGi
YHjM5llzKWO7vsMUsv3PIHDJfWhgTCNPdB3yuHPnLn6gaWrn5PsYuQeKnD7pCwMg+UenklhIh2+c
aVU726eacJt0FDpJPODaomQ6qWrSGpZJvw6x5ub6yKIpqo3n7vf8OPqaGq42qvdn6RQ4e0d6vv71
303UvawzAemNsoGmqFznMGICx6hW4q85FF+1oO5CYr4geKIg344fW8v9oBOcjMKLUvE4pI7mxaup
gtgs49TnHHR1/G205HVFGfYtu05IJEJGlVuA7byySEyhuca52qwUMs0bvLSe82iX2O9NvW0eI78J
6bocZKhCWm7WEMwxDBs4e8boCB2HquC/ORKepgUhwT1yem03sTGeWKXXR+dMt9QOmlt7jXghyvY6
36bbGAqj1ek+NmBtOON8gGHirEjsmqGryCO6hQHVOzugM5E34XxV+ix0Mg/CyLFGYD0XyukUAL1Z
Ofgal5EyZajEn2w3cgqYwdnbjKopPSFdn/eIRIM3pnhDeZneLDTsl23oMTAI+Zqqbt1tRsDZICE6
ldnOcigm1J18hP8jbqH6LUgWZX4e17bPgT49iRMuneS4UGlQPWTZtw+j5mO0+w9yJUJOdhnUMdIA
dX77UAwJg6xxoYxEPlw8Wsd500zAo3u5wKHzv01FA0gvriMbOak9gHq0/upmG8RMgU6zAbZF7xv2
pxAdPUp0uhljTkUHKi6CKV7ChftRft6Z3dSVm/uqJ2YHRC3ybO7iyvpO5OkgcNRnZaknjP0g90+0
YU2pb+xDeuDdtNCF7Vmeo4gtoR6rbCF19KAWCotpnSZHjakIN3gE0hO3jdDyfUZ/UlrLCezlR+mM
4qE1o39FLwol59JpH6vGlLI4zK6Bb/q7/TimkteKqkbrzTknMdQaGJGyYGrXdBLUQZE8hkB7otjQ
7mdIFD36f3G3946jOLxhnE/+AZLiyA2GwZcRzHI4gc1s99Wo1iwAA3cJMuArI/ijlwGnLJUhBnOC
OQlxfPs/egy2rK4ABuWzUsQS86LOyQn57dgGOVGwgWf6StwX9kQWA8m2/582X83dYmysi2Oxbu/g
FkTymX2/0V/x3bI+aiAaVoP9n+lyjq6El3crMZpU4y1D83HY3PA8qlNFn3YQt01JZJCiZPVnJ5sm
6Qro9u43JP2zs4a54Ppzeh4zJrmgPnUbj8hStGxe6et5KxrA+CcBoqHmEXzrqCg7KeH4dvuW2fkS
5chGxzADoR0QPqRR9lNitttBEqKz5g16h/B7iOp8bAngBWUCpwRva6Nk0FPVvOV2AyGfKfxUDoUl
/wl6SqtrwEx6AGlSg2mMZgTV12d6eyL2Mgy7/8hSv+HdUT4zd7r8l7U10q1OSz9s73D75mID5fUK
+faOUVIWZb2Nxb7XoYESZwd7wdvTmcBW6pGb2d/P1BEsg6JGsvMHXToQKs8nlRwWfIQQNsabFYLW
3sUslOqnl+mqrXQARWWAJbtef8OgXFEQGviaEbJF/qA0b80RIthwp0D2vf4Zeb/mG4SSfZVsMO2w
rSe4jlI5bbEA/tqCf8hAjzTCEBWnpYfKZsdED9gIAQhCiTUKLf6J5svvKW4vgZ62bfoVSAnKFHp4
kNVoq9LTSOMXx8R10VXrW0FsubbrgbQigze5iMzWh5H2371nNsa2fyEfVqOwN2KiPoHgPyX5d6jm
eXrH06i8kfHKwuSVi5hkbphgc/ALSLmc8sZ6YxTUyDrjiuTMknjFfaaAKRD2uskkXMyO91DFS+1a
BJCJfEtlRnPtv0qqZ9MNINulsB0NK4saGEnoyPJmEu2mfFiJdFWje7gOOOAPDXTzSZ7kqUCEHavO
24LmRe4H0TZ/cnIMnzQqjB2YULNYqD0zld1Uhs3DLv0fZQBUaPPXlVooFaFAUwulV2PYyztkApzw
1vu+YvUJmAKG727jGgFpKMDnV6h2c0cwHdA6p0A+IcPJUobQu1V5yDw7I9rMWXllEHyQqZx4QFY5
6LC4S8G6dL25f0S45IyztuUQe8zbIWKPII3Tz2vd/4Vb41ub3iKph924kwHIzCDd12D+gXVCMaJN
X0Zr7hRNESeyZGZCK5pVVGmjbZNezhfNdJ/R1P5AU6UKP+JIXImAeP/Br4ZLPN9dtlJuTg6dbm6o
/j9kOi1LGtc2YxU+3mbP0glllOe2c4qmwXepMDq5Z+WL/Mv7gVf16KehHoFYc3ubp5dOet3ptfdp
GRr6BaXRV9fX5FZo/VaU798Bj+NElvpNg1GzDbeIHnIt0pqlIfOQzWctNuKEyPVhH07VV3jNQfwS
mutbq33ko4qgmKETdcrmxq96BVvMZnoFU3BcMGvjcrb6xMB1WWqdY0EAXBgAl4j5ycnZJZNMBUMA
RSBpo0jQWJHlA0npUwHEe4TZrldWcY+GNkfqV4HCHWTFCtmRZhVxw9HtbsQwk5QawdH8njwrqB1/
KWM1RbL7+Zu5M2zcGf1jQIv2X0CUgUsRaCb6zwOHpo5MRuA7cW3s+E2dIP814xxhHECeJMWCsXxr
atcCjRIJtlrvKgQKuztW5dfByWqvERXocSRQrUtOEW94wic7E9lR98M6RFJ64la6VGlsmRQsq2D+
n1uD8sha/ApUGvrobNG4/Eec3b8IR9HdiPwEpHWH1qG5RqjhxrlBZOOoj5+lzuWx8n6QFwE4olBJ
LSsFLd6c1ZY7uxdx/7KyoiN6O12EMpAy4kpzYyA9QkGBnE4qbuBN744M1no1zLY/mSsnlyKOuLz3
PsG+tmdkfgU7VeiIMOLqRSQO8oazCiSx38SbUY7jnSsezx/wfe6+WcqGfBNBiXMpWeleOKj7OM8+
6Z9hfM010K+P9EIkbnHyTZH2bJYMQAVgCv+7HzxWsKU2nUR039nmnmIR/FJagmpunhR8Czb3W4Se
uZojPwWPPQJKil+gW/N7SoWp7pFMsb3mrbxgOOF9JHwGhDAu9Dcysve9IFL+tADIQIkoaV6CKDAp
JVm7q0wjF1e301uECafuLNIFHjeZdTQWsJv/fr3ISjIVzXuB952ED0ZDX6h0kMDENcDORMz2CTCJ
5oTUPMJBp/zCcYNXjKLdjV8aKZQtcloUyKDqAAoY+sO7MYU/PxSgyaonEJBrvpS9ZZIwdi4IMQUK
xjbKh5qECjkATYZmhBHyJvWqOoqwHoQLXYivEPoS8ZI70G0ZIRwlN6KTSvkARUBrtgK0ZoavTxwz
cbNzyLlXF5kjcwoGLhouyRme+H+Ui1+pQ30bIz+NatZxkhSAxv07v5yN02f3kp6KcTbdXgcxvck3
o4QIK/CIqD+/+g67NkukQME6xLedFcb+RcZYPjQh+oWHs6muifXnorhWtP67yB9PglCM/wt3O9RE
icUiadMtnM+2g0lBNISs9Y7PAQNOFCY6NLWTTKGSMzsCi+KVQqpSlsveoYsuEBctk7qA4OYYfKzd
Nz4EAm/rqyEfH2GE/pdlW4hjw1yttqfsnDspZNq12kCu5gP/3gHbXvDktfq1dBZwR/+MEMgXKIMu
j7WKW6D/96Aru99Hm3P4NBznhMT25C3Bi8V0XhknfrTw5gwcNvINKcqYAKYmOnQjIg++mNNNIpFO
Glsuk27HB1Q7Ob9UB1+ehBkXSDKkbqRSeoEhxG9pxQilJasyE5qI37T/hnUYSSJrayfcr3JKfwiQ
nBIuwo9AJnWIZEhBJ5qtrKl2+CGIzst6b+kUuXbO2IMEvwZ7DzHCsW+67kCXrEn0ljFiCZhIXY28
7uJ5GbZhItm75Z3y8ezpvyXx6xyin2Jub5BKohIIstV3a9kWf3CnXy0PeeA1vWV8rcsVwXe9rjOh
YSN+GADnK6CKqwgA6SSpYelu1TJPaYw2lsUCVr+uTOFAIW3GHOofFOvPcwrCvCNKNFLEp9ALBlIb
OA+BLT+KzaFqJh6y+wH+6qM9gfHg+UHhoAWGynLYrZoWCubAs6oOt76riS75/lD5X1zlLadAFDpD
QSD65uAEEMK6Ou09sIwKnIfdfkfzp2OgNn81VwrWOFW6F5tJaP2MSVyFGfNgLENmuT83iD/EouZy
LXNlfLTY+gx8/7wSdrcUrLL6GZBCWjNUPfhtgCdmEDN4kiRqr50VjGGlx5Hew76n/LZnmvO5vq9i
dnOM1c3+qW+nMWXaqSVY5rhynBpkzkbXXP6jpGJ1H1WYdVRIXqdcuIPsn1vOIombHlNAiSc5vxmX
02yTm/Hfph2qFmho3Vh/39OE3tbN6te5nZ8xnYjsvCqHc8rzZ1Tcq26rx9oiROtSI0Y5VSDVd4Da
jMKIE/Hhe9DdYYAWK9QMyUkNWtB4q74Bz1AjkLJrGKU83TUYQMhIDY8CBzXUima9ocJ2M07ijv7K
tjmEz+v4WlYYZCtMY7+2Q6deDWyzU3xL2Je5NzaPdKwSS71Vp9COj1DKQkLHRG/tGi7CFQDrOE12
jjQzS9VliyD8W8C0lSRh90tzqD48G8Jd5CGjXh9W8KF8Vlv/Pzxam08rWjVVomSAupLYIULxC7ra
NklzyBy+3OV85PafvSAwFVE7aLj/OBigELpveW1wwRkShhMOURVHBXnRdWQzn6wgbfNL1deb8/LT
OBDSySeXMM17HAILy/NAhc1tUmLU8XmBRQV/EQ3YtLXU6iO1DCO8YIuBYT307+u14xdcvybf/EMq
d8kMGJLwvsEG/saWwXwaqwEqzb/AF///F/e3+poWp9DiYklgpBZZQaKBHpxD6WpQJ05GDiFd5X3U
2fs+rgRIbhrVduLt0MVZHNpAWETsXLBIsJqe12FI222aozU8afkbDtmnb3NQWXkx4kgVKmG3+8SG
3bL7YeeNE9QMI7mkolXXMIIsBAfsq2GxEjTXX1bTfHKXwlpN01DHxKfsvZyDsQUx+OLHI3/ArTyd
AYlZyPLs5D0+pgPZ3uUhRqTPrVaULaZTGYOTW7Zqu2lyTKh0INbapdBRfsaMIiWuR3j8XowniMhf
63KRK0vhbRAHAri873hmYvpHjTohYr4UcVAP9PpXJlggQiInDDJKvtwIqDwZgp+G7iHffuZUO2se
EafeDSTu8Ye4qK3SPIl6mj1+Fuy8GUX254aufFEFXaHc8OTKDmxqEpo6soW3CteeXZpAg17MQBia
P6+tL2H5kaNZotx1dy9NXL2ANF0a3lhCCcXkp7ZCec4MmuwRqgk7pcIPNgO3Ch1r0kRD/mf8LeTe
NQ5C41mbq7IjMH1fh0iT1gQCcEiN4Y+bsne92IdXsTuY141SH6lh0peVDxGfIVlZf0GEyEUtLa8k
5fTW5gJCghZa5n+MdbnBqeNybnX4F2Mj7k7tF/b6AkvAQzgbpkJmD0medxJVpFH6kc/fFP1J3Ymi
dqfo1DM8vsKuMST5U5So4re9Bs4n7W/JRYnTICuP3VQi9Xli3rKXC73WDWj4CCkPFvZW2vThu/qs
1PY4PqWVFrea5T7JqrkVrnYgo2k9IZxI521u1vP/lnY4bfrQqYzY7+GdGzlQKVzj0LMrUbfo33nt
2ENwV6abp1pcu1TE9PxTn1TY/hSKGzejTNYKGaMjtCAvsKyDjYBMeN7oqDx9PA7YHCIoCMMlUzrh
NA0nZOfjHw2jJWhyg5/8xkqzKo2SDensKZelFHoPKnofwEk+hu9ievAZeuZSzVe7FRJmXk+gi/7D
S6pgG8N82cS+fCxwozoRzP0pUTaGiQ82cBW4PX/T7Wi7XZbbzWTex7p+LK9+Nq2iSQTtd2uj/kz+
ougJo/wa6ijEuLUjWzfL3bbjUvIsiuWdS/FrS9xmivEAbVF1FgvuJtz4hVbI08kFsY8WdkMu29Bi
pvU24K41pCNNg+rWqfD37Cm2qVFN5igE/dFxGrBzPTEz5fxAV3TikNfPCAogbHJx1nt4Stt15yRW
aK3MROn0iikyjUhwqNCJJVg7V3DUj08Xt4V2gF9n7ETWVZMszxCNx3kzuGxsVgn8/vgTH5MXnpnI
XJ+zU9oqmNDtS6vCUzM2PYbF/5LGeU1KdjmF+G0uuuLNCUfUhQWmHDNPkGljNxT+T5f6n1aa+cjt
lW5D+J971H3whTENgDi1j9YlIBU2okSBb+Ud8ZLrAv5uIJmDcPnPj0r6+6cHkgdJt2HKexTop+d/
vusnGvObhLG2BUpO313IqC1uRR3UmVH+HsRr/7Vr57rSTnyGTvPH/xyk72nLOSYFyQItY0pfp3Tz
qaKER3mlN5TxnkPyy6w9XBAEPWTafmQzZbxje6hjk+omh+h3Ek9baGt6T0T8HjGAYhCVJidkdQAh
r/K4h/r/gip2SDPw4NLRi0L7VDmyYpHfGEMlrFkwv0ZsTrAMEkgCMvDaA4kbA8Tsqny3vT+b3KIg
gjchRLY3fNgQT0GKcMbTbmKY2KusqrDR9TDwTT4rmIDZyXaKGhxGyWe2MThigUa6YqmCaQDWxs4X
/v+vHHZuLQoFTGXRsizoB7l5N7p2eJCEE0hgZTwqaAhwsNMqGU0jDucjJpXEH9xbZLxdWX0x5+6X
2jknfwJdQED6ki9qRjBzf8q6bJpb7Uo3OEpi/NZZhduh4cy4XxJD0vSm5LBOeIt6sSNMGaF8E/Cy
yt3vvsJi4oD5WS1jbnKZAs3795odWSjwlh8CgU68/OqGRZg8WWjUiDBQbdsWIldZym38YryPO9lc
cswRuTa1uk8hDPUfwCQZhF5je2tM0Mx2xqar3F6dYCfBXy9G95tOk7+Was9apdX9NvxAfjTuZApH
x4xO8Gxq1JDWdQWHxFOFPC0vyJn3iz0KgGz5zDcIwgXF9WzbSlU0s4Xh6NZ2BF1+bZKoGb3s7Uwm
vIhcJHVJTg/wCp3J/U3bHsf4Fv9uCO3kvX67SC0thJS9jQwqfEn3lHSKsxXHheoBmuEjesMbR3ua
a8H4zP65LAG03RY16EB7mdh7JpxVc7df1buDpF90rlCcgDXO4aIl4fh/3NLsB/wmbrovI6PMvJm8
8o6trTvjasB1/hTpLrA9jcmDmojR/wVwx4Lc3tq3ix79+TuzKekPU4jqTikwCKHLCL4lJKAz8G/5
04HXk9c8N1+LlhkFTx5GLT68s39NR/MJ5N47mWJynucN1kIgM1A8un4cmPQALfWdXr7mRxfwZ+ne
qq6LB3vseRFYC+DKr33Nb0QrgHNBCDY1gv4f3KpyQ1/yoprf0VgexGlHY7lCMtPPsWOsyd9HjYSV
Ko04uzZqEZ40kP08jcju9LcctLG1rO+j2xyJPyiLa808jYGggbeUQl3cOpENXVYlv5KJ2vOD+/7c
v6VgaUmpgOqjHMyfPr7be2oBnhD0p5u7aIm6JUic2STllZkYndQltWQeWDFNl72FWrFk1Erspbtz
dGkd0T0oOBIyVdi/yJsJ5kRBPvpbwoi0QX4WHw6FbJ0WXK/JUnixNr3mH1K0AmFBkVh1flyW7lxZ
J8wwINg8s9BUdh4e2CftCOJrEfLjkIwC9x5K0ILpxpd+ugyxAQGoLOh0kJis4GGiNa1UR3DBU4rw
IRMQgisJ5dUAHQWzSmtOyvYz7DqCvfg1sraSJEyg0Ptkhdaz1x6Imc9g0LMWXcVF4XWrCE49uFQP
o/MxBPFXpEqJtAo05m72tTY93BrxyK27Z5epy2uWEfDVB8Axgjhw/DErcxrewYB06ehYx7A+DlKu
J3EpOC1EqdNeQEExeWasZKY6Kv49NS2Pk/NdFNj/8MvUuobQ32SlZK4pP+zSgcp0XIfiv3ZpK6+U
V58ZGRPfHBGP3+Q3EhzLekfExPvmocblxqxNu6runzPn5qcVJd+0moLNK1fP/CWmaJeBsNtRSlK6
/wqqLuexhb9S1m6DMNQrNg3IUrZgO6Fe+b4IkVXl5DyEa28UCJKrW53kPbVQxakgoHHuj5LdQPKD
P5i/FGQhWBCQGwO4SWlOQVZwID6MxDjHEPKd66c4gN2fY3/qAM4MUYMN74zuVKnPzMLX4g7L+8Y7
Hk1ToCHivcWXyhonxa0uA3u/9LOmkHxigh4e4P20aKlo8rszbzca3kYkw/XbWw34OdBPm2oG6hEx
2DIWZUdWoFZzoNHAPOOQSnr5oyXFGUPzLj8K4Yno08PkD//dczHTT8ugMXhOp2YH6SXQth2uT26C
eJSxtvkULxuFEHlJuAoWLvEkLsa0sWW99Z+tZjjLz3/2SPf/rxfGfJunG5RQhNxJGDNL+Z5cwYE/
bNMmOqY6Ip0AJOJrl/sdN2VPmF0SorvBMYiQC+T6ggxGbZK+LHgVl/kiOxZI9f7NovYmUJPWljCR
iekO3bz0DPhqse4OqRsKeb7z5voKzeQ06p39XIL/tvuNRTRcNu8nvmmOcy5IcJqNPVdZM0hSTmra
yC+zabB1ZVxNVrbGDkOHgI0aQcnDCxbMnRry1PbWB5JHjKborBWHYB+jVHSAJWkg/i8cLHGPZNxx
fVBKpyzOD56O9dkVFSeooXdghGwJTuffSUJbhfXqQw0Eqcy6AgMUCeYzbZyyve2ZKlPa8/XNu/3k
lP3rVm4h+HRWIXKXRqPCM3uhGM0Uxd07/Cjvmgyl4QW9A/p6jWc9EDNKKWAhH845U1eH/3NrRQPh
FW3ICLpiUZ8Nej3T+bVmbpHech6wR0/EPLL81Q5/eKpk3RJxX55yYjFZK+/g/5/KbLm2zyEr5DT/
L99LF5tygBIc9ZR1je+v8OaeRc6rZ3mYFG9+IegT3SeN1n8BPX7nLQZCiye1sTeJ92AfzCfLkmul
4WSfGvVkdA2VxX1iAJmNIvxxzjpkcwYc/J7TZ1tD8RD5HqJPsMEBhcCvNu1hTMA7/P2bsVaubLGT
NCdVGFlwTR/1ex7rAjcXYgDrnSNXK1aAUSTn/a3NKzcsyciinetagxbCE7Pbbbzg8OJYVp4Je0hD
KJhAPv0rBDrW7h9p/9KFYljhFkRep6rZTa0wSC8Vkm5xlBZf9csSoo3gJfBSNwKs/i5fnxgcsyLj
2jLLaGq9I6BPNCU3sJnJfEnSYO2K8hEehTyrdyvRSEOejHjbjsJvsrEP66gArKzKKAT4VpW2volD
CJeswGsa5qJb+vVbOJdz+fY6XlrzuaxVDv6jI27jzhkcXBEuipug3GGwAs6j/etQ28wujzHg3pnj
EmqCewEz61J3otEUC2EavxGm0nvuFidbfegE5Wi9Miz4eMDk7kENL1izyeRCS/ftUkttfA7eHs0t
tUxwvoYrLe8Fe5JaQsJjA9gzXo4ko2wy6h1BPbvLEBhOq5KDw/NJLiPRXBJfej7KlDMOsUZ2KPcY
RqDBCPqkeEoFQMFiwmbyhRv2YZvbu/V4nNmRxvnQasyz+3HQwiDCnAr4Kgi3OyHfIdRDI8NuxXu3
3vxfoMWmUjla/x36veGMM8TuE49MMs3P4R05Hu8Lr7l3UvWjbJs8Mzz6wZxSE9T5N66DSB67IS+x
YmUXLirruDwFt/oj6XAKMAwRzF2+ryB41k4Sl4QfeGFFpib4mqUVecf7rs9EAsJxQUxrq3vc3JSV
ntKdmRRojdeYXN+ppLMGsGkejrEhPETMhcvSTLaWQhSy2nY8kERded9syjzjrpeZG/xIkGzfMaUT
eN88tZNa2AEkbhn9fxVeInf4mPvM9i59T0ks+DcTMVSWDsBGJxzm7LDrV0IX60SaLjRTSJL5rmWA
y2oqQAriHZlKQhSnT73YyG74U5jMl5KRyaJbWDo6Mv5M7CX2+15ePm2TXFcJ0OxKwnhl6/bxkDck
h1P6eftDARnWBnefUavOoDar39AQyI010yLfX1bpaCAly5QEg6N2iQTJ1FdIzagghPJfAUGtTHr4
kroH2ywDatAQaVx33P8dyEw28Id4vZyjCIK/HLJNeCQUTJCAITBgfuUBfkIEKHwkKPmKkgNaSYtS
O4tZrQV710hdmw15nGphbg4NteA1xIKiLwXQWwETcIprxfSK16LX7Pg8iYulbVVdmX9X/vgzSNci
N9WxxD4TEonC2R30zaLNSajNQX2wftENamSlbyxaplZ29uiDoJLR+jguen2bTvgoDYpnoV29AH9y
gbCMjFh0nUSNjqki2Xf9hSR1ZXlVDasKn3ujURkVo00t8FVK/ZoIAE4NXZL/ullt0sp2OLKuBodn
1th1xNNsufF8y63FrXlsDoDfi9GG6465TfbLQYgigQfzNRr35+HLIyJJqBbgSbHRvXsxhBsSmekp
bRNmVtitIUacTgbKR8v+aOvW8nXp630Mp1tzsW77CPYahv3N/3fe83qaKZmXiQu0h7TnI2QhG5zJ
IvQ2bAA3KgrOP4VdJ7mYZ/FsoMNskzIoXI3pJk0ysNk0112xJiqPacFKHkRFjhL3Uef/Yl7AXY9t
d/9DatLMazXyY9UxSZZ/NwBKt2O7n0jOn2ZdbfjnQCcl3mbXx6j/WY9vo+tC+oiYLpohu23p0G3R
zMUEFArkGoksRk0Vyz7BvlASXEVfP/ttEMlCTilQQY5wnFVtGt5BKoHVm9RxPQq36V788iMZZcfR
I8wj4nVsegQL8wF1POlJR1ccXqzxYyLEfaNS/PsH2pVTYBgVvEu7QCyoZbNeMhAVwAhP0YINJQdb
jefbb7K0VPHfQ5EkgsjPFVYc9BZVh68in8INb6S+E0C7npSdwsjFczn7VRLV/hptGbMveoZTkH7U
ORFlXrlLtr+OHXd3MxnzxSxnEhgOR3X4O1QUgmnuFWtIM9EpFm6flWI6MRctx5NHhPQ9Y1HZ/Rba
1n2xucK0OhLWJMV0Y45h40lTCWzz3J1kMFFrPy7eypWZrc87ToNxD5Hmu/NQ2wnXEAKxyTg8oYJp
Nh/UDvHt5TmOoNHLXaTlbDLxAnnicwR5DUGoqXfxebAf/NwzR5tksAclIYjm//WyIZOveQuUfCci
N+4H6zHtGMOttbfYscCBMFQpjFC+I4TSbX68n5vAbdZuFf1yv5uNTwDPkINbrbnGBelaFm0DIL6F
wPZvEGbfenyc0j0UJFXk0tZO9+H9coXJhMbknN1eWbxrEiGMIQjOq5LjqEgmAcgJEbqA/C6W7tbf
lsvK4Px7CZ9FCko2crSwnK7HJd/pBIZVehT3IELQyak5Q7ySWijwl7ZE3Y7QNC5nt9AHFyU5HcwS
1Bbv3lSTeJooAJDamxi9Gl+UP726h1OFkmeTKJ1hPJ1Lt+cVvt72rbqmaEBxKJgpJZoFmzjuLOKY
OSl7B9e4uGgCdaNZdsFj3tp5iuaBJE3sgJGa8FYL/IC1MjDaw1XqPWbDywvumm6Q0Z+OJjJsqP+8
UTxN+p74kclYx4zzPmrOGsRP2r9vlSC9wpBrEiuKIQyhIXHDpUxwZLuc3p2b0+Ng/Hn9GLroa4AB
O69Kh6WCEZkuaiGhZ4tjI8kF6ibDreJ4xK8la0anWPcWZKAvfgWGY5wu4Zh0K26OCEIctV0nCSGt
tGcgIaBhBLy3b2v1ExI/K35TO0ZTuwmarp7QZriPxls6PgdPRrwYwgm/7xVDP2a4paODzIlzhR6A
5PLuPrn1nR80K/XIGmH30AowrefVSHZH51e0Lvaos/70EowY6+dBSV3heTOqGgUhE7NcNlo/vtAU
y3ivZgjEQZEC6P1ZWfCeWuOP3ZYgy/ZZIa9YpO4rIRdAYIU+fNjPHsG0rWtihsB13641TLVMaOf9
uRvYONr9S8ksPI7TtxNVdHsoSEX+lSGNcjVPVOBDl9BGfxjBloNCifRcQMT21kSJ5aV5rfqP2GJ9
YLLV3JTM39NomeumRhsqx/lZV3D2hfFJdeQmNgcNTwV5vEJWl2Ay+gEqPylF60/+r4VQZftSFuO1
s/J5y7SMPITM5PNOZvXlR9xecDhnSwLSEtvqvWoR+9vWZ40e+5Kvtu6vgZWZzlDa9bRrP8mOH9DK
4DCxqXPPJHMSsPIakWpPGPX3B7NEskOclJlqPyn3TOYvSncXK5DJz0KzeNcp3rhiqBNo9cullfRa
FjE9Ykq+JIosk1h8Q/YU6Nx5M+DXMFhg1JCeljQx16DgBjcmmU8PZ+qqgQsjfiv8NwL/XJuSvfjo
xRD6YiQxMDRM33DgN4mraVmVK2PVACZCYhEptgxBjBWo+Lq4khmE0l12Ev5106EDAfzd3BG1NU0m
Aw/LmseYJXCthdghTmkUT1J5GmibTGZcxvyJ3elhzvcQGNaxABcYCy5uP9GHhQoEAzGgGHG8ey5C
qG8b2gOwxltpfvBGs7syJtkdA22BvfF7Yi2C91eV+CDP5moQUsKq0VzNzWvuU9GMw4A0IC5OKPdY
hfNSCas/BWSOR7MheFFuCSQGoODW93LqZq9Q2IqAjxs5lUbTLqA/mV4xImbTRxjc4Of0BCtZCgza
oUtF7cB5KbmW9Qxwkln7gYKUMfymdjxSksqEKxcdG8qMXbAn2+a4ncw+ACpFY6Y0wBU5ZmBPW4ct
hxyeHphZM8+lTdwzFGJHrBkDqNkD6Sleya8MGB+wj2iQ+bCR6vzbazZMXnARl4ZXwXVo3rGfUB8N
w4XDzjGFxqwrIayElAVIBhN5fmAfM+AJ+ia4Dhch7zMRKMd4CGiPIVo/QRbpfjnXTzlxiVAchCr9
Zhyo8b9LmTzMI/MUb+4y8fZK9Lo5pxVdOH/ablZp0o12C6PN776Fxwlww3tqWv4PGHQAXXGXpmND
Oa0NGKP3CG3k2rfiAwHL0bfzDxBOef+8X1Cxt0Q5HokDtyPsJToqpMQhuh3M1MGjRxX96cKFpCGl
2GN3wQzYcayIbBrpFfMox16RE3W52A7VqCWtLm4DCDquT8gNnZDbLE1XGHf8VWrL9e5wPrhdsrdb
xWhngUKXitaxr6A8p+yvlrS76aEjBLPp1VOLWa9ev6XzEzwDPqS5DVIj24bRvd8LOigH5KRPqSWQ
ZeCgS3fJiLSfPdx1l6idr345A1XmbxO1jqUAWeGzAEV8hMGuOBg19JKz9Ba9gcV0m0yyqEdLQz62
VME3wLhsACHhwMN3VUCdiVhNkNHzFICiuSUiE/ybO3E4s8WpohvHUa5ZB5ocE1xcohdU9gJcmvVL
8k2QrPNNV/tH+m3l6DNTB0amXdS5yZnRWbqvHSPJlxZF9/XU/b/L45FH+ufhqdNfmURSGeiOa18Y
yKkQqxE0OsPhjEOM/C+ZVMssitFWMWuzYoe86dLU6ZJrOKJQtodWz29DzvUPuQroEmtS+lbUZddD
yORXyZAtuhSLT6bGHMLnvA+s6whOnDcc/Igl0SZsRfbq5yAINy01S0/MVe1bBPfUZx5PMMJLnaHi
Yl4SiTJj4iUCyacAGsPOpUZg5zDYALCRIjJ/DNLm0L/NuzaQlMy9t+A5CnDz/oE1KPdTaCjqYE+A
SIMdWTzxxj9Z8YV5kcq+snPnp/XlXP9KBXldNDNI6lgT39ad2HraJ9OJhYI4NSPS6TXKMGo/i8dG
dG6wUyDgyeg4mItiyYTRfGY1lOz+FPjakjDEDeXFb6ptAw6vlPaIy3goRwes/SgOJ+JSLRz0Fm+G
rKHDUS8Z0quLMGY9rNaA0xaXVR5E+gTwVWZSWobvdBcZKfGmxWdz36iByX8RICfhuDF9GcupLpIn
l3u5hBXvSNRjgLch2K7lm0J5yPaWB7qaFHuIF/Sw3tHdPQgXbxQr1Ffc/Sn9F+s2xzU1cgz+xDii
vwSRe3TOHC1sjYqRg26vGzaibtdA5P/uZkj3y2b7G+vRlc828xznvccr+hlV/Ye5dtjwbVo9Xnda
vAp67kAT+a+7PDScb6tqbq2bqQArt/OU7uJkLYPZEDaGrSR6KpYSKoi8aTpWrcn9HS5A7w1aQJ7F
H3VY5bVsRsZjspvmHn5+96nAsCkVQJIPd8Kg+G5L9RJ3649+e7uwwW9NeKmluUY/rMogdG1KAJ/n
VXHzclMFEoaFVp6JQpOqjSLEwLGnp3oFLWyOD5f/xoZjY2YiZ0Jcdy5r4H53g5oMgCpEFatp/EPg
JaKdxnh9ce18kmmyQCY14AaJjTwhhFke1ioGUslBLPb1FGwPFnw15jDJwqw21DFHnwAKhEyEPD/t
Q7sCXQ+CTfHzB1zSWPW1fWg13jfsoLzKmqHoNKj00nhv+KQQoJMHJSG5g/oGo/l0mGbgyFPwnM5E
cZG6QHEIJ628wMYSpGQrMb+l22aDbDYbMFOB+CHINugmuM17oSDoarpT5gNiPpBAh2BL7oNu374b
Tp4v4wafGYr+KwY61BVWDAIvsqtscTisYpzwqBvV2MACpAbeWMf3egWQCXqi6b7AYzG1baCxpIwg
1eC9Syzh3NC7bGSyz4Ufm+3FUmPtz767kqCPu92q8PRLz7vmliNBriKEhshtWl+mbRV9CoxUvlZh
DVqW53PKMe9/2H7ZhDF4yQ7iruoU7mMe4vdet0fxyfwq/DxmJhBZBhB3NcwNzOUfVcdKJoPFazvT
5ad1HCUpS5auuF7YAwj66DL/S/kMbTyqz/lo3YdRgh81XZe866jTiUCpcJszcL4cDNwF8G5EqsZz
bjNgt919Gfg7WjmDa6pkqQy8hLUzVGIe/HBS8EGPCESSzdjvkrWYmLp/kz9XbaxIDvwlxQ7dTu8H
AgGQMrxMmnq29beFT9VaMZ7ITtXHKbKy2skRrbWsKjUpKtqPwtUTYJU5/iQrNoLVm80efw5blj+0
S6IrkKvBJaM3CBx1xV0rk+7NufPQJK/5JMo1l+L1ou3YPJ6kkGhT7UONUhmTEhgNfrnNZNucNMGb
IEFJhsw3JVVGSrcwGTst2gyyhoj4g1C/MxTgywl/qhVq4LaiBb7P6FLrl4+FdAq37Do2nXiUXsHs
r0f5CO2KRcyVtwDs2OWcknleo6qowKWOYK6bcfq3SXvVM6mEZEUVYmWFyty+UhU3/k0wbpVOdhIM
YbM//XQQQMKlbzjJI8F1uvGN1PAskJMo5W576a3T1StuNIgzWsEsBkmpF8dw5bC0w6nTZPKLZf2c
/gunhsQ7YGzllGc29E4RBmobBaYTc41k2YLqqeC5s7Z4p+KvUdOUsOBuWppEdegOHDoyMrLVMzDA
P5wqF/9kg+0omJKvKmVvNQIh5vg6FZDAteD7yz8lmAhJp2BwanjBePrxNIWY6WeB69PYQidK5nrP
xgNL3XPVKoOB8xfOEIEoeY2evjOAOGzDcMOfJHObKcTkz/2dxGe2+5asKvMG6qqv/tV1lnGRUTUq
ruJXWV5rl1ek6Vl4A+IS7vuJkMrq/vDWZc/rS8PK+/znQtn3cJjK0M4PB7oaDfPBysXF4qXO4twp
a006D3ejFfDzuHlSfx1uM6pYB04/b1XtRVls7sERWI6SYUlnP2QZkYObHbBJJs8DSVvEQVZ6+kvh
4qqZ57ym979Bmm0JVEbrlGBWIWeaF2drt7yNRce/NOY0d3NAnOL8oH36phFfm7r5ht/4yrnq5u5L
/KHHC51/ddUGexZZBV3Ae3n3BY+aBQ4pGam1/BY/GM3OKMxD/+DoXLjqQaiKEbPGrzS6B5O7/kec
Q2SDyf2D5mqSCCb9OYBbOwgvw9WFu9tLgLjCXSK6JcpshRmr3SMwfV6iNW00TjTY8/biEKl8KDW/
AZpj6EUW2XZ1L2VygWjXE2HW+PrciNMFZyQ/cpRJxcVcDldoZl76iSBOkgip+ydZAiwHIVj79av3
78RmEf2DW1JBWAwx8vY/P2u+Yn2OraftBMx5fZR0cd3BoJGVgTWet3aOvhw+37RbjRyF79EjTOgq
d0CtPRn7jHEkIYkqdR/zTNlvX1KqlzyVle8M0cguJcsFQb8cUHuWNWwxsmwNR56UnnhCrwIZ6ckA
Tgy471OFNfKgNDpZ9MVHCouFJ4BzexkdY1b6al4sbOTU8HsNu4z/OHzheY+IZbo/eKnY7qHBRVZb
ZWI67rZZx12PFXlzx0SvXtmIvBiFwzHBw7Vb9xQE8jfGSpDgpKuSg9UlppeNrpKzD7iS0i/VnA0I
AI17rrfYnaeGhdmae2SQFGs8seQTwpjBD3KIWVHDxASiJIOBmJ9408xC1YdKA/qdssZtL+AMLChi
Nk7Msg6gc8Pcuv/c4XoBRIMH6TWmoTb0Z7tlkJnxqy1YVJvu95Y09Db3H4jtredmas8sQvFQi8DA
bMb/VG4gnMSUPxZGOuCjgmOS3DMJ777F6L8B1J/PFqRlrfJhCZzV2PjgHjQ0Qtozljrx2QdAb4CD
YS+OObE+UxvpcCg+l1aYU2QTmQT9vKYxSXooOvAZXrhTw1LEuNHg/QnRUdcoa9aodnJ6haFExnyy
66EUNH8u8Bb3Vz06kNPdWw3Tig2zVkUmuexI4tW6h4gJQllEipXPEupQ6u44WYouCa2HrXFEwviM
PEwy6NnqXQCps+BICnIpsascwF0QPf4WROKR+Nxlcqm8ET4zBouH/62uHylBLDk69JSqotY8yAFR
FTAup4n4EZ9BHwzBIfU9sI5XfJV9prkyjXkLx897gj4pJfib3lvL29f/bpWjeGZg04mKiyJmbVwp
UUEbRrgWlN1NOdudMiZyMJLmBaXrqxDahnXva5sWRzSIL8fD5cvZfuZXdDER9P+yOaEJaQ/vFiCn
QiEAyw/iIT7lvL/7nngimoFfygd9ewTZeHEbUCZ7J1FII6wlkhm3iheJZTENXDtHKGaGGTs7zGao
07R8RlRcRVkwr+1DKLbtSa3EE7VTw15Uvc+PQgBT6in98QkB8EEwZaJz5odFDTBb/eQW7anN0qRD
c2KRyBSiFWnwYn8s+ce4c/mwYJ3y1YA6VHzIGMA7GshRv4+IXv4QrzOmsXDnmNVvsgDTTFLkShrl
dLseoHL8TOVFXiIeiQQoSOJKKqage6iQOmb8IvJc0mf1YxcaPLlDT5xB7kAtiqYPZ8mnp96BddXG
4a3Mlv2hv5nwWIkRWgkL7Ukm+ztPvVj+otYpDwYIchnD1ASCMSo5BGh/wPl8vqDufWvvWBamutfu
R+H6n0bZEHVaRpRkekygVUgDXP9FSjL/UiwN1qDMz6T6YT+MAw0H2iw22yHo9fC0t1mGUQvF16b6
AyIj9YhSkuAoFhMUjQqFTtWou9HQJqSwMIIfUvodYLay5RqRaWm60B9Hn468qgiZJUkUz3iSD8qY
rnouHWbAYc6nGZ7X88fwEJszDvauwN495JJhwZa8JOI6s+03FcEBc69g/srFMpr0N0VmS3xbxGjI
DOaiMr+Aj+D2DKkDwcH6jzzlLzsTVY50uTM3j5/+jHUQDGJAFAetzoaulH5xByYAMGayEXefxJ9G
CZq7pABAlZFLHzgWu1gAWb0s3+lKzHWH/rfB0uodOp43m+vNWbUIX28QpzGrFh2EZyTVYTBsDvCy
PcqnntVEtndkYzbmq01LRikXHpbBSqOyV8vJwFFRi2xqR7o80dWdDyJIvk981ykr5ND0L9fPO3S6
qNqnzXTcWQCK7BCYWuJzE4KyfY+UUr+WCUSaj1d6J6/BYA0Cj81Dcydomj1KP3+M1wzYWQV+lyBI
Sh5Qk2l2/sElaDyz6r6cfqosGBOVVckFTaDzZZkLnRQFN7qJG/UAkJfuZ4zprBpCuyxKu1VMpjFW
7sy+CI/BpYgApZpKVeRoScb++ASNSWxzRBY9bas7gARcoY4i5dnD9B0LnVdAenksxCaQKi6NMyuU
opdBsQj5J9mzTkmfqwvO+XBJx+D/EqXHGpX8olV/oG7AGIC6fumZbW62K63d1B8OWI3AWx/CK9bS
6ZepxeET9hIawyXu7kTGzTMQY9yvESmICL0bTKu8zcD+reGsXPYZqSCd4UP+maW9aXZNpGX7r2xY
vOYdHO6gTxXES8hISwo3T9Ai6fOqtcfL3nxTTLK3m/Gg2fvyGNDgCTF04b/5XflCt9NJyjd9vOQR
B7KMRQYxZ1TMrBkK1hoSQVEkcEqcgeGOQx3nscIDvrAByJdSHVIx/x9ZmaSMgkV8vsZeUi9eTxru
4Kz8WYIexdhRtN8+Hrdhboo62LCMqbkWJSfpISFkmdy3kDW15zzGjfnhZQmzmZfsrAuG18BZYRky
9UjOm3cal8sg5MW2/fVBSGeyNGCm6sSzwj5Efci2FP07Jr4ZhMUjN1N5OJkqeTLscTuyClndSOnX
cRCv3Dz2u3UQINGswpUyJv5DrWxnJpMGPVvc23VipAJkUwkwgfSKhW+2qbCx8+9wmJiGGdl0QPbf
D3/BIrF71ssPEw1me7MrkjbAnVwEZ8QrS+XCK/g7vAJjRKF4ypczX8q55rX2YdmX5QNu49O7jHoV
jZzLHXr2yRqWlVyQAiZjpbYeekwX9bx4WiGjmlnSf3Fuv8Y9a/5WfEXlqrT0bXmTSBO3dcXV75jV
z6eUvMxWOAxfsK2CLbnGUsJbn/rI7AxZptSsxIfZhamLhlmWCf0aOZlK/DFASO1LYSjiS6+FZByw
tF/UYzQHvuAy5ULxGN0LwqbB/9uwrFv7co57TnracESn4Ai3RYCoQXACSXgX4dOTrN8Qv/WPwshU
fMumcb0yQlCWskRx7gekn0Ph4PitLs1hb04o3UXUI7f3mJsVXrqvJWXmkExvMNo74TrHrUHg86GR
Ch+F2bj4vHcZftie+Hu0FxWsBPoxAfrIGr2Bo+GjKCvJufMLrdMuoj0yKJqStUTuO9g+jWpts+9q
wYEJO7rlnzirEjABSBaQ/Pebyj/n/6ni/aSsVxYkK8ChMH0LC/Xq/GFVLpMOisk1k9Xc94Od1hbs
eklC0SczceYerZObi/snsq9HVsQTZKiwfQ86453sBfNUJW8GFYGlnDnKT7jLMDvFWBDs+297k9Cr
oJZ/O/prORb1n8ax37DcpKnW4lIkmIM7LmZHcGsaJA2aaqANkgYIrqpzW4PjigtkePLUeDqejjTF
abyjx9nBMy+PxZFCYagIvC9SAfOLW9yFYJFoxdCQAaNvMvHYiIPIeFGonITZUm4e1PxynxWEmvTo
Vg8nZ/pARzcX4oiP5gn+ub1rIrCSInOhhkPI/48fSinJ+NQNxws4G5Xo6VmjLhE0JNgTTMqwyah1
AbnCV7qb0xLFENn7bA9cxDpKkTJmAidBWSn/CT1rOGdQRf4x8DsiBhg3jklo6MzHDr/cCcs3ykjj
mk7fgammHsOMMuOk1m/UGMoh5998+bVwHLtuusDcwCc3+NEE3/hqVVcvGsG+YMIQzrzF+2UcV5Ln
Yc7xfS5TcQmBS2Ioz6VFHlhqn0C5XRgLzSYyFmV4nKqnRNIjXFJXPZFDDN+dl9w0UR9ZLaW8yzAB
aIEVKQgWKK/cIgMO3hEpyJWrUGiRtugU4oV3s1PquBdAKJXVe98FLCTEnPbv+xgWYnRS0H3My64R
BgflnxF1HTBP65j4nC8N7KQnxLrf3GOxlZIwwIBFKh72qzlQZ8hRRggvzFvLOdrYNyrzBvpA2bt3
e7SAdXxithzxihoYb1JSdSySEtJds+XYNhuE4kTdGs/5eTzr9+GyRC5KUGwo+UAt4vkmz1AZs0ZV
tRsHpE8q7XxdP81dkwIsyEgGcIV+NnukoeYOWjrQyXqoR3VXzNcyr5UaZi8iVrMdPGsEBpfdqKjk
jDNK4BDuxRgaR59fsjeIpcz5Renhkz7PywN/ONeIAM2NUDDnAqH3RTXSB69bqd+qfdU0JtVtv27u
wU0N6Z/BCUNYJ+tE9xHNqnX1JLwCtK904M7l8eNy4VlQhw6nf9SrOjv/MNdy5kTfFYl62fD7Gk6v
RyprRtR3YWh1MgfHu+SDYtLomn9wh2A3UzYx7bgtGdX53i5Lp4TvKthm4nvXT/zjQRcp+vriFHo3
CNwI9mlfkJLdVglVC5AYACk1SPNljQuJkDVRaedDxREiq6YmPUJA8t1eOCTigAr68UXgHC3ODmmD
qfuqoXbyVdKpYnp+iUAUYhml6NBhtkVTiYjK5WwCZcf2B6zPf3zsA0peGoAAlNbiVF80RYUtJgKr
erK5kbRvaSWydeKXErnDIT09kFiPLHiqazxRlPglIPbS/9H2DflWgLFQMeQBKlcjClFBPUyf91lz
J5C9HY8c24HpoRU2awOJdg91WkS/+NhY2xuYEwoKLdAWBmrZd+UKAGUZBncbux5q2sTK5zyaX+km
UcrqdkRb+BUZPgk7dFdWMXUGkaBhQnyuBV8HvCPadw0GSalkXS8MVNxfBhpxpJk58ZXWtzZi8N7D
5Y/BldpcbM8MXuru/i6bwyFGKmO8/3Nva+ENJXMnvzTHeSJIJEXeNDmvKsOyvxRFinLHV/OQnqrN
51BA5EIkdPvD2BDKrK3OyK6akt3kw5nM73A+6lnM2sfFkSXRyTOB1HCNVF6txd6WzDYC73Z98zvS
jOjRAUAJ5oUakzNkjOSNdAS1Fk+cpsCQz49DOZ3ML8foG5z/E6tTVG9rzX3VnaP67ReR6NBSWzcO
yQtoKT0CDpyVxqlEYGqSN9xhYrBDZy2Etj9RVQSTA7kyiAUJ7KI8zaiKqdqfjB/P/V1DBLSoFvuL
YXy80kjluK3XiLI7eQ4BIy0bXiJbRf8O3e1lcnewPJT9LFA4XarmkRRA/MSy72dqaqQNsexQ/0jJ
Yt0i3+roz7fZ3oKPFy60peyh6FCR8osIAomi92PRYPgiaZb3yMVT1LEMrAVqAtj5+gwbni+EH/yh
W1ELaufVZZySRMJciG1SxwAh9UEsITP0RKmkJ1oAWoDsgYiCPUNEMxNu2PkdnoSYRxL4G1NK1PKN
QAsvCi1PgqnP19sgXqROHVi/gwK+K9bxoAqtFHKyTSwAMV+7sbHWUl1gmHWZuLSGzel8SNhOV2SA
9etW6ZvI1Ba30JXOBxuwd9Uu9VEHd4hirXDN95teWHxeYCOFKGRkBDN7xh2OwikTvd6cDY+Cc40v
QSweAuUqTPqDi1VplVq9bAJT+deYObvxr2F3R3X9VpL7r/8+LDs+93rCj6RwIsv2bdQyKnKINf0I
8QZf9ZDMitiSdZLdV8XnCFQ0doL5PgW707JyLFXDRzqhAs7buuFe8KML60SovJ558WX9r+H10w0c
8EbSVmyOXIbqEQzhCqbHZW1HuwkyLEhbo8R40ic7xZkNuWoEf1SKWLjcxXtnyx2A/OCEovqUo4e+
EkeQm0zW3WyH53Lsox9dATi3Kw91Ya0t4EsMHSMgdk6JAghqdQHGrOJr4BkoYr2T35XQkKHY4Ym9
no4zpG86mWyCoE5PHjIWFhDfhBUM56ry4OauT5Pg0Jp0u7skSHikA8+w9nZc9oq6UV4wQ75Bhz6J
2dNye0cttlGbGH/C5jrQJ5hzePuwpIMfYtR8EleHUb0zPuyovTEI4YN07F08Yek9jrcexMAuALNp
TJHGoQSE2yIdEFSbTDxqtr5rF7WuVa2nYTCy4oHe3RdnTbnjNUOUUEJKTlAdmt9ULDbh/c5gA/Gx
10pfNPmCT2RboLKPivndfjPj0i//Bsyxt/KSkZNqrqQkIRzOQsxcJsFN+DVXJIvmDZ4sxmPXZ+rm
Gdb6INop+xgtrI9TOvhQPwDQLemv1msptsXVnsmaySTakZaeuDiC5NYApycI57nR7yKlJ/ANxblT
cXFbwspoyxIQa5AS1frro/FJ+PMX8O3yZbjNtUgxsCJrssBlWF1WAKxg8e7wQmN90T3TD3/jfySd
mjOIzqfxKRFXYtmbYUXKrkITitDDr7j8udMhHzn7ugeLpJeqE2AR5yCw1mtHG+h6VgV9ZEzrttEl
Rlf/6da3G3MICGcRTTsV2yT37K+/2+DbI8da+98x4e3M8Tc6SkhLXMM56CPmT81aA9rRGjFwc5LR
/hDyyJzMygSM1hZeauuCBvVgvknOkybu1dLwZHqJd8NFBoCMBS1Fg9lOobNE/Tm98Kw+UoIu27SI
WnWgZ2gEcGnLBvdgvXXBQ9dHauDDkAOPQRaCaYxI/m6Hn/iT8ydW/f4ranZEc5ChBebflR7TnlgD
TSf/JOPqNXv5l+fnLfuVMgzMO69UXuhcMsfQopWIlriiWXl1P2pwtAX8sQH/tcr2W8M9LGL0+F5q
d4Nqlsc33Y03Esp6rBuAK7qvNZ1wRPadix97RS2A3/zxejGgLDFNedMDYu8a7XWjD+knmCVB5lQB
RIHR71et65k1h6iL/g5WunB0qqbJXcE45DSNEr6Xz+vHUBdeNVokh+9DQLT59x0WU98FiZdawrKO
kj85/ypuMsKaHgkwkExcW8JaMuzDxYgwvqZ2hL/4BgOYr8nwaAaLoU5TUqLcZAmOk8bc6fWX4oyF
ybCScdDt/p52F02/i9atWmizb79mLpIcfYv/fitGzWoyuusWQu+AHodUiQHvqjmZ8ah5RfTrkf0z
a/FvNkCwyXgCt7Qq2j+fpZF5qPabiWX0NP6wx3Lhmeh59Sz4eykGx5n/QzUqqDjoCgStYqXPpjH9
m53DftnVufy3eUY3u8vy9H2qUQF9NEPeIRK2KunIaX5wlwLoSmEwkRNXdqqFU3fWh1PZvtUasgsv
6Pc6rGWzeasYjK53owZEJQn0mMvOGI6YMUpbIj317jAlR6VbtLAJB2X96i9EI5xyIy2AfAvj24GF
uPPpA0nmWg849Wz1RxOTkeSEtvGo4VXqhI5NblH2sSbCvj6IxAxeqUrgOwVInOsSjiGvNTJRLNhY
qrd9uVz72tsGoxVF0X3HE8z4sxBWOWW5RzaatXegew7YFp5I6raUnkbUPhQO0Hvjx0/JVfxLLcSO
yL2IMHcKy+RNe5V/IN72tXNXlVGXueT76mxJ3QyOBcXFVOCzHjx1Ha1fZ/zj8siKywKF6IoPfEhl
0HbgpD4PQg8e/yyAxIjWnqHawO4iSWrptnzEZh6utzWbiE7mTyeqk2aoyMgzJsaryOYa+vCpWyfl
l+zKnc5sqSHwnHqQm9WunoY/rDeY9JcZw900680wy+5g0H2KMkL1NA2IzfyIFK4yYukWmm0MiSOB
aibwtIM36ujAvhqPksNANJat6tbzbHnwZQugzX+AsloCha5t5b6pvjHhJt03RQxuCUPjwE/lZ5mq
ZPjo9xHi/7A5uHPuhxH8yUry4fOYl9Ji2NQlDSSDqsMi1ikVtp5KRsm6M1sd6FPHAkuVZ7PwKVyP
utNZ2srX2QK1oUi+wiaZUSWDX9/R9sDa+9ozIjTeoRuzGszm92TabEXOwKbZ3+uWnrudCof0rzZq
ZaYcRXAtxyBsPZuxHPd1BmWFzqwBbSs0anWX34Fw3TMikiZmsIbnRnourWM6ELqSA3p/o+/P/S13
2JMV0+o1ydaBonXseFue/T9HuKOVulmhlyzIY6mRwuFyjJ4KoP32Sh5yNgvdE7Lh+j7RKe+dbvFG
Z5q86k6urTtxiD7fI9lUIUwsviMnmb5M1+LQeZ6ursmf4tML9f7adppNGyaq9w4FdSCjh/CVJCvq
Vgk2eEThJNG1nbt6/9ANaCfWW8QgSrhuMxZZPdBcA6gXH9Qiawgjfvxr7t20FiZvnok4w34XllGB
LUfQffsU5ecUWy5f+Fuc7fFEWFUX2CBuhev0YEdGkudHRJXKfHYZzWWeE/wQeDzhq3tFkNPTKmRs
+A7DQEv5wlMjxGoQpOa9NuqavokI+Ac3vvVL26IKoVTDqLifPDvD2LWfFD7AFzVJUWWsfzqCR+b6
QXp2vTY7MLg9hBQMwF8oCLBm1qHDcvAcByeHxkU60OEwxXztE6sDrrslmn2cPDrbqZki3lBtA5CR
sLbuvFua6JfZ4Y8xWcX7EQMK8/zJbmtCYHAZVGSLR7Oa+jAVdCuebC1qKExzb8WdO6ab3JoVk9rL
WAeavU3GRDMJW3siBj62oZuq8RuE6Ckx5ROaEMSjqaUVJJTSdFnjZsWGPn9qrg0gcIIPYgXzgan0
KPMRkZR6GifTMcca6DiAPe8IFPMkfWGjXRBwgwmbDl6/6/n5IsDZ2IU5nhv6liKNfo2njGtgGQTo
NbR7rFLA/0A+UJwknn9tTukEAhYpS5t6YffaUjYz6PwTJq4QpQT0l6alUZccaUkHszmvQadLlScV
ccdmtQ0e6RB6YOGB3n63jxu75r3jAze18SdzfIz2zSNGdw59m/MlPNdigDGAcAZkdHCgzORKNfMT
Ab2RWvC8b3neQRmxRN6E0DTpkDZkWK/ZKN2M2rRtmeegX7zLUYwLd22VUFbkMiuFeVBUa3mtolAh
doz6NNhmQhe3A8TobXBs/PXzD9iMsFtoWf5psFFwzi9TR2gaJJZKjtedwkHBu5LP5QSDaccbJdtR
B92n+a8elQP4ohcGikz39aJ1rLR2pszSsgFDGzDgQcM95okMdaZGh2LRtCasoSU5tb7M9RSlXVrK
CkIOgS6XifEWU2AAFC7YIBJq/rM5FbfCQnA8ZvnEraiAsqr3CN1Sbvv/A3l+cNmfgHFQaSrR0Q6r
Aq/nByJtX7uDUPOa6BzhA7mVFqLfrFgPvFy8jOLTsw0PbC0aoPVvxLsY7IHU/2EG8iq6d5I119yI
z017DqDfyJSHr/Vf1seMQ/b5Bw0t+odXb3+4mqjaBguk5+sdcd8RAKxpXTeH91p0hUZQa92rJxLy
u6B3i2tJjjJ175q3D+AySIGtcgsUJLuMl9nstHnUWVnPs5gV++YST+ijJHeVoHuWVfhQHVdZOSRp
1rcbeyMyvBluXle8t871aHbt3m+peja/4YCPq58YsuuGgDdvkXbG0IJWCJlm4XRQqgs/m7Y5I9bR
KmqfBmtMU7XQJ1CRZqOZ/ZZJBRaDDyD7zSUd7cSUW+vlXs2c3iQWdHtt4rxWZamW75ppliTScyPC
Ad+Y20NGC3z7hfd8ziwMbA7us85A0OuEsg33DTlf2Vx6fqNazcN6WIqllS0400lK4dUENVbKwOnD
BJeRL18MWMFYzZA/f1Xi00tGi53twZSTs8FrAFvXiMsu7DA43fCIAx3tzaCmzQOIJpb7H0Iw0UCB
db6YL8YjPSxad69MqWcHBd5syI4GXLmWL0FLIgRseVaqTL6eKe/TxnNbxHYslEzXwYEF5AtKvFK6
NbWLyJ14eqBAZ5gwb/qgcUjgWOd3C0YF0jAelqWUTmyF9fg1NiAd7N0csJI8eYhAR7naUorbCZrl
JDWOsLY4nfVS1PK4qeQ00jCIznYpqrkl/B3XI5rtfcpKjsNeWnkib8GItc8yVByhJgQG5McU/QpR
UBKdW3b624lC2U3stlV97+DzUEBhb8gwisREHJ5q7w8Y2v2MLxvsJlIIu8UwR+hGBDqVgYGhbPoA
Q+rbLqXiG53ecRVCwgvHJcT+Tj036Z1sIXgzp6xFLW/Ni61rUXzwyo56vDnPunrmaX1Mzg8izYm4
pST3R7hp1SwXCvzpBtwLpmU6KIBnmnI71EgYwpoB8v5BuqJLIj3fggfLcmcKtk3JfGPUsA2u7EY4
HtcrFu1izsPM1ZdPVkRmJNcVmX6tzRNur5zif/PiNA5D5ogCFB0vjupMNV4LA/2bzr2g8m9ugdlG
xQEDoHmxUGXxK1//G23fIKIIXqUnqAeT5CVEdXHvRlAMs8cfSzi+s/EO5oDRV4sYNhWleuUpnn3y
Kq58UivInsYHtAkCNSkWQb5BCoVvjLNh6PgiCJlhogbFdS1Z25XXcOOD1BEu9mmgfDW/NtA2Dxh/
c+K2stWcL1WBO5LidB6nfuW2YQiAzkY2pR2obrVhjOsMAAtCXsfDBXkm3LMxzR2E0i8z9Tgd3X+4
QdvfGD5FM/Ij9HpQD9d45WrD3a4Oi8zGyjGhVR+e40A3X1hfuhFko1AB/x1HA3N0E64+yFy8/a8A
Jbsxlzt/dl36SiL8A41qA8PLnRd4Jj0ZdXV6nFuNRCBfBK1Y3Gt37Na9w8L4FhyJcLASWokT44ww
PqTq3HtpjoCLFOVWyZ8h0+8Of4XO0b3gvp1mZjRTlZe4h/T2+Gdqgcq1pOqpibWDtlzcZt4hcWJt
fSnU90MWLy3Yv5IQw94H1gb5/Z+Q075gGXluCKqN0Ln66+1YGYhjgqDlN3QcJ0TxVPa7SloPhuoi
FM+K7kBcN0mkbFWo54yUKPXZt0A+PEmAbiwt7DiJC383kZtfQCeMt4vNkE8o0uZOfHxUvgjGfRws
P0VraFTD3iVRWZz41suFSwrwZabSRyaCGs0ncxWyrxQNLNCmApF5SMQu3N5VDIJcYE2bFIEvaF7e
kLdmDbewp8I/8D00+7zW8oSl+cLjt3r1niBSrzogAa7Jk6U7M0rks4zx0ERMKPOdHYzCfVOckjo8
/hcIrggLatUJPkVxAqhC/0Kn0ENvuURJ8pCZ1Zfkm6h2XcTrL77Zu1NAZWpv+BtDD/+tLgdgu6Bx
rx79jDioHoZ12R0SytXWAQz83DuDL+dkeWIwuf0fNWX8FfGTn9N1Hz4NvYSPt8L+vp0xmEMPgStG
y59LR4zN4NsL+w3q5cd0+VXMuSD1f57/1kGleqbjHPl8Si5sQDQDHgSuZEkC1t0mVfqFkhynyte9
WDpXsSUGzusHShEkSjY3xP5A8muuhhTbzkbcNbKNXIgzlwr7Ue8PvHVxbN1qVp3l2lSDfa//qkSh
kDCWGo/MreBUE2nlg+eQvpzwIih+1nBRWtzZ0iKr7k/PcvIfbztQG6LeXJHjWzZR4DM2JKfALFTH
MyTLaZEvAFxMWmm+tzDRY+q0ZpnzhbMzt9okMypQj5F8K4JEzYBe31Uf5hOl0zrGzrmCxVdZRT7i
73m4WO9OH4+euG6O548ijN0OoC1x9OhxJ9Um1RtzrtK6gmWcjpcyM58eH119xBbeNKdUS76BhL6b
Sq7m76DVSZowtB0F+s/DkkS2NvfBqJ60lesOWV5JBQSRskaGj2znErwEHl4nCpniPPUSQ2nHPSa/
5O+quhUcYy7jI49WS+/Uwvn9ecJTw55kv5rXnHezX8nIz7eXyLqr8Y0AtlWthxdC+e2V3stJvHZX
+41J7DeVLO2fFnE7OReeel7F6uoXdAXGymDgkR0QIUUvxqfM/iBMmwP+odk+JIfRShNFXKMeKWlh
5/Pd+NrSvCwhvd8QtB8o82wvHiIXxvAkGWvBcWwj9vsoFWgmbNEaYCLNzJHA96g+pEpA/k+wUgeP
bjXK51HDYqYRUM+txm4nQB+DlgVURKmsxYnHHAWE/MVzrW7svQsLTuk+njhG1f4byWCrLLzwV/IM
ZFM+s9Pc/CQ4FMw2hUfrPpE5IeBJvQ0cDPfAFVU+J/nmWUV+FPV07to0RVuOGaCi/0exkJ/qMGQm
Gn91/x/HWP8Ez+Zhyd0/9iSjrF1Y/Q+rAGgs7TDwetclQQWFprzon8VhBRQgLBF0+D9eL6Qu3fqV
+TQsQPjC/ZjBMZ21SBjIUfhaE286KqFr2qYohpSvF0ZU0scej4cYbkyCwepl0udMpXB0Uz3kHKki
an1FX2/2DHyrdoM4LTCBPMyUlrho7krRSbScuVUCYgV6jQt5r1SKJpzH4XDQKCPwQiCupGYnvmJh
X3xmNKbHVFkRITttiRAR0T1yUylcPRfYjQgq8MwYukQsGVTKkiRLguj/O7HcUC8Zavhrmc0ruLuW
oaz5t25weCJrZjJRiOnvs5+EvFEdcbpIyM9hnEGwX7ZS3fZm3QHR33CHlMdDP4SmW1iMtco4M2Lv
0/HWFzWso/5PjzLxNjC9Cegrz0k8r9dcvyPvFjwuGBjs7fFeNd1/x8CGXCrmUIiB3NSdy/5sS0jH
aZCtvLxjuEhETFU2hwfOIJpYdsBNOgwbrEXdOnfg+v95IRWGcwi+zNBCcpYint0SR2eQRHl38uOZ
eJpNwpmS9W6IxbvrD0h4w5lPqglPPOaChiEmUqD7Yq+Na1j5g5C6OFs9dpQ7Hr6Lc5qB/PpP0CfJ
EkeEHnCgqEm9YPG6cemufW22Y4YDg2vg6/snjjRKW84zvZDAAf5PRKvGC/p/nvfxfIEwyhVC92RH
iDV9eXSd7OMsHFICCkYVaPhOPmnlw3b3LB9oo8NmbK/eAmtcciRAg5BWGesIgrJ3CIjQVNhx0+F6
GFvF2Ogk6Eu14Wi9ZlgKsCNFq9oh5LpoXeq74+GtOUtE+I1vPZnY0mKmE0sLOOTrQ5emZWS/wxAa
kg0mWuyyFHB4NTad1hnHh7i1WrxfH1WniqtsZMQOWKVFmaOpGPi3nIvQqeaCCjCPHFhm1R/7Wnr4
1W20qqWyLF1Dek1kIxUkal22xnfs8rrRKZUDBX0dm5yuV/iEHpT7hEfBMwh8QRWFEvF2HiiULG/0
1UHDsvRC+9+MRVG2e/1DE2oBH5Q2P7YD8Dr2GeXf5xPxUb5Z0iTQjmdul8I3CjGN2KeCIoR9wB7N
XtSnFiD3WGHcF7JjSaxJm3aKHjya1zBiDjFgl9X3rtNxeWjTwVilBTOKDAe1jLjZGhJzigg9pQ8f
NKfqMMBDId24JilRZD4ENq4k7f8JlOLwXr7YSgd2pMcDUO0dEv5anNVViT8xKXJ49b2/bsUHMQ+P
O7xl4aqKBpfBhFC8ZnyQQQPfg5A+226E/UL/BpmoyR+OdB0Guxt0SYCTJ+SjBZxPQx6u9t6KjlhL
ZsuJ8S61wMxHXTaA5kqEElNQVhwob7Z4BjMwwB0ca+zYhqy5CJERbzmmA5L2IhjJCPL+xITeq09s
fE3F9qS4XB73U05WO7s6ktzU9TRuh/wTrKjMi7LGzqflapqGGV2tBFjBO2x0+mmdeyJuPPdyVw7W
nxb5MdG5cNNPdAQvH0gcJjueD0RHtGJrvl6ajH0uCqW2WM+Dev8T4ywEiHLJ/X3Zl/eTe4ERVzqd
PKxXP9Ds2CH4TlU4JqFCZ7vHG6JU0U8CJKrtwHcxZK4BOH9FwyqupAVEJloYoxv3l04LBewIytNy
tRMzzQL7eijARPlC53I9hUYJIZ/SyD2bm7IwJEEiZegIp14DWpCo8U0Uy+5MnmPZJrsMpuxkxgkG
l/GH3rZ2KF6vBYprSMOAhDqF9jt8yyXii0Wc3iAy6wY2RSS8equIC1cB1lA1c3qh64L7dzhajMr4
I0kMFRaInHI5ojc701NANQeXvpS4xWxsDj8ohl3R9THASZAsoc3jekWNP+CsljsbzlySxZXKoNv/
eiHu9prDy3qK8nlrv38BTZeRqWohbDQhZM8qBKDbJ9LVXXrXDvZbv0uYngXRDuLSucvF7WXIy6Ew
eYBEfqA9yQr7OPoLcCiNN/dnYy/u+B/2bEif17v1buksZrmgqb95psyuQE327JYGa5dLgAsbQnVz
sPhbMQE9YkYPyao3qHnJaOni7MrYSGyW999RZKjgi9jCB4p27Aql6rVP1svw9vDb5n07jpeFZsM2
P2+ciT1Pk9QS6KLeRyNE2f2tfgA6BtWs8N1eGEQy+Iw1wqgStR9pTo6gLAbxpakq1yaGX4LG2TTE
2yanM/mfmm2d16cQAtAkEXW8sUL917ZesefwDVdATQJiSlP77RU+mQNUlSAtz2xrP+a7CkEovIgh
7wTkQuuotfEijznYPbTqFOtv0g5E1tfJBL0vejaA6zC4t+r1Aot26Xz+52VOWscHlccgoDbMMD5o
squ/usSWBdpkPjc2ARj/Lcf2OZLgADTl2xX0oXQzHgpbC5O7taq1gU4nIqxf2axu2VbSmKsKttI1
DF22udwloenmif7+QWIVw+Cdecm1nZ13tTvOhUYSKFbXwNypRhldD6bRvvCX0XiOZMwkJ4wgBkkC
JAh9kshMxPP4pNwQxJOOS8u4GHN4dlJvdSCvktXlAG7e7s6pFmoLJs9Z4fWAGKIxW/BqX9Ucx2wd
OgJM72hG21R6tvMczihz40YlTLa8/2XyjdJaNuQqpPZMPu0X2PzejGtSqJeMmpaZAQFTLWeVjzro
VCEyJo8XcydGPlcNHv86C1lBRjLgnalb2OJLmQC1vChSl1gLFUAvF3Wt84zb7CwpMoDvIjITZIzo
Fdu6vib/cU1rHf9rKdWvqyxKMcRx00pwDhGtPf2uCOfEXTThqMfiYWOKFUZ1Mm+FwdsX1OOtr9QD
Imn3BpjAnr4QVBK0pnfVo61g73GjJu7BjXC1VsY56lJkYl0TAZ/O5rOBZ+KhfrUMg/ZpV221Y9Af
FwYyORKrHxJh8JY4WGeGGo8odrFq+MWcufXz55MP/uffcx6phtw40LMR1BXPbGtAlEVY/G7OXTJ5
DozutKWoU0AhPyYGQ+OJVJdtO4SihDHCPuEDeb14Otm6oWWGZf+7uGThmez4u6OKpSklRhIvqrmh
3mZ4UNx0GCI0BDmxbt3dLGIzKzUEqAHGOwQwHIcgFuCv7cArMuGro5pHZdTXBkvQ7V5mRqI4imjq
Ts3We0LGZD1ALWr/2xbRCZamPjLMzRdhKaJVVoyXEcdsH5Ybp34FAjlYe2Fil4hXMSrRiCVxqPlR
uxAyC3MXg1eRQdehpLyOQ7lfA2y9FsOQc1NGW5fyQNU4Www+NACz3DZzNH2Kuk4KVGMwDcYJNjqT
bF/reDIgZ6sePcTi2IPqGi/DCE9H2bTkC4rpR1S+4GOjGWaGvZqBFAbIfrwF8H3QLsifNGs025J8
9uevW8vwyBkeHCiK1ZwtLyQCzaZO85na9rX0HkLmpE+kkL0zDTaT7phyFbwpE/XQBq+I/0nPyYZl
LnUNATtoNqdz+bK98arWM8G6KWNjO0NGgVwEIu1uVvdkgdBVW2wviaobWAd9n9GXKLvnBO/YWfyT
vqoQM3H9GhGYgkjpBBv7Ue0O2eTl97VGXL4CqLP4QLxYXNZL+rXZbwRVfJxGHxnKOduqTrPHqPK6
o6jgu0VO5/6yZplWXauLzz6UTiy1eduVJ8CHUDpjxCYB41uGu6uWh8/W+/g1TJFS0FXO7p7E2WSH
e/PWz9KiDJMJ95Wc0OlZIiLXL0p6ySBxh2f3PLA4FotIH4tQ3TnvqTRdUKfQjUnmqsQgC0Yahaf4
8fxr/Rme3qYLhguWhkPHb80eHUPYwLVUejDYJo32g+vb/tH3fCKFEtBvNnpINmwiGJOh1CAUgB7h
YISAlPZxikXBbNg9tNf4N1pF2QR+mVa/izSN/wy2jRNuZPGFhoBaveRiHb6vBPr9iFrcT6fjlOjC
H7+LDSw36nzs7C6z+UCEaJ8ba5+Y/qNmOfRpYg5Q0s1+CAwZ2fgoAQHK8jG5mwThYxwpuFUW/1Lx
4P/zs0SUPvr25lwKvVgd2ShhG7SglXJweNwsll2hEjV5K4lMGvDHdU8N+OoqyfTf2ydclxS3jdXl
Mva+LXZcJu//1w9GeZ8lyFy0ABFtSkZiyZBqA/J6nXbMyIhOXddSfJUgiwbnbpnC91ebfdQm+CN6
ytTPF3fXktFAqvX7rJsAl2b6qeuCV9Y1N8jTdG7nEF257QlOtbjL1s/we2EJ3+zoYi/I2QQ2RqoG
Pkr532xJLrFrLw4glWBmNfcL7A3ZfZhDzCmyiJhiHoqngEZMXaKTtVigs+yhQ+ONkVjxgs7wpdvo
5KVcha4k+ea9Lv0Gs/8/vv/IU0J/9MpP6hQnDyCBxUCzfkWB+i5KlOR9MzkdSF/8xeb+e4uFesjP
SqkdzYvMHAfpNd4Eo3r7q5SZmk/PctDY1EMgRwcitJzBqfV+ya0tGmamqJDSoaLunZSkB+VURvW/
fcc3dFWMnojtRX5mLJ33emNGD3wZGkId4qagu0t3t0T8/uVvwSkGPgLHp3k0hmRsqzToV9lvlrVi
H08/IbDczFJM6IB7+kJnJEt+I1kaQQnwe9sQrC6Ol5gd/2xQHtuvByvjclfWK447ev1GaLKR5lgH
3K8jhDT9giK5mHoo/V9Oz43SsRmoVp59/4WHvvjFpQLqIYHbxsZ17+KKQyX4dkMCy/Z0Qxzgo5zE
6i5cdLxPlT1XBOuKFR8CMnprKR6ey+ZfXT3Ku111jlWCS+rO+3nxFbnfNaay1CoALk7YM2tfw2fn
Tf3ovaejzn7JX9Yerg6Ft8xgRVr7ikNjASXtw9h/bgg9YcXQBbYFWr7eeB8hiHs8B4rJl/aKd0oM
V3LVj4Uo7Gsse0dF3YQZT0dVqeW2YFTCe2QHxFKgTURsQtMp4sGIzZMWZo+FyL8bAcOC0+tQpQok
b2sHqUxd2XBue/4Auhp0NX3JGM3PKOEpxnMi9AZcLMYBo+t2nS9gfOJBjCyqP1DfC0DweS+y2tBk
l+WFwPXz6lyW7IbpEU0Lw9QEUgR1YxRdXg6gvlHnkSnh7d4H8En205iGYSTdrHVyR7lnNxZMb8BF
EcTwmL94MihVihmx2qkje63pmo+ShMeS/EvttLuoL02NtjeO8KF/oiOADxg69/sj5h62xau9dYnO
PO4VqD4Ex75ZMQFCjPEhGQT/Iytaxe8HDrTAgvrrt90gNIRqC8KEUgt1ATSXlh/E87BFC01mRmmm
aUG4ZHi7Qt8SPgSklHRLhpVTWjHE7aN6YcpIBstT1Ox3V4wOrj/+YOotQPQEqVLREdOFaUtgHUaf
a/KKfDKn+l845fawy3T0KD2VpgUTOKIkweehcU0tO+FcFp8Uz4MiSo0Oyu4HVBeSWKSgkiJASyI9
f8+S1eVnjS2grnlkvCjbjor7BaGuXrCtLLItgB54y6R90i2VgvSxp4S4C0Oary19sgpEKWmqUNJU
UIPGctwinfnzvWwv2iv5KQ+9S63/WiyAC3VED6bLsmTagv0HcitkKP5WhmIwrhq2P7szxpBb5if3
OSb7btoJr1EwOoyTAOZNwAOtV+LhtQJuNuxI+0E5BtP2iELY/rSgzAIJqCG1nXB5blDmntML7L7F
GoSCny8jISGE+QO8xPFEJyw+ONDCcG0RXTbJtV/Zn3mD1yagZesV3Ny/ccDP65VuXk38rV4nEjBd
KD0o98dN59qK6Jyc6r+BVPLDN6zjAuyjPGYy4qsOskh8ybiPdIcOEQH1afMCe4ip4I0m0j9YbCpu
ay9zT4D8MMNIJ9qjKtTNTFrzVlH6qQwIsR4ipAwDEHR66i2FYtAhih0orT58MufubOv+3rvA0erT
DHUjoqDf0sYF3tesZbGy8HHcDH+ha1bDsdliKgSzywvoHRw0RDlY9L6CQ9rPeP+eMvhNRLlq3yBw
0mUp0MZ2bslUCTRO/zEZ9XAehh9A1pMxnTwzYhOxJLPt0oUZbN+LlZlY4iUercJvfI9RyjBpUL0o
p9UFau8zyCt1gcqunHU17MizHjrGyietj5nBiwX5DZEHfYvaHuQ0OAZ3zVbWwqu/NUHWii7O2JuW
Pi2RRSUs/iBmJEmZ3v2bDq7+1iLYjxdJLcS9kuiwKpN2gkQ7AY4MFZpifBCoxcApJRrHbf0mUXt1
yuD2jiBv23LcfSCXAn2v1iheNTryQeA7xg7cKowvfnhtf3IEpUJsQRZCYqJO+DKkspWms9hRVolF
noKeV3unYJJYk269w5vv6ZGQe3h0ExNuGnWbZo4+zyjAVF74QgVtpa/+Ig1gZ+ZLY0VKV8D6j1Ls
p13M7a3bPNs+dHyKhgFpRZ6VjPaXY6c0DMp5/4MpI3iSBESMW3NPoHHglbebIj6VFESEjOD+jqei
ZHOz/2zThHnaeHYml1o2cJaTzCKdxHIsEaSiAVqJiQeZBPYCUngp6Zq0lZ8mcv6z97BWLse7U7Np
Ca8ApD7I6t7ZL+NL0eT3mODwCmaV5kMQtoGlyt4rL/lQP5UNVA3PDEUOwB+zwbMhEfdj7KF8EnyC
vWLPY4D7KMDa22lzib1Kd0xzAHtSbqhgEdscKlrJS6aO80tL+OuwLrIpErxfbveKlk+dthMpM3Fh
ixR/cnvr6m5i8crH6zBFzT2P6wzix/3uQ5McMYzL77HoytsyN9Zl9KZme1dhfGBWoI++uAlgXvFn
Sbf+3W6lI8oGySRtVwFCOzUpHTc/QP47P9MDfPM+MbEl11iK/PFUNGVTJeNRooudIdNRO1n2hc+l
XFvtdgB8xxHGzUs2198euk6LBLtaEK4OKrjUISxi2st9zdwNwYVdSYSz4zTcCvIkTFOnAjv61ZBH
YefuN7emdiGNHn0b7znYHXKOG+Satk9qs6NA9WZrlQ2rATLAyI6X+H0rM8yjaIiTHa2wvoPFPaPE
tWmIWS5XbmblTQ0p9zp0BUyrPKFChYIqof6IVS6jFB6RuRQceXJ4bTkokgFWzKeDOLij/jI+iQeY
Pn9vjpuzzN9mBx//rOzAM9iUa4OEj61rOWd/vt3x2DPEhQokYHm0v8juiclZvBd0E6yorXeMYpnW
SrmrhOxHXjnmBMOh8FXG7FNUFWBj1pZJAqRSiMjIkULdyfKFZSwem8ocbaeSfEIM1QAlzO6Ci2aS
Gg1SaCoXhebeA1uC3F4D1lVssAC9k6JLRIBQK2Odd8ia5ASsjIAOqk5RLzegI4UTO3a/ZSDIvzPJ
09U8OvESYSTrQhjGHVykKV6g5i2kYUphdMGIkcWarmxPJqZmAxWP6v5S6FxSIt8gBM/0X5vlCBkL
fnePUnCid4/BzsONucN45/ZlUj1k5VdgyQUuHYIQm7zZ9PvjfZIC6Oz56/VJaOawICCG0ve6O7K+
CyhS2XEPE2zUzI7xLsGH16ZXe6I6Do8GqiHOqeTG38Y7UUWutv6hzhNZWeFxy8J35EE5+SBD6HlU
xA/TXO05KTjc1BWQHS6rKKqWoQJYKUotxw9Blp2VChEee8ZOUwndc4FsRFC+751hIscNpodHXgXc
B8eQFUk0mTvAduVoFsQzvE9IdSOgtIrK9pSSWTA77lxgTxbpT3W34wYqpddqYbAyQ7XvBCmjX4W5
0TNjFE3CfDYYC3AlMXTSlAe73k1terX9iBmez6j0ApbKnT3BW/yAsFuzsESTc/6pYGB+QBksz+KG
GBr+vkisF4Nx4ty65/3xwWM0NL3UqIsm7pZJFalF51IHeSAXzvApnRGpV86zFBIh56L2Ubiv9Y66
sivi7/6tXQ4ka/nruQwD2BHY2JETlyjXPzUsiX1Xmkxga+EtugIT06foaaGZWQWZR2021aePo+E9
w5BECmuWo68fCOpKhfvBCuqby3gM5gq9cJSgM50dB0W/yWrzSOO9faWEK2evJ3P2jSR5N+xNDcl9
7OilIzF6eF1rQ67buSgNV8jGlSf8nUs1M3pOlChvTz1KnjahYgCkZBf3I8bDYCX84w/CtdVeSID3
kFAKiKOHn1oqCyAYdQhm/GElDJrCIIE9awcv9ovvlnNwNDRiDjyc229c3LAKrCsihNw5dydO5Yju
i/AqKDH1G6aX5nCPoebm16OKRU99YVfyO9lg9yJ9YEIQqQmHwiTacvaVxoX/yDhA33Dp19zxgRvK
CWEno2jyJAWnrEWQ/5xu7qb6X7bOqAyJnZB5NFRTzSWoYUfNa+7hENfWtQrKCDH6GUxSCqvyMuYZ
TRQ4xrXgEwCuoCxKbVFpSjtJCFbJjJCanNsGIZ6f1UZoS/SSPTcVId0G6Fo6LqI1ttkjsFPHoEB1
Cf6VCd0GviBLcsjYk53AiXIIjqdDE//3q/9EYx4y5C2Em+4oydETtQiAIB4BIjWa9donynhI7c/s
da52UKYzyo5ShW/2WXbXCHSwM5Id7U9boW55TnPBAzuRdvt+b1y1/UwAwjwJPof99givIdxNxDIn
qKKjCDECvmcK3g8lwx+p7HpHfHg5702NH7GcAHF4MdVA41o9r2fJ9DYZLs5kPShW4LvmKw7NAmKc
19g9yBhyxGMoqZMGxsE7XxNRzUzUoJlnVPNoyDEqf4qR/8BY+RpAUibviYsDXQGf5atpcjp+hMtt
cYSdBRLy7vx4Zf0idjcEIrsQw7YYZQ+gimVjUAjezehv5Rl9i/SQFbcINuWw/ZzbJH2IwZrPXvJc
gT0/NQkyZurvuIJv5qhbjt1X8mof6z/syfacgBXFoYXrPPA2tRK1E0szSLOyXPIBfktioy7+JmLm
uQm/rr8rLITazN5FDz93m+Xnl0ppMkgQXGYN1OcMPnUdVD4uQxuEr+wiUd7NZBqy1QHIjqZaqi7h
BS/xQQk4qoYdZJGWQ4V2UAVmzzLuniRmpVDMyN8lFXX9aJCfNkWW+6ocFvTsUFeEdGQKJgKu8iFG
Ir0DYCkOdfja1gKMrlQluprIOUBwWdcJDKDD+OwlJlUto0FXp01Bzlxok2qtuaH4FBlRUnWg1RPv
tNwawztCfIS4Nf87rLR/iBzTWC7ZCE0uJyZNPiHOjEu4v87j9mWkVvHnxHnHhOtnsgZduW5N8zfm
p4IYeyBKA32HBRzkmufRn/54BiAfpZB63bvKoZqMg9ni+30pBGTSIBn11eUBGxdhIr4X2Azw+/q1
T3sY78THp6YMizsMlSS42IrKzpwXgkJBWxLiqcCNNQptJiFZJO4exNQyvq+U36fEhkkw1PlfgKsm
/Rp/dRX1qA8Yso8gucDSQA+aiGWjBf/fD6fiT5hBCW+0n2BdGNe7pWTInn7xZsEw4DMagAO1cMJ6
UUWmsQggvinIlPTCMk/hb69RKIH/yyytP5jSF/9M/v+x64w8/08u6ElBlLRbbvvT/ghnOfBLIdoI
p3ftBtQWkohJBVQuJF1yZAF5V00qrk0ttnP+QgFHoKl5ReuyezlNrWY1g+B9sE6hLSC/3ynBJrIw
DBTwn0oC0jrI6ak6wyY2c8hN+zsBehZBIKBBF58agslXGPBtyDoCzwoP44a1F1j5kA7VRSJzr2QJ
lcNj76Ld1dVFJk4Zw54d6fNdVglBn8+aP62zsebr222Bg3gudP9misIxuTd099wPhIpvR3E2CkfU
TubkYjaYLXBKY07CPL8AByOE0nVMlGXTUQHarbvK5svZhMyy06ZOXeV41J9WkQ7MqrhP7qKqJ1ry
i6p6DUaeCRXhAnTYM9utKNEb6OMOGrNn4beV+vqel6kIcqEoR3DTzxOOMQJN2V4KdTfvaKnqS7ZA
R9mhB7+btLShmCqvXCIzzqI+me9DVzpmumRgxDgA14/8Uff2n0YXv9KLOwBa3M/j58iH0pjiPSV6
R3TXpiy62mzBN8f3WV3fktrzzgnq01UAuSZrfIJSR2KqLU33Eaywz99U/AIzMHlRpcqNbKsJ7WLH
cTVM1NrOJQdu2JMMSHx7pJoOrDZIIOhyh+XTMscl/HL1n29a539Wl2xkh3kHfnpT78U5YLBdKaLp
l+oXSHS/oyCMgiI5wz16RKtGWeWdChc2iYjgMj9mLc/WlCXtFK5sSJyOotQNrlfMLdx/BY5riiLC
ZQRh5aYSsMOuA7xsTI32GvhRkjATwbOsl4anVMaKAtw2n9NNycdn6AZ6CRvtuGP8n4if7UvBlE+Q
nGO1HOpRqV8zHchVQFx/FOSjDZgQux7KVBr1woGNfHKDWfzNMZeseLi+SU+gDfBRx+gxCrKLTiPS
DoKJlLVeibuyjnk0m4YCNcGfO44ktKV8bKvMawmKHcOtzejO3MYz3UKU77xbQfmT2i9hgggPbcrp
hbXHZ5ZKPnsxJJXcjOkUxptvmd1lii9uWNJxwlWiOxzFcNrNsWLIDnTf+V5KxBSyEnrvSACFMpLU
qznE4UmO6thKNm8/MVH9luaHHwcTHLhQe6J/Pd0binYwSAZIgqgOUxPX4OIVPHOncy3BMJv+v+Fs
DS2bXq66SlIy7+JClFLiDFVWOpr7idON9oJ/4ORYFX5+5xFrJSM9Ic13Os5gC+45ac9X64QCIFEg
RO2NRS7oSmz4UijmTlPE42tdGq8UGb9euJEMVaBghpnYnFcE97+gSwKDyOetf5f01xz/PZKZN+aP
dfgWXNwCIoky46JRCZtPXfXMgEKjux1qcnBnc34VBuUb3ovxbLHRC3KVYbKM3HyYlaH5DlT9CbbE
F/Ky5yRAAJx7XKgf1tIO9/GRJKZDtV/Sp5FgREm7Fm/rURDKthTURB+vwIeDKdbnGLdwJmM6gHdb
fwsrGHhGWLes6CVWWkihoRdYrB8eKQIXDlwt7lQX3qUI1rVfJJcc+skSXDAZsacbwU0RC4ypDfar
mgAg9ByURDeBzvfa7lhAz5X6efWWyqNi5boRX5IqQHUSApcETLG1OSOEzbs/xzbDRuRibMOaPVnN
VadHRHgTWPT3kX1iIhk4aRsP8poNtNVoSJShrwQUvwd4tfhZTXc/6gB+9EFmB88pkdqO5z16bzMt
Wu9BknzGxeTMWoDt9cr4FzuRv1gX4NoXxhfpXfJsi0QgHrWxa2+RtrmMbOjeddxCSuULFlNBKw8t
1ZNSlROYp4uk57mFoA3KQ0nFOgsPAOlJaBz3F+IrTVySh/kVag3JQkgEQpxZiCq7qk87v4j1mY6L
/hv6exrcSAP8ZyZD9wTdmwocoy58HN7TdGGlMVVbzeEKS1TevpHSW/GyvIWzsQYUjJC4sk14TQ/I
p/YPTq3FQskCT4YqZnGTJSmvX/2qHUW7tdeeuQJghcXofQGZ7IDUqR8FD/Y5K80DEaA1x+th0Lxr
0okgRO7DJJQVXUZWBtjyC4v28o+WTV0HJNMMMWBhh2T48x0TaE4iLiRsY+IgsVpI45YFPUs8CZA4
FigtNbdxdQfEJ9+vTC6T2tjAiUw1UVu6UFho7KWC4qveols60XD/HjewKkXI9QWY00To3+dT1jaJ
qM72L5YyK5csFEBVpc9SGBf8e/77+QwkmwGla2OHzShdFyCq0BtWFE6Hr3BtjnQCIDUfjCfkUHut
e1FhU4Jwz3QVBCPSlMgoxdzv9rcR9o+FretSEqxg6AKWlAKXb45/Hd69khVfYcf1wpeGi0H4tteJ
auzF6ud7rRanxNHbPZ8xI4ZpUKBJMIGT3KBa/nv95OHh2yWGJHY+l56+H+s1A0LXFiOS/B1uomL+
6SYUUYsfmsPeluAwfrXjyYaoOidAjCE/DaRq2wsj/2X+1lQONouWQ7PG0vaNdNjp5OhXitSAxc8f
sDSXLZWbBjz3Pps2yTbsqCKCY4V5+jpaNPiRZLbgTI7+BycQFSjqgQgzUGrdMj4HpA2YXjrNOA8z
n8JaxpuKs/DWYBe0g7ij6HIpIkMpPe+A3NdObjGF/uZcUeF8ya9wrNHV5eqxAW8qFibRTwradXcq
0Ds6jSa1kEdWkgbfQhtuE+oqvoa+6wmWPqwq3lIrork7n+b4npeg7iOTcrT89Imx21wvYTQyRzDE
R9jXrlj24EuiEROu1xBCf32Wj+eR7LNFhN4/iowmspI/gQFsuthsF+7qodjmDb1tlOHq6PJUYRdg
Emg2Gy2Ilvh0mh7vd9GFdnPdExMvwoxRxpwOWgUYFuJ54vQvsiff/SXqrlZBScqqcC3Pw9Ls8I6U
+gQPqwb8UqGpIlGSPzQ2FHidPlE9uTRpW1nx/O8O1HVirZypcYZgMwxoZfOt6nFblAIzK1p0ocTU
NTKZiULOWpsrOsoBOZSPk6vzK9isJjjAe/zIiLpHmY6KZ6F1Dw5cO8GbswbF2MOjfnGFalNqzGca
VdCt8R99UBqCyPkqymcrOhMb5jU+yAAJJkuCdklodde+XfyOSCYNi1Vwl7MSyprY1n5Ed2P7lXHF
rv5HgCRxofcItmVcH5/uwSDYzaBVp9F+1C0S82kivL9XK1CkZH5ZicJXpPB7Np4yK5Obl0L8RbAw
etpVijxWY3QF/XPhdheYhue3MGeiviUjbw9MzmEpBI9E/+TISIpdC3gIJtCHlcCXXbsDRzsFMjAS
eHX40pDxXEo4ZA2W2X9maLyAmi15j1g7ZkBllM6kMfZDEsg9lDtFP1TMByomj9pZ3wws8nMePBT+
p/iuLRNX4Gscz3IuRygRlMGr34j5ea9LOIVVI4+DxVK71cbBv1En8cZNKPkj9U4Fdv+SezJAgwUu
JlqXu1e9iQ1brsb87Q30DStbG6UcfkZUe8zv4ECyN5lQELgXUOqvmUhdtFrEB/GHUtk5dh1oJZEn
Qt6/5aDuqIpAsdaXIyWAEzdrBxdfwofqPx2j0qIZZQCAGl+YSfDct6cQNp6+9Z92F3aSxQ7me/la
4Wiqpy1j0Va5EaUavjjUxM4UR7hmISyUTN9FYHRTGJACy+VoDv/XV2Q7HA1C7xjEOs4nqP1g6up0
RtXXBQoQHxMydRMawITsPK9AKj9L4q3KfbHLSbZeZowjd6VLDLJ6/zwAukZdZj/cupX0DgI3xziE
2wDbQDYSYTD6gQN4DnYD5pi/on6l+gWFl5IolDST+ULX5OUiZgDJJ4oM3vPsA1Q3qW3Qnk1WlkFO
rqT8yRtEId8+t3hPx94ywWa/aU2xJS93kd10m9pFTQoK9dhb95qlEw7f8FlhO9mDllpl+GI1gHbd
1PRxhzAHiVne++cEI/+7wBIBSOcnqlJXde52G7oVepMlmiwZpgLsrhmUFcSdSEaUQ4pUC/UQZdXn
69dimg7Wpx6SYiR4aohHB0AK9eW5bvMc5mgGR7eILszWOqFXxcKeZYEStO/YhZy8kD39Pg/mO9GD
Db/1CEB+pV/f706bnzvgLCzhA1aRlektslTxqjJLYBIZkQ+UFJYysYPKdP7LcHOi8aRY+xOTFPN1
BsIdRz/xDChZzUgY4Kas0oRUABiRNjKQogbt9ht+5E4U3YLITgusM33u1ECiQhnqf8xm6iqeD+th
ktldrxUx3YefEr79/l+BPsiTsMrcqvyoolwCmvIHufcxRyot4LMtT+Uj2Ck2XOwSQwfMB/aNTm4e
SZYsVjLtFT0ILC92eI+SeDYBsrqc2d6n9FiYTt1DxNOQixN28QhLDWBATbVCWc8K5DBn/sTDSiIc
pTfCFRNyBYqm5TjmJMT4uVRJkrfDyBvoHOIYQvEqphYBqsPlnptk+KoJORwIrEaFgCHBvAA+Ol7V
VIS3mL0gCrBwR0p6j2EC8XBihWBklPB3aBZ68kjf9rVVuqFuPig0Z/yGbNrzPi7xRAsNEIRYgCrw
sKuoLkmTjlLDZH3RZL1DtZmkXZZRP/kUaRGUnga6go9I0ioKnWewRZVlGPgWEXoX1xWpO++Kav50
mk0BFdKCyD9FmHmeLGcCap63iSD335ATks3UKGfbHUWElqkDFjozf65s60YuQ5b1QtxcfaQ50Bdc
ow1qqN79MjqICjkt53JX7OjSVMj8u262VfhaBpRKUkKVXWvGL/C9EFWw1BmP99G/8ISz5e0Gvkei
5Hp6FaseTtS/gau69+LmwTtoENKhhSTMJ1j9wqd71yYiKHvLlDwcZTInyQtq4PJwVYB4AAJgpfui
zKQZIclWTRJYtu6MAdsO3eC5r0JyoKptuexlGVpQDfJ9WeBtRSvdLveMxQqM1LiHQeov9V+JGnBh
uC1OZaH054nzLT1saN65S0RUfbwE1zs+rknINr4aRk09RAv48/5BHsGf5SVfWDgjoucL1BQQ39q2
qPfvjsArdTWr1w17quBUyoM3GIw+oNxtqWlQZMbCF7/SikTEr7nkKeXVQn5XTba2FCx00FSKJ3Be
lb56i32cC9WN0yZNd46d3K1ASUk12s/X+heiwa+o3T3WbdpXxTeMGLu7g0yWduUfBTDqqTMA/iiJ
lsOgj0T5Q9rDoKj/Tn+wSnZyHtdQIJxCVjA1YmHl/lKC0xwSCtazygTjit+WjzPFbkC1o4flONqC
arpF/W62q9ZXGTnPKjvbZVm7CA5ru3JvQvot6Tn90erUEKdpwFEOZK+Dq1EcI9kU0mNJaLNaJssi
dEW5utYpIAdMDFSLhqtJhWPPEOq797mYH6+eiii1vHvtBEKN6VDA6v9NCImme5xsuikYwnJfAjl7
0oBdFX0D85frSEX3v0pzgQV19O8xcYhVNfDMx8rezOq+1FPPjPeSiab5Ty0w7b6WoOC/0yYjSsMo
cchwdMvU0qH+oQTVtavc5YjdaiPBM0Vvk/M1C+uUtdY8qz0G913Pp9iXI8RoRaJYOXbAUboQrKaF
nsan6fU0acp4uP4VgfcVlsq5fw5FIL531lF5Vso/X2f6Qg6sEwbG8ynieOJJKKqiXTdZ/N/tcwxa
mMmMI4iuiCSq7OatEMlzKXD18uh/XT1l/FIXi2NiLqtdNb70+yZiuo4OFJc/2kImckbGG8MrBO8u
GmzFUboY7VMgSKON11zzW0l/TK0PxqQ0tesqyoqzoHmNIUnWHwfEie861GyktelrXgUw59X8w8vQ
FVtPUmqzgNc20H849eHHBcgXZHz3JJ12tuUvB9LGJZRlabs1RHr6ilV8VSwMMcDjchoISiHuhQ6S
/6uQILmmzrc9s4f5KTyYf0LEY6rtLWsHj5hR1yoCRUz09pGkqSGlqsI2ddxIpeHC0p5hrBs9JpAk
SiSxxEBW9N0fDkReqg+dcml0JQS/apSQwoc/uwcZRCdG+/ii3pajxa4WGLeEVyJPQPNTBQFhD1Ln
FRAqZ4dcPImtPnR8AuBzYdeVHzxNzbdmGHMD/bSQgMWbPQWt27HnFgW6OerJCwmSUOBavdfK8vCs
80MKyEsZDvWhJplzL3ikfhqdkI06oDjpt/nRvKciuXzCoyffiU9kwzLqToqaYghJWb2AoWSHNt/H
HAOGTIk4IGwnAvbwixLI5KUhL6QnvJ50INDZWJL8Mnhegzee1HwqBwrGNTpOC/D9SAIcw0mG+plM
8+SPI5AFUujmzP3ZRRbllqXYNrFWZef95vydUzAdAkaWS3N3GrdxVOx4NFFE18Dnlk/9j3kkKy6B
QNTWMhTQr+ZZdZUtM3F9pQkfRfkUoUJimVFgj6ZjLxafBFGuwWLp1Lk/Rfq5E3tioMZ2DKq99uVS
Nn71dgPCghyXHkJ1uWKq3Qp+njrsuIDejqlTsWQAuTZXwFsuKKHkUYs9ui9Es1I2CGX04euEy9Em
GjJ7DrjF6pyqhwOGd692EAKJG2VUzk8Dzesxp/JLNhPRzzQfj5+MndmujFGXKH1dyZBpUgTkfcXr
KSO2W0r8ksQuR2kzgqeuStrvduJir8fBtacQK19YVTJMQMqLEoHrusT7nt8HTvqxg0GLDnh/syfZ
5+cLwqBut6vugfvxdGreWnhBHSO6OO/93R9xS4CEMT3SzwWMeAsm0ACN02B098MHzsa929DCZ9fR
ua2xYmgqrFdyFbEGjbQlv42h/I1giDrWfiKlrXlHPnfFe2shl5FdTmCUHwGPazfBT6qoankch9w+
UhfJbjXnuOyiaH5T655p2oqcQha3NIEAIypfuZy4/rXW3ES7RZbes3mAiwNLM7crm4iZW7lw75VF
Voqw1PJTgzsaN53zZ31y34kTYc2MdKl11twCKSreR2uGTOrmeDLkqbirwh5Bqd79fHc0LwWhZaEz
IWdJChuoSiTvmVn60Xbp2ZtdKxGhzBVrnKM2m06SPaQ8cMvPbIJzyabgr9nW8D/qzWmuJZV35Ouh
yjpNGsktMyuSekxZDFZF9Zg2V7oJDOzlMopVyRZT0TDGGnYCMMhlTEhxX30sckn6qzhCpJVl2Zfb
buY+x/rIhQ0WdcxjxaclZIUpmY0zF7JfvE+XfyCCkPlVv/LbJnHPq89n7grLGqVAem8n2jLfFy1N
fe554T3dhTcfuBFh3A0YVaf6ukryd8I5eMP1EDMBuLi2NxNoLWdAfIgs9QB9qhnyNBxMMbF8dtbx
fHqJU3XBLgnckE+p1dBDLGtUPpRzGcQlycg/Cfc0yEJeJHYtooD5vfdtJvZ2t5GUSUUdb6+gE84S
07hLtNaeD5tv1yzIm0fkMk0B65v4zT70IWzBrkEAEt1b+3SF+VkCAmzjEsWI0oD/SB0dXDB3I+QP
Jy/hl2LUb0nY23Ygcgo+JF/GyaPIIoKGs2LU+y6a19Qfyc7MI/OnMZwhY2b8uyWDfuJnlxFzIGuc
NVWME/5sQI23v9q/5loJSrLNxRkDG/QdFnPBjIL7qOSPv6pFfQLkCLXDEoHkQvuXYYteQT+3QOUJ
ekRirdMPS627oOBFSSLE9z0yx9ahVk790Q0+UM0DfTVQu137NzARgW+j/DQTatlTNLeHChdbSK/9
MO6Mvh044YR6RSiJ3clwn5wTaphgy+N40JGnc4t3MvckSufbd3KxA1hYTNORMqKyWdK+vdeXV2Qv
y0/nyh2oCuIfEJWLTiYw/GRA81JfJEL55t1Kmft5aWq/8nIr8gpievVaWE0AHTUrTi4+O3OPnwnf
joEOwCdaLjLYJsYJGmLviiABoOEuCHg7ObF6SPRSTfd8Q1Pau4guSWFWkZhOvL0sX6GfjHolOQlM
4vB88QX0dLjF50xF+jWUVvI0dyirvt+IwsB8SORTAt/crPD9D8Zae4wCigQtYmtKUEI/oVw8/kGT
6/Zh/gMPVDHCNcRkOgkmmkFpIz76vbrcwPExU47B8fuFk8aEDTM0yrYwyoZIiQGr74H2FZ3YQAT5
yZTBZWmKdwTYk4PaSy9Ei1F2rYBi+sVhheJ70KMwdoqqQow7g3npS/83Mql57VLk3YNjBD4jjGZK
BiSFvGhWH3nN2AO+w/MTn3owRcqA0Z5uC6MTgMXF5zZYui9xocIFb7id68KVPYPHizDUQNKqdWuV
REXA91Z0JIKVLW8L3AemV9oxTv0R4f+JXEKkRQ7tHQdQ3rMAsl2kvx75sjri4SPJUlZhpBS8AonI
h27HQ72NCydcZ/dXIGwnRyYguvZOQrGdj97JbpY2SkgqlsjysUomOJx3MwIuzO/TDDlYbZ2n+bPD
jfw3j9m04v6au1hiaXiU1+ob6ctbhe9pJtJq0FWovrjJ0rEQwREXk5B4olnCaR3UXzZgdXf8WP2j
2PZd2zJTOCVXj/XSRkQQtT6Dq7O84c8zV2yzrabYfAbd6FrYUF4a5VvsBcgNyo5FuwVDmN1GYQ14
S1kK2LuYP3gMt5ZEpoyPhtxnpS60i6/zSGKLRXC364hgZRL77y7NQGmMhoIZozFvHuhQmEpEgfc6
+EOAXNK1mqVbW/A67jH52+Xx5m8fN4MNEWDa5yfbgxqwrliDO5gHjrRmQnV/yOs+Pkjh9j3KRpxI
W2id5go2BqmyIuYGO59IX1EjAuSf1twF7cH4u0LHjetcTVfN6ZTIwow8UQIGEX6AGrQMNVfXROqd
zG9SmRv/YX1rkvlN25gsH9UysRGaUMxw16ue4RShR4vLd3FQIMC0hOXsT18rRqV12I6fVBoBpSta
xFqxMMkuAkvroBWKWw3BcWgbylW8pSog9+Pow9CfNBJyl1A0Sm19ZdJVdDN9eZmpVbpZ1Q90EFiG
jJNy2mNsjqaRVnaaPtnBtFRVSABjgC1itRecu3r46P94cdSHEf3FonSXrVEkGX7C5sqSJjPXBaJW
4mEFf7SUpx1wVQWyKyzhmMOROMP3AyZ3QYl6UIppvQ82HMPJRYpZzUiF79UIfg7BSfBlY4p6kpjr
l/+sKEVz+2U3FamyfVNFedQKP2xX5luK7RNOrE+V6I4+yPRx/gMAPUYc/GRHk1ZG/zIpdlPlW7vH
R6keWQbtlOc011F3ir8JC6TAumvMB3AtZL6HtfTIcW4mMAivrG6MD6YXQQiVGCa8wKp3xQIOaljk
c2jDw7whlI0wh7TsBneMxWkAxo6lplyYMGwH1iYH765K+XkF1XlJv54I5MGJBICM9OuzoqQZ2jvz
uRhXV4zo5bX1kTNvWHU0fmYvMAqBwo92JWyazTw2YdsbKgzvyCtV7a3obGXn2og9GjaoxJlDQZFa
uoQTGFapD/L3IkKqRJsWC75p8T4pLpCxhaLuxIYthEh/Lo9/VCWzbRuFJJWHWnryqnwU75dsy/wn
5GGm82dQ3ICxo23vEyt7XPupQwdwI5woUX5U44JuKtbMXuds7Yi0HOVYXu+407ncihveVaGy4462
HRqPt6qlcYKfMpw4QmRJGVX3wNA6kBZIzrt3tL6tVKATCB96uRtvqsh3xTuurwCWTB79uKUf7tyo
x1mY5D2AsqzujSOj1M8BIZYEPEGOn2R4Dqhf5R4WWmiYKTz08bRcdA5wB7ZrLkIv7bpI4kYGH8Uz
FyQ1zlxBhkRlY/rYlNB3q3SUd1CgXhyQIJCQr3GPEVn00pTt3lhtv96DIbirEn/VFksHU5Ed5GFB
ar3dfiehN9ekDQaSseZC5qrd1qRxf0fzyohN+vliq8EeiQppxU6taHjEeNVy7KKWt2hTYFglRLNh
tft+lcgoi/69LJQ0qVE7bR5NeIxq0J4ZAgBHr2LhVXxtZcOaYDq/977y1QcSwBGjFK+RvfvkoqEM
my+XJyyrFjsFhaKPUvRZu/A0Ie6jDQxFzuj7Wp9k1IcM1ie1wtysohJW0LZIJ+CX20r4ByNTZLhP
abcg6uAKwgpiRy4hhjD3mmQez2eRBaaq/jJz7Cq/WyT9oDhdl5DBGMOu6+T7l7ZzudR/nQNYkEeE
Bhoxc0Zg0d2HW7GYnFOJvxyovi/ZE9mg1nkME9O6hH2ybCKeoik/epJ7Z5cjdlI24rW+xc+yn9Qz
Fx2qzyzxiakbTa+6ArEonmIHm9qTLXfpmnF9Al7StMeDKKPwfyw/cYw4CtzdAPd8ce2+RRfkd5hy
xvcNvtpvVuNHWL86pgLElRxLMmxWhs0JK06S8jgVbb1LzZqwXg8flAh4hPN6yfd9JxMByfvMK4yT
DF46WzaDJrrUGM4TqyNh8CznttRkRHuRcFZqyZ40UKZixOgmbP6bSuKQYRo6YW8hep+69rWwMoAz
UrJaZw8dgDtVk/8ln4VkF6QidP8FcIJ9YLRry7BYYPHGyVaBrM9YVFkfI4uBsLSkUfuzDh0y9pZN
oYWpEKIP46RHYa/loDZT0M6Go9D85DrwAyC6jDFUeXGcho0VNkbWorBOOtujZvMuNi8uCUJa6Fxw
wmb5kofCv4mBlqTAjppe5E3a83jTVAZCxCwXrND+d8IDv01hzMBqt72+NpMd8m2ajTcqet/IKpfK
+VnwDxM661GI/1MuYicHIqX/18yJotoh5qftOrbZyqxwyRelxq+23hiqK4Yc9bidvf8Q6P+EuMDO
F4zGgWE12eRSSqif84C2/D5y647VoCIoNKsKAh1a0M4MtOpXRIGkwkWVtQRpwfllPn54jr9RVufN
URvYseuPS+aazf0D5vRN9qhaCFdnHHaLkol07DjbDr7ySdelmP0cWOf66dcaCSn6nKzFXIYGKtV1
+kGRbWROsxVIywvDLQ9+Be6ieqTA6Uq9imb/DQD1rEuRNNanydRzJt4hMKuaPqUMKr/ECzUuqHri
O3SfifkdisR9ax0vMKyz6Od03DewjAVUKljMwTXb0XmlXu9N6YBjvDHrwfeN2iOuJkuSVswuRbtM
/4KsQSvJYMb2xCmfuDgogL5e0WZ5BxWp9s45HvCXoPy61OV+Zoz5wfrqwiwFUfp4MKquJXI3yB45
szTXLhEWZAKenrNyv0aJfEEg/AetPampggfcmmHcLp5cmwEOvDpbHHMkhxxGYgNuxU/kWG9OJ+oZ
ww8AHKQV0I+Ki+6nCxhJ+th14l4EuJU0EbGC5gE4UBzIc+pPHh4vOQYGtJHhiHvJXXAi5ZuX04bK
ON05j1TW02s1u3MnlPX9VRmeMU0sP9V7dilruXQIhTm1kh5mb90adLyh/T54WzQz1fyGj5Vf7sl1
AcxjuVJgzpVrkKbrEywI5rvvpSAHaUmvB5awkotojCsIN5ty6j/H9NWWuwUmgtycsBPRdKKVZXbc
bZsJGw6I2rbhSDptkzLD0A69hEiNmMW28ZRpR4doGDN7szaBeJqxgTvemGPW/MjfFveE0hGQ+RM4
/IGKbljN70Cg8GZfKuuUgxmb90gbrXgxv0k5IDsiEcrzrihuVb2iIjGzjgjerQ+GSD5bjeDJqF8P
ZxJzGLPwVkyQfGE+YiYx3vNNkpqk4qUmBxnNSYBMq7lWSKY3kMrQS3+ayMOb/Eu81K6z8jVygfGM
xagxEis6xHyfljyki3vJwSCiAJEGIlMJZS2sYnHhb2Zl0L4E2y8uSUywYCtzJ+rkgEH7yNUt664g
RWE3T6XbVo3+I2VeeXrr9C/2wlhSEzynEjrELhAvEH10sw4gvkySx/pGo5NojtYfBptIGQCQXMqg
XGcDbuSilkig9YChJFeetI2j9+cKOU+Qe4lIRgNOLDGoh7uBwJ6VeoChgy+msAnKSWC8cvnGGzKp
9zbz8yf2Ij96UbJR6cLwe8GyESt0bz9+QxXcxv1eoP1S28tXJCTBkaNA7RDGjzVUkbD7cFnuY8bl
Qj8b2kBftGZim4C9zvHfkvUXMfdCswwkfyi7uzKbMmXZXnSEyUk5/9L8PnLUNTFw+nvgdkAarb7e
Glb7YdRGkwiLez3aKYnMOB6apZRAQOxspAYtDnbf1MtR29BaGTQFytoF8FmHqOm+lRCOeYO5sGtG
Mx/obAZEP9s+0K0NYfIlKyZ+e3mPEy6rgpNeUGYnjueVBYaJASr7NqAdm3xbOMZVFnr+WqJc56kB
wVqA1Jx1IJjCxPAdLAbNvWpkZvo33gfxB5rZEgY6ELuyET7hNK4QSEvkKp8j9fHQZrmkh56ST+jW
M1PmCFfNaq2gFrN2O9mOoeCd1huDoY40EtlQyQcY/E+/KR67F+i8kxWb55E8ajBWffciOgzVuo9U
95ExpaSUrHpptCTaKOad7eM5SlUpamvlvNlPojKBW6lnswge0M7RYqPBvCMlyaFaj9lQS6vNy8Yo
h2ijDit954ZzHgW92GbX1tqnpebT4Wa9NRqdxPkeqGjsfuq1NiNUzRU24nX9EPJrRCFEJbDZm8YL
HdeB+f6ba+fAY1OuXVcGt18sUVSqi+8s9rXwQMB6JGtA3KLALP6zf3tsEkuuic47mrkRRc/zeHmT
48hpOPHtdGyZWihnm6hZD7W7j7r5KHq0y9ZNOv3eFD7CIGWrljEbv1COhGH+4s7Ix3pWLyxI31f2
sIAcJe5mPKwRf66EtA4aDVs/ZEZbzOOpPSYfXn7rq23lVJ2i/bztVxaDpc3Rw0VVuBWc/fdo3fM2
uNnpUqW5AoiSQWDaBYUwjwp/GiGTspu8IohSTguGr3tkY9QUsbdu28jtVmWTSL6l43D6TXQhqUIb
/EXHGHHusTB67ABaj/zf+547146wpreR7WU7ZR3n3hrZcEHqV0aotrnM6TMmlMVrTcaflUtkH97g
NGKPqjJnR2Phj0VfqXlL1pMwDUS2ogYKcaDdmPRyfq3hNlxhbp0sfItZ+7pmL6X+cuG/J9UHxX4I
oaZrDzKmotrYyOaP0iG2+1orUMKWx1yI0ZVIlVXG+jKSrNiKgA19ZGk6r35jC4yX0pNv2tpbsORc
UMdFMRLcfC1Mj3X3/GaWkMk/DSMca/hEyOabq2Z0xCBiUxpxtH5Nrr+kng2Uyvnk/QHl8l9wHkCY
x/sCiOd+oZ10Nz5dCbX+6UsVbUqNX2YcDpV6VgURuPcLAX5pNM99i5Yh+zuTchanJ75r2lFtvw6V
ujdq9S+ZkOLj6OJE2csn7BhvE2I+42dtmxUPIIkH/0E0X30Fp1CrvvUZLAUyRLsTuvv9GALPY8nU
xzTkFVZHnc2ZQmyXbPBFzMWAAVWiiIeM4XwSFLcm4xE0Hlap7wR3wSuzZt9C2EIQrtqlCfVvBYeT
KjozOtL8Ukd4L6x+qEjLfRP1WaUN/7x3fJwmDOa7tC+6BeLL4DYL68VajMEo5cBxSTWxZ1qgNa52
L6GMxM+a06mNgPFFqfV4PmPsf6OYne8OJUkXP0CKzL3LYgI6TLyY9/2HvJh/j2p3ISwhbHrEd3Ci
nN3KDUOr2NZtKskOta4gPeWoFd+GbYCe5jM4nxToe4bzm/fzmVF+8XZ5vQi7jKnk5/wNwu8uvGN+
Kl2wJKdw8rIz+ooWIO2zA4RwTIBbIL5U2yuVfgm/jpT3DIDXnE6/lqy0KWYeRQ7oaPgGan/EOnCR
I36pUfwVBoSL4wIIZLgAXO2wNM5bVsw2q3XKmHvtIQqAFTFo0z0EEt7DVCAGXTAiq62oZEOZwPAy
oyfGUiScu6zj5Riu0+e6Djdko2R7pKSJdZYMYiRIfUZvEJw+1OdJ9wolTcnqvby1R3P/i1kZBO16
TbHPAuZcM+tVyGE1nICS5kF7/AcqMD66g0oeN1+fK+G57Q4tnx/dh9f13ShN3yVJnQxDicJVXyLl
wKAF5Lf8zRXvOl2lAnTLM7fAl5q3lll8qiFS21yMjo+2r7p/JUIpzxuoqXXRr7ycrPfZ9memIMAg
5Ce+WAcou8FgXUI+Lh4uahb7e21vzykk7SCgFZK0Au5cR9VjtXj4y9IbB+56NEZ2oAjJshfhJUJf
zBfVnkm2j7HfhAhUAXOAjalYzrb7R3591box3aKKMMMMZeyiufuO8ng0SO/rKVftkvrltScxqkO7
mGZka/WERZNxNJ+BBK1FkyAYuR7GjbT548YVma6P+yIGyHFl2pYULyx/ivZkmDdL8uSGuA+RXrq/
TIX54pvwAPUm05VYrff4Dt6AfZi9v+pvYm5YvuvWA//Vh7XSwJTXqSIhecfum4okpm5aHIeWjWVH
gsquK/R9K7HL0kzqWo7TbTZ3oBYXWf/Yc7+qK+6oSfHpeMdGwct2+kHV2iLt/mEfuizX/9Tdko3B
r36atxENBYEdJk94h2FGfP55UJ66wEU4dMuZWXcJK9XCrfXPGKuMIDDQMcnXFHDb0eE0EOMXLEHb
QrZgUB5NVk8rTS6RidfA6xvStgK2UulcYwKfFX0IynHdHs+aEcnRS2cAoF5MrtlwPD3m22rJcm9x
M3NwQuMm12fegNSP3FTBUIcyz4JiK+tkxXwTZB28kA7uYZQ2IRYhDDFN7+I7toNOCRpH7ddphJMw
oeC8BbSJB9FJ20YWw+z2Uq1FOZWapc/i/EpAsWbJM0cMitCv/HGxVeFeroLvh5BKyyeEKUg/HeKA
kIwedzVAtPkEBDCpFRJXkQJSjg445uEHbiI9IuGy7NYd6iv/CvoN2kUk9ymWK+9wgbkaj+vUVjCl
Gyl1b/UZNgyCqeaWl3fOUiE6MJ45hpjN+Zn9WepETnJEAhq86Z0h/Z26BwQnHKHGkUHp8enHiriZ
UVBUpsvEs1KLCx1T/2CQFMNWjx1v+ilTglXUSeHhfEuJlQwwjQhvVSy+lEtd8cRS9xGWRWzrc7fZ
hmyYOOQksXi2Q71IhQee8Eui4dkROSRtznl5wLn1rodpURj+qH8HzbA6rnYKcnjNEYBv5LD+Cl9g
VlDePaN35UFQSU1AQa5yR4Vs4biwLSL4ALGPEE4jy4AtIbO/dJRQ4UmKsT67D8LB/wNx8RYSZlvL
N0isNukfXYE4je6Xs56VKZ8L6cd1B0GJh0st4dxeK2NCwrAT91VeOwTcHh44oljeD/VHjE3wcT8B
EQf8SJFr6IJS7GqLGltUJ+MVhx/Igsjp1RoQc8k4Xh8miuW2ClzNTqTguBAgMZLnYU3aDchS7kzY
RVme17JPBwGHqpFpiPTiUrO/B+XvS4AMts/+yKZYSydivjV9vFD8SqGoCUzEygTIH1WXtnzpy8BN
dMEprwAb+qEivNv6Q0DhQOHdx/4WBhBpDJLBlCj5kwNzQknOuTQ6iD8ibXf7aOc1ZMbWbQyT+GcY
cLFhnIiPmrpmYvwkaU6nEhANZcUllRO4RTv6ZPYe7lTeCYcBSR/dPAJDsnhqiWx8c0en1RFQTi5L
8WVLE90Bw94frK21wHfCm0TK1Ohe6JRSxE5Q4cfCrEeqegfErY2GcCAszgWfIw5ZFW9SdVZsrswW
rJhM+zf4GoL26nnPRf/rgh8WhVUyc7nkrrdWKKhtA6maZgoH5ZZxGXKQWgjV0JMwBMoI20kidAte
KXtii8Z1RGZWiabOCM4NdebBaWYb/MVmWWcXSxrh/vTHgYMtYnLhQyxi6At9AcYAchdJPllyvPd3
qpUXPMfO2VFnbi2Oi0bOK7pCQgcTorFRMIKw6qKCI2Zk5x0FTNIGDMh8Wrk20JvJYMZ2II2C6Ylq
fVg3ER9QfzwCz5ADDc0LSkm8YuQcHjeytGPqS8lzwk013M0TvuveEd/Zu12CKd7xJPzHIV4mT8Yt
NWllnngkGOwo6eir2d4KT1TeNXMCo0PcoHC50vIYoA6B0J4fhoA8NevP5X2e9ctduuQdzMRwohh/
+7sv73p2QlfZ2hUGshkgXsktUtqhBWv03/pX5A1RimxpcjRQUhSOpct9bMSO4uDe3KUKAcDqSlQZ
5fDEz9+oeLTXALC3k4BP6FzuGCB1KWY1Qu+8MKE7gyFFhv46j2z9kTV2XUhivB2LP/TUUddMn8yx
X1yEszTRLeEU9xCN2J4DKvRZFF8BAtra5rrXkR83wX6TSZeYZYg71LNkyqPO+cdjdDk0Wme8RBka
9M1e9H1nTVoaUY24yQRIMXngCU2G/TB+wrtxk9pBfEPAyuhopv52B0+hggqwX0v1TpgYlUxgwO8M
M47ooG9tMKgupcgLvg2RDaXmqpKzgthiK7qaM3gDKxs26P+6TYLhYXIpSw5XIDgS428u/yu+uDNs
gewaJ2ftc0nxrHOjiaRcGg8MTkmytVkTDkxgu24yxHUidN2/cR3KoOU9br5ZSDMeYLF8ZXRnWF83
aDsq+HxdjvdUSmBvI4fp85enU8J3pzHBBFPHg8Vf8FrxkrLl3Eh4cMzShvBtyD0Yxv1hkfyZMAO9
oVLm6ZX92bD59JxoecaaWqKJzDcnhwtzXtHj3da7+SMlSLIDSuJYzdzYGVl7dcF+pcFhVSFN+8cX
nRhdXHwnkareXgbzL70dkLTlhvY9jUmwO5RwknJjKWR8RF0/CFy/r62acum2AzV/6uLcIJYXfH34
zTfIS8HJy2j7bkqWhCvX/lP6aEEecagYSZC8qFe7HtfpLetO12oVvaORhvZk/H0c5Hc3gOYv4KFm
8Sxgc4QOgiVUmjxFK8JxX70GFqvTMIp2DfO5+pFxYSPbRRdrdk4caPFkK/cl1pzWdvi0QqR2N2gd
pJ2Vbr9a+514b+1FUKwTmfT2lX4fKaER/xs074+pV9tj+LnwIQ2hvDYnJEkOWoJVZknFj8Mi60X7
Rdk+73pPZtxTOn9l4byrNon0BP+GMSRy07bakE9hnzrVRdQeBrCVfWL+ZwrEwa7enROB5QVPsN0O
gyXfGvDOc5pEVNt0TEnnZj1mAdiML+Gs1gEtIaQnB8/tW5sSMot+uQiAX+0Rc65cNpwWtFqw6zLS
4w3RVndUsz57hGNxYQmtcilzIzCMNbdQ8xv8Fvyaz5k1r9mam8h3u8p37NdunqrxtITcFY9rG1Iz
PFU+JETcVec8LMZFKdPoKRPU09tSAkgZpId/1hTrQyEhhoxZpclh6r9HUOS8M1nkviTPMStIGZu7
llRtl9DVrLcgxuwCLFELJUSKYlv39jmxM+DFLLpQ4CGj5SiHqItO1PG15kzZW5t/rBTDeKZdyB8O
2XhOqQnCyONomxQcxXwijSSLQMr4F2zh6DguuB6pLiC7E4Cc/Tu2FKde3Y5+rxAyrvqkbAZlSRQw
IG2f6sS2mZdXRBNr1ovMrkU7HlKiTDV41hsCqoAIPib6A7j1nz6CsBBE/ABLbzlYK/gwiRDlDopn
fqJdF55XqQzc2he1wVWWt1/1THbCm+wD1o0KpjaOO1DJk+9w8+35taDej97kcL+OIXlkbt32wCxa
JsCWuLbmW7vJ/vAV6vwKsJvv5hdjS1pyXC0zNRjYnQwzhTL2Apn4mEmmNY6HQ0YdaWXRwzgqiKUo
+ugd6fsVLxTseyCW9/mgsmKM2JLp3Ns6pnflzU4BEA0raptzZS9YzEGH19WXwmH/bXQF14u3sIO7
qSLDz2zyknkMyP/hXjA/mmlJ0kSUkdgvCumgTpDePRG75lvhbiMnoQftpJugAeFDuMuC4pf61JdJ
p02B5Re7lAVvUpf33p68uc0FX1+lUL9d0+6XOO0l+9axXkoskUjUgBzvKyDMTEcXnty66AMrJWbO
NsZkTkCsuiT3h5DKaiSA0lSRW15UtgVz8y7ZKqQdyqupEYvGydToShPI5k6ciXJS58u6gIhlOC2n
4zlJ1u4FAU2Xi7hdKB5GO4cQP/5mVd/dAWtGjO3IclgOaIhJNYjBICLCbo6tYk+8b/uAXBNPgdQZ
BvsnEkoy6RpsLOsNbzStZc0LQxyOsspdgw1N68xTRu3YJshxCfUgBUtIVfsqQ0MVwcABTTNSv47a
8aeD22nJgl9Te3q/Yb+bvJYRMPhJZn8qpJmG8QNNMlugVpDk5hPR7WGVQQKWDDtvzW86p226pKYx
xIO7XoIqynOY1TIw+YnWw5tu08WC+hpCOrVFtUaUdYpUxMTlXH17N07xuyFNb+MHzdnObJqYBeZS
iquoOyypqg5fQC2wmhcNa/50sKjchByFneJjQ8VUAtIW+0xL+n+bvRpJt4RTJe0Z/QEH+Suo9QZ+
EwVxXPxuXKKu9ZXCIKhmCyhMeIoACnjzVxO3hsWKV0/sdMi69YE1DTSJUEtrJFdE1yuYhwlFg74W
+KBTtDqVciWmehbx6lto5ptvh1qSw8SCMueeSIsRIwJt4Ifjhbt1+XYI2oSvbKq+Gt5y1Jzc/CK3
pIAjr2pamHvdaIjsuEFM8tPJirEZZVeDrTAdZpGHapBzmjtGmF6SGkzZy5hR8uY6cQw0ZfSLyqBj
IljQH5lFGVX5mb2jlhytfRqDshohdsAwtEAgg1sP3G2LjDkyQE056S0u6nU/vQTdQti2K9mA7I4p
+EIl1fq4kXAgcoi0hcuOPews52VtchfUJ2Lhnx1x5DLRAI45WbQy9WN6VhAZ4oz9ibySSkjIt+8F
5ypOXrHOjWl4ifC+sSeJnfVAgRjqH/rEVInAAivSBvnhgH1v5SLBPMdBCu5+sULTn9pQIRKNAhRt
FX2kn93PpU4VJf9TIzmFuDuVORIp94VlItEhXuFNuEIpyIjNHwipUqCfzx1wLXFqm/7ECEJJKUsp
ZYBFKpOIFnLmpdMHmnA8Q2C/KoqAZbpS7qzp3QVpGuX7McY5xpXWkLHzClUK6jVW/wxxqZmUgg5N
quazbbv9uIUJqfp94qAZseCZYJ/Ou8aP2LRjAJh795nGuypmmz03y2aANre7jiw0xCP5mA3QPKcP
eAChPOCHaMeB4waFIcmv6k0W95xAlUwehulQ4vgneRTntZV5zK/tQVzQXqRSUN6ayy9b6ouOqRHZ
nekWhi9RGDLLNWHkzhLnP0zqMukZg3rSAbhFBPBRPBpfBVuUaBiRk+cUTRUg3DD7aCNjmdAyFMCA
2EgSnu3QTcHgv9mTO5I5iY7mehOtxN1jwjOjMQQfjzym0mEspW5NQN54HGWs2Mp7CfY6M4uBL/46
cg38Z+HF6YfIcx/jiuecBNkqh0VFsYqC4mk2KyLJvEYYOOvhNJUZf2mTsESAsaT/Cbrj4g58v+3a
oBb0l5b/0rl0vEG6bJ45mB3CoqOHrN3CWG2og8bpk9LC0c4B9BFCg+XG/DBfEPrbW5kquAlO4nmd
NCKHgmjS2WsYlw3g3LCPYRXOKRu/q6unWWWZ1i1MAuKuNLbpgOFk1ivwa2pMpZdrneN4zyBIw4KS
tSpT2SN2Tl8NtJA0iBGld1M4Ps9JnO91ZPJKFl761EDlFekOJ7YfxX/YQGmb4ID3mwFvt6Ok4nR8
gnDBjPtrWm2MM+Nl9J832Zo+z36kehB8g1pwzmvp0FXXtJGkXX4gfZuSfx8pYwXwNm9SecAmKxdt
xUO10ecVkJ82LZ4IiYt/xq+iLVr5rq87m4Js973RliAnFXylxUQUY3vBvarNt1oIuNvNyicZa3Er
ttBIy7QHJko1fCrE8PlPJjjVTiBR9nTqwJ1tRGJQZP4YD5eTxvaQ9qfpQr8YzI86yWiGyhGElE1v
pYC/+xkrZWgo5z2fJwoxNWRxY1k0mqIaYlH3I3qOzGMlRU1d5NXf+dUuthovKmxz3Ru+M/syL0cW
Qs92RPC2xAkRuFjQpv8It1z7umoWxT344ZKEmHi1q8Cix3CwpDi04Bxsiac2U6pvHta5Aaub+k2R
dB1qmpAdSjceE79hIDZQ1G/RlvfnskloTJA4DgyG5itIDxoq12EyFoFrfOSEtBvZmJg1Y1uAWfVI
aMMwVn1VpwkqAzYqbb2XMV6k357KRLI4AGuaOB+nHEe9yWuQYBZd/r5bNwzhqwCz0XrbIuSJGGXA
xvX//8Lau+Gkr60lByna6Hur7waAbZjXqhYUYn1LygdzlziKqYRMza8KPL833hK7kcXHr1ZHOxO0
HMtMNfn7BvuYrS10zhv3NgnLAbTZz2mcgNSr3Jn2no49I+Lu+TyY9wKkbUfFY1+V7ppKfSFxKBfe
4ADAFL8swRv4tsWHBg7QldBgKtC/qhEqmtciU9g+We3gr0pCsvrJSl3FafdcuUGC1qZpBCc1b+JE
YGAIPJ1SFK1ocYuy/KT+UYa5PLWCj/7XXDH5KTYkoL1ML3JI2/aNODbtyJn7bqk9lDgKE4KMCEWz
AeiVass3aw5XZgdntp//D9shNEucjZ/JoByckXVKbC/kAHL/0x7VOs/EKPpVHxOFJsoL8pBGKQ4i
IZs2kiwHawtttv1B/yFjGxT6S7JrQmSRj7deIC711QfwIAC8+q+iG6d4xbLQzA9NWlReX8Uz6TdA
VdlsoKyZqpFK7w8gcLqM2MkQDMQlrGYSK04yDDwImFn9Lk9rMgGkUKZOGEruhdRF8cgoLsTG3EDN
pi9y/z/sxKu8TVdStQ7BQOvZ6hd1e/TaTlxyi+8QI8XypUJc0PXG2mdupYfb37nOWkNlSpHWloK8
S7SVo+ye3dLBT+xFDS2IWafFm9al3tEV8Hw2b+Wv0Pv2unUnXCZBA/eciaEHGdBctq2C0up41r4F
QcnnS5oVQ9QRViImx5ksTtszTSghLueu4MdkAiOVOucZXx9Sf5Me/KxokPzYCWaJWZbr4vUFwOfb
5hk7HRI89FVLUDJJQYkobTF3O+Z/xwYB2fGIB/F323voGEJS5KOcnpnYhXtt9WnrQi78XJlMqv9U
J8w7DwRWa73HMciLzceLts0H/pP1Sv343sThDXRBW7+a2sw8fxPThgeN72bOI1Zrp2JZOl8Lr+5M
rPKkhShxVnkotOlz/BoATg0dQHi6LKLmYds83vLivQSjPibGzmFTT11utA1xlCZ5zf/gYA0KT2WH
A/5o5yIKSE/b4TgLwLJr3yR2Z7jYMh7RxPdefBUQdlopEtM376g6SjwCUYFDkyplRmkqY7U2Hpio
1vjh5Ti9dToyp88laRIB5C/SYNL5AnTOYybIWUAWDpL2r6loc3bZXOMUkFpc99z4cm0owQL2JS5r
rHG7W0o4hlc6GMlE22GJS/FlTC1Xh1guXSH+WsjUXJe4YJPhFzCALQ6FQOTmHCJIzqQyDvNa5fa1
pbUfptWS0KBKa+aOo9rFm6zKiHx6Wv4jGMqzwsZGxK7ImIPRqbq4E7mOorlZKqAUW9zaaoUSKNln
FFvrlhpIa2WQBRLJsNgBYr9jmJzg4WlL8poGmP05eo9z0Uji1HUk4Jr2cEV1I9BD5JmLGfJUjhy3
bNkJzY8cV4ZJXCDcfyaLJC3+kd6h5PlpYZ3sg+0aBkUtOq4TlpTZJrj3U0R5KMVIHU4DenItVJTz
Z3+jh5qf8Gj6Aq/ARfj6KBAwNjWtkNtq+yf2WfNurpPl1L29qKBihD3uIAdZZt4u91Z+9HZyK0tT
LnJAhM/hMsZbop6lXk0QMiyTlfxJL02kMmJedUOAUSPGWD1DnTYkB5FYxkGhPZdI9YuOFwXCtAMd
tVfk84K7aHgDE73+woo5Pe20oRbSjZ8W4Lg6c1WsSss8fqqC3PeRk9shdV3N0GPWZ/srUhVqSQvh
sVLo5u9L5km27z7a6G0enzWvVU+q8w6QZwM5qcl32sEjv+T4DSxnNFiGH4RjYuMy1WqQJ/BSj7aS
bfGMI2mOwrQF9rrBc6MNaiwoB3tD+EkeQQaKr8liUSm2xZjGiHT70iWqIKVztZ+3jnY9FTIMAi5E
9PJzhpauNy02VASqrwFPDs24DvC/NhO3FOj3VLU+bZ2N6hDmRK6lh3PSF8+OdiBMCEnv+rBNmbNC
ntOiN9yyWMSeYJxCzXAvGuIW1jxnCQgMAAYMA7rqVAUYu9A19fgnlwDtaigD9dClMbIyrEvBRoIe
XMcbdtpf6xZSF+4cZHTY76WyUMYYWAzaY/GPNi/DjURBsk4Yb5xNZnMlsx+cN4itnhm4+0NDfHsb
sJJZzAAvAxEEbfD310Oi8zwf8sqTVwcBOWBVb5OIvFjGxV2oGitzCOnGSfP93BjdmvX0FpfCd/A9
Sp4LP1GM8w9f4s0rUloUVcRwksQqFv8/cNzbcsnl5yzVbw01rW8kIcW3u72daoHpWKgpfKJNEYpj
67EdvDnRzrUgf265pyXAQz73//h2219X+L8erQbjZVXI/NjRUsNOG/62210py79yh4klknzebwKt
CaMT7+h5KrBPcX3MVBvhcJAZRMtDetHVHv6GIf7xikAcrJ9kHTUAHvE7dUPRBOCCf9gyot/njLhO
PfTCdCbdN7JXTnosImKRxdiiUrpbk+LUIl6BNzFDnRcCv+xfLwGNBXORaqyEJQ/9l1ExE8jwdP7/
9Jv7MpPuGz5FHbCG8OeiRom+Bf1AiwJQY+RUXgl7RlRd+4UE6SUq8jbya1gRLxGCk2UZo1+HlhoF
ngC0UbwLlmfKl/hHAMY6MmzWh75nTD1DHekR2rzxNCa0D/Cgpnm3P8QTKmxHX/P9O45rm3mVCYAu
tQczas4MpzFBDGqJixZKpwmQ+YxVIxYyv7miVk9/KDr7acCokkAu22NjbMczQhuoTe2DkTdXcYdU
nEmj7QKYcLFZx6Eh9tPQR/fwISfJKeORr4wN08NcC6ThCvtlnMgBmPENGIR58XdCpX2tmSDpFeUE
YryYPhRlJMqfY3rPHcSW0uBoFX0ylzWXEAq4hrYttqzjyswT7M9N4+QdxlGwsUkSzwXvAHnALGiz
XppiwV4o9PFL+8Sitn8DAViR7PcXjB9yezc6rU++Gi3ZVlvNW5unQRnBY/7z1BUn1y/oNIs9R0ec
azUTCymdzV/rzgrbJsDnyJX2cj0gJlQjtQw8cNtFondROkQ1twpm1LWXEI+j+c8c3/bhi+UBPwWQ
eOYnfVxVOpIzHNSmYpZ8Fn3wo0cupoEbbFHldHKdZZu9QUHT++3/2pWZo6ONhYadWvIe0MOjgKZD
8xAeYKlom49X2KXQ+4EJ6J/dGNIMiozNGTxHo6Y3MzVRxGJ1ssXlQfVn1KApRPEryHeZYAN7MNCV
upxwG4QCBQlrW3gP6MHOx679GjcKl1DChZzCYNdJ5WlmK84HP0naurVXyIuyR/d8454JpOvHdxaS
0LU84Bi+7h2JYaaag+JlTmDMayGiyPoFajJ6h0HaILh0ZWEc5U6owdlIMGA8CMA0yIO1gw2bZrWB
4Hw/Tn1AB/BhwbcJYjGRxhNiosVQj3S306UrvGgzckI/nu68Lc9fqVDGmKNHV3k/tktBTIQwrZY0
DjZ3dJanrF7ycniuwky+0U9K8ewkGXccOtWtuRVYE5J8ULrP86WyPT885Hg7Jkp8cDZUSMgGPU9y
EYQ6EQbU9gz6+9dg57217LBfqHMbL1gtfZSxZiWwLCNds0INCffdoiZNpxXUi22pEE91lq0beG+C
/uyva70jHZkgJodEo7jOwrybhMuMW65uLddB3JzZMKfvd7dbbUD3XYCOow720pMluMEGpyaA6G9w
seSYlDWQ+sKtQKsVdK49z/0SUvkZ2ju6unmey5Ac65wTWutLq1dPKsigR2I1yKBbOi169ZqkxvYM
+z2iXSLYgMDK+ZieAF/r+j2PpQrAfOAwp4ri/y35upaK5Hdxrqd5FXjq4zYhycfHh5lQ7LHWlalX
u1jBnCDbMSDsu2WoSHXYh+mXoZQ0aYfvyXjTPx9zCQ/oTs7mYHMi1MBquAD+dxQP/fwBlH8umyjm
6cz0vGzplXFrRAjPmXKW9D8kmHWd2b8QG5FRR1hM3onEI+yL11QWWwsbrBASnCJvGfefhd4dVY0A
6T1F0/E88POvQ3EpSk25V5RdZjWvkOeHrx6E+Ze/1CkGqywtsM+1K6l39xuYS9FzFSr72wqP3PJW
gjQ0nyJmD+XM6IXK02zwjFlUU6vaP+qZYgEhE7/2irTtXGY9Oo2kQT/A8fuLkuyUUFP09NL8Yhhq
7/+iC3cWxg93i1l4CWEFY50mHfoDr2quS4fMibXI21p5sCkVsdwOJST0A3T1xPceGKqlFEMlkHkn
jrcXHzZlbZzMKbhjMDEP12ZJZAjQoCb1I0vKSFwpYjWag3e+NXjf3y7oDaJX6UP4tk4OFxYDNk6I
hM6CVDiSCO9NYCxWxiLwxWiGYHvkSHKCI5rnZ7j4E4LNLT2cOs6IN7KIO+atPlsPh0lTdnLUYQd+
knVTziSxf63xRBz7myjMx/mCAWPI19F24uVUF7zp4VRm/3YonfDR0OSBXQx2Pv4r9Zi2iAImCiJi
BSV/SuNkO97mIwXapkhc4WVCYBxPgmeCx+G9VIovY9PDHqa+4I8Dwz0h81IV5n/uucjkiTpR34Jm
lduLfH2OTsqZ4Zdb8A2gmKGFAfImLvjpfjRAR00EwctEl0bzdjcrJBXBFxjhLIHiEUnnhy21asJ3
jvx5XzCs2OClxlJ2P86aNF9Vs6VQwEdgD56pTx7u3jDpJhH3qKPlYiKP9l7WxRrZHwW40+xiYCOD
j+Opxw565qCce0VT+TZIizv1yK9x3XwI+7nm9CaJPHWX+vrVagsqUy1Mup/cQIIz7VEkPLavhsUS
m3zi7LIF0hGHJJq/Y3dQFeKKXxcww/nx2T40kRQNEZ6HByVgfR0I621z+YfgjWD2H2/ajNRVwNA+
O01Bv8uH99nfN2LAeMSpDJdkFDgVC/SCbIQEhBcxCHvojZfvITIuin2LeaZXy3M0e5PaCDp+TEuT
Be2ue6Lkfvxwqyrel+S2ZYoTftejHXT/zhVI+Gj4nngyD//cagVykivsoBaCK/IJFxs+qaaXZgPQ
cv/NjxG7DQbEXJu2CFg/vQxuk2BXjc/OTMdGBTxMbLRp/ziFSw0mL9Ok6JSqNwnP42LVgquYECk/
aGUQNoWRm/yfvhRC4ecgGKjDZrhYVZZijnQ6oj8va7DjeLLJAz86E1sq3WSVJF13y2QZtQWj1lkp
RynitzJJdPahgG5Aer661Wjt6M+WXyDwFQQkL+LW525j5XjyXXbMV+wiXd7bIw+XI5ThTuNJ8oRV
i6DIVnY3bIt99MI7FPcOTaY+c59r0cmmNDC/nUv38WK/HGL0XlI5dewX6zrDwJ+PNmqCFvQHFVvz
Qdbq/hMv5NV+h//u4l++VuH/9aMdUHPBZsRBHb+2p/vzrHsZvDo2Xn+f5i/rU/eqV8I/zIe/TkI1
XRHy9wJLCABmRhfHAtImU7vny842/GedO03oG06rC0eOgeSelCKw3pNd4qraF+UiRyzVY1KJT95y
HL/eyCld2y+e0lp7IdiqnVQ9TFjwu42j5VxtcqG8wm4+6EL5QPTbfj6Jy0UT/x6765qp4uKhjkOc
cs6JQ4SPuY3G12nJcyz60d0JDDekgKPc9d8fPya+X5+nbHYeg3Dt49cAz6fN0QrJw3fIwnslfZ3B
0YThIrl/fhl+oD5Ehn8grzXmllb0vETvH/JtCFp0FOjtFEZ14RgNwWsDCFdBJrX3CiH/i5Yld242
Klxo9c3JLGaebqnjC1LpVzCaOMBCQR9rxes9PSQaYfTaPwQDQKSCDLuUau61ySNVNri4605fvYd/
GCDiwMRw44jjAZavu7MPOP3G0rRlJTpgV+5neX40Gqfg3de5/oehHkq1ml/EGEvDxoVuOjRfbnO6
xZrQcaoaJrO9IlwhTSwWZWpINcdJyioD3YwwSyKb2PYCu+dmmM/8FHUNI6ta/SxYRUUu+PSB0gn+
4LTaBwiOqBQKMHIsD9LT+xTZwlgmYRM/G3jm3ueafE/Sump3+XHaBnkgj9CkrNH/gX+2WfS5AguV
bUClq5nGh1O2IWJHyTrCeJR4JtN5QZsrs8PexyXTOAqg2shHgC/zzzZ5ubuWv+LoGUo20bPy17f0
QeTpPjLpsIbe+QXOq3ZjWHTNKJqvpNZRTtCGS45OHOuNPzBMNwYdgzfqPHMFJ23+tj7BSlv1dp63
S2lW2ldO68XnM13IBnaFP95jEUYGkMdBZyP10x+2Spavv//Qygg44n/O8W5qvI1XsHYY1/yLrmTX
G/7vWCfOZ66qK3YzsLYwWnp5PW03144r/ehvhgtChniOW+tF6EpNrAaPYwgOYdb0UaVIIZuUwwcW
TpTbYTfVx2E/kIZKjsCt5lyBKvB/XFSzMcj2T9X4Pe+BkihpactF6l+nEcA/r5FSVB2ut8tNi3dD
iiECUiTcfPJsVefMGy7c3bovYf4cbBBQkx4r9d1lhu/movgfg8v5rERJkv+t7HwLt9+Bjik9iLcf
xzCJ/wRrnhiVE6XKOtSY1laa0ExEF6rBvofPpcGDbeLZqw23rCDwKQ00WMpMmUkM0DtgntDvY0A2
vtC8uQb+2CtQ0kt+7B0OXK1AeyzVloB+m/mnf2VXVRTzp/4W5F5TeqBaeNITryjaqjBO8MqNUfnw
SyVv2oNIwbTpwKl3nraHPv0abocGoeNw5zNEzafnyVaj3c+KoHXJKZCGcX9n4iJ2x1vmR0bJeCTa
UHt+sCH9PLSW2pBesZo5KM7x81z0UoVAf6fKgkjsns9aB6C2G59EsSpA8N82gLedxl6ise0z9qY9
u0EbGGFOPnThYIHQt13JqyJ2UyUTEoMNKzB2TRCAYECIuoGVQmFNf8mF/O+ThyWUaYh3DDGnyI5P
TQl7Cc87JTEy3R2S3G1n+c8FRueh8S5PrCotwRNv9hsnQwm2h+favMNq6vnj+jKwiFke8HnYGAMh
1uNkTGVJRusnXqxQdpc+blxigKiei+4tX8a9ZemP6BSUtzlvNV5RqvHoPyJibQGEAPSUZtxjB4TM
YNycKDsV+2ZKwKJZ91AVGXbkNsKKRAetXZq5GvUKqSR/Aah/+PKg9S4B0WV8A5DJ9hPdSfHqe1kK
vMtMhvFIoljtNZdQ94PjhHqpx04IBO6O5uJsYTtf3u7oK5BUSM9U2j51egHfsvYhby1BI1eda0qu
GUULs22RrmIJfkXnJg2Ty7kfS4OiBc2KlPVZZlpNBQTE4lpV67Ohx+8tzk8Z3tyuwdYZsM7B3do8
c6NxXBd5j2DIEFxXEVy6jGSjO2Bui0ueOQFLbs4XxK5YvihjTTptUZIq+1JsqwQ0q8J9kBZl+oQJ
sGd+ym92VL2Yo0AEWQE3dzvF6iCrtBKZJBS3dueGS1NANy7wdddIsKjkLHHUXK7KhOR8wFs5a82e
bwjVpnEEvsi3OKDKi0xSYxesH3KMQ25V/z2rqtWVB+lG8zsj4iDm+6qF+datsc2XF0/lQkfbwMun
rgrAyVHdSKNMj9onkLbWMeaUvA9tOI47vDI7objYwM9HvAbkrU7TGyjfbl7K3cGlg0ZHdUcjnL58
aMI0nTuGIH03YZW57Zjfis2pgPVmCo+z/OgSh2vz1paKmZ2ns9xVgaTO9etMAu4AEWIkPtcUjesp
cGXx19YvwBd5IjkkaMqzLP/29X8qbUHgHUj81ndl4bmQxwjPGAMz+pi9yvAtYaF3qdlzDLseZr6f
q/uq/bKMKPd43JK/8/NUqDAWUEIfyItgaGE+2tAFDrzniiCTkefMyXgPOxkNvKfOj6ngxY/F4x88
RYHt2lj3kAHyAsGtxwhiZ2QHweDJaFpwy1AkfmL1H81aTfvZW/CyahI9GRW71CWsdGHG0UpzDhtE
t0p62w8eiLPDdsbWhgPxk2+UPYCk3OFDt9i4lFLKRtFh+Z+kDFR/4aoITZ/EMnajk/G1c+aoSHHT
h2afRletJH1dKeYRnFjMgUzI5J1gvp1kltABdF5XulWt4QYtNs0vS2AdhiM5fo5f3UoImR+EPTrN
QWIZ17MkAFk5Po3QMslQXhFoRir/WRVeROJTGkSJi6RXh3fZPu68CKmlsT2tU2e3gGTt+5eNJd//
M/r8jITy4SVnrHGWZl+6uLUDkQoh3doqqTUj/M5Ku4YZqrUIdm/N+DuPhgywaJDRU20zaNMNU4Hy
S3SSWNuBrMVMuZ4QXKSHPBv5OtD7c5bl9AotkUEiOli0vcymEJIBYuXsDfiJ1vE74m2IJsLFBLZ4
+wqCPMNKmHKlM8OkB9/4cgM+SMxi8l10CBhJIgbjGhu/iBiasYd7eztxg8zAK9GMDmNCEvwYRVhE
seRVSZ8vP4VJ8AcsHwFQ/dEqiO+/vtzx4Nv81inEZAQ+XP6BSTsGdkS8j2MHDpH8QTINzScI46Wg
K7wLBaL1t0u18/yhWvtFDDSLNpWly40FAVEq0HoH122hHxm1JGvXRoemCTopj/uKeTAyy2yQej8R
nytbnLb4/RPSd6PjbAaAMDELxc/Wr7AKquKREsOdJLyPc2xbyOLe8qso9PLIbuc4atFnhop/JcN6
uO9O1Gddlsl8PwZ4dQOTqPLYnBzWechIPU/iNp6EAV4+IMEFSEhky2oE4pD5fsNqFL9cnaPU1cLe
ROSfzmcOt9wl91a/UdOVKcXHTKUhvWnnYQ3MsD2YYyIP8hAGkFIARbJQu7QmmyVLBPv72L+uepHG
P8NGkTfLhTqejouuf4DBZ5sa+QmVD9olqlrnxEnlpactEVD9b0K6u4QJNHesonl6Hn0klV8R4Eij
UsNoGkA4fz0ULtTU32EpktrYkhwV11QJgZ7pblebq5Ad3FQ+BFxdvUoW8NwjzPcb4JeRS28Z56EV
mBtkPvwIISUOhImX2WjKHgTxbrDy4DEV42sBBpbFPDMB0f77ox3zdkCjnXW56cOcn/cRmGpSgilb
AMZ+SAM4ldoc6eJIbGIC56vIe0vvGQIPfhJBB5NSstJ3H5hsjIRUImw33sUoc7/kl3lhXdw+exG1
UsXIrNS347JxZw66921nB9wp+nGWdGLUSe3sMao+IjTh87SXiw4brwoW+QUlRnI/MKvCVqJUFtVi
iVJwlb/fgTIUYEgoMbihJAjP7adAal0xHcmA4UgokKy04nTx19vMNjEUbs2y2qN0HICPcrMzHYD3
snMhHa7v1t8IxHl1cWUDcca9yO3x7gtV29mG42Rsh+C0d0yabkS+WkIhLMdA607WakSgjFgKbyn4
HVke2ruALJ+QFVjd3fpib5qrov+UyZkDyPAfvhBR0Tr8PQC9SEAf18tn3N9ZFf6AB/EHALifS5QE
GgDHgVU2c+osMWR6Ckd+LttOg18ppfeYatA33nzhSvOZvMs3soEiWMeP9Onf+Rco0mBVDuwMvx74
FCWs+nK4S5LHr4aHnhtoSZvngJyugZQ2pAZ7T23CKVjrAG1uO8lx0bt+bohJQJFpT+cq83q7r66R
lROIALJ1rVagf1alhIO7a/8LNBl3VlgcBya8EyPbrDTaKR5fQD0bj8TV82z+N1+Mm8gWHD0BR0pa
dF43KJqFb7/o/gt6GWiO1Sk8yBtZ3NvqXde4SFd3yPnmQGmn4PXpaGiCqHon9xJxN0U048kRPSzF
MEZcQAl9D/Iw149EOCFq7A5YuRTfXU6IKdn3/NnsLwPIMsIK8KEpEFIYGVmuf38uR0z3do1/I9wl
xy/zCdJi5hS+5jjfvkgqaTIYTIwm9DIWWF6769dQMQFNsMcZXCv1L0gGMzaBPI2u64PSOPhOUpQA
OOPTH0XorOt5+7YMXx56aMsJEJb+R/udTiIBbEbyMUeraFWncD+mmFaX0ztSPOZR45Ik2yx/uSHQ
C06GsjO4ghreGrFRFP3GmKYPfbPp1lGMzFd8DQJoaKiA4HFn9ZTvR5zDRFqBOV6D7k0Pqf+PRBu1
fNhKn/NHKWCEemUvs6eGP9z91aLsc9XbYmfoLpoZdBieKp+NppM+ikouoeGMYIGhoysKZHaP+vZ2
AFDJotERBQGeaGdTcT+GP0PF+lxX7KHRhjvwvqbAD4nh4bGw9MCkmk03JQ5w35iJQO4tqWNr0JJd
AvP9/8CRYsyEq/gkV5SauKfMBo6MZPu1jyDcQh91JBgjVYO7fCjAluhd5rpoRkS187uo6FaQViga
kjL6WpDl8E6PMLkyga67sTK/j5C4Oa6jldjPXoVW/aR/Qtko/AI5NyfblWqrSdIPFCJTQT5IE0V/
exjz4SuWewXCsrDisbqwyaA8alUOMNUJvANArxFTBa6LJVfhaxtYSa/X1NaIUoKEOyJn4mRvBRQb
B8wvgiGvxch6LW6a2M1mRVfcvbe60oOhi/A5/rlKKp70oUmDJE6pnIns8YOq8e3/vaXvffPVRC+g
eb/rExgc7eIUZMWsfcbYVgp/xCw7dqSbnq6v+dEUuVKC/YK7PrSL8yysSh2J8hFiz76et6IMRX98
BRNfOW/q57JHmT8FwkNZd7PQFIIVDDUphVpsg28YaiZW6jMFDpgSSziRGbaNb55nFGQAz5HpV90I
jwkSkOf7jTSio4IofifUj5XhGJ8xcxFC6e/VHKj+dbB+GPu2D4Bl8ubT5MUkQ/mw8+Achf6Ankho
rVqD7q9FQn6ruy8YAL0C3sK0HsCEZnbk7Bj8qX7GbkSMPMVR2hDALJdnkR6YE3cE0LPn2GEEnjDi
1+lUrZyAjxKZGh4JVnx4MnbIm7qE3sZNLsuuomGsY8yg6LSoIsqyULVYXzWjm47MeXMVW7kW3ocB
1+3tHv9L9pzEzISiY9upIIuG/FOWXpgqP/E8VP3UqnDfK9W8FUupePCsp9joi9lFAAvpMfAVK57x
puBXyRmSQ1GxigLyw5BNaGRBem6x335UOinx67V+wiXte4LIZXP0+8Zvoq7pVQwSOYcCt90yiQkt
6czhaIimmeR6ofZUUcRFRaC8Fy3rpuUC3eQ8YQBdtWjVUHmf/gn6JLzF0J9OM9bNNiiWzU05g71p
xp1V6wkCmPIAQKhOm9YQZTv8cKh/GbauQyHpAgGAQIOzthemKAZg8+10V0wQGsBv4H6CfhlYsDMO
C3wGGr/tQVxKOPKxl3JagqdWTxmGezm8BWzySMprxq2nsIffekNsNJKMNP1t2qmtIPLHHvuDhPCh
FXO0iZfQcVlsEKYSz1kesa6RujTztlWdgUNjsGiP0lUbA5EHUDWa/d1odntvWUAQXb5BNc2eyF0/
5Oj8aI58+SVfpJERjF+3VAJ7vipihhEyUqL5W6+fzC9bBzh8Md9Q4dn19MVNZRngtHxYqlfSCYh2
XAw47UbKnb11vja7mKEQzyXpvt8SNj/CfS+OmfDhg9z5zWvpmZTXF0AMxrLOOyNxBUUPwQlsG/ng
DnBRO7lfUaQrIIOotMmoxExWrROAIEMqL6W+YXzoROUSS3gSYutd/N+HVFBNi7wH6VXLJn50+sQy
5kHXm2tHmPPOMVS500jo1vtDqTgZj+c/K9Kk6Sp1xmtWslkWPCVZ9SCu7CcexmfvneTTMF4GZ2Fa
qhDVXypsreuUqn/skO+q7wXGs1itxgj2l2E2n3x0kCXzQcBG0X8fPbYoH512Q3NmZu5jl5lbdloH
S5/MRth6leBfIySWbvGBBd+tA4a6a5GX8k3vYurfzEmBi3IzRMHVQvZpNm2kJpfLn1rZeGGw7v8k
48p2oBGaatw9UXDcElzWYDtCiAVVmySgJbIr7LuZvvuaId291b6poXaHGb05EASHzoKadlFRk8iB
ZsyoaZ8Sy8For8kguSky+OvybNTuLY3hFL4yvX7xyaE3Rjj7+dmgshMkU26OBFFc7n5rUbEnCtI0
aNsCQ8U0kL+G5Q8KKX5SJr069lDYrx8FSysnQNefECjNl7xJAMbsDPU67E/La3PRYgrYEPIp5mcK
SVhYDTG80JVczzQNX2hY86/F6fAELcmIeH+eh9ZXv93dMTwFR42WHprD+oRK7Uy7W8r7GvNm9oCK
YKmDNclrIPnpk+yOTLVTpVkdtV928IvvV0IyibD2wC8tbc9GSMx14XlKfbU+zdFpCh8aXo+gDEa1
fdfLAJJuFu7OayD5c233byRMm09OSYVWc2TzIGSLF4nBPeevNvOTgh52KwKYs8utYrNTRHvoi/bi
QkduIvg8xSJYHkdHlaJs2s2lIAbzglJFb549x4LkcEPX/z6Z4JV7bJeSKr2yg7bUVhM5/W3fAGHg
UBYbWy3HBgsmS2MEGhMXmspTgopSCY9Oc+iuCVvDzGvzglJMEaai0AwVHYJzE9tgA2BIu1wjGVvl
OLXj/KzDXlY+D4TYPT1qQlJpVfVjPuDUcSKR00euW43wUmS2kIOKbgv81z+3vgPn5v5tPvl0Y4TL
Dq8BptmB0dn2LLAYGVGsnw1m4NSIJBUYIxAHNRpoTVZlMbtowdK6246NysySTnLdj87kyPhvUQqe
bfes5nU5G2k+u3Qc8dSi9mKAhC38eetOJfhG8vgfPdTfmVUTuEXn2GkSXqAe/RurkM8x6IGNrz/+
m+B2WROK+u/5TSiq/n8eJnPWVtQk6CML+O90HbNXsPEWZ5bMHGjdmJQwcoC8cliC5UY6ZOgkeEi0
38aJzMmo+jY+yKRJg+Y54RJOmvdqHWtdSKCNV4s0EAPh7D4joZvlDIPF5On6RzlImIs3CA+eTips
vLQ6cvrYWzO4bluDIWoo+aqC8TdQqvSh2c2mF+gNrd1MRQoAzjZOYXtpHBdvtV6rWD0DVtzfwN98
zi1fgzkC6VaPGEJ3To0pRGQ99i9lJXBR5WXyxu9nQFARqE/A6kXpe/pFUAh5LZsAgxrmji6eFSqY
T7mt9BmueMPQZ5VPsyPwpFxFRrgj/S94i+gGVNrNwNaWMNZgf7fYF7FkRLcpddO5CAia85Fz4YAQ
AN1HzINAEHnTmxLbRv+TdyiOT2TddgX1NeybPDQB6Wedo2JLICSYFQOxU4DezxU90yWvArEy1Qfb
SJBbbhN6L9IeFEUVLJB9mIfODznocJles6dvgiTjzMmMdbg9GqSMUUMa5KrhVfoZCFII5F8WRCB/
GPj1Sn0l8h9LqJYq8O1MUtcVpR8qCieFmNNcE1RFsDMK2StbqeDFZG6QBSAJkFBF0o3eS1TEdB7K
bbp/ULe1WJQD0GXurNV/TKVR3UOHjA2YkB9kba8lVpZJVZ4yQtpFgp0h/jUKMqsHBqRfTK7hiOlq
g7LYJgdwS0+Enf6P9uUd2hVaMHqEkVEA+3EODhcZ/XhPrIgMhriTZn5+8PqOja1114je5D9dJnMt
rOuAraQRRYp5Nx/rXray8o/NBixRm3/IYXjjH8ZV60Z0rrrhBbkqW37wwYTyi3AYbJ0bxlYFQYCU
Qz2mG2+NLTyOjkb3mU9/K8Bzlv/I4vHxzVFhDHz6rQ/9Y3Z6ydLq6aXY3T+WIbPdZ5rDBApKI/r7
as/2bhQdc1cwH4KE4dPkpwezfz4hgM216yX9n9HMbSwEQf5hpnhRHfIOFucMyV25W4b3t9W5xsic
Z47Ilb0yJYX2CZE0bNuImwNbQw595mWdbMs4LNm3USq1LU0ks/SajBRuTBGZPrttLUxWL4OlXtMB
cB42fkTnEwNXd6lTkNp+j1O4tSoxbO7seB8B/8LxWtRSNsv9n5kSwYNPTnDI4iWt0+2MqKnIW+Ve
WwKhjt9nrQ6OgDIgXKVEuAqEihfWu4QH297EkyJZ5O0uy1plp/vez8HOvqkltJRoo00/VcyYbUhS
BBXJAl5cHwIpaJJdc0blM9n24qUsy3vaF7BTbjGgj0QlJ1T9s9fskmMlS2OsUkRlscNwk7ni/MEm
BUHX00fvyJWLJ8oHK4ksmBtCzaJ6S8h/nM4NFXDDd8ABmr5g4QOvco79JjI5uhk2tj6851ARdXsv
V3ilJUF2ocTzX0672yGypy1tVZHuZAwsy12cLp2DMU0ZOyrhf1CE+8pUBbEEBwo8PQrkqMc04kgI
qtazld34n2capk9F3bNsy57xDm2JGMGYf8lJ49v045HgZA4G4DZR3zCouZTYdt7s+NhgR1QLqSyV
BxaQF6wt5OnG45hKqTAhOMnSGOLZpz99DQUFlUMoSCboixGnsgmxamPYWIO3z6CcYn4sjbzww2vz
V7/WUIsTQq6Mn2eADRRZ0TW36W6aln1enRG2fXjUYT0z7Wj48pzoBFcPdxBrvobMPS4fjVjQLk0t
hZlE80tMX6WJAubaqe07yo7SMC3mlE9reDU2KVl0ro9RLhnr+wTab6lvIFDJAnwjeky/4R2/pBpM
37lgwNw4SuiTdFdU8Yortc3QIO7De0DTyFYDGpF3vHtI69DT5vc2C5ZKVBKMJ8HxyUq9J8H+l6Wk
bBTTjXMgP3Tpmw1ddtLYlox+9lpchLEF0bFaiJNoPMbP/6ZLxsuaKYMajayfl329+pZs4x5kttV0
VqFQ8sUKFrjEAYesIK0u8O+BXoKNsOfueLFsfJSb8/L/cGCoXbscYbNess+4jspn2q8ZI6CQDop7
jbGIGUUB+qJzLhg8bzUd/RjCHwHwEKd0TNqIAYRLaEqktgumzSivDoZu9YarvkdnCk8fv+lRlWeU
X+3B/lNeF0ub5Zzi7N1aLN96YJOtS0ED82zWYp6UreKNl/O5LFh8AVJw15arc8FBHWc1KVd8dUIu
E+O9tYNLfUZiO2HiCTFB5+m8pysJR9fleF3iWVL9FwdYYtSE8U0/4AR4ij40yeFuA9ARiLt5LWHk
Q9pSldVoc5p4QmoVmj0JSPW2Dh1uDeTw3rF2SpHJ/zg0n34l6SdYJMdxfIP3tXMufBmPrB+y4+aJ
Vi6EFbtv1gsbz6tKYUySS6UtUYqWvUJvT02Hy9Xs7iL/+ivv3U9FUcCq9dMeHawUCwWW0webApt8
zzq4OAlIpCxK086+xM6X2VIMlYIpdHWXrLyNRVgSUEGvL+KA8QO7QaMNlbHcvY0PHgrAme9pV436
5JsBSFH9X7tSDkmZ5TelcfhgRibU0R0SEVEDeWJHstl1651Mmmu18iXK/fq0NCSd9tGcYGS2zbG7
6HyZFzUk9/Y8psf90ULlCOFRd7NLEH8lr3d9mZUeuQUYvefbLxx2apUBPGkyNvW6mdzjA25ACXdg
T1SDJHarMOUPmHaqGPpXlvxfpYIPzN8mykftcoGmdI7AQjfFVqKaAp57Cd4UTsW0nO5GO2va3WFp
5QET26Xpwz334LhX0H/P8uDyjwU9ZicrONqb8CDlYGjR01XsMVGlTdy049KVa7nGZZR1/7/1c2mk
TbhxAb1lLo+VUNRGAWCfSspJGMSTh2pDmUt5/KBGoDD1wkIc8e8CRsHNFI/fCQQWVY8GBblRJ1Ed
+vIw4q3TJ3Xq3s55DCeuQAaN9p8GMHWuiUk5iQ2K6zksdvX6nMqj/ZIRXYDlU4qFqvEJudaWnWrm
OL7PCWANapRPkMTuTfX8Md7JP4mTvrUmpS+K+7ruvell3sl2N2S9qLHI41CVeECfsJsAnDvRmdVx
IhbCXz4lls+9fb76m0ZAm8xclE/8+/d5yZJCaDTBxlGA48AP6HWJsHyNoa0Iug+Idv6DeBQO7T0R
dHjSXPgLbwG7WVapcsVo3saVldF5OVTyxkhW/U3MdtGutQ8QxwJRGmVFqJhFKONVR7Fq1CJHcMat
FLGuamA9rRAaDWqeLbzj9FhBv3dVVu28KZB+4w+RvQcZ1lKSvw/gUNxx034//tIOQpt5JcyL6Qbz
NjsIrT/zFY8nUsuSapcY4LFLU3ssmnG0sx6qyOaoNFdRywZSEuq78WiKorbaonH+Fqhu1s0ygjOr
O1QltQCHKQxuj6iuNMLzzCtmt/Vy2aBoEdFNF09vRFGBAcgFKUip8KV6ANKkBt9MMObBFCyrhOKS
8PT3+owTcWGftIriRrUDqGIKWw75joT8ZdXBtpCdD9iL4NKvCVVuEfIPvLxh+VWxytXOeVC7tA7R
NLgzzo/M33R6Iy1DSh/vRPLQVn/2zzmASy9ZNrdp7f22usXBg/cznILIstpX+ehWV8I+WcbqdtRU
7Av4G//dfP2YFqNCYCG+HXxLoOEqa7+MOZno+2Pi+C2uEDASTf93yXjcI3jjZXSfJGujRn6/TeOk
x0C2Jbc4I3qZBO1/1gTe8+yyjvyyKSo0UnZ2GDu0wTBL4gV8bB0VQcpKVq8rq9Pi9a/DkfQE1+nY
OrG0smL86huq0Q40nqN/qGvxt3qkrbOiK1W3R600NW0zu6R4OTHE1XNqKOn170fMznnIi9My2vPX
rOVLN06G/vnXavuvs+OGggf5vryxOBAHeZpgj2kPdwHZ5jmnUlpNr/nBkuyzwaSYtRTPnue080Gi
NJsifr3J+rK5yK6gysav21bhRmDBqoApT6TLkb3OiEkFKoBSeCCHelscM6NMevzpeGwa6nf8RMBZ
6gievuRuE/32SzZ71NaShQB1ypthrNn0BcVVKtIEmKIo3un5JAdrsEkR89lUpDlP8z77bVgo2Gol
lRR27DKYgyEbMB7039PE5Z9VkgGOyXyPKume7i5P44voqYYdVa2ceVXeWCMzSaQX1yruKQ7Rejcs
FqxPk2Qwacf0yYZV77Yy+G82BthJVVu4CtR94rF0cg1PMXHSlKjZ0NaGSww7dAZ+9/vJWmVwy4Wr
R7l6cyB1zVX69DxnhOkURhTKgAtSZaCQqYM09kXFIsCpIp+jTU69eoHSUfNxOEzR9CtGGZJebT9N
ICMK3k7dSuqdf4WJ7qgC/t6jWQtSKtHyM5oJiPp4Er75L1hdHJL8UUFQf/BgsCZI0zxNfwoZELcQ
r1uj/f03q5QjItZKDf3HlNcvPa3R4rQw4+W4aru/aTwZrDxZCajezxIIzqF5iyXrAqCbTumAIZw3
uGXwYaScj/fv0xxRkSahFAHRZdlt5HvInR93iBCXkAJ/NfQLaQ3no1QRnGg9dmgfHZ/GMwaMWOmC
JF/Y/ZiQPXl2ZluzCV0ld4LAe6PfHrTOIcYsfPEpoJDVZQEtJw4Rc9Ya8+3c5pdw5mL78eGZElys
dWLtkl6LTZe5q/pgW0VO2bJPvTB/gJ+1H9VKDg2xVfvVAou7b4oy5IGrQli9dUbhcL/ACoNKkeuF
gvxuonxMLXhpk6FrjELoNf76vMq3itgUy5bHf6Co/Y+ZPXxWpqAiVQ9kKgQ8HJD7YKC9a7WS8LYh
PPK3IUOK71UB8vQw1ePt357JoRFtSLKbr6uVMFfWb7Z4gGBKaDUj5b6DVQdIrBsf8Z0UNgJmgas5
TPd3Uwre3/b4PbjkY4Qg3n7weyM9VxIWp7RN+MnFYHhOZyBOknNdfqI46tKeT49WQ+zGk4ZUwCjN
OD38spEYBvBpNRCksEiHwRYbEy0Ga6PwORK02voIq0WLjYoM47lLAqN9Yk5FL0zrJ0zDq315FJKf
r8GYJpI1LETs+v/i7eqS6MzIEvVYBZ1ZSJzydD+OoAYaVm5VuZLMktW0lmeUxU/zephokRuf6RQS
+uMGZWH2QQgc2Q1csw7TkgR4vzEz/gKHgrXQfnTX47ArXXRPQckByqbeZyMt+yZ6xZOA1R3MgxAI
IDoEhoRD49iPhdby7Cpx0fKxpVusCaikGxD0Q0hphxfa1MRF5v02eZeL460KOb9hIS1b6++QJKKO
M7mLdSb9e67nbz/d1E6k4Ws4PXxBdDv4hJXeopdBjDOWUDwwcX6Mv8FN3hbN+l8xa3+khQVi5Wen
keMxR/l1WgtqPSYj8exBFBzygIQ73YSyYD5Jj1SOEm2QyMegs3Yh95AiQQ+oEiM0Ix40iml8E5+Y
xUNwU+qoCGcpOt8QmyfphnOfc7THvxva6T2OyhurkBsvK76gJOMMj5CaiDiqLO+74+GTWFZio3ZI
4BnhSs1/GtkzGoE6F+QJ1hE8xsSfYuZt2MOGPDQHAMgx4YasbFv+erCYZh05CSnv/RtK5evx+zuW
V2EOjUOWvJU3nXs5yZE9iRNEC09FN83WcPX9oCPo0fG4JmdI9JqFskIrTqf4x+uzotqo/y6rG9xV
N+a7NslCyECW0LEhR6w59qsshfSPYRNmOqyIxD1ihvYb6Gd9MjCroHYreg1uDcPxPMQcJd821K00
6fDozndARVoZLownflRsIScmzhwkInycHh0u8D/P0FXoVyj/0t6GcMAzze69cWOSaorUhu4sIvPJ
1QVCu0qSBVuFSaMlcIh29XbvZfZ7ordYL5emA86ySRhn5iFYRkw0aEz5ht+T8odYlcW5OMCyPkgu
O6+bR+MeWA+5/5NkftivLwqvPiPIpvAJ/zGEoyYkZKVaB1EnIVQWXJ2TyN9tP5YkJ7mOhf2WpEpl
SMZFnPjUyMSCMZOI3dNJmw9TSqgfwJvAPLAf6ixAe320d4lzW7AZlx0JS+O/YSS2bVTBOdzLupmH
l3rHQ8C15FZeAoDyF0fBalnXjzPp1OS0xDCarxdp8YmAsM7K7LdZaxish75Hwl1OmIIJyoU5iArJ
g681dbVXSc27hHoMDQQdC8iV3nv+3K270HDEX9fnDtSXi1NCuF2Xtv4Zcar2TZsWrn0g7yhxHg5K
iKhn0l/UTSK0XTSuItbQnMkawhRvLJt8owBwbVCrvNwH17eyf9cuqpu2ydztf3LRYwU5+IVvqRZI
Y6FINOZl0T3b9c7If6CCsaVQtBUeeYdMw0N6bxQSS/3IUIn7sRmBNN8Xi5qYX2rSEMGgwaO/8Ngu
eZ4K/AwwUvREfvS00Pm6DA9M8YA+tpS9R1sbc1VdNi1Qs9lwg6BZug4CcrBbPE9c4Tsiht9LuuAg
VzPt/j23YZazwEhD8bi5F6bcwrZolhYdXlNpubkgNgcfF9btNUw4RSFSu6lpOItnMZEpN3OL1yiA
fmZ/YFAM3rhw1ZOrNpanCabTdQG/tVFha55jNtbFXo1AVxE2VJ2ia64sOhf5WQHkYccQ6gmBR8js
UydnS7AIxtboBjnITA5kPLb2p+LeIUo9ErbeludILML50Jf9J4rN2OhZLag/UCJM8zCtQ7/Jn+as
QYleohlY5kBVuahzFF7ADokXwVWJB6JLlyQV0YWQRWLu94J19WtafLwUkC7dJoe+gBhPOmPA9rGn
oE5ZAnFOIX8yTC+fVyHQHk2Ia8MVchJwcLLjVLJu89hwHjtYkqPrjZfma/co3BLDUrvSuzmfQUeK
Lkt1qZ11gpxpSVEL/AHGdKRHGWnvph/plSTpHudB2Iet4/ERZjw+uHJDf7K7UA54xsKOITbGq+PJ
fLjqO5FyfFPS2Q8YcqN4myqjbj9ANZPhLWcx7lthJLVdRZOv4BD2bBE/Ivoa99ePTQLq0ytjqgm+
7/LBaRzxf7ipVgf2BEYKEw+HHYUA7VnakzjDMD5s4yTGPia4HTusD+5kFBWSeC1DArWc5dlSEA0Y
nrdc7OtyxedmlmxUYHw6HWAYCWZ9s5IdToFsEAo1tH4bFAXBYgA7tndlsz4FrRRPrrWWKebl681B
P6v63o1EPUS0R9zbTFGna/AqpXdNnbVH+wRFF3dQEn2sLBBNno4hbu9I1mT17TJS+m/VEQDTys4F
1yK+2c2m+2C/9b/oRbi2o6aHBfJ2TNlarXBmKkNJ88VPT05GxSfiNM0e1dzFKhhLxB+9NHWrwgp7
I4CpXkl5b5M9sLyDn6+Af2esj2wd1wCd8pR28z1qvvnu5JybMasG/8JopA3+Qg2ZK++t/M2aY1em
3XGUYUzTFFYKtRVxvPeC0fEwjkdzY9vqSwC2COF+5g6zpANXKwy8437s2XgzBIxEtwVKP6E6PRJo
x/07mu4Gl4P3G6yw7ZdGNAPWzmrXUEoy0Wf67qEy6VvmNHIFs7iXRHsUhNvgJv4WlSu/Z3l1dH2e
aFGRAejFBmYqmfDwjdMI4GdJP7ct0bbByhtkZGC1hveriiv/07jtzJcswYC6HVkesNFau//PuzUS
g1D3sIMh1w7BDwZbBH2IepTkjHHXmJj3mbMxGMwAFng9maKrflN9ysTTClNniUftxfEcrE5SMjXJ
t8pmGhsv450PjII643tCT8wSMMDupsIf5c3FggoftacRGCZcDFO9clULdyl4ff6Na4IGtK05KKSx
HU4hHI4T36q15PYNm5fpr6ldu5xALuoXCWd9+HiuJjrkSEWXvCyJUVGknsXfa372r6bh3GPzg/Dd
Cg0re6ivjOT0SyGGV+DXtj1xOJBM0tvsfb8vhTD9zagJDvZuN9zmmZ93WdCzYFE2Ucp99YqY538t
H9wbHdP0a68NC+wWJ2gXGW+qonyPa7FULTOK02Avi7qFQgLAxmHBdnd78QGK9fThukdXg3jc7mAi
SQCDAkRr74Zsjl0xuVRdbXGJQquLnLhvnaxE2kNPKuiWMr9wfce21abMdfVOlOuIIAMg4faAi1dV
HDCpdmyuKK1s+rPOI/H0uJmj51tuU591UFNZ5nM4OALnZDqgmG52zSQ/Fi5VUIlmQHu7Mxw9xTka
CmoPQMrHZs5TTeB5Nx1ljNjJenKAH8EuQlo2xSwgiYLLQlCl5bfbYLBlaDsAZJc74iexCxNce0Q8
yKl8+ueBBoQE5v2DbAM756HNj4kCT6GpvbJ/3u3nBNfSzf9KNs+TISLDP7CBTB+R+cXHIuOc59ku
ZUf54O4PfrmkcDM3jvEzjv80Z7aAtZ7xUMDO4Mwwdyqwhb0NtlNaZGE+Kauin/SBoZfwLN2kqd7x
XrKitja1s1GKM8tdyG3Y/nKGdG0NQySL40n9hE2j8tLPdbQ+u4od14b+JqCCyKYYqf5pipZ2JBmX
DdsIFoTc6Q13nzURmDVDUdv/O/4RqwkVxTVxJ3QqWHKU0AyIAA6HkAOXOlED9ewA4zZ+7G1/ANrJ
2PrKmw5N5jT0kk4ZZwuvsGXES+q+bjg/MVEfP4GK8dEZnFf1Nm1vJ5TzxZCjrH7QkxrRU/ytz592
utFyOAF7wTvChJHcyJcPVhUxhWzfhmGF4h4dk9cqdzRYZy6fxogda1pNV9TNQEzY/qs7EnSkvUoV
pEtln6WgAe7LipxiFDEp0gnm+Gj/RCIkYIpCNCQ3xrGZwslVnm50I1i9MrH5sLX7YIbOB7VtMObG
bJOgR9owmbmznwAKYmsv2swAW8UmUOiE+2Ggf6yyrZG7vgmo+Jc2aj0/SbjJds9UA+6zatj1D7kC
RZDm8W+y8xBZxSHlDKMgwHrKo6SQx3vXQFOikbO8T7ad55vjiPt5FQY6W7JT6qvbdOt87mH7o/Si
KFKNQ203GHEweVf+ufacfkAAMGKjOijziI8iV+hxv/gmzgSKvwZwmo/ebUTIkMKICayVeu1WjYUe
oXWblnWSlpVrOzk3SddHSkw1pUFCmPgWCiKfJ03qj6LENvMBANUQdwLRYYxz7UiuI6SlHO4TVtGW
X7dB9GAjop+b8Wzql43AeT66lAL/v5yqcMBju/NGnRJCr7bQN/TGTVwCYBgxBWjKT+a4a//954y4
QoYp3U32gjKUIaI8CORmaDHZoJmdKAfO16D5xw1kpF6g5BVzzbZKuowjE5aKI6IWxkbbZth5SDzV
TXf2s2jXxQxQ/MK5kjLiRaM73j1UcR1IdyjCEpiq+wJWmvhDnJJD8sumRd5kptqY3kCcSgZhffJ2
35+0TYhWTTGCmEJ95m5urPVSICH5i+E+/ysf9wdClzE+GiNQXT+ST3J9mWhtecjFlUGKM3w+AFjb
W9HSqgJAdeEPVeExtjVJqgT1jp1sRMOZ5Sq0GBA1xvUzLkfc+4hbMLe1fG+7TGV93I3zQqoB+/Jr
M+w3/h/S+9COAsAWRtxGiNTYWQzfUTZMLvq3K5vUEq6XNM1Zw5aydP4xGPp+jpOloEWrNs8kBqLt
BjIu4yTRl3lvi1y44wms2RgMEtLaUcC7PC8AJI64DEAqqcO6Djq8SqJwartE2G6tAZDgoMx84JBk
UPVPrsMQO1Hb5NkBKfIHm31WAq0yMdAZlSKqdEEWP6b6lkO3r4CxqFWa9zVjPPIsPiMqxXAhdrmc
qpyAp6HytjoumDlJqX2+dmUOoilvcofTFtkp4KBEi7gj99PZv4kV0k8Da9BhKb9BduHbiLX6zuYC
WCcflhW++Hn6cbEJ/hTI38jczx3YSXZMlcjBjZia16heTWLGl7AuGn3Tk5xY++vtLxBYzjXnOO+1
2VVHDsRSS1yeiQN6DERQrtnxVUMRI4jcUc4NlY0epi4ZhQT6NOVIEqeNNOyzLwzgGt9/ioe5LIBr
lj7WRfeXEziUZ9hXgF6KM2ierNOtgs8fAvpOrnSB3iCdUXuv+TytE7pUEmGQYP+2ZSR2QHIeVS5e
Kfiqc+ziMgBTOimZEVUODtWUrqvm/lZphwhT5fXTcGaH8ere6uk69Z5/WCTVFk0wFJNR9neGw7sX
GGhqz7j7PO6LYy8xaCX/L4YvsS1uHc9zHYgYqF/jEcaw6FrLAKIAUb/8SKioBp67vlw2DnMnYLA/
Eo/DHZLibag91B6zAUOL/5MYMkaWwvO9Av/kuX8ANPfL99bxu3pCJeYmS5GgZRVPDCgr5LjaitCq
5xagpRrNbUGX+ZGx1xsqX4SYR+43BnnioCMGOU9E4OhIJcVaipqfhVmkcmIuMJcGYGPbUhTLc9gx
VmEKmGQsJiXEFnS4LbfrqMh/Qmyefj6mbMwrHv2rjXtgz00Y6KaEeRckSQiFX3EGUrGWEr4/t5wl
4n3GaLEqDZ/FlSwpgoHsiI8Rq/4CA1MjyDKJ8W5UbmOzRcDgrLVYc2cE5TsMI4B/0O7pEntT5HCl
gUpEI7evYZLiU7MQ0YVRo8biVz2VXqEYGNl+Dnh4tNijAk4/d9iQQ86YCCQcoFByWAxj0EJjUPV1
1fIEBKlwUPJsFWqd0bIoea/tcMB0ZDPO+jluZAF1n5x8R6ACDPSa+g+AEJH+9PLWy/OnV6xvM7VF
1B75wlSNWXBykv0NJYf5rZPLqxKDVQwZMDdhoQm73dLmIePBib/O3sSZQXAqv0Ppl+/UqSBuN6Dw
N2fSPGkz+7wQIvNYpcGe/1LhjKVjkl68ZdYP8sd+nKQQsSJSGXIN02aEr5RKxv0Wa0l0Y3RS+UMi
WICI07mOr10of59NI3fwtERQtA74dU2EzQUkvVwpme0n3jQ5uJLEdTomxBcy/vTIwKiWd+l2Kdyh
qkTJABsn9GSQJnTzBKD4DWDRby18MT1uRtKeR05OsNSEQmwCN6qllOuDiNJYW0sDfU2jN+NJnVb6
e4J7kuafT6vAPN1/EM7lcpkFarkL0lLP4H5VGLpz+qwhsg3VM7iqrjh0NijSPpXZB+nrvK1MG55j
9UMDsAGjg6Z47mb2iLgnxiyiDyJqsCeffJqDMEkjGYt4xbAP4VrUKPBSGIFC+0epOdeFFjaNjZee
a2zNPgZ9RmQde4K/6gQizGZ0QSxWcdd4yMYG/mByJTUMZi14VpHmWn7KJumlA1TYqqG+l4W/iBZl
OQFLEM1mpMHyUO0DJWoJxxTLsZoIpaXm0+KK+S+68DUmW517aq33RltaWwM1eMpz1766kBRo5W2s
M/6nvsNyQyVMHF7h8k3e7+vSQRPsx3MFwYOSQMscXhueB9Ermf9hqXlLUH3gTazSjpcEBWRkznt2
TwP8JvpdMY8Rr3LsG0AzyrQUd7bSrt8msw1RzJnYSezKLao0grcf0KPsybpS8Gn83vvpHUdII3Ij
tNEqb4xvWZDR+u0p78nEEvi+WqS8YZKuHWuDQDyfvqYXC4R5MdcOk5ukTBpJTEh+PiOOBmFDdJc7
02Iw9TeA8Tj4DgUKIr3j2F9Zby8VYOviSLv6Wk7eRU2UkURmZBYegKUNoRQtwzvRevvd0cYGxzjD
W9UHTwFXNn2oHX7TlMPV8IrMmyHGEUv5vrgPnhhpkkI+mBYJMLh8Lj/tArHdOZ6dWpk1vZjCzAdo
MY4WB26py26x7CaKXyDEt1E+fJlR+Q5AO43BwEIOldfhafazD+PKyim2dhzq/ov/6kJoh5NHMvcX
EMxlhjG0nqk4G2NiyJh3pqqATgN/Ag2I98Al93X8P8o55X2HJhx7rm3pBY0ZzXJp+MNlSnAw1ktw
dVMHMkkB6S20zSzcfBvuYRaKxS2K/oYc3XE5j2OxQNCJGgtFTN1rCKo6YggDwRCo6u43Ple+F8oU
I2LFutc/qOhEiD9oBjEqM0IH4vmFid/J4TRBd2QcY6J8yz8qumAKPplsbu7jG/4ET6zYSQlvT8Rr
RSL1aH7dd+i/K6Vq1m6a9TjYZcyiGpqCMraqbVNUpFfekHd5NXGQXF0aheSZ198jZ40tNJKSw/g+
gsMXgZG1HuwhMQgavVxhQ/4JlSpkDw0cwwVNsWgr3i1vvIiCnU2AEXHQA8DW8dVRLLW96x2GK2aZ
PNNWEjORO9sw4t2wz/ZRAYy2beY7Z/VuewAtJlPW9ZVNDR9vwz/CDh2vXknxhYBAa150XMY9x6K7
NPXDAXbIBsqmK79wZR8JLxZIF4yEtpDmUTLEWGxUxX4u/R5m9v/Z+TOA0ZWQYIUKcGsG6rJmKEei
0dpuYc7f5zX1fHNQS1Kr4toZ9WScwM4nswEG6MzkBViZmNy0OY1pbPMp2jSCz2jtmyVApoAU1YXs
Kw1mMaSK4yE2+rB/uW2/Qm8pUsAcJLYnwoAsqr1PxM3YIAnv9XejTzYRzdoIGFI4/AmuWKcTZsjX
KvPZqXHdBQjYY9NcT/AvUWSiXoQCf21f5GPRjoGyPIY0IR9eabCKyWfIWWKHJ8ksZ0kdSi5B86Vz
bRPSK33sV1OM4DxrBDEXuN0upJlpE7P8fAMYoiA9W/vSJL0e+u3WMyS9C65g0t2onn21iY7ktSdE
3PEoNxSSTF8i/DpyF+l5oSvRkKno6//T6rTP3ZFsNU3P6zWeQ4M83ZOYbk/dC/BJDB4rMHESp6ei
dDwpPBMPgk64UdbQpek4cusdiapZMTI9Y/rllarb1zPQbSQKdSf8CQG3EUBfrAx58JhnvSmj9y81
WAQuK6m/rlQihxgbZgfMxx0TWEU8JSe0ZevYcAFzqMJGMXwQDl+cWICfm3oUPBG0TYwQdFLN2T9/
/REG77avwrZf7hPvZxIfhN3Ot+Plz99fAAe8g2zvk2CorlwOF3VU+aY8wg+0yw9yoYFDt5tubWmw
SUAx97VVpuF8g1oGvV3qIU3hYGLqMjWnMtoat8zx8gL26OE+v9/PfAi9/V4Yt8nNxuSj5yQYyqgR
aQ3hdVjqkBkTto7RHC6Ui9q4apaxPNr1H0pGB7A4O/Otg7fd79UfZhAWHkiLYgGNffZGBcz8FsfK
n3UccdUKhAMgPxaTFPRUnuMAbWAgamc+IXivKjZJUJBCjk3nsvsI0LKObq6dJBgUHbG8edeMMUt3
6TEdaBpH6u9QYJQMTvZ+Wyto6ctgxx6qSkACFVcb1dMqmw4/PZbR8O5V7XTRwKTGbl0AFlD9VWSa
qPh3xbJ85VpNMTrkpylr8diZs7b11maOK+Z85TrVwgVj58avL8LndbS+Ye3ca8ldjOSS3e5TsHvg
UEeGej7b3vgw4QNZrBcb3Fl3zq85rsn7W0aHQ7ZmWq0HOuTs9NKmtj0cRv+w4jKypJ7uixN8fbz6
wIUxcT8w3ewzn0M0HZJCUSawK9lliOfh3fhrUEdS5h7PHJbATp8fuN815X70af18J6D6OaPSYoTp
JNVfALF3xAzQm6rSiVKap/wKFPI3YIvBHWOWy9fhRqDdQfHxaeLKhhU8PNtpfV329B6yP/ukdQMr
TtI4t3SPB3nDkAPG4KXid/gaYM9Pjk4Wtu7pGy0jKqnPMOY5BW+97VORZRHZ7vtlLrggj/W71WRp
bGiwiI2XehyVEDZGWT6bSEqfR4AB4ymaCTn/b29zR1Sezao2f3CO4W4Kt0TTtfK0/RIxFVRYh5x6
irUdaQFV/fg7ZyfEQChDGCgCvva8j+P8yNKhcFgKXo8UPXWJmml0qIqnKWd9Ex/9TZI+E8dxJBs1
prUvSL65sIKRKXAJgKh7Q8IchDwnEcmaxYeKwZ8bA8B0Pal3fDN49xyck5VP4Bo11R1RPX/dJQeC
cnZOCCg6DUOKJbCrQ5nlKS+6i53482LOneMk9D86YMC9UoDtn05pRQ3dAIQadAVZNrfTXqsGVEgU
B1pNOYzsPhwq2+OCuNAVdtsb2D3wJp/3VWWX4W8HOS/a8utwFyzxdzBMudPL99vqpSBsilpmCa6t
pf0l+rS9k3dKmxnD+doAqHP50Kb3abAeCBCNZieC3B5/z+qJwPBlD+PSqvZeRnMcPeAuwUU14DEl
hSyXwk5Yn1hAdMC/Y631l+O3u9tFUBK/soI/oygGomG8aF6P6C9M34nZudEUW1mzXO2r4YS5RUUt
l6+rYgnOdXvhS9BvxlT8iTWHNXAVpigS9fnAb5ysBx9pCpeWBm5L/ehvex4xQxRLEAlUxcK0BDdq
00+hY6IeAbtmAJgn05amZHvKac8kSyfmaC5lCTnC0XO9njwrXOr9NfoRfdGIrOoA32+C/6Y+RPdV
orLA6Ysue7Z1RJQDQ42EazsNMqfORtgA7/2dJ3HrZAY6apH/fkrK2Fbg2D6ggSYhUO/h4vQZI5NJ
vKYyoqptwknLVtRim7x6M9jBsVqv6w8QLMDWZT41/s5R9R75L8hN2qVBejFdmHk3+s2k3H3JaQMF
HrdBez84LWi+ouTj+YGvjUK2YRRyVNKgi22sBE4YOepxIG5GtQ74iuYpVgLrTAt+vm8X0p5a2e4m
KO80lxzK93t1LMBhhgNbXD3HWVu7QPG6BURsotF9wHt4+DrqWtFK34h4iETl69eiYmy9SfjDRo9b
3tRG/pAscczikco5rccbxNpPJ3uxIDAqsSK4jJKwpW85YeKPY3dW+jnlbGH9/ISoumbsjfA6qXH5
xqOyGWkAPfxMg1I1AfoZc7RS9x+skX2FdHebOQgqarg3k3OufkpP+WERXWwy81RwxPgoo67Mop5T
9EPzrEYi4OLPsubrkEVQpJxRi7WjzQd5+MZZF+EQPk21r3eH9cMGzVGiqJPqY/dPxlzFa3Qt4Fqq
tkTaWGYUn4SvqylSr5/h/lexop1QF9JhWXCk5RA2oIInsQDmtkWwbr/TEvWybpqfvepc3spjCAET
bQRzC4y1hhbbzpe7f7whZMdWX3NMSTCv5Tk5gHWrPA+1bmqSI8q+1XGmL9dWR+yOk4kqGkwjD0hE
80Po3NEn8XljZsqNczsGkQerMk9l1jGhdyrUrubh56lpvjOABNbxz/zjxf49z6IUTFTQBjt/5Cgn
Ldo6KMEu64p9OC87v3KiUv9cAhC9K/baBhFXD7+JKO+d9jVS3MVoC1w8t7N5zZK63CKzdzkS+nmW
lNykdNfchx/Wcq/GsZRX0ma11UAalg0KKurk7S25GV/b2NLKBUMfYMtHGmqCaICmjReX1zin0HKN
10o39lSuY6IKJBCT5Cc0dnklreljNgIUtR9SrAm2Jtx8ibPfZutRE+SFTwqjWD/xJ9F64QjxPSL+
eX1GNIKsYMzN3XLn6dFKiKT35XYKCpWlCGz0FYI3D51BbdeNVkLBU2WnGPVkfYj9LoNxTctvQ/UL
LKAjMhS+TB1EgE/MBEaYsVzLXNFihPLwS4bK+OZsGRKvyyv98QrNkwadOjbwaTMqpQ15H0WuIp2Z
GGyfEwXOI11JmkS+4+hX9LCiWKKg/QLVn5vNhFXy6fcXnpqi49N790D2kOClEFjqQfjh61WrAYb5
4fSFSUEC/x+bfIsGHmJlYUk4j94ZQZoZ/N6nCU1wg3F2+UgRTOJcpFZCXB6UiCDb27Ftve8yJo6m
LAApsKgSXWTVqiHmFm48Rj+HI5x+64GhvnM/HESiOS6IlqjRejsYMs4YH1g/SiHVfo5nq5J7Mqde
IALdP4AC+sF1Sujt04Ieec1ad7EYUUkgqvvC5/3VezsXSnO9ZsAASARJcqOzcNPfLPhMPX1ycSjL
TQpcFjdNLJIZasHjXVn2ejp8Y1zoyidcSGJt2tr5j8lZq5MCoWbocn+fxzUX1ipPU71oimbp47ht
YcvzLKLisQNfBfregkPBa1nKpF9w37AJLrxpxta7vRKSD+kOIoUGVU2aU1E97zpOGBWXzN7t2BQa
boloFab9cdnAul7X9xZLGV7aHG2QTtXvrwu8G74vlLF9rg0I7Boa7ZY5TxwL6JykTY4h2yqSK6KK
vuciTg0QHXIwP2xGTyv50a4fhzeekl5/yaEV05Ii1wbfISMoraRV9458QICJBx2eOukoNoAnyrJk
nJl69k0IhIO94hQOQeCmQquOQOOI3JnL/EpajZGcyDoKQ3Zr0FP/V0UEmG9jBXZQswe7fJIgUlWt
zvDMNWTuvfvR5VvWVPm911xjzDgw2gi29bZ3LGe7Qgj3ey1SEmKvescQS+iljaFYPyEfRfovwDJ8
GI8Y0vdzKO+iZWXyb/lw5q9HCdjoJubhkrY1RITWVT3lnKD9b76nHB+lE1tw2UMlK9isHYUikIrx
/zHUciYDiyZ+6BLjJIea4JtEleRUz+8EXWhRAAXjhx7+sWqQdWEdEA1EiidfhoR/4/ZuKyayoCid
oe44iMyZi/RfoiGM8nH3NTMZnKqcOT+OxB3PE/KUtA4Lj4xsrdcFpBFlGd2yWXemWu/R/4+U4ZKv
3coXe+7SWY0ZnFlkLnHT9vyufsM4CfQaxK/9QLXQ2P9psWKR7LIOL7ARkI0lDsp9XIZ2dESmGwD5
bCumtYeSEQFnz5AzPxQR556rwuuhBwV0R7aR6l6TuORy/JWt+f1ckXojCOn8og3X8zIZwOfmza2u
41Vvov6lJW2TQFKF/CxunGK4PVS0oJFgiybyZsfrZlA9BKbIpaDQkSeX7fqm/9X6JZG/PuRnCXRn
HRge/DDIxTYOpgfHaoSerQhQj9fIAyIEtOx1xRf0L/WIkDnsx9NVFqrsut8gQT9YN+JwuMulF2Lh
F440GS5NIjIn7QRpCsfCxGni+FG+BfA8c/GlT3C7lF2exciBhLezK+u92rjbwqSYCHEkjZRU13tS
RrP5a3qealBDauA/sL08UBk00LVWmunkZL6zhBke8QMDboQCpK7raoAO+erBSpaEGeZ78r08Mb4L
aUeIugDPKzWRiQ5jKz8FCMK4CU3QJdjDS3WHbcBXpfGFTHf9vUt5YUOEULID1iEfOaKZ9MFHUtEx
D07viQhbDI7+BUaNtA+TPxl7pSZcny0H+E8/d3w6Jd9pM8VEMv23IFpiOy5opftoTVp5UJR4H5dz
tO1gMKgFi8efjcjQAujY5QF4zF3exHkT2iN8IrPX6BKAgH66aXNtwRQ3z3E/t1oc3W+ZXaZsPAR6
oYQRsK1Ip/ZmPPxt9hJdfTne3ThkD1aoo94VhE1LcLsyTgWXWb6kRueVly8DCCuJ2SId+r+QReI3
1w8TTrEKrd98Xc0mX9BzDCmAQrJ1brGk35gUAMQZAbgujhAGLjVoXVL8H6UrXp2Jt7Yz3ALaM0ty
vMTmduFFv1+4n69NhwiPgOglf8AsXXLx7hXVoR72KFYEIjoxtmFJHdwE2YoGFjVrhZ41x8MVVQwP
Dzs5vyXcXOXdAjppehiMFRMeePCzcdFhtjPkIGhlFOf8cJvpUuHUi7P/474pgXGKl02dz++OLSJe
1viKEj+SsbfamdNd4N7ZLf3Tr+VfZWoPZpV51a/AEB+zHsbiuscnI9NmRGg9es2G9qIPaEjP4EeZ
2aDDYAQ2GAoyiFsnjVYGr/Kom6c1GKxncMsconbrdENIo8poZFwrzoTV9dYO5ubO3w1Pud4o3fHE
PWZLkJnECJTskNQr2gi9IehFFLoCSKdBVCOHya2cKviuL3+4W58YPCwBFLUspf3YY1dJFArTLLc1
ggWlxkBeltBhDLQdFcIe/bj8kePBorv4OSshwqDat9I6hqQQBO+WvnVErXgnu2bKYe2MaIU2QpOP
aWrdOMZM0qgTH97z9d1xmWpqn88r1uUOH1h9XrROjGXq3+8ryPF3k43F2OWKbBfvXtUM7FyPBvw5
deAf5NXhLw4lmm1DqA1DPB6YreDZ4SdzGesWzHY6X6eiN6rCAMjwBiHHQslb4G2Oks2FHm8UT9e8
+qMIjcdySuoQoXua35XiHxuYy/8sKUPsvw6LiyhpaiGttU47FOPPz5cnwGSEVcKVYo6DRjs0ve6D
TAMIeF5yV9HHVayKcanOVo8URqRUQbmylVSc0OjYydmrp1s5AzSjMWUbVgmMkbfgU3uwOTZqDch/
nWVdLfqOgKoDMUffV1+tRnQ8yxmOnVQrMxqlcnKhvPeLoeaYNzNEYDtM1Yx4iIihrHGW1PIvXejf
evmwzGIH/H+7ZP73tE2tfl9XHpKFgGuNwTjFknP8d10blOwiNtBlTPfa1a0GQSRHk2Qwb6JtvCnr
zEls8cQbFyiFAQJbG/b7i1wSZwnJA41qS3vQK9hDKaPEH3IY+tZIgjZOalLTBotV7N0sMXf9DzmQ
hE9u7/31fUVYAHPD6PRlRWyJsEk+tAW6W9h14SftjN8AF6L3cjXD8shFFYbLGdJBjvEU67XFs7LP
d+5J010Hf/ys44BLXrEtpLpkhNGRGfBGCUUL3P2lsFoWar/yQg7UoHiHXHpeztn8DkJq9z0MlfHY
AmBX1Y8IrgAky/kGmCKff/c2LN46Qyte5agTWE9F/uL8vGv23cTYgnqa6T1VihOHrpZAW3AJnDJU
3bptZOCz6Ty/uNA/CS+zVvlW0LQ4g24y688NZUQGPE1421DHWQ2j+PzSRm+Ij2G8Sfflta7QW1BX
HusTMTfeLYtJJ7kJi83eYx15LlURowFz3sHAykJRqZnptpqBTEEW33biAwGxgAMW/PVEPmtuuhcK
tLyiHB+n2htU/CesLhVZkDiqIt0vUaKiwyKNwaKr5EiB9OwwfgM9ccEilD7arLCSlb73VYFCoVCV
GT9iXXcycpzYMvAx8rKkKjYIhS317R/Pgv/NA3EFom4nyFN7L6ggQidH6oOxuTarONV3D/llULod
LIlSlJKQXi8ahrRJPmFVGnDr6wFTkLZ2E8XVEslrRwmBrL9Nwue5KaBO1jXGMV3Oty28pI6a2gaM
52+5nrEs+oThbecAwPprez8/HJVcxl4kIswDFfqgHvKc9mTE2K/QsTAehSh9ORvRc6HalxVaIkqt
9/OvGw9/aCIXPjzU7X2WS6I1A/V5lCjwfyzE5tY/tsWM3Ak/g/BLZwDLXnJRB9cK7+UiHh5pk4aQ
V+IVbwn2U6GFUBURqT3SKO/JTK2z98gTxxIqa01k3RSblOaDPV6rFkp0l74lqMp31TgRtacj/dc9
RSbWdRRajrYtoRLsbj6La57GnkJ+Zwv4wL1fzzBsFIWN1PcbEGbKtNgjVstt9c1qH66RHiqkfh0B
hIdRkYRJSSbXPrtk+8tflfShXdI4yU2X4fwe0CfIXQ72RSleixcg0texoZeK7AIp1ghVxx6vfS++
wr3lDecwl6W4Lml4MXdQTOZMJh2PkV9elkVGO4boexPJH5MpAmeGIkQQsSI72VDhx45W3uLOpeH/
03DZ6Rh3Wgh7nVhguwBS0xgauO8kb8qNCp77Vys+X0eUCQj16b8GguKlzvmMk+CiqSbALzwO6QZg
FvTDryl/sXJj/A4vH0liPhjypjN5vQf0dvEDtSKr7xM6EQMFF2PBemkKqz2b8jD4/m+BhXiVZc3x
RZymJT11wSZo7UtQt4DsRTQtx30Yhgi5gcHOxDvfVgAH3ARVTAUNzg8xd7bFvd9ZmT3oAns5blaa
QUZPimaHQxbEDJLe42+gddpJ0FKchynu3yVWBo9kaweFMVqZDHWVt671n4w0PHu2p2WgDRQmAAfe
2jUB94ZHYMofGGzyPUIZlVfFkfvRyaapXyzSxXKPQtfI71okXok5IuVeLty68vyysCLuCZRmQtdi
45ncDvFy/g+RGGm5ONFe89RX9UopMf3XNUJaoKCjIM+/gTQG9GltWkO/g6yzDqUqzOBWaCk9WFeY
twmdpvVTqs88tENsXMuYRHTaca09RbD05awjPIsVa3ixic2YT18DfiKB6S0zNqex+ExUl5n57aAM
7PqnufgY4uX1xCQ1jxIx8WJjAz45MiGKFK1dmn3B+Wz1qRz6RxWWRdPLJ9sSjl+uhbkjbF/9uAOD
dsRt7VnRk//+oDzjwABKbGPk1neWQl+DJa/5rH9NEptKImhUGhtjLwOsRvQZfE/WWACdo2VDnqIO
no2aEX7CwQ5f7QNbg5/ZlojvjjG149qPXJhnT0IxJdO2bMaItx2cf+n+QUhTy+Fygbir72+2WI6d
yJTYFi5sPBmNVbCoj/r/gmY9zOMjWoHYeAoj+iqt2KBGEq6nMqkTEhld4XkAUSsYcT+Io/GtiNUx
ZMXAUd2fJErkylLimROYPKSiOXvFypXnaXm9IDC2rZc5dy9OmuZURL+/o2bCtsUHKX+FrgndD21c
FiRcGYpLTTBPdlOvx4jFg1Qd3hUVpZtROPiet4p1OdLPbRn0W5ILYnL1xowtEWdddveZi+HvlckR
p9/fMaO1K3+V60066ItShidFAdbsZkIpFwQZ9FOuhPaSLQbnjNMGtUlRnTgAOgYsjlXTKXOYuh52
2Hw/AzGLf4T1317G4k+qE/RauWR+kXgyVbg8+IZrhe09DihhUb5A+NTg0G+mDeTnmppeCnFdFxRT
mbmn9MQzmlvDp0ZXTByFZKca+uIaPTUqN30DEKudukWHjxi/N0tFXQnbkoyUZvAbx/dJnc5oA4sC
SNUfs13p+WnP+MezOk6U0DIYNmJVKPsXmRXhKS5neKRy62WxJHdRbFaLX3ymQ1gVZSxJY4fjgLw4
s2AklQmxknyW64L6AY3vwV7YDmsCHTFXsWeP4fMKrYQgw8VdkiXjryPow2DxCaKsRN2RxExAqrVu
JYWmOK3pJtF8keNcYAA7uXlBWPNtaMrrwC/OD3br+jZ3Jru5aYsfLwIwaS9Ql55+22e5m5HLQVZC
wnqzSJW4T8m6VTJ/ESZXf2zM7DoI8ZF5cQy5kfWiaxMDUqNytz7OHT3jc63IxLT2LV2CE6E7Q0a+
aGhcYIZxPZExhNFiobSg/NXM/m65CvuVxLuQIeNHOpOvARfK096WQwpBJy3Ip3oUb2/T9HfvyX6y
4lMWNhduAxZ5xRaHhD/rl31wpD9M3mS79ejg2LzQKFltdJJ4p45I6Mdx0hCmLtSQr5bf4cNHIxiV
OWLcggSmny3pubhvHN4nC/ZjaSV71HolO9Jq6k/tRf2JW7F0mklIbKX1fMOU7g/xOixOYFH7DmuH
4AHxVUjKRZjp4ZWiDqPwfMYcZf5TCbaX8jL+LQJ5/Yaoc/UBgUNQ+cHI90bUdDNv9iCbnyZeJ6ix
0BrkgHF6f6cOYn9kWxBsFAaUvAgFAUYt7RN16wLZnlJHw+B3getQXyCagilIZFaRgD/7JtwrF9Ky
lZuy3TIAde+0ieQzfp129yOoi3fd4sGkmwGxVMdEHvjmqnW2ULHM+HvK3YG8fdadqfjuTH8iesn4
Hbw6FndZxLBx+bab+UAh7pTnKXFOBgqtbCibTbplV1+4+PdwBvmJyMDgExG2/XG/Pp7li3HzPviL
m0eoRlrRDHAewIzsxvNCcFYQ8/dbBqJpEPBFuZua/+rFgkM1Yw2QXEFpu2iJjySES/ktVNBVRdNK
FlsNbZBnd2/dNMkeakCQcbrOjKIEwWXfTRBUBDQUAZUL1CBp78x1IYISSUwDbeDtv+TFW97BXhjA
gbYcb9I3fr9e3FxAhzHyQAFuh++YUjiOjmpHoh3DB3mwwgqfih1WAlegPmZzEkrOdLW4za4H/UOl
OnITLskYydjPh+5Qw/qYaCKtu7Nm9YTu7Tq5dy+NOlK1ihULTMrJuUZRJZmsTQ6y8F+QxAXM3USe
bmV2XBlp6NOmNlwyymHLesMdg3BZeQhkjEwvsL97z+Ib7II9WZpEDd95zkuM6th9G3f8WyJwRgrU
5f74ZzDyB9tMoZUqW4+LxrkE6uWjb32oTs/pCSqIHwqVrhCu8i1WwtIW56Kp9Wa22tmyXe4hnbD3
aACKqU/XXkMxd7OFWlUCSYGrYPqRTI6E1pYpB6d1ozMp6tpuDjqvpCTWtROScSi6kji4njYgr4N1
pRVrjIO6NatpaMi3hzJ20XPsjwMLlCk7v2jzcx0u/RuvvzFrSWmjqkEn9EhvG/Cy3i2S8syxQmcS
TuSt1uQaX5gyT8ohdwWcQtILcCw1cbp4ZEQwzAOiOZpN10PkxWJJ+Zx4SOBy4ECLVOHtRxzAWkOR
2FF/hHvjWOCArNDykkeZuk3A78cXIfkqNXxi1GK/kKQ0yK+sQcfa7Ww+70ieFcC64bPG7nhypQMj
2j6sChNR9RUbRek83YfBVs/28OhkbB5s2TbMuPw8cWgrmpCu/WtuI2q8JjWB9k0tlwh9fwKloWJF
NqXiHexA9VfRECs5AD0iXxvE1zsL/ewLck9HzwZxcvDAjU1TltOm74gDI8cx2wCuB1HC3tI8eTo5
ieLrQL2Ce0WGHSGciQ0XhfZrCjbbXWbou1SbDYMljr5TcV75YQubGaXxFDA7drGrMVKGKIHfc8cr
EArebvj9z50gs6j0FUKx8aKGciJ4bdkOoiFvOE6wi6ib5dVfrLCWPr0aW+SHizasq5n4Sw+AApgR
kyGWPAeGciijpVcFyI6mhd9BzIn8Z3tz6Ez8WZ03jm+M8y2sTyr1X6VD6WTqBwiY7/52FX1xwY1u
PMibtEjbm1XSV3aIT9sJv+82rXlmtUSXFXaR2im4C1c1KvZ6HmaT3DnSvWNvrB8biF6syoP8MCtO
ZtTEFEtkqret94arTQfRfxy5+MGX8TSrVPWoYLVj6FGXoR3UaCT1xHCpPaG38PmeAONVQwTcxDk3
2o27yu3nU02lt3d/XzROA7PiLfgSbzb+bWufgwF6IRHNIWo/3GhU2rzRnoiU7Eb46KuH0jA6yf7U
duTo4yxej6IFLd5w6xdthyI48hQ60pwAOKSqmwu+94vTC3iimoSN+84P8JcQ1rwBN5Y4O7WGNFMk
6CLCBZIzcK1yG09XEPMb4GlepmaHrQery/p8FQLgd4CFAhy2wNHoH9Uz2zZobECUO5bJJmLunj/H
stq/GKXTsnZTedG0L/xJrmONSPsDHl98TRdH23gv1ti9NR5jKbwQ/A6E2ilrtaJ5cPz22b3rqnF0
C47n3FvK9MT5Tdz/FgBqbAksLAcRCv9YI0ltcfN1c+b2OWa07HplR2s8tuIARLzsXXYuXPZF2Z10
DXVO8nYJ6f4vuTHJhzKVU5KzMifqVm9cQW5mG9o8BrlGK7gXj5b+TFeO1HBKpz7bn33Cyad/91Ub
Gr3nubFj0smPBa6p4YUjoKFsBnZGRUKaLjpCrjc3xzqfDLBFfU9ytRnjPgVgx4jtg6bwPyQcxUaa
qjPCMfsKu3V3kWnGlD7Vu2GEvEW/oZskAfqJOT+aGmKHKwx/E07tekeakMx+liK1NpfmF+3RUfUD
yeT934faq2uDhyiFyLnyQHkk1Fru3drofoMNyp3A9EwCTue+W8EROLr+C+OK5+TPQVMIGcIOoY7g
iGFEQ0xoTCU2yuWRhKYhpzhJfww0BE5Q9917aQu1hJi3eSQGThSZ26fdTTsFjc9G/TLXvSSe3mx3
M0NMnkqsc5yjYdEnoz9Uo7vkJMNIam1Ia3dTuP64QEyWri216UYihrTBvyJusMN33jCDgEJraOwF
/upIHilAykILi/XQVml+HR8qAn69xOJGOB86ItuNjpto5w2pf665ejikSiFhqKBtecHHsLh9m02L
QijNG+9GyV8/5eTrabqohPV3zEf2OZa8X1u6r5NZIldVTPBn9PZi8IS7BnB019dcqYiCqMrkJhUn
OOXWCRE3KCqRc+9PTcAJyliCr8xiqr2MIFabxyrQh4FgNw8luDZsv8uVA+rXLYDV3/ic8LsMPjhX
u600XrV70RceajwpYvbO4IQkmTKZ+J86ZqVsNp0povUCrKB0xteF7GgpswjENpa8PWMpu7jOk4Tl
ZR6HKtOT7EP7js6wtd9XsGX+RiqJ7EympCvsLJ3C7hqDaYEdRJsiqWfojuX4nqMHgTwkNC24SCtN
Bs5+Q+BwdzFwf5ie0rSUxC48VfRes7j3mWkcVarpf/bEsHBRnJLeCxFO/YrLXhr1Zgt9ZsIG6l4H
f2LAR/i15EG5/04TUrXwr2HjVefGDgPZpLJuZJN3pbjxs13yZFs9v1+LlIhJaiu1P5Kbeg3055ea
lfTIC6AZ5uVhU9JiVTZr5g9gG0/i/Cade2af3numNGeuMfN7WDtjbf0z04+0/5Do5y5n65hjBNHz
ZiPWX3DQMtPadr++8EGHnykhzomxC5QtIGZ7R4FhrIwqdOngZwrYSmajomgLF3GnrDO69gcO1D11
qQ3Sq+CFiR+jqWHPNLhUseyPJw4uDhQtuROoVpssJT8wavoNlr/uvcvr3BCezRshS/OPQfawLycT
QGwF72gvaxZmZ5ZETz4M214/Izn/RzSzfGIQBBoFNfCPu9hG45VBXgzYPP2QHg44z3u21RwNJRUP
gIrF0PTulH9Nh2i91S1QRZtE+w3l/zD4BGzl2P0bBrHuyuKod8qC2NgTvo6DZtSpj3TcCOdZ3VMr
OO1n2eVEWp5/YyOg419An1giVINMMbkfXyCxeYkZ6hldJ6VKXC1EVzobPyMgrc5iAlT0zCBLUgDD
lgF2AwoFEhIdU9iIGYYs/6GRxcVtNT+XDVW9k5ptI1ThcDtJEViddBKZKdhE1ysWurj59zsaSUC/
+OuSEUnOwW0vW7y76A46r+gJZd8Hs0fHkLHZ3SgSL0K70NcN1Cp3GYLE+Ko2czpEO2kL/GCUs1gY
FO6jkHiFerKBkawlLyQyjNlXtjTLVKUQe9EnuXa4j0l6ONtrs0E2NJIml2pqYbMQqycdzJs5Old+
sqEglbuUxq2U7e+UMYQeb+PZKyZ2YMY2gMEBt8PM4hau0fDsMvUzb7yLF5eQy83LgtwYBkTfQPf9
Yu0psNBa9USgkXMjPrRJ9vCAIEt6Q1HylGPp/u7vDceOTgpZNoOQep6z3gP2Ot7oh1ln14yxzAkQ
CuDsRtdDJpj6DABsvAQOhaVUrDyZMQ9EZOv330ty1ToZvlIxvcuUyRYAHqNt9sYH+QMa8aCnfSyE
q1kt8Fz2Vce+Rmg4d4MhhJ5IBuvVvk7YbGGHTDroQPLWUvuV9rj/yQVUqvRgqvBFohD6KYya1rPx
QVC4tbGUhKtg57TlpRhsiKSTfO0t7H6t+w+fyCQfKN/nnprhbI6QnUFePUmaxEUD/YM0gxip5hlI
PErc0YvFw9ZV1rXYJrV9UVAgoidYzZPoTko0Yde0V+1wNTEXBVFPXvxsW894MfM878ty9qTFtkSw
MnXxHzrzchyVIXu07F1fItmHVrjGQWieY0M3LISc7q2B56EAQhkVFu9EZDZvi7lHIgbQ4sHco1ny
D1Yg8uxyJwJV/mg7EBfDaeJ/my0K83RXUG3tU53f/R6O8bRMNwfgauqSfzjn5WGrZj5Bv6MUgAQa
LmUHkJvFNm0MzXjOYL2a1/VBQmdgUuuEpAhBNXoWX66wJj3u+fFRtnSKkLGIxVoNU769HtmZmQ0U
MVwaLK8ISIS2nDsY7X8h/2iCIxKlrzv8hmDW7dC0ewO3MLQJRU75KwGS8qcQKzWhEUr4fMg4wOOi
erSzvLyfT/IDIulhRyGOFg+vwCCcqIdQ9F/hUgklBHJ6GajBFwBNDFNFs1Xbmp9WFF92h6kAxtkf
OXwvpNNChdz02Z4gEKIGu+LE1C2eaNdBGetdZZJezXTjGtI+DzjosdMobn3eIePycUTdGeeU9JiT
EAWq9aa7Iw9RXp65UWFjvlyIIyqBLUNHLOzYO9bJk5RvMZbjY+f2RNvdTjvFSYg4laiJEYodgGiw
XZgHtqmU73baaSRzEYrpZqwy+wH+zWjtLzyQD9vlmVCoP9Eq7O/psfYCQKE+W8pt+M9zSH+/Hbp0
Wx7NTEFf/Cq4X4Yvvk7EjzHrjp5VTDuocJX1O8NZfvGjYynencaA8LzGftrlaT1NlRBo+lte/lJ2
2omSZvv1+irGXM2P+6WHHIQcstBI4I1NCP3g3Sxft9spLD0HasgfjAHLLWNrZgfRcEDbHOv17TYu
1gUOTHjkPzWQP8+iHraFAtpizK0aigRZ3Jm6jvNjhI0jlfpNBHhAWNj/cLJmLbaFVR8Ww31rG5+V
zUxCZEBUPPtTHixFlw+3Ay0FopSurmDIT8O2G5Asdrt/0jlOKNUkuTquWeZ4MvTtsOVvuLax/rs3
CHv7uWI3kwX/GRg6H8jKeR0LEbAJtTuoHke02pgfPrL26EjKoDESxqCuVKZmZs0VWKnvWj0CAWZ1
LT6uJFdgfOsgfPTNH5NgMT++Dx5S5SVwDaq/Sx/atp2a8LDFOFThkGzvz//iC5i3htmAnTUiFdGS
yK4lwmZ/cGKsnh0yMeKFg8u8YVoaqA2mb4lgAzDKBGFQg4EIIooyHRM0HTVilN6YoTgEVdcH5ph1
bKZSHciRafsAG19janV07hNc0lC/6JNXTb7307JSwx9cursHDjybusuzas+l/Th6dovJw7hJDITS
MgkapGsc9pxcngUpdQrFD8FeRWm1q5N17jIQQ3G+ZHiCii+P2nMVYWkEE8yIoonJotA6XuQCeLIn
mL2xz604Za3yHjy7hXHC3cZn+UNra8eMb1yuOcRcog3qSbUprP+t9KDbNH7gvvpU4vfbrXzgNx8l
5z08LOiTVjPV0pds0YRBNp1U7AuyG0FXdbPxH12s+LPB4eA7YLbrxDQdgv4j3ztM7otyxZdi2Asy
TZSKC8C9QUZCHKDXYDYCurdcSKUlhxpvQ3zcnKIKBKvEQ75HuQeibF1l+VHi0Io7fOB0OTdq66sz
XNMCch+FD0u7tFAvW9kARP5eyyGsP7W7QmjwJZIew3AfBetMRjvr+ne697EM3K7sID4Ujg0Oxm7V
Nb97I8cSuauLzFcp4oeHZEYrPZGi1Knr7MtyL1Spxx7GD7LTcMJEkRksvsu5HpLgCXeEvULgqaTl
/KrKZ+rz+S8JWXhJTHXy3LtSlc8v83vZKDxAOCHJjayyehM+buB548kK3XsjDQxxK1NtRhrmLwdX
9W4r1EToVmF7nqc///6yGOp78uKD4GSv8BbO+/v6pak/bajr9S3Nv0RiIizDbfG00/9yzsq9+iL/
hIVW8WTY/SFn2gDNnFgbAC78DW3bc0Yb3bh7isxxS7wn8hzF/Rre19ct/qHykYcVFV5SWWAOB44n
48oqwbiPkiY4OLm3JsdQ6IROj5GUF+sUmPDYA3Z5JCyVF4cQXWoyzsCaXeFI8dLJwT3tiMd4RhB0
wD38U8X+729y5YBAadkKLtN9/x7hcoKqIzzRPiSh86bBBPQKD6FeOQuP4VxUf4a/2K9G7CkSGiUk
s/+hrC1D6dltSzx8zd7hVTXjeGpI4CXdCZlv4glmjeGex8pwWyOnyVsw2HTmHaiW2AkiD6DppkEg
3kZVHK041K9+FPFnxLLo8wgfMoMrcHzEPsBcDXkJN5KhbGYCBKcLkm0CrdCcIw4J5tD28ppIoDcr
2bRA2RD/dCnIxTYytqFYuci90zgWiy4ztTjI+koPq2zzpWEHpTeT9BucIGywqtibAZp0cX8Ge4jP
hAYtLXTnVndDbR8WuD67fQUvK4wLBNrKo/k5qITMN+VJhrBjBZm9A5LKobCrfMdukoYJQvfP+4tF
BVDxf885iICmch/qgou8VLg7f+RHQ9GgNi9sI8yzS2yzlaGXFyx8lRfCTL+9/lFrsV99MrkPn8bv
1YtpCDP6/shmMm7oGduDFK0OXEfVqQx8tZrHrGsxs5uQS2aoXdwSkxh7XxOMgUpoCuZgjPVfN5Lx
BonOeqppMlo2XG4QcSKaE8cUzilEgIa5GzxFBmyqg0ifKpqupDIzfLW7vAlZtoopdMaZFaLmXyt5
8E08TBUr72mxEQDCfDpU4BpaeF+vYwhjvfIYatr5eyUn/cGmikvTokBlyCeMNOWBoe2C89qVZiZp
rhA+esVRigv8C6r4k+VTP+eKj2PcTt9O8tylqCyiRTCiOlk3sZJB4YKqdhkJYk4mwRaY4EJ+1zCI
9lYbt4LwN3jsS+4Op4K8d13lKvxvMRdmRvIpBJ+ryMZENXv1UmmRvLf1HXI7cLX8VSIQxsmEnyh3
cg1FAeGRxXVIAg5NU5d1IFDfG3XzkaSdkTSCWMM45E1/jGY412zIb0QwA5onofXRfN/4i+DS8/as
kX3t9MUEoVoXS3sOqx2fpi72swjqYI8Gqp6sYfbsbWUCwOdNU18rxaQHTorEBrWi/zgMIEIkPG5w
vQLlVvedrNoumYbJLvAHELcpFyTMgDpBypXZRsZlhNEejaoERvrfrWBJ8wos8Bh4WIMhVKrt6CvO
5esC2Bbim830gPlPvK43NSpId/Iv+BljFFnQiMdiFrYx74BeF5ln9e5l6xuptSGIN1wScMkHkhER
+DOEf0JMwM4fNYFj38yCGeosTtHUkJrYpqiDCKUxAI8zDybZ/Wya7ugo+zzti4ANEOh+iehajQE5
gvcp/jw07RpZEcfoQm6k0QpcOOsp+r2sTqp1TO+MZA1+GqlDF/DDXFGYgWqk3wM0P0j9vhVtjieI
SvL0wQAyAzZj0vgnFqJA2L4mJ8zxL6z2CAOQtxNE2eUkS4Wu7sA0ytlT5IGijQl38P/6sucnaiQa
aznS37LjH1v7nhNQGHasEoJb5L4EAtWvZ0UWBKfHVZCpL0wsc3NfMU+L8NnhfJ2o099cgVOptWFx
drrLwK+2Clzx5XRfV8umBvzMwPtdVxSmlqaeCvuP1K27UhTuPZVd9m4nwugRqtySZ9RjCsN6lQfg
rThenJVUBcOWlFBTYta6AGF8DCTL7B9e1fXng7vwOjMdS1+R+sqXRJ9s0sKyQEa6cAhcoibBvk5z
4NhsYiqdtmmtTwIcojV8JKoTVMki7n0dsAFthWscE/bMNHK9Wer2/hkQmR3MizLhQdyPUFK9s5sd
B5lr8WA3M00MWVQxHJT1MRDPlQuO35ts1aAIUcABSaqMYBsSPh+so9Tcb77WgRORJ/idU+qwlYc5
fNa1VoXQ/dshlJOr1aN1H+0YyfN8p8IklFLBV3M1gq7wQqfjkxPvP+MmRwiAaHqHOI9p7TF+0rAE
Seuhe0jq/290W69iUKMV7aExghpmiEWmYsUlaGDjkAHpaJyU1swzO3ib8ZGEo6Ue3Z2atyMx0j31
88FCKatnwABrsZ9C1rDYZHj1QDNgwnv+fhXh5H2cwHpO2xWi+uslB3VhZz9/CxN4ctJdU9OzNTe7
CLU+E5Nwb/QOXgeWOETUdohMlA8moAms5EHsEjQ0wABI7KaWJdg6ct6yqErJ3tOzSaYjGt8T0N93
DkNlHFQf60IlPuYFQSDVIVnSEA2EvyTNEa1mSM2qIiCbqqzxWVOPEP36EJxxkvxr5Hhupe+EpbTu
oWbLcYBK1DgzGufGs32XPIwAdXYLQJN0nd5yNWIgU8hvVRjgXerZPmudOaGaTVrBf49OzaDI+S6F
p6SOtpiL1Tdgnwnc7A+T031as8eCXYyL7dG/AxPIyR3Rl+pD9wQZeaENF2pjmhO82ABg2kKZxPfe
16enH6/SZ6ExxOphYBVHYY0ZD2qNC7utqQFG/GEeBC1540uBwhtMMdaR8/Qre+t+E2YlYRtSv1Ra
v9Se2FJqqCLgXNeDAwB3YJwlukEQ/0T+KYVP0PEp6dkmhaCh6qtJ+zL22CFk867IvuUdrpdKBBiy
DXT1uxLACQ3drcM0c7Ttq/lpSP01LZ8oNIkm4gJbhbLZxSveY8YOX5YPbtUslACXMw96Olx32dDQ
dBUa2uqR3CajFSXbYL5MqUfHMvTScjvaPv3Ri6YnJ6WAeNe8MWLxC98PQ7nN5F2lHh1yRFqyYiQJ
+5DMH4CwWU4LIwACNOuJPDCXk6MmqiYT44pEhLdbs4v08V/qb0KP8c6h6AQeTDFZx/l7jwIpl/cP
5oF/qUqlgJgiVnJ/NL6zccakfqT1II3zHNmiDgl14v2K+PR7tYQLEL0vk08XmtFvDU4H8DWInJVn
A0uKsU/nqHYLUfEgpUliPgCPw3aWZL84qD0jjf3rnx9QGhdLmXmejs3Jb76PlZaJXiRs5pD8x2Ut
/vRhBqcM0FFuoeJWUXm31xduPceirMbmMUBv/zXLwLlcZwU6LF756GIAFetkNdgBPzI2fE9qCc7N
EBlRV107yrOC+iQI8N4c9q4pEvbxUnv6xXxmKipGkhpbpwDOJbilsmX/O4Z7BGJTtaVl+NSCCOz/
tRwtNzrFa+1oFOJm7/xQVp8xy8c8dNRobf56KOyhiXmNb432JFTWkFhNSoDQ9WmBbbqwOg41WotC
h6K2j8yr7YnZd2GWurJXdyWyd4HakdpLAmY0YbhHF/C1F7wav2rDPp+b+NKJnFw4fqPAeWcjfLB3
NSzUyvlp3t/DV9bq1luKeb1cTKIp2lck/ltfRZ0vdiP4LJciDQMDw4hVoqcM6O5YQBYbv9J2u7wY
qlMWVmbxhRbbgn0DqHMnitHdfVboZFzMzyuIOcpzF4W+rSvnNaoPThHdJJiilW+QTQCeD9Ci9scm
gDJ58C/iCmLs21nF2btGw2CxuALgnsXNPM8J1zYUV7VTfgJz9WiaPPR0u28rD5G7CRaX1lxJ6Tii
48XGU1TJ1PfiDN3UPt+Dddz/91/YQIfyO2+ISDgW120SdAiWja0zRLyU21i4ISVKGleTz7w8hr6o
Re/4xGMaDFjIW4+gIsdDOw7N4UdEV6Zvi60CBu8af1IY5ZCk8yeV9owhtg4NMNJm4SlMdBhuKKRj
MRpNRf2AYvLe6KueJMeugPOQkPOvbO3WNQME/UUEKOWUcXmORdyCDA+PFWlG5Aw9bklfJVvl9kTi
wC+QeQKK2MFr570rJGEDzatMuRtIradhy9NZePgJz0g6CybiHsV9Ez0iSqqxciU8hJ5hvwJ5sQLh
tHzaAsNmMwKhCqQmqqBD/YQRL4FvqnsQBHHUQKGac4b4stP8rGezyKDCJbGhlQIbWphCkmRrfFOw
+yd5CKXvTiHPmtZow0co/MewU3+Um/QiS8x/1KALa7J8ZPtNs0vvA8pKs4jqIxYZLvUS+SReV4qm
EAcG4fbPMyInEcmYU6Jun62gPhwJlxkSK2tZC0HQ04uTy53DSNCoJ46CHpsT9jOCPj5ykhMTaAKM
rpEKioDSFRKhuHCroqRa4F8sh8OUum8vj5uTAFNNiE6A3TaiW7pkUdL1dT8wzbFNRHHEMjsJE4mf
QqgIa8tR2/RsyvmwWUfAWCiuxfVTbuLLszOiULBcbrpmm8vJYAQqzOLSkmpW7WWBRwwjgTDWjT2+
i+cBPY3rQxABDrtU5VTs1lP9/Ocn6j0j9eiZH/fLD7K2Rqgc5aIuqMs4hJTyJnT6sR630Wb/zwKh
uUrkD7Rnykf0FO1aWxvY8OfIzEcaOJJYZZyWLow2pcDUPqxmD/iKZ7XASKLVE02Rx6dQ+e8QosW2
uyavW8E1oN5IKoy1ANed/+RrYvpvhc72VIFe5iNIEg9ptHwV6gX5altyzgbziZWOVvZ9g+Rvi+wP
FSwYcHP6vBHJKCU5GcFX3vmbcMhJTKh/j9Pft8l23LiFNDcNU34KaV3Y3isoOfIt7VsClOz1qIYN
mj1O4XSEMvOiqv5m9n67ewYsMrmWWG+dBq4tgAT3bqUZR6Z8dFxPdL/g4cgOJs4NAD3kZjsGMEj9
W0YTwe4SnmK2M+kBC7aogGo8l9Uaa53vszyyVgkfScgn0BzwlVmsGI2v4l7nhu4bl8667Hj8jqg0
Cb7jOE+PVNw/XVz5aGfAJ7dn8jmvYGOUHKJQIAnoJj83VkniCmO40ac1akNXySaXMbsd56Y9HLG4
RUMivct6Wcpl5kTh+NM1+cU/2+qo790eI7wyKON3WzMKX2x7ah4lp1IuGOG1hsJ4jYrB/72QoW8f
Ho/SpUgMVQHoIZIm/xU7DFzEaXgKA9CZVyjVFSPhiG0R1eOMKXadExf9le2WiIzKMgJcfZNaXLqe
TL8LGnbZSqIsOPVzD8kysB3kg6jMMdlku4FLqvLsgT3q/v/Zm1F/3y0Vb5th3jFH8SVHpKMFd5Fj
I4JWUK1xfbqd7RXH1ImwY5GwyNZpIBzbqNnxz2lj9dqgcK9ChDnN5uglLtn3nUAhNcdBHPoCPONr
B4OK9LBlzhL25jlWOw1JMB+nNRDIv0rp+QR30v3gBBTXgT4xLPYAvRf4fW1BmW9+cUBTJ7je6stb
xNhIpc15sb/rXqJRfoiCa0OXDDr6npKR4exPIl520UJkcHhcOrqeE8SRkXc/sPI9mqUbT8srqlst
6g5c2enSF5jgqgPQ9oPNv/m64goz3BaE0ysStVwLad997ip7h952wANrmgA1sq6NAMEDvaIryQpG
Uj/SvsIyMQKcJM8RZwCoClpM2CVJ8iLRznmz1iMtdURICyxnzNHfx7M9BSqw0aomww0UeysUkYWl
h9Wuc19+aobka0XCfN11vWmDqHju+Ujl1z+CAJuQgQPRAFYgenlF5zf2hgwr/WKZCSY7PQYGviAo
k1v/Tbzr7wQ8Hs4DnuWXQvTDYRcwKA6nRXaUmWfsG8/gVwM23IPh4s8xgNIOJUHHupw/ql++jEzY
RSoHPLGl34V5QXxsLmCgYOGJHRtUc9xHdIwUcMMnyJ23l3UJ/dciQMPGBt0nJDHJKu1+GuJzvrvh
BSi8SGq6TCueXOAPzRRX1ev+ZfrNFvcahTD8odYPANCdrEIpPT9RCXwS+chUmHM0GS0yyBDthUVi
R2POmWFc/aeWtDKdAwCBoHeES8BO6hGYVbEeysDlE7iIOCw0o7cYyZl8tzVG5mi7omEHpuVsmy7D
Z7yT5ztvO/iiA1mmxzIT3pmy9QL/6q3/JE/UBv51DmPlBo4E8sVZQ/weMoY0qzPmoVtssSkKwP+t
0TLi53oSVlohFahMLlCm3ylFsB4Wybmhx4HAJgq/9KVtf4VZokEro+X2YlmpzaLIUj6ieOFxdc0r
aCYh90k+nT2UyaINHgx+tB2KN9CahQtj1UYecOUaHA/p9azjrniiZ0GYvCSZofVh6M4ZSVAwsue0
Yk0A5Iugou4xBRsIIbN5E0RTXFsMre6j3bIthME7186NJumD5/X1S/zXh3n14W2wfZMm+NG/XVNV
YXjHs63KGtzfupCjbtE1yuR87pVrkV7KaL8Ru/XRCt3EOGzpsILKlZACI85t3D7weR6AbHcX9zEO
4wb1XMO9p1hHlaIp8YqF58KNfcNqUMZe02fsIF91eScTAGQMIp3yV2gLiIrroTU5Hm8D3wisId5n
QaTrtdPS0zE1PzmSh4BglZzlp+MBdgR0IZhvWaHneu9ff5HXRl9oLFQQXp+8EBLfqkw844JRyQwo
jgSK/2qhVO8OrP0fcwVdLODQcfmP3m8r1udG6dzzsBc95iFgd+JiLqyD4zMMe6JiOrFtby5UGZei
yaep3nAqC4WJ1gEUYE/lMOnSY/yEEyFu06H6p4kir+yY6HTpTQSduL2FjI41lKoHbGQsqTQcQ/wE
V7InXYxbVt/7NZUQAdVsq2/HR/OLbdPIm2n3h1iEmd4DDsRZuOZEodR4z06lSwrZcC03gMmjYJbi
9E6MVRgR4Fz1Xm48v1n7is8+FK+F9y9tGWCQwOaoCVGOg6ZSOP1Xw8FZldgLDSOqBqL2w2YGHgou
fCVuH5kwfmhdB/psHhmPWovg83Gnv36dgsb3AByK1U78fd59V4Rvvh+877U840WhKcbwlYCG3CdU
84bMwCE4IizDJxNtH4ga/8QEmt2WoeZNhkpLfP0zS/HiwmjaSpsOxZxma4ZELGkfwEqyn47VB0hN
2LBH2NOgOwAcIghN4YwAZn98sIJBZpcZp29nAUUFzY2I0gHn0uDwSUl9h+qgLA5S2T6rWqgD5MIj
kcqGw9Np9bixw8ZL/7h0NeN/eu3Fdp89MJIds5qF2OaIAK/Da/rRfpvGn6rBld0TI79zdZMOSk5x
t57frI3N+lUrSc6y3tLJSYX3F3OwZK2mclxfIsNZHUBiFnXkzJIt7XXoVwHQabRm+jFXWg3TkWtb
c1qcimcVsYUZbowxLOm2i9EIktpXtAB3pgbdI7kEnzatGHFbuKrhQWHjpdMg3hjbXoW6F4LC/T/y
U3K743z6G3z/d0VeTdxd8MogP8qU6yzef4BoOOOvIOCduofUcR16uKaDXCs88yXkYIIM2My/d6Dg
Vl2nPw2eWOms61wbHjFa8lj0eWCwGmuQXx8+Har37sPn+IhHF3BfC5woFthSU2zlnFNJMaU7XGGC
WkmFH5YJfFyzVNTzqtm5HSbeK8i+mFbxdxscXJ8oZMdqAyFCqh+FVorOPZAULB/XqSbw1kNy1B/4
0E5wrWkOYKs8Jw2JBpLs1tV6IxwblZs7mdzV2TjPidBwU4j8fUz8setIi2kmWbzcgqZKiJHLP+rk
3FruVLb1uUVipOKqRYLKi4vwdvb8klpQQjxeAhpGPaB6Hvlct1N+ki7v6+z7HMwIj072bXa9KA8+
zfZSjUNUV+HkxIYjrBY8WTwz2VKqYWiyEnTtTMqjZd6IMwQoF8+n2I2iPKiZMBTqcDX7wP9J6kXH
TMhhM/KE5PlbV+W5SmDp1oGdF60NlQ2UvRkheTONMPqSrkbUuhiQxwKAmSLU6rYudTSWWa+86VVm
7G5rTxViL50XxKXPfy5gYDuLvj5RF7HiCwukeBW3mnoVjWVHuw1BVx5dECPp8ICa958eRitKswar
cL15j4UId8D5TuFflUwT1x+5BV5MIaDKq8PZbgImtaOhVlgyljfwQNHTil6YHRdluOD1ge3hWFUf
VtaD1bsIm+CV3BtVQ+d4+Uk6s3ENbOXPNrs5w98IPXdnl/l8sgOcUn5CmhGHoHcTexm3UGZGI172
a3zzFe9cucdCpfBkGbl+wDU53et18eR7iXBWjIg4tyj89Myewp5cckY6oKfOk0y+AwiyZXcrstg5
/QGXRV1zo33Ni2twY8gzCHJMpCnDenx78teFk7zBuXASnCPcqd/0FF4hjew0hwQrrwprTaZwDD84
hByj+ni7L3RNGfgyCIgCHieevXZd8z4VQUfl5GMoyw9m83i+9UWiKUKAcsXqxoB9zmznMEuMwDqm
IehMuTt8zkvEyAEflb9HjUyJG2rLIDxMlLwyAlXeaX9ts1sgDjl6xvEFJ8BsHoPfzn7ZW007jyFz
Kn+j40DH92GRYrkjaGJrcGz/GxXy1wK/2wm9dt5F90HxO2BXHdLxVacOjxR8Jf8tTwxL+YO7dRLF
fGogkWchlMF117Q/0RMtnSSLIAVjjlNaHEqdV3y91kS+XO7mq1Oy5ykWSbFT6uI6XV4MNk7esy6C
E9YCWQEsLG416uAjz1wm+H13r1QxPla+j67xOUxW4DeTO0Hunma2v7zJa6zzVIhSWUj+KpX32nu6
eBuHIfhW+fbg+tP6q2B2TaI+caSZ4hsoprL6NCpka/bF+Sy14zbzGhVhpD4E+42Tl0GwC9oJ1zVH
gFW95OsIPO6nm4UlWCN29V0Br7thWBeuDbTqWO96GyzGJox9Nu3iW3Gy99ipjA2IvHvK1JBiSyXl
0xUwXdy/XOPGdWttOScy7sYXJf6Y4/B6LhWDDUjz3DtN21h0BFfqXZaXyjW3YLh79gky8Vtxy5id
ZWA3nzQDprt02bmayTvWc8Zz1PhpeOZ6ZtcD7CSblW8OUF4kZc8np/2yVcv36VA4C8CkOay9LqdT
iDLu82ozvfVapaozNyI4KvxCIoj4IGGdfWXJAb76V1PAiWDmw8My1ZrU5kdADzuYGsdLK+6Y21CX
ZP4cwottEcOYp0TgisjKhjGvUY967Te/usLy7zV2IAOYaf6+7OcD8mL0W+lkvMjMWTSsRBXEPQ56
WVQyekBzCdC1jkxZ+3mehBC+A6xZ6gl2gVRInrXk08r3BlcU+3ko+xOlhrIenqEz48h27I7+tb6F
aY/pgW89/Z0w6uNs0vUGF4tO9m1X8jY6j+qYcynHBX2GOTs2jDBetMLZMM3aaV5hPl2H8/VbeOmd
ra4edypuzqkLHYs9OAz3+pE+IDRxXawM+7+krwwN0qoE730ln8jMc8pJxzKGrB8rJikUwRsd37hQ
vQBLzgGo/TE6XYfrwso7lInTRmmV/+vS5id5M2fJgCiYHGVxX02Qd/piHQwkRJyJFH/BI3N5Ri+y
X7oGTgQi4KkXb+zhLG6ojKb9iDJVhJMtZl8GzlAz/QVRdh9kZy4lhExD8hH/ytCUknte0fscyEGo
2cQE0Gx8yPcT5Js2tkoA58ltbHj+huSN9fBXV3UkIGeoPLz86BmIpEQoCZvldAoEJR9h2YJgxfza
kyoBWrE/TDia579+rYkA5+KRJKn1Qt1V5flbu1pler7qsZZEFLWyz6/7DEAuFu+RkUElAW+n5uaR
SBsthUlo+6mI7xvicru+E6i098XhpBpoci6wBSANyNgNHS9JqN9kKTtkdC8zm1TUrPpbF4WM/Y1j
mXkZTTGJP/xCiy69I8wVGk97cpBm6EZCT0nj+hNrYY/XCvcRehhs/WdOdifBG5nBx88dqtShKYku
ln4Ct/TOfmB+GYgKhhxdUKTpIJ04yh+ohuVE+kv7YsNrvPC6cldmEz9sjeOXc3EuJa7l8dplS8Yi
o0hqE0mt+l5xBCHhV4mZf2GDa3eeeOWDDwUl+zWopQhemQRXXARqEM2kiHoF5KsIoTo3XdCPaF/A
HFPHi83qggz5INt8SPMcK4o59884ZvhwEXp1J4d1dopV0YPtEAp8Vu6YVSttkLu836pR4Fahfd7a
2+E8D1WQhcw/WKOm2mSlzOe09uSzL/iYwjtRGTTJvh8WPF8O0ATswaFwyHmFfkdKEh7ev0KXS/D0
uOV901ALSR6ibwgTTTZc1WAFJsbSsvIjcl6muQc2MiuWXdKKlYJOcTZAHkmN3+SIjNHvp0wEweZH
2ZfT17VZ5umU+g3prD+vfzh0Op1J420EbqsoLoda7LAf4u0FAsTZawmfxnDsA5Dkby6o5ZO/96Me
ZcvK6tB9LcAxfgv0a6m5sWzLecrUftkoVvU7bvCd+NwIoJINQuTt+Rw6P/yQyzdGEzr/FpKiHyoB
SXZ5zMlSIUm/AdGaBYAI0ECvc7SpFk4c9J+gFYWoAanPZAEv/QKshS1zuaNho55g9zLAOIbqqtX+
qdJh3rPB2PwTFaT2+IwLHWkBXd7VGJHiHeWWVjxXhXxngRSKxFEGIqaBgOWqeje1ilP4G+Tfi0uw
3z8unSq2Zfciuhjbzt/Y6fC+4NK2rj6BiKPl27YyAdB5TnuujQSlvn+oUkPytILBetzRpvxBzStj
JUlElGDDXhTmvteAl39mKoFX2zbVmOqfcG9HJ4EWf/bv9kQtdKVrbZwmKVGyG9d7LDc2ZS95FFa1
EgwsfusuyPqi2YtBBv8ck0jwpq+xqh3RiqhYiCnpmA5sk1YdRSZ8LZyFtb1AnUcjWFKE3CNqJJFk
efKFq5sLS5w9NKbZWtwuAZFL6fHUdHFdEYsP/VGS5YjEHU/nsjP9VT1iS0SrfwfekTzdJ4An/ban
XOwqtoY1VpHr96qZc8ByzM4By5fZ7zHRu7qQdxV/Uc+o6sGb3scSbwiK+tImvTVCVTJYkpwewa8a
vpeCu+HU+9yT53BnurFMdnIghax4zys7MJyPn8CR2aeamWsa2LrhraqqwtOd8Z3ZdifRMd3hpLXR
HqXZFPKuzOHocagm21tNtJMDWePt1Ra06O+okIOff1WvVtq8o4FVJ1vvYqfqmGX7BD1iu3Fd8l0z
5j/3oF5/TT2s5jp0fZ2sGPHWnUljtUqNNHgWLG531fZtYbn7UA4qWwrapxgfDU+fkzTGzpsMNAKB
HEVmKGsN7JeuRmdwQxLeTXwwGFUzuolG7V6/Ke/Hro4KUg0Sahdf6FL++k0Y4bulSsxc6nR52B1f
+h58zBd3NE0PNzIU03/3uTjo8W1qU9ueZU0VyYid5hAL1wqe1YMPokP9IHpZLc2QmRBRGt1ocnIa
Y/2iWLKGtTjrqLalB4imdSI/zz7c3uazxMKJpvj+FtxMzr1jQ++n6JqJS3OISL6rs82640mV3UgC
Qg530stE3u1IFYC9aCS02i3ZgsgoHtypGhlwP0LVR3+F0zvB5qPVYYKdTocNxOGAr+xC5yB4081h
wwsSZJ8sqRr56tRlk0Xfn3NlPN4bJzf4iBMPPZTBQJCgAzaSUV941p1iTY7d0KfOE+AJF+gbxspd
QAfYRpQSX2jBs9ZotL4H2UFalT08fv/bT55EPLNmI6cvsh0+chd10IYFgGFzCGKta4q1EdJp26Xp
voOOX0WLbGkaLXVnQN7tiWH9JNlXEwwIA6gJteRzQcvadhJRKUEYc8q+qzGsainU6eS3xWXw4tlU
kcBM4dnLCfgn+j1DCqzjg5oU8nrk4XFZIiANVBOXtAO+16V4jITTkPb3S6hkCMfXfx5p5tB6HHml
FQiqxR4ixqJ92RiPDge9LibU3nTn2ff2Y9pT0jvVQxcB4wRstqIB1oUvabXJIMd/z1e19gUnN1tI
dLahXO//Tf/Jmgh7cfA72XNii1z3rbucNy5CbOZ3JriCRbuRfbaxcJ4EL75a3uQaRnicIJRSwoCm
Js5tzz3oQpl2E6u+giKRVusMiMOFyu7FnHRaeSCNi7fac1AYpi6jkYPMIw5jzVa3JXHX1Yvr0Liq
bdQ1SMrGofNBWbtHjrep4qjnR+Wvlu3oiABIH5T0zzEGjuJWOX0JXavtBdvd6vzRLQWRZuzgkLCh
6ryRqzG1vas8Jg/3oLpu+yUv3OfLz+QO5mXUiAQd/QcJ2CzoOBhKQhwBmCHS1FFz9b+XhOJ+Pp1l
UhgHxrs4LHAVmzKsdboLI1qUP4pKuRnYFxrigTxZT02QIdcJuS4w2BjIT2AITArXkGGWW8O4BJ0r
erpNGnfclFbsASlUkpy2ViYKADCzXs12FIGgADeU9Y+oeC/ndAU0+MflnMIiFepbl+1kFn7R7IMr
Lo6DQ14ZcuvZhC+KpG6IboOqUjvFRcQilDUM3Bc2G3EiyIB+dueS8LAa9rbOy1NuY14C4AbNezoh
t+mL7vvrFLllXpNx0ejj6f3hi4cXCaWpU1kgQCbohWig4/YfvVstLaoYCt/8J094p/lu/h/n3elI
G0RtmECFGiy2iw59XvCk0V0b/xoEwGdIvJAXigEUmFmm9MmnFj3phjVFi1ty0nBA+rVWTS9w/qD5
UQDJiQa2VMVDmbzPhni4iRxnVGLscIhXK5quxCYpsf9p52/dSG0zixLC7VW7wRBFJbF2xfER4IFa
Qwt+6eMwKhHQ4UUXxkcZpfihzxuFsKRCSSm63DyKqjf1N9DH1L9Ew/rJrMAq1WIUg2jvdkXycwII
DGrPgMpvaY3HxAbJVCVgxa/PWxbS6IF0WUF7fIv71B+QEMjBLB7hZJr9isCLdsl0pjokedt0F9/Z
H7NZUbT/KX1RZ7rFZG5eY3Zw2xwubXEdzJwdm1SQ+/d3hLoL80WmRtEZd7VufPY5B/5SMZwMCSbe
TzwuzZgjdMybhZ3u3+2KGEeaE7cvPXH4dVBZIyor+Wf1pWWxN0k2q+AakB8Awkhm7OMVY4k+P0ht
gr+mHpFWM+EjqxYwLUzqVsp9c7eTTa3DBvCFMBbZrIJk2n1esME6h7Ar8HuvqkMPm+noKGN/sloM
9uvBeiwmG4CktnnUn3y4itWNkC8cR+nAeCPfQICYRo0EPMoK6Td72MBq5d3MnHY5WTnPd1nfeIyc
9WfLs9Cly5xTrsNw3zJtCDqkDdPZWs4PD0c8xQNHdfpBdlnQ6kRFO7yI6rszFKeaRPR7i/zWrl3k
q37XV+ZWzPCr6IcldRAqFemv1aZ0LgmGDXmhK3/9KZwAFJLakjoTH5/iuaFxZsWPtglDS92W7X1J
TRjwm14xTlcq1JXkzn0gx8prE9LfvBS9EU+OaAwiLgGOGbYJSnK+nj/Wk5hXtfA78O7VE3BgQhwW
TRJQ4rH18zNxmFQzBkskp5sjqOGld6DxgNdoC1oWFunbx3UZqOsteHfqqk0AYIfhMhNR39tCS9Xv
PjgnNaornf+00cOj9SJJrAsfLb1B5UkjU5/Unp4bXGvGsgjaOgWBaSmsd+5SHtFWF3gPozAMlvPG
lAfCfif9SMOCCfF+dzP9capyyjcUOp7hkMCHVFwYaYs313YA2RhOrgYBS7yFLhRbLNmH3eq+dIm8
zGCudNKdePqTeM2S/rdT8eq9D2IbNqDfIpsBBPS8dUXBf3l5pS5+tMvSnOZGvq03dAcfWQzCDeLK
NHOZ4BORruHgSWL16Gsde2vfTZBGOMu4GuEit3sRAoXxwLpR1OGl7fMs7qfp5hOBGmw8wVb2rC+N
lch88W5vV+X0gwcLffjpih0/v/LoSKCbXcI/ZWlKJxSqOkrDFB4S/SADykt8excmg+SykEcpS0Ib
ZULl1yttzYz3UiAVFb+FGtxbq8ZkMCBfDIX3eCHy+kUycMErpV3fGD8Jq4HU2DYQGvIo0qyRs88P
UeZqFPR27VRGcoGjjVcrW4jXPdt8qI0t3Q0aS3gN7Hy7M/LrpPO2ehc+ZAo4orYuHnQA16Z0Mb6s
DNhVm8sOfjLxn87jiuYWDDZskFwwwl4fcbfOfJzULxR7Su/As15ggNhqUj7FqS5f6/XgxECPgUl1
8f9CtDUCx5ZH52IlVdJeGxmQaE5BeKFXW7QgAC+52nn8UfrPd6mFJTy54tieQkH7nt75vonAVKqy
PYOPVIgPX2GL/xJn4iT6MKL10aVfBoksyASfmvoJyuae5EbDYgTHFKcvcgULUvRB8mnbuIR+MpOT
TYRArA41Ba84oiSjhzTus6JQ2t9VX5lpdE0Xxcu8vPeL8xKzgXy1B/P5/Dl/9ZBFwpRlp3R81gMj
YECWEQICwZGBc3KRDK5iHbOdtyiJwxxEjiH/v0tS8OL7Gm0jluoYxKh0vdvtd19gtiF98hPqAURb
LPtd55WLS72BahBiHO8uS1gnC7dUjLX63jL4ZxDRfeRseTOCTcNrjX3bxcE7BT6PtYJdjE+JwKAQ
YG6DSu29qJabSmaCePH8+3pwFcUjJHJj03oyYXstNqvqjQtgv75n7UN/zQp8pvYPYr5F7dRn/cK5
+v0i8n0oJ6l7e3etGBn/KOTip63mKTBqjrSwKUWXq6YrPWevoNeEKrbwgzA3TTaI9yFtGj47K8Ni
Ki37yEep1CS3v/hePJUnh22jGdvATQuuooties3Ocbth8f4dRz24G0RmxtDLD6KEBf5zLUxDxvYV
SyM8lnPfJYwXGNBdXWRQBzDGxf14ppWhyGAdVf9uXQjWLFZfZKVaesdSNekvO1D6cIWmIZhu6im0
9/gL1NpEy/1FL4QHiXQvq0/WX3zdXP+khliTFDBv9SfPPoySlmdCaFFc9//Wza0GOxnWoPN6nE7Y
M1/b0gSBjdswpdpqMIxnadzcJIW09yiTAd+teptG8ij2zpb2bn+UeZ0raeCKf+PUGWpmVb+laPPs
cjb1NG+IU6NGenulV0TgEnV6+5+w5q/PEdMRcfcIdp1oOTw7qk3IHRIQf0VKDibRLILJQXUSUL/2
BNrA9VSHNXryHNiae+V1vGo/JV3gk6tPRJR0rU6mfZ5CxDPqqyuC7loxpAkGzDU8Zo/8Y8q6BGjj
Wg+1bmfUMDwbQdTzR0cXQBig1ocRVvnqT+jj646OyQeJocjMKYnKjk/JM8NNRpylsXdb3UDBa+lC
Ew/zKXLY87f2UR0T1zdU7+K8rWereljM4G/0hyr5MZ23AsFM2SW878oYBO3gy1ob2RzSS2MaS79E
DtoLqzEY7qfYE7e88D2tyf+/KSOYOzPopcDZxIiGci/UjATI+ePoGpc94YhM/01Lvv6t/cuYiVGb
9Wxv09UmzAoT8/LgUChJ0dZZ20BXcgvn98zG01JiniaOnqlJxtEty7jIpku1f2kvE7z5s+0lRRRQ
oMwPe09MzQNY+8WaYIa1RmGIDFEC26q7114luK7q2W3nHkjtAygU5MO7mAsxEyJB+mQr5qG6BaT/
GJqIuObvYGiOYb15T+LbuNFMdIgOdOWsv8eKzaeElINAGOqEwgmdqGeJUmUKTO/T/VFNJwqsY4Y4
uN+T7AVxiSxYN7i8GfuBY+39i6qm8reVW0MEoxG08DJKkVzwcxZoJY1cayEYsEJgOLRplMPU3Isv
IcYGp2RT881UITf+CDYs7AikPgF/COTtQoH3WhfbgxGpWUkZW0STIGn+5rp49gEhCGTJSQcYYS7F
34w/VLq7VX8SNM051fFurPSPIqH7hP6prFFKmcoPEghV9Bo/VBYKsnATRJc2o6U2w+jG49ojR2Sm
tHe8WEuTNxrkosS0IlEYbdJVoP4Zaab2mPaRMYhqtyYKoGPBbOs6iMc38lWiH3cwlw7krn1dWcoL
RwLym5JtqqKuiqyBtmXP1lvtESe4WqCDi4f8ydg39RM/Dwe2Eskc+44H9GMrqu6xSfdx/lfIiMua
qU1L33CO78t78anTlMDxS6pqwlHL4cWD/1McENzHQTHGT/3jQnKfK8l3F1dBGRGjTDGbMtvKIrFG
rba4iiF6qXur504BkM5NEyesO74H2WzwbhmLqyo8tAN9Oyj3LBu8mun34d1Q8kQtgF+S4Jo9khYv
ZvQ5t4Gd+VzFzBKIlRKqixoSk4MTSzgEVwUvcJ07W6nkjbrveYYEjxmzG4Q0lF/nZEp/P7kAhbbt
pfLkwcUnpHpWlPz3k+w4i17Dzwx5LX8vgquJ+K5mVQO6LuQTta965fO3zdl6l+H2m3ywq4V6s5iI
H7C6h5UC2g4zxIuj5cic3AV/kLhqAT70mGnHJoRp3/F3Ca6qyIhyGOktqgtYe02YIYDwvaUFnTh3
tKwD+Givn0rHMvMJk1bD8FcTFWvOJp5YGbZRzuFb/Rn4/3YYZghKFsADy2KktBKypc2IlGSoh3EJ
W3mAkkOb9nYaCAN2Pa1519vFOO+/ez7wbq6upEqRowAj69sw+wp0+DTAQi+G2fulF6gMbNVwsMYW
maxKsAfdJXjxd2NustPJ/Zyn49JYyXYwGqyUv5Hcwo4+b0PLQJnRFggoGEprjDrOxJkdfPsSBWuu
ABJCjYRUFrPzewBM2jSXEZBaxGa4wbHpGhVJqgQeMzk84M7Qv0UnZxAYT1QeVB7AORntLsrUNQt6
FWxXYist6J4XJutrz+S6Or/zVjW9p2FDYnjXZ96hBXguCS3sXBRIc04ZJCd+z7mnfWGNZYAthOcc
WCFLSnT5v5a80RwR++1PCAj+ljJZTg4xe52OODGN+AEBH7xUYPMePG0i9Rsy/RGPA0oTGP/1yqez
DU+EkN3SPG2Z4u2mLijZJAe6Fl48dLr+0CqAXXmGNkoHxHo49pWyL0Kyxh7KaUBvXglAlQZwj6Y6
AumWPPLxy70jNrL/vHjn4DIMCPrXIVfyk9T4yOVty1zWx4/yd7ZKez6Q20kO46eU2Autsp3kPC4W
aE6j8nXC9eqJw9aanf4dd0gvFgbDMrfwZ0sEXlLbNEUboSbG86fViuqOhz97OEVn7/LhlFURXWEH
bZGVfRKo0UMzR4DBIu7+spObsFQr2KpAMB4GP+bYG5vwl9w+8hVClAFXsie3vvcccj3vE8wP5Gsh
CHPeySJVWFrdPhWIMXUXdZSbbxMURwSoAxKiZyL+clL+3nQYIPsmijE7kUAWOpLgCVm/ThatOsRa
zfJ8Vb1e+65oCwjvpB/fhwIycVoaM7rfFvLUYFMzVPT3643Mw6nO93YmNvexNVR5z3sDaxcKzK1W
79UiMqhqo+q3u7QfinajlRL7cMu7bZnwWDbNFPb11TGud+BI+J6u3oO8MqW+4fBFlB6FF/VEk4FF
C1FoCryz6sjbTi15N2PUNgRm76cHbBsl2Jz1zp2LpdDh2E0P2WgoEYOxpJz/osY7kBl6zg9LxEg0
dOj/+rieOlJKKaPn1yLHf0/TSJbfGw7yRi2VFOg1+aGvuxjBzzVFNBUBuyecTCWLRz9PZ4lUe0hS
XnD6BDZabPT4hR/OULgUudX9h5/vCVirn7pUuJibIJ8WSPdmBsP7On8/dcY2AYXcuA9kBewd4CZS
xhe3Bbtt2eBkQjPd8bf57lGJSR9eFWfJiobIEPOI1WmaXC3qgDYxFoksYsqZUiRz3Uu5f4xCZo3a
KWPeWQ+PU6u0/NYqBY8NVc4JoEO4kYFTIY8SzG6+ZmZgaWUY36c52w/UvoKmeQNcW/nyKL5QMBaM
VNSmQz03w66n5S29rvV3DFP2iLBSAieGYj6s5HZZJilWgXsSa6m2Ht0bNzlSiOJJ6wkG0vfp7NPw
DQmh3qjiqZvVekAJNu/TBxdr66H+0Fda4jJsIddJXVdTnzuJQ7JpqR+P8pCQtSvuprdP3WBytUL/
h1d3SSCZKkZ9euQlk/OSMOTJn2H3MeljYvFNn9TAY0yVPv01a7MCfAcgFZRYU6phZ8hKd5Mdpk/e
9YlCKGTRA7hjBRRk5HARE8Fm235klvClg++O0l/0TvSNPCJe8AJ5A5mBu8Q88dImn7USyZBU4Zx7
TsRl5jqpZNOnF2VBlLVZtnvts8rIXNgscoXz8At4fvBebDLPYcUh47NHLAcgzhdlGRwq5mo4cBE2
yHPcG9FG8Eeh9y2zbsjjZBA0TyewnDGRM/Z7c1G06wg3xKFmw/tG+tCKMuKoC4eq7NlOfXovZav8
yPVrYGTBH3Ynbvd9BcUmslifAOIqpzXJVAzFzMY2r1u7DCycDwoAEGy5N3Jrp6H684RMRIQnyNb0
Wwj9sL0xc2RKpKe2dWUJEAC6iSDPw4jtdNQL9MDwEWI1PqcmX6Gvc4sjAbZ0Is+XGOfpZFTXuenO
OPLXfzGUpYijLRHvCCXZa4oXBexnfq9zBrv4Gch9vmdiQ+1NVqAnAMYc2mbK+x1KBpMua8a+dZa2
pDiTBcbAllJsEf0UCxrVC0OIJTWCOT+Hm9OwWAw0R6GyjUkQg92kXqxD+Hl0CsasIO6l/1R2ndSl
hXJNEhDMQyQCyiBgUkzOlVKxQ7cnhfYCYB7DAuDEXNWY/CGFWYc30Z2pZbr+JaO3VzEvIXXgNVg5
hJkmSKK49P5pk60crKE+/VxsdCRWpv9Iz+oN8/A+wElDBZFkxALzUSCRFy+AxMK9aLPE6HB4hyLo
fyv9WjN48YjHg20+KNhyb7AUuPF28787e3ioDz6VzmbbpequNlD9jVwbuzYRyNC+UQA7Lbyh1uiK
yEwGY+mvFUwo0orxAMjdt96B9aVFzjnETkc0k53sVZq4VNISxcJ/nUdZu2szgYswMoUJRc316EfL
woR+UGBBof3QXdA3ukrlABx2rjwAtBFi+/bdyL9PQ+mV8SnCiE4GyFJbBEvMy5EWrMVDQ9gIwH4a
BM+voKw5nA5RArmow5C9AhSLDMPXXiUdNCUgF0vN6tnrqijHze7VOpdEbQmrCrFslSSfNuGIv54m
87IoZbqM7Ayzjen5KiSZQQSvdgGh76B7zDS114cKuZekxSGdNwfax7+NMbPBF1VJ1k204tkq2ysU
eK8Wywb2SahcIBEsgbq/KK3BSy19KtTvWk9UUaHoyDnH0JDqJdCbdQXBmiwtWTb0cvMmYBHpZm3a
DD4mayKVFTSU3grXiO9Hzwic9gHCQoRU7t1rLr6gfdSxT0RbrSI8b15By7ZMadH+azxKfpopNoOc
+fHAybmPCChrULiVs1LGGhvVQdjlqRUJU2EDAceAgt+zDRvqc3RZTDbj+AZtdPgou4bHZdJE56z7
pXhwHXC6xjoiCC2beYlCMbMK2ghV4gIIdDofM7+4vqkELaVPwL7T+p1LwVS2NO/I8l10VOVRUGBU
JOAkdwPwl6dkPgQrsg1DzUYebiimsg9yx3iED2Ev+uDwDDGf4YbyW0lk8N2z1j+d22TYobvrhS0P
JIG+2kK0aczxqT/nl55zah0Uk25r0WJ3zuOfcx+bNuNanC8k/QFR4VdcrrKHHpsw/VAac2m0GoqM
ntorzE9UTk3+/Nxwn3Wu48WCoklwPa8R1RW491j0lYOKXD8aiFxdWkIle/ONkvoghxeRxlARHEBS
gVVDVMFwSgBqRk8kHJf+ia/4DygbQkDZFTwWEJlX/ZO5B5ZgVgeViG6HNipFz4xvHalUjR4pOGP5
MQ+7rtMUQakeT4aNPHji6jVE+L5kXO0g3ZLzLjdqzVs03ZKMhIaTEB3GH78EdouGbclHUnhT+DE5
+7YncgWFnpB2Nsgc3BBUee9XcGcaLQagWuvBnIwA3hu1ai/RFcbe92KdGy3YnhUlt8opuAAY9Sw8
ql56bRd4Sa1n7f7EhRSrDI/SZr1Vd0Py9L3ApqRwE083rORUHhx0bVuPraWvyHCUTX+/7/BtNW3C
FcGQE1BB0t35G5iLQEwHFuowe6nMJ69XBNuYOO9U+bzPVz8tWIfhOMkrgImoE7ILA+nBVUp7/h0H
drckHN4qC5x3/8w7HtxrBOPI2qEEMozfgi3NlJjiVPv9o42cHZxfg10PQxpQhE8Bl6vl2kcOuLah
sw5XIt/bH6i2u9ia9eEg5yQv+/iJ/kqwEYkFq1sOqADFxzJhs+SQz/BDKZ8pwb2/52oBvIDLexPZ
PlwyDVyackfu7s6bLDBNEjBkk77nzYCw2DE9Lpp5xoRp22BveSAauO3opc0nFREE2RO0LgiI5MaT
rN/rcpQ0kOlL+oPN03CTD+2KOBAoAD0u3oJGxg5RSBrXRrUBETxQRzb3ZbVa2Z6p6D9HJYQS4YrW
6etKJy+fj9GftX28cN2ihwNcYt+/IYjtupr94N1kHsSxuMPr3J3/mgDff2R/SENMNTkz9JoRddzT
0Rei3iCnqoAvmxHZQ9anah4ep1IMVYY8CwVRt05Aknsd24+1/YcbUtfIrbAxvo94mbgG/toBvGEu
iHyvUcuAR3ZbuYV0mT6sYttbKPjo7WYcPRZh2ssPVV0qsVph4LsvF/2kDGBAsfGeg4568bveGHBe
AIjZDVUwG4c7VKUA4diiNO3Qs0GkBr+dCU1h5tB6pA5hmiW4L+f5sexAMTiNhYvLY7RWYNsTEv7A
i6vgSXy2OWBK65iqXOGPo5b0vZP3WQoTVK4H5cn+HfK1Ae6LM5CkCuz3EwBi9tuD3HSIDD/vLJlD
h76SqYw+OkLL0aJTTDlYzP+GsJF1Sx202JVhJCjb+eH1f1H/du01nEOZOjdQdM7Sz4rbj93CyZBn
UYk91bEMEM3K16ifQPF6PzbWo52HflyaWCCx53MIVXQOMv/d3ixMLjLIQikijzR0InHVC969iHc2
EG6qKfqHsNbo3nTkSQi7bGqPqWwQ7uZXSt/smMMk9JdPMCiVsUQ+jb+mMRORHJ/Jd2A21f2EDn2N
OGVJodfJh2Deo7Wb/iGcoZtio2dk4O9OYrQelDArpnkkDo61b70ztQo2ASabq8Tyq/jfH2pWqZke
I+gTaBJuKfIkF/vT+vrbig/de+QuGxQBm8pgAAN+fxmud2KXRYED0k2eMSxWXoo0534Ei4umUjdz
k+c5nydfy7v8hLSTLfDEOBTROv99YQqnp/lRXFzPeFPdd3x7Q/aa+uIGZBBg8NYJX43o4kKaXUGb
OFGmU0zT/m/6nC7AGiYput1977BBWzSxsLRbBuCKTn7STEEQUHgvacsd/VSEcD55NR/udM/GPnYg
hAK6u055IgwcCJQe6McxHxEpBjTadcOWqYmySVszqNO9JALKP8loWntxYpjKGIVaV6+L3ew4nw7B
ZbcRW5pnrB4iJfeWLtUVeNL2pBvn7VhAw4wAYWUTHiFwezo0A4KIPRNVQZN+LLNF7i2RKEsj2GrX
8V0bgqlraTfd1iyg6vWyMQkeELRqsYYU50puJb8TLpuTpIqOUwxfhN+y0/f0gikQ4RRVCeB3ByT1
p2lV8qzPsivw6eGeOKaYjVD+l2gkzTLFRGH8U1qIdGCaq/VpjENyuX1upkpOOrSSO+FmuLUZHMdz
Ls2PT/sw2moG16fxvcuzUgCYciMMkvNRg0jiVI0Ge4I21nfK1aAs70+NVqNJ1ZlD6wI/qWQB479i
cVOhWh8cTofBdn03yyoq/7k6W8Uh6nzC2WA+v8ezq9xhEnEvGg+Q6+5i5TH6QmpGD+ovdUdGfpIJ
gKi//kaXVLT3eQW5a8FTyUlr9IxIeexdH1Bvulk5TfooSe3k0GkkSzR62ekfXBdiVX2NGkEfLBK4
ZwEAJ8iveZSZ8kFzy/2VQc7WQDIHVVFOfaZa6ArXwY12zB+rWw8ORCOIgG4+mtZhgVTQvDNyQr4y
xG8XOL7GWlr0XXFyKG2BjJwkLE722ZFyh7U87iuYOQukc5iX48GQk0Z4EfJ59+7L8qkHY6bzNCFn
hPee3vNx80b6W88jzeWHs3OAGRufVLnVIN+ItXGtr2UT0wSLtL+jxF7r+TUlumc5iLr35KCKlGRi
EcdvuG8q1ffyZgdPRPtHRo0Xn2hWwQmrN9q64a9Xy2DhEZMK0VRuww3wHRqIaIYdHBIFeizkVYie
hY9r6R7snFL+Et6yKRHajCLtN0qlo9dTN6MSVxyLwtak9R6hOn742cXT4L3XqGZYqb36uV91OdO5
x9NPAZ1GLJwUU8LCsUup+hawbq7kNDO7sQCjozJnYjK6s2oayouPtobolQbXiugLaa/N2YxqaoqX
+wJxQzj5ZHEM4f7aEtkvPMgwwr1NDWKtycWvCehzi3ssO+YuFeWkgeVEmFoFBeAXUdC6LRu564/K
oyElaXyBDVypnDaRdBv7WUU0DAtHiiyxhuBuEjtYiRcsnqKgqEXXpHHTzxOpIK0rzFdPtDK8z87u
c64Rfb4ZrqE2rqT7uiT01M6sGsSmTgIqKjEJMr/gbJNggcVDqap17x5KS/1ILBW0PoyVGtUfI6Bm
339k0aKUnJw/HG5e+XHxOzCpZTOWBcNtOkxa8Z9QoNpYsxepO6aYf8v/ZwtLf08d2KpnROWsu2oF
YnYWjkf5+OqEQowC/fkAKIcHET08IlSaqMmI4E0baT3C4evyWMDVF9hYZUS0u5HJLVMfEQWRx/5O
p61ha20o642wAqwa/kNtyrB+fRQG7iGWurwjoUpGv5jjg1UbKAJUAtcuPgfLMNlECyfdrGzgMh1K
Wasax4WZRkCIJ91nBKNyNpbvSZkdnaWlJAhvLs2EDyBtfstOAkmtJF1Rf9GBHBwWC8LmcYw5/iZA
oDnNzccBpurEpfog+Kr2jPukhQDnldvfxlBqOSNgWvAwQsxxh2BAOjpo9HoOg6r+mL7VIBsz2Kue
T+TOUODK+JYKA0zpX4UswKBXqYNhhaTf3+G7ol3J9TgvvvPuodMxQ5Srfwz03/6BO1ZhWLmAER6R
El+J1WEBnkO9e9EAEQNvmSWapwrXUPBP8PJrnknQyYNCusMY+3Gs7qZzAKvXcFmk0KBpldWOtDle
rZCMdDZbURxWKvv6Lr5lQYxWQBj/2YqA14WLJXpUqhQ4zMAtzvf70w905tw3grLiHVej/8N39JA7
q9i3/RBDO2cszDFoEMntpK66UAohbqOdbUtPdxm5JqFbrMG0ig+zkIFqWHmjrxPQVTWadRDlnlfY
rpUwm+nx4iPdK0ebasEjo0KaTmy8MKzoYjbkrXRAPeOqVTKjvbYo2qlSJtg7qwPdbnFp3ILxh64W
UF6jIgGJr8zq1srHd/LjgUF2BVd1SIfLIKh/zz+yXpXQFaDIs4tKNmYg0bk8ThOUKGy4jpDIyK2G
nyKh3CbGmNgDnS1yxZQSWLDMc8SJLXAbL1al0OCsbtkuVZuNSjWgi5Ez4rp+IJ+zGdcIEFy8K9LA
qGCbooRVG+UBdkoQx8MqceDCykHwzFmhL5qRoND4RbaGYp7ySrm5CYlasbGTr58gEAsKBSeu/9eE
jVtwOmaayga4kTAav40CNaVid6GHh4lzpCibNA9WVhJuP/b+dNWM0ewPuVzaxqZ4rl35GWEqbhnw
7XKlzhklh0CjJfkVBYiw8LtlQwmgs0dynhtYiDqPbPGtgBEO84GN3qTRA3NHTK8LVNKP75wjWb+8
d9Dvttfd62x+BmSVeeFy8w4dsncshzmuo1cH6fX7xHj8MEzzQEcf6leE11wakgQoVIhRmTP4e3W/
ty6ZPF2Uhc6CIUKWZBBsZR+BPh+Rm3N9E/O7gh5vD9x4skWnESEmoFKgf+SviJqzUjm2j6PLV90S
ffj87ZGtQ4XPQCr0jvOGyQ0Ao4Y7o7tZF5PBqJCIcm+K3KewrELld9ne1o4LvlGQFWrALp54Pix/
0jE94GsKluJSohD0QBLgySZx41cLJDAYsirYIJBfGsGKu4o9k7HWi38RZHd3REr+LbtaBtvzXI18
5+kDDiEd2ss+5pWXQqD17CKkbQfsYPiWjANUvND+o4GDziMgG3GtGMKc/P+jk4S7XKkq2HTja6ln
LyWGPEIMZCWIBqoDhmBPFPVUq8u/mA744cm4UfPcgq8YZN8IMcjKSWb3crYGTv8ImS0MgaFgwH9X
ro1MWUIOyBXIFhsg3rfme4XhSrqDW++LAus4yeLYixN5lJsI87JohQ/xOyzpB9wGzsS2bryfGdBX
GBZipvHQnXIrOuOpUnPAsKhjXYFM0W8imAA1PIhmEKemz6S+H8WcpvWjAIIr/da/PXbNYPcBJBZA
8oKJhdpzURYQOapeiOaHllEqxCtCrEA0Wop3kjAYfjF0NSStObf3iAzhm0yIrW/88ne5OmQ+9Kq5
tlqwHDONLX+K8hgA3VieumDnpx0KK/cdd2qys14aj+j+4JuBYVg/BbjopmNUkqF40rXCMTo3daOM
pT8g9wQLtZlsKX7J7iM3lEr7/BH5R5xsdzqPPDE+tnCP4fQoKEsXOtkuvtXkCZ2S1QyBZxymynEU
CWJm97YJfsa0lam0ktRfh7f/NrH45LRFeCpARDGCmZ8zpKmWpJVtKKGVAPpeoIDs1xczAHA3UH1G
4+bSkwBKrDqBN1gBr3aC6Je8DCWzwwGy4+9906uWI9aPIj2Viq43STkUwB1kWM7FlgQfpMX9/tQI
ak4wl/W+7bWTJniA8MoCcjRzpJznmdA9CSluIze6urCRwe4Sq8uBvtGQdAgVl+H4Fo87it5YO34P
TvKGs9TbluJdVxc0FGOrZNjdUyqFPWlE4SCvdRjJo8MlbPNl7SKRNYbrYKTYMxmkAvAgFOTSy7dj
6/sJX+TCL1dyScMsk9iDkT+4OZSTsAd4/CkFGv+jo3IPQovSXvatVTnxqcBsVxekzPSSbXmIFx+9
b1/evkK5QCqK6yHO9KYKEOHgNkzGHbW2nWMpFtvSeWdu4f6AOUnWZyyH9irbC5wZUNXb6AMaVrcb
KmL9t7RBCBB3yDOM53ELsRp/4/YUv4pzLYzdZuG4ewm0+nC67Wc1BK5AYgwjrYkobIh6578iyfFQ
CkLZvDuTrEx4RiF+61OVvXp0+P1POw/v43wn6FwWClnWNd1pi6buci+oyeCN/BiZdyLIoGAZp2QJ
/p6vHOaWsjHXuHDzBY0W708mBSaIbgd/69z6bCtwDtkzMyBEBN5vwr8lcluE3VxRX6nODKdwfyQD
SIgCPe6T1jZAT5JG5F9+26Qr9p74T75hNeE9islF6en8eKsaeJy0o1UEkaEn3IWB0r1gy2BH2bU3
q0klYHNRpC0QjjQvQxDTiyv3+LdHJqbKkLZOSk6a9IpQo0knoVThEPv0BEq7NUXvHwOIBZKekIVL
zV94F8lt0Q44h3DB/UnZa2nG7Yj93UbIwp+vCLR9HmSLwubmf0+zZnBiCOb09MNink/+qwGGNCMj
deZsIdxJ6fKXAyQ/mzUuF/p5l87LwqSsx1vkBFKZTb4Da5gKHCD+Hr0EcjoBHlJ37P1HCau+rnbI
IhpKN7kRhrKrJ+XEH84y9hnSsLTGjxdY8LAYrR62cq4eGQrM2FTZpTNeNOO7yU0n0si5CEOGF37I
r8GNr3K6w7fuPMOH27r/7D+BpyTQSYtxQzozSpxJMoXE6dBqgKtoGm48zz823MP1XXhFtpC1YHuf
Gtp6hhbRAQRCqoyfEG1pHg0hTayBE76vMeibnpamwuUuDU0xUjPKzBDbtz7qHN0xq1k1oaZAcBRy
0pLHEqVqNJUUK3vT+jonT7ox1ZQXdDM2riPuWZvpByG9om4lGUjZmtU+jKTwXGtGwceICkx+RKjd
vS7cZD8QkEl2CJErdk6rKnGaEzvPdAABN/Zs/XmClhzT9zfy0FDZiMJNZCaBnmYJxyv3FJKL28ja
0JBSjce5hHkIMTzFSR6iZxqidgW4OSCPcrVagZZ3zuC3N+67EcG1Y5z8OdEpTjbBQEnhQItCbOHF
LNPSvPyqE9VGDrl2J/kSz1YjpKmzJr/Fks7h/s/maqHKjXyalzVwxSg3a9l8tBlFvHZTt2Zqo95X
kRnWOz5NahfyD5S8MuLhdkUtDyjzSTUTcvLFGOjqnyNOHz7I8NPHJdZr7cleNAyUF2/MwuSltvMs
WD1yHgsTom5X6cqJWqLhHMoBgMS+9283QGWwNV+L8mqZ2j6hywQfoKlER+tkAKS7Lb8Uq/Ybzd70
w4HrJtmySoao3rRLQQJDmOpri/vbkokCkyZHI9Lr8JztctpiOSaub50/cNSEaswMsZRo+ckeIurC
kzxWfumHXb7ybJt007e4/K2HcmUhl9x8Oh1t4vjD13EOdY5nUOswcKNnsNZmk9fTuPIHm5UgzsHi
9P8zeMVRKMXNR7IT5NVFRUh/XzwgmIim4lwODhbOQps4Rek/4f/RgPujt85X4ahDjYn56u8jSCy1
KD3ay9Vddxdr4XqBbfObqTUQFn9N36MZ6o8FLH6oSdXAJuZjS2dZS8PBDO09m5YBz/TJ7GZ7e8vk
8uCbVYcfG1xHEp3catXBIV1SN+OWM4YctP7I9BWnu+V76Dg6a1qJmYm3+GOMsG0bAoYWvN5OYEE+
dH0iY3mH+v54egoL6XNQ3QNnGyqQ7RRirfdUaMX1cuwJcu8utxk6IsHY3HWP4CfhV4JuKXfqVGlo
aMCsbh5QZ93PSTRe+AFPOj2pqMgIyliwKzs0saHTzuT4xqci9BG73rSJj/AlDwxtHOVjZbWcdxgW
9XPCGRi2+OKmNP4t3YTkm2Y24FUfdxo5b/uYVOkgclt+g+KZyferVXfo5moOjnqj7KfUcD/jJrAC
/TSQVutitdbhPwhDuLt36FHGXWNUPtfaUbQL3qIj4+vZFftEcwHS7O+Ihtf8fhpgHggvLSsrPtyC
AtLMOSlyAghpPSwM3WQOBbJbEXQKT10CRrsGfgDtxIq4Oxui0iFzTvF4dvP6AjiN46wWi2wwUcXz
OASyib3odxWhxJaPzw129BZ2+U+UI30jS741wylpbYyANXgy6ygu0fbAGzdQ3iU4ZR4a4JyAatj7
i3KKYgJYWKuiajpmdynRb58vwMmfu5E9Nmm0KqqOtU0hAWLpkwE0gW0EMQ8X5wTYUh87Bpdwlh6A
IrcGzwj3/T+7iOnyN8ubIG+mMCG6PBlldn3H8XvQ9rlU1bB04IZVKp+jPYRYcGwODl6w9rQyhUCN
7GewAcl5iZF2bbK/tktHC4EEgypjU+tEOQl/QKSZKfq1o/ZVY+m0g/IpgUNUJE/Be9eg4Yxwj2FZ
eFouR3acPkA/h2mAm7twEuJRGxYx7tC8l9a1KTSwq50wFnz2sWNJu2COp8BOs/46Now57N7e20A0
TA+c2YPmQjoIONgpavVyhT/l1Pwi/5P+IxbpYNxeZy6kbIUHVYAO+JJmg28pRe5vpnhs4TZ5Nnkk
2ggEaTHHTSUaq0ZB7AzqKcqtLubfpPdRQ4RfOH6N7X49s/4xcXW43lop/jxfG1nF0yeTJMr3PsUv
mSOMUsjRPOZbwWF5P+kpW0gJ6tB6nYZcA76YTjIzEP8xBSr8KFWPLvu/v8hexWhFR1uGIKS8IFcf
21Y3IrVOusI2JeFsaxXP2nOFadjgney4Z6r2+McjYULmjz3TkpueNQQXbHWu0nECUXr5x0QGB7nE
5hY8Ugv1/Xn8CsJyNzR84YhfUC+wq9wqlcC5TD1hXwePF4oKoLL51CIbWIy4MG5Tinh1u7wsAQ/8
tFMp6PbxFDBC4BC0iP1+t+7MhKNbEx4tucOUCPO/dqY+QxGG7OApUHPbmCSe5oMiWro0qh1jk1Jn
z0k9+KFT3VJ5BV4nIzQI6XIfAS3a8mzfYRUs+0xi36DyclSRePSbqKLwXwrzc1bGlKO1ujG+rrWP
nBERJOAvnfnO5KdmfzvZPLTM1zTq2XOYUvnNOOr9bCuGCNtLA2nQAUwR95YnnGeXjsvSCig90gPV
Ks/gczPvNTCwR+EnGgZuUrJeTq4lDNyVL/iFU7PMfz/QYMIYdqJBs9cYm1BaS2FQjYHzp8j0A8kP
aoaSB0DRDgs/jxsAimsoZSzrD/IXyHlHkG/V1uAiNNgRq7eBdASGKGLcBBZ0BmGLL3ZlQfA3Kriz
f2Oo16KUDW+noYgR4tblu0mYRiuBhegMjNSixDDDQChKn2usOFbUm9A49Oo5Hi5JXc0PZTdmtTFa
v2I9zMVYTyyRM7zbY4RWvE4fijWFN++stFqIFDMYjOU0M3mfYUR3p+9KB4ETQWY1hAFK+my1dXZD
5He9sAnpz6a2FracDLpCLASnpVlhL+PZbVljQUWQnNPxfoDHr2RXKXZyfLQi+73ktggbCwFMJIdX
oRqUlHJdMhH69iE58MAzIdyYK1a4ZHL0RybnMct40TieZsGoTRCIn97ZGmIAe9VAGci3uuk8fd+b
+mY8J72/oyUO2xjJ3HqduQWOd+ZY3okoQaJePVnoBRJRnDkPELbVMOvE36WQdHZBtwQo1oFavFmA
ywyeKtPB1SkQ8T0qjPCx3s1y9RHCNAqH/8N645KUW/6fwiBq7zG/Fp9rcZpFX1o3osqzCmDLIsH4
BELL40hYkZjXb3evBY/8BcLraOCvJfrUdawL4VqeMGszacM4ZNCtEWhEpAZitMp5nt5gLCpHVi6f
XoR+aLDmZ+dRImpoNwjhFlzjN17qTjX0T3kP81RTtr1MEmwA+D7UxS3UDzN92pwM+uGl/TiguE5F
z8fF+v1jRHxPDBtxgxRZEzBGr+iEW+ZHoOzTwJxV3CvLqhqnLtH20g2m5w3cclAGZZcGKtWVC9fQ
Xh3uY8kqevt7xk4wdBo2XteoMdu9L01p+Okv5ewghvwae3XoS/7JOROTW7BR+FZil4JiC+nvtQa8
n7+WbOdSdRDSgH7IxwRhTSUFNeMv6xOqRonEA29fOT/bxTuPPj1lQN31TfKoo34w81mjihlnn3qx
cjOFi43GZ2vHZvsqxztSmn7UN71WZuSK2Yt6373CfRrdlyOn2sP8aG33cAq+79T6m61eZLQ2mTDA
rgPuE207VsvsCPYZin+rgiizp7n3ALZTn3zOUUfo839B0kCpxgoSSd4DSU2V6f/AXkIk+Sg3x0iP
fnMP+GMtQGv1L4yPS7jH4qaD28zCVRCDBKbO3Woa5mr5e3JF8kE/6Ip5LRRee8uBgJwmQaUMgF2e
fvjtPFIsjRZeZPAbDHP+OFhqIcKS3erD59c8Z0LIK5Z9/FwGNSr7Ui3W1F5unp4vKpx/ug2XOBbi
Jq4x6uN8627PQeSSfW+nkC9LBo0i0c4W/nbv70CK3Z5Os/UkRdXbPS5v5kPcm1etfH+hR4t52vZX
tjnpsN0w8gigW5eetqhruxh6X1/tF/glhf23Z07HH2fDZL0hkKKPoj8ExWSa9v+tKkr9Njq7TCdw
Ai+JdKouPyiON29jV4Qf4lECNr+gMKjhq+7/UAqCZ1W00i2E4cIvzUtvjXoObNd5l/EH1JX11cxy
q9mvEHUO1JJH+NPJwnVxfC+n0tWjZu4s0xGSJiKKp0X1YUcVk4m64MB4Mx0uLy6jzQQnJ/YgDM8d
FlF81DoQXJ+fRFaQkz0vMQm+0EELrCtWhB3IKp72qs/WyMakQ5EcndMsXPxMeia4dm1R6NdJHh4g
BNgDBtPmvHVApUUpx2x7Lark/f2J6W/RfYDAREFuq1bXO0iUz3yz9bWMcXpbXyJhXLtBfBKaET0G
PWreSDphgyJ/B4P/WqMPfnIYIuZsjN7NpiH85MIQoH1jDo8hMqyW5jiIcrUtLaA1+ZcJ35HqUCT7
mYq5XpTJireBRgtybhYgD78VkzCmHYW2yx9neaCQwUJIF9ixCrfEfG0oppH/HaSwjGYJU9UW06iR
iNfecg3uj4H7bbbBEPfVRI5ovaK4C1sjUwUj0GQQOJ8x8qCQwC+pKCxrT22bELJlNNFPAJv2bGlX
EMW1vZGSoeGfG6/6lR/VcBDONIQQHj+kqk1Bbh4jG3TEHfhkfWqnOTi8hNEDN5FgrPPJiG+Qqums
aUqtZ/pVs45kob41o5lU7wCYa6Ozg24e7YGTunpT/UYkILgZDl2gBSW75N97eA45QUB3sXm5zPPN
kcvbpkujn0ey44YnAVWOZN9yU7CEZLsyieEIReHXdzRRkBw3qx0qH+oqTX6Nmy1I+3ny6v9a3/3t
0tZNNetmtFgj3qE83XIJhJGDg2N2bl22P4qjIvqR5MN7+E6jsi+SgnN/UtxYJUJL3jlbmaPlQ/dS
FLN8M3c6o78EUGhWTNAtaIvYK/GW/9TEUkrpyPZUgbfyX/cfr6b+DDSlayfuaEJhb838KpfNWzYH
AaRP4ZUGpZgF3GREovomU/kc0smMwFeJWnb0OFndsEGWQl5VxTm8muSA7b9/e3bdcrLFFO5gRmRO
ycy72EsbCNUC/jnAtY3kN15Kes2ve5OA6pNuFg3QjbNSAMHpnE/vCWzS7tKbZepIXRz/rYoNe66q
CNPHxzO85vyoXiqXdOBBP102VhgJuW+oM/W0e1/YBdGoGofYtH+ClkEhYGlphBDSgZLMdxOdnNAn
dCMbl3gYylvfIrZexNEGNPMug0GT5A2l1CgwY6lhxs5fwVPW+gHXth/XEa7KHYtcXh7zGWrGhWIG
JbazlsxTNHzTGTacRzgwoGkdV71xx3zl+po3H5vepurVQaM5s9WFs3B54Ofs4oHVnpThVGbnqFr/
Vcio3dD6xONADWy0oHigF48R3FZyGCtn+hDGSQsw9a2Edp748XXeEssoBVQSVhAtx/gyMDx3ISkj
bxzVNBWEC1wGIEB9RaZd0c2XduXxSr7alp2YPqNBIPLeve5+QmoxNqIVCT7mos5Yk8fJ9ujI1/qM
WMYLFz9CP1+M/CbEboOdtwatYkSw/uUvRzm1yRu+PwDXjPdVQk+ck0U8JTOFcbU7CMRe1MuI/02y
sINhjE7cyePys4tDvxyQHDa3oDGeJWxvnbqVXtVIoY4UipwyMfjBH6pmiQ2Xx4LLvrhcEevSw3nk
gwxRR1ZcluS+Su4OONTEUyufECRhd6pxm/d0RmQSP5ccYkANJSiPwUu78GTfURBM81lo3i7qZ9xl
HkAAZFdw08TSOHMD34MG6JAIqtQWxhy4wKC7K5XH6nmR2Tse7CvBdsKTBOSU3xlpLtecOtmpskf1
PyBCh7+cWRpVcCoo1QREQfI1pV17rI4Be2Ks6dbcDezp3O5dqM53KyTkgzRGSVGl0HUMl/xip7Sl
aCNAujze7jqq9jQNqZ5/eq+w1FJ+8Wz56NkbvaOpPbXHvroIpk1uk9vi6/iwGSEgbUUVNYIhBKeG
ogk4Or2zsVwLIjCYSUtzEcD/LG/UR4+oqnHaIUyvECnUEQ3w2diKQIOC2gunzvocaE1sEgTs4KMI
OjZr/ac97m0A9l3e96P8LrQNKEGj7E8zYbM3FwjFQDsZwZqfTNFk6MiPlClfTOjpugM9Sl3pt2og
uFH2ML2RHSMboNxqORfMM9rEQUWOhABoOYHG3E1UUeQDRRQ8Cpg7b9SNniTZEvJ+E+uL2N+EAaMq
zHQ++mhN4aZGA+ycg/qdXrLwAQhEsch6PXvFzTbaGqRcQOh/g24/fFh4jmy1q9pOANiYzwjja3KS
08tWuNPH4aeTMm0bbCfPMKXLwCea4A3IAkvT/5cMkn/6ppZG+2T5l0YFpoaJLShBXEdjP1ONUyCd
ju8VZ5hFLyR2z9cUB6bCrUfxIkxrjq0GFfjAlUVW3DFosFoeE+TcfvJfwk73ypvwhi3u6BGrM7lZ
OptzLwxAQ9as7xe8yE/1i1UjiYHW4TMVgGPie2He02zlolqVbN3ck5Dpvn4OrZc15ACHe7xFBiKn
6+qv9AdOQTs7NrnrguT3Bp3DXKrhY+JEvkc5uFcWDLNl6X9qyLKH0nT0XiwjCQcvK2pqA0itEjj9
WNNeYr2MvIQxfLGxkk94AAKdnjGEsxVt9Y49k7TY/xnwXzcS2a0D0vJyRXgmr/TU8LxR17r988Qb
bYck8oXKDz4tVENgYdqLXfNW0X+/NbtfWHF2PjfeBUNNOwaEWJQ+7rDwtNvLq1W9RvYn93kUgMBn
vYQWtwI64ouNf6w0wYgErNY1xA3sQu/VnLg/6w7GFdCOEC8IIAq0jOJnncH5zyGJeEbzQ/wJ3C6j
r38YlU4fJt8Unj7KeFGMxip/AYu78NrLC6QxhfOkgKksEJK3XIUfkJaEbpGhbnXH8wbq9qxYzwPP
5MELFDotmPfpZXnlO5d2HQE4/uBLUuEMjLFjky7h/i9OYIJDDMqumrdwhBnaViDwxGQ9bkIm5Ukg
8REV9nWlunb+oTYMSMSamjG/YIwzX3GDPj1xFPDzw7tEoVKRxLRTGujKT3k25CvVObVFeTS2ynOl
KDwJX8D6h1ZWwOgxrUovkfWiY/Wv0F6aavrokI4yvt/jIqiDLdsojcjcpQcFWD5MuHAF2Exh9vh8
e3z9qDcBmLzjtVDMoWcFN2fcyZXHYjSNaXNMhosyC8sgJ6SCX8OAhJo1IxmzKh8HkLW2WpYsxYuw
7Hu/o4wG0c88EoqMHl9dhNW8C3GQCzv/U9HpnQcffsRlrROaiE3UhDrqtBT3aoakbwinTVfo4Fl3
/x4+hTZEq4DYG7fbYkdoOSzzrYERTT39bwrBTwQNADgZuf8BNpus9tTw74NnkaRTg9KaYUBXlJgk
qytgj2fR5WMxW2QnmDYE1ii6okISpL9UEx6czjDzL+WoitYRJtBG3HzXLNVwMLW0wEE17m40ZlyR
HPPVydp4TQ8sT7C0Yt3vERP+0X0QVMizLmCtsbZNeSCsH3c/bu4AuVgf2rTcZSIrgsuQ9HrLIlNO
c4EqnZbHF9axKEHC75LIJ1Bdq0OOEZ2NmIexDRxTP+sORB4GewsZSUidpHpR3RPIrtX66rPZ0qEf
+cbDkDoZ4SxgPf0cpK1/K34s5M5pN4s4iZ+5Jlom8wHse9ObxcVfd8nZM41KGJH8oFP0VOFaMHYH
zBCXZrUglL/4aZL8mQFzKH1Rk4nlk0GsD1XLIAPQMHDJZBUrQWQLJWWbs5219T4D/qDFXq2x6FUL
Xq4o783dQShv1tI5PLCa2T5dPrWM7InIrhppSLHD74H7AlUUycY672yi7YwyljzpnIAfbLFFW+1c
wPcgcOw7H5hMy+l2F5ZWPgLSLRUumQsaCQUoL24TWmNw5+kdhPD+PW+r1JGhueaZCSF8OlGGzZqj
erfhYmLaODKV8ASk7MWB9WRZYuVcb7WwmyntnYSgoJt3l3CW6QHmfUo+MoL35LeeECSxDcRLZ8hY
vLy+hCLSmpc2o8TI0z0Ypp1cQQLqJjJe2sXkgbCnzzOwTTz09JrP4teM2msYFGEJwMP1LeYSsDw7
WYhreDTq4Z1UFhtM8nSFrzFNjidz/+9zeT0CvK9NofJwh/Gf5fN6p8JqYBg/Jmn1Tu6F192Ce7Oa
0Bqbl85i62lTDdoq1WrcIPl0MEo5C8DMybFTZL3Rp9eoHRAnANqf7IBjtNUYAIsnp+9LplC04Mlw
rtr25e/iQvIL6De5oomqwH6Lvg8ru0c7+pMJdvHcGPJWrBUjE4TOn5FAtZaqUdaWGmWrgxGP55SK
SId9QB/f73iIlrwzQQ3g2JhkROZE4TLGRQ6BG2Fx3lpWYcKtkQninU4Vvr2R+BXwIBLKM4C/UT6f
1zITUrDO3b8DiIML6LVibPL6/HsZX8YktciCxV23j6tFRpUIHhwg1UzBtQQZFOKKQDoPxQfnoS4H
wu+GS3L0B6NnvxCp/0K6CKkvj+WJdFAQntfS4x3gwPDlieJR9Jqo/+WnAIsw2J08yFf+DVeGmCbc
YmBMPt+RuGi+043eMZ8poc9SBHJzrT6AASxho1U7c4VntOIGi4SLI89C9CMgD94CIoqhDJPn2ONX
5GYVtJdDRlJ2DYRu1N+/QcZHkNnlwsnYwXzSo3BDlf+9UYnFUMDcFEyt2zXc/sYTHVKLV3zqVIkS
iAtkOL24yFhztbzlKTSJk554FjLpwLfZ6bt0ygrS9kaaVg3i6pl4nKOPGVw52uD+lKMXUH5sQOhb
9ZV5k5ts+bb5xcG3ZGlxW2zpN/ke83TxU81bVxTp6sMiizyVk9+9lwLJb5IBpgQzFe51Eh3Sw4d9
Yr3xjZ7pymk2AsFeGuWpcTLqiIX0+GNiHhvRbBh2s53UIRFxjzwBKQLLATypmMGuR92wN4inumme
qWMXquCiYpsMVjq6tnilw+ozYdJZlnzWmBTVSXHMDfwiNi8YV1WW2Hqe4Zj2NSTsA6NY/9/bDWNa
NsCAb//St4Axoy4KthEsR8wOeQ4VEWf+tRhV0s3zztL5AEoMNPzhpRLQXz8LiP8ApKPh/FtDan4d
+5BhbKyW80551E0cwHTNx6uuDX9wXy2QKjCXdTkJQIksCSA0O6gcrFhx/XUXAwh6EO73gPKRkQrG
rqAQQzhzyjiUooSBSE/EHTL/G7bS863YDUzQaKcPwersSmKNEGhrl7yXRaaDY52GEZvtg7+dJ//O
gaJg0tFLOPE4cLcc4gFyPy/bl6cwPlxWbFGPTs2tGiuhTEgJOcEXmo7xUluOpWTVDDD8AoVW1gMz
kY4innxEtSQJR8pYr1Um3iPaFl4nmsVk6caIb9NKo5ykLfdKqrcTmTqp2+UsVMbzyoUR+734Oeh3
RW0k4EdpWnooywh3yWNzf/dpis7VqjqIxVTh72aBy9s6FPd56LH3mWK8I7K1TsYYt0tEm6ZygGa+
eoEc2sKXQwlSK6f1vFm79Ra9FhJ1gprKtMVSLLTisraPzPzkX1CqgpWHVl5+FSJuFNDakvPHWjab
ho3gLJ31XEgQGfcMjttu00s2M3PQnyocCAFbtkvcjv4vMHeVfAXIvxE+bm8SkeEqb1BE+fCu20rd
jhNuIQoGDaBhQN00CjEVdbmPVSvvBGjAzZ9ykhGl3JRkox0h3UiQmnLWiK27f29R0OZFL7zvebud
sEws+9J4yZW0iR9y3fRC0HcPia8pGeYk5mZZhWBWP5MJWv43rVVdYZzRvVro+sjIN1rAhHRIbgAg
ahzPcGXRBe7ZQVcaSD5BPiKmaykfxzU9MJjslWQ9XeAqXIeZuAPont/4c3Hyl5DLfx8YyqCRXCDk
3O2mmm3CM/gFBYgv6ULQHkxMcXS31fI4lw9mC0RGsWRFvZDpggjiE9rMq0O7CwEQAywtP4sX9sqp
zpBTjbKLzxa84r9+jSDKEHwSxSyKFFautykY8YdAhhZJqUcGB7fNForYVIK+sxRlaIdMq0pMtRYj
Dlw6U6xKpblraSHhEAY/l6yqQInC6f1pBBOQys98wbukId/UZHdMJEVlj43YCa8lEQcW12mzustu
5UMZRhyR1oqC2RvJ4vU96jRSH8cikh2NjeTfieR7qA//kPK8dydkHwsng7GLIur7Py+5Y/fO9Wjq
sCE8s+mnfnAZ1NaAAtPagcH1ujrgFnSkTYQ0UfqWq/qhpp794cZ5IEn61wAv5FFcP2wMXILpOljP
uSQ6gr6DXPR3ORrRV7fzMRKxftxCZIvkVgBSx2QL6n9NkIR4J9RJ5rZM0QMMWYs3CLuodFWRvOl5
dbE7/qPhEDQj5mVJJRdPtVh/JPy/i6NHPN/p5HA2aD2OGb2nvf51UVEnSDQGhEipW9e98VoBOOi/
Yr2yU6J6z5+RNl0dIQh8aM8d+6HhJvU0ZvDlCCjL5OF2ZWp62x8oTfWpLE5tFGAoQNMVXxGpJ4rI
vzOxFNZuI3vQnLGUAm1MEYWLME8HA3ozbexc769QN78EakOFfCTgIIJf8/6LKzdqyCNfIpbxhRmm
Q+iNe5kY0g/idFUfv2o7CoSqTbtRiuE0/wG1Zf6SbfUlI9aCK4d/mcLP0Ow+3+x7KZBe/w9BULo0
mDcncLQV5SVAOPAThPtzgh2k+ItJsdxrptyc1csdMkPBC0CzoMAy566YurmuOCzFOqqew9LsNwTm
kCVRso0B47vXPEQA/0+t9qbIbk8mjDfz88SfDc9EqNwGOQsjK/xhjiGHhK/ZuERkti+UNap0j8IM
wrUzT071gq+xUJNO8hWbLO5Mj4cwxPhIL0TXzlPi1kmRVjk024toZIJaL6eIbW4afpPtwu7VgVS/
p+s4IHL5f4NDLtfwPZxDmMsQ+h9TYWCAWAIhJEdf73BsSHmcZ/Mf54uSTV+ryW/K6zYQa/d9wA/6
9/znyRlaQFBowfd6B/1ranExXtuER1zw8yUHtMYyJkTeIrUijGUBthqRE7sS3H99wlfdG/Dp0QAS
t48kBSwSDK3vr7qO96sP1Z99tFtVu1N5Yem+41vTX8eIJe69bT/1gbC3skgBM+Js5fn4GhyCR6fA
cUQpWPrfzkADBMWJ8k1/6Q2Y/xkf1KdBKnqGwStwfugbmXQHhu7Dg6S2jVCTYbsLH2ZtAYy8SJVE
tMLsIn+CricH5HDLmEwnMawH5WNUeX0Xivfq1RRwpHWU7N1bDwtCS7mGKaQGtt2TiyO/IenXm2IC
oizRJFoDxaf6NDEkOqC/s83vXc93Jm1CoTDICo1SrhBNCNtaTGxsZ6wpOS5QsVCYC+OtWzWi8mnN
K8ih6BjJr1X9mgy1xf52kqv17XI3kTzH7xNDjm9gSXmeneuXbNkLeprFFtAAl3ZMSV+6E02IxFWQ
HOVy6ucTREZA2jDilkpQCk0tT3z5EmWPmB7sgKnryUGSEbj/sLqbsiVKgWa2obKNTKwzSph3rAzX
zwpfrbkfHD+mO4VlgCLbOMW9j9cvQ/dEERGUa2fsPXG+U30PMn53Vm9BU7Us4tQU84kcJMWwLyHW
u7Z33SUV8m37p6DffJEy7ll/kROoA1quTTgy2OXEuHmoW918s1wAQPyr0cmy2KMuL9tBPuruieEv
FFaM8XKEXcrm5OghQYTm9iIi4nywJdWKRsA3gJ24XiSXV/Z/u9Y7lVP0pdlm3hXc+D2lp9EeAZMz
4WEHkIfYp3Q6k2prheSegfF3BBF0NylmQ98B63bSdW5MfGXZ+Q53Alz3E8dZrIic0UTg5qjntbw6
JJ4uasxGdNyqWrd+1N2zxqmHdpsOJK3fym6ZFguY8daZX9ptfRY13m445jI6TqBIWahZW9N1+91R
UA8a+YfwnqpcXUAjHrbkThyLs9oziCk0KRxec5HaqBsdl6BZyB8Rqzoc1ml9cbaEEDnBclt9+6Su
7evykToXIv71M89iaOmKCp3bTERzXk2sJqNYNADPzHMaQEtgUhV8slNWlIi/OmU+9dLHnvkyBmF1
IPXCbBW1cYLlHwqIPGl73bh/HZGijrjUI2/IhCXZKRCA4QQSyhaOnUB/EMzqUaDIhPbhRJHtFBpe
ye+BPKLN5afJOTWb1LGo/BjFDRGBUo2pZcp+gHMdsM3MTXOrHE4a+5JkPeSncW7eoK67wcLq4nSd
mGGpwqhd7Z2RMM5Ko8nSgACZl/yM8Fmk61bsc/NDy9QUM9ycJt3nwUgNm63EGJQShdJhfwwO0yxK
X+jgVNGL7StCreZ1201rZ1GefS096xIPJfsAwnGAr8/zLuy5jLyrzHb/Mf9+/LNY7dkEJqhsg2O8
cSkpWKSlJJuPrQAYE4NdM9Udb1aPyUJlhD+Xqh7sRIcCcuBZdoTzdo8iLKmy9APkYfZttsRJLzuq
I4CjwYzv70V6wbgtvVNRyWbvEtoVabzX4VM7nSCvL8kfrBp7ON/vlNCVA3Q/aSqwFPw3mgGsJL8w
szCTmwOUyb54ZjW6nna7HZTIT/TY/pSAKfYeTT3pzctqUa1MSm5SUqjDvTTxrF8hZDa19ZTp2+89
Mu0G9JrZpX+Pw9vz8CHZBfD5IVQKdhBTB4KBqxpOQlC0nQiRPmQxdPKCZGAcV+kNcBanRsPZOgXa
Pj88KAtSrtKto8LDu5XAiKUSv/6Ipyuxd+NJWIvQBsJd8psucf5YsRIo3b1BixWgM4cf+H6j36qA
je2AtOVXDtJzZCwKF+MblMircvzTNP3bv6oHbxrl/NkTdc+ooF0mOpjlE/MFWQJKbcJbXeyVxGhx
XvXNxgCl1JImo0mWYB1R+sj2/I+MqUpSe8lTrQsS+vluVWPQW3De8nuLtsSV7VbVM3KbXFyUdnjk
kd8pXGh5d8enxdir9RBmahZ8TrxkoOXYDi7hcdoCFsFybxORQxllhB81+nMDt6trDr2rX7dIolXS
dVnfOaSSxldrP+Jshrx2oxN+U4DIjIzuZEF48a0R1hYKbRkaqI2UW8BbtYGRKZEjGkItIGzHiBgv
PRnneOf7lOpkaV49z3vm92a/7mK3xQYGjpRQ5FRFHH9D/QzxvP/GIiH7wwd/tBnL0WuMGVsV9C/8
4vX+/iXuJ+EGGXImfjR0JIb5DcjvGu55zLNxsUPoWP20xpLDhNAaP3WjoOx6pqRHg5uui6TYN/0E
cA/rPmXbOrk/6LiHrP2NMu2CR4HHZNxVr3d21joAUHRJQ5/XwjGdG+wrt/GDTaCTZg2y5RMFuNuT
gD3KM9CFpVypopctlIAY6RdIf0szEbY0ZsK98dtGbXMXRgFi+I4PyEm7nqpDIf/SynT+uDix+Gzi
6pOAAM62PeQdKXbp1Ylm4XlI441xaEOxDZ2QCwnlFmv9iB323bRCrFey9UOnDM+7uJLKy6QGjZvU
SVerzNJWdZ2wkN6z3arsxgTkiEy8wt6Jia9NQqmIAruYllEhkMt7kOPJSBritYb8crRiNVZao5Ei
NcR2ppTILFfSYXJ9Y8pTYGGHctH+kH2aJ3Mnz1cojzNLsmSYA+YEomtkhtwHXwCPUrpQ8kJ/hgSp
T9xY+3glVwxLWhOcnUfCtoFzCyStMCuevC9wes3+qV86zmESrvLzBg0SfWh9oH1lG5PKEENdvc5l
6luyqXTLoYoHqPnQl0wkx/s4cESgocLNctj79ZUIVYRkVc/1UmgOk+oZtZRVMnNS3syPSPJt7pCK
SH53uOPBL0RvLBXZABSxEEGMPEEpjgO0BVs+ouILWQ+Nbh1vn1K7sciJYnoEl0/3kWWJf5N/579H
IkZSHXOB5SWkKdKxQUuvKXK/4/fgEhKoJP/BJpMx3N+gpGuXZmVhj7JkrFjcQhIpUUYZBFCxRb9u
FBWl83ZevGdlCNr2qF3OD5qkHSTQPiB4xbi/Lrib2I505v7wlEYexsv8AxlwbdNgEftcEwdW6hlh
0MGZalbKUECwJn+r5D+G3NLV7CLHT/uwazNQOb3htzRFl0rEbQgr+lMTwEAuZPEVP+d097o3e0/M
GX62BHv5D/K1e+YfmC43K+KAOgVGbpjoMrtQkQ5lc9HqQit8N6VLIwXc3MhHSL7wisH+ka0cMyya
LFNX3rLr/iBPAR1Xk3KmvoIWvuKgXMNKJl7dBXSf7stNhVEaehmD8XPBQM5xj0Y5P9L3hBO05Aat
UB87x0yO348PJWhKXrI7zpBbyWyvgjGq1YRtmdc9xckgtDalDlFTPnNeezlNWBlATZ5AyOTjaDf/
tlCWTVQ5PNhG8MqSlfJsdEH6Rlo0kCqLdRc2S8BZnHF70+nr/sGtkHA3+uX1jNqVwsjMM+TnclMd
jXmJtK9VEBYh0YJnm1Smvz5ZmWxETrEWLZhDL0ELXnDRl3JuO5O1nYp49stOrtGUMnRbvU+vFpuM
aavewzMJRuARq5mzrP0UMGNoOzhOIhkHC/CIaY16ePpDMDLA/YIb+1Efpdl2mb+Qkbn20KgW4IBa
tG1MZ7EuKECHVg+OQhc8OxlPqzc2ogt2v+QAu2rjkNpgtQwLc1t1mICpyPefmJ0hzGuBSOx29vw7
ogQ0eEi8byPLitaObYS3fY+w/lAYFWbWfeXT+H78CNLm+TmO5/n2GOLBvujCmmLQ+jaBW+OXAR3a
wSiK16okiu0Japyq+6U8EOVa2GOmIDQGo23l9FUvlKURPN7ijVzcyOlNhNDEk88RIYpwy7XSOLW1
xPTXm/mTadiOHJ+mMpPTsinIpcMdzraOc+DaCcX7eQ7ZSjDOuMEXzkIkA7RuwGyIcYzK0stSij9L
ptMQQSh3rpShQyFXmrxvpF7cBuWxH3AfTgnoko3MA3xniNcMbo28FBzDrhfoanDzGRcboKWcSuWp
qYdYMexFQ+v7Un2xBcbY4Lcix5bZ1I8J2CtoSgqDWf0Ob2bEcFjLpUsQgRXSsvPCdrW9gHUciOlw
sYq5aVdm0LX6USDtB49tksgo3767jR9dqqWNDbT/lChaQ4wwu6+lvp9j7mN4XcM7hjOh3AcQxJ7+
6K7ysPNqBTE9LDXcKAHtHgiGRg/jZd9EzsTwS7bVp6kWwyn2TaAH5EjUvIxcrGMKiZR8bBaLmpa1
ry8B1xxFoT8/r//r9zSyUp88TNnWpsXzOym9G3I4wUsBOMNtQXDjueaAMCr7A22PHc+xK+GKCahj
jVqKTeZ2y/0iZnJr9SW54pNPdku2FUg0Xu/feOSGeY4wXe9z4kYwbGkNR8IcY8jPQDrZvptvGEgN
8jkBfYq1klji1/MduxJldZFZ/KQCoU25DPnX3NaCuhrtEmah1hJPBbGlBzZyHJUSb7A1X1TtElTG
8Om0FX8ZmhhfVPqAqx5Um5rxsQVQwXkXCNnbpy6gu8YPNxUShSNUcCBL75ZCEC8QmVRf66RtJ6tc
86gTQJpR84mr5iIU0NcRdiu8Ag0fz8BkUPInQXUQmoaCb5nG2iXEXNIXKl/mPAPMntMKrSKZU9eE
P8ivgISrqKi25dI+rUX0zLaCzlkqupYAIFa4UUtxDuJ3Kw7T5DCA73Cdm0bXkau62UIFGsBOgu+E
tTNv+06MgsVk13eYx0e5WNsMmgqushcsaxu3fgBzq3tFaFfuoQWFTDMSewjXolKBCyuj+SlA4VrM
rLBRqW05iP42aZhenccSxj+wwpdZzTmB8xiVmgkWPL9e15y/zUnpMe5lSJwXIvW8Dyg8y/oQGpcQ
65pHYPhivk9gGj46al/N51oEfo68x86MBct+vGYBlgXFz3fGa9q5uThaS/Cu6PfoymInsWtpsqB1
OKH/4s/Tq4lVPPyu7woGLshTHHkmEyfXPLNGYzJOYi3idj67jPzMlOLNyVwtJ77GgQtpkimP4ETy
f5Tn2J3yUpF83mWm7cSIULuAQ60tyUno/SEAR1THoFfKmwh/Z335hlquCVdq9JS0DV3+OShIhUTJ
B+3KcXzmcBlh4FYRhMSkItUcAlMLeOHnDVJMXCPXu5/Kwurfsb0zaItM+3tPBL0V/IAIq1LWx0Pp
LXr7zl6zp2eXaWb+M5jXVqyqJjSDbBfZgQLjLS8OCCRXJ7ge5JHnu4aMN4QhX2N4mtUeVqdVSuW2
WVw8rUMJgaFn6CSsOyhgLpINuF+2DGywbC+EsDkH4P8FTbSflI/5a3LH0UU/HqNi2Y9+3k5I/amc
lecdD5WIg3LShXdttlueAWCFaEBloyOl+k+APV7XEYI+EtPPjF6S6L7rGMV1VSa2i94o2usNap+y
a9Z/QEAyl7L8le5KcqW+2Q6fyZBcdpbU5blJiWo21D9p34xetlAw7B7kq+lekrnOUQT70T+RAGxD
fXREthwuyFyIq5hLPMTSJ9luorWa5DSXXyqM19d6EHB5CidAvpSuWjsNKMTSDuU14ue4PlrTZoiz
6zhkuf2UkxNTuhVsB1pwrjnk+FipvtDfvpMMdxas/JE5SeNp+m3vg4Hh6wGra6Wip6JuAnwALG3O
AH3KrjqXbjDN4QX5MknOAVWqhfp88aGJdYOJbXGgeslryLCBB2iX+KxJ/57U2NHw8VV23qiLCpnP
cE3LsrPO7iDT+JHMKm8MY8s7gB249gZDCSNMm3kDGvSy2VR+wZhtqIUBg7aAA7vIne7E7f4ueR+j
vnpZIB6GhEmFTiGf93xyI8AZFX4IqH7w5gjqGfc1E2QJc93mH8zZosAoT62vMiSzeW1sQeEmlN/p
TohY3qiT6Xulo2Gue54hPxjK6fpWvq5DEPK3Im0SlVfAe5+jNyxWqLjlDeApY+ccyrFOakI4NDnB
KAnNw8FH+zxLrnRDBQWweUz+a6lynhbK6UXwOT0cai9k8oqxHNTHOZj3p+7FOa150NAb1zDeIA7i
S1pMxnp8o+SOx0FTEza0R5UPtMLQAg4GS5hjRoaoXuu4F6kghsbq6WAvvzaMyTO+Fw5lSuLDWUwS
7OSLY76XVH6dONIyLyRmpYEqxYvzZ+a/shPLaMK/rBBVnMkcmfz1kBNdMTsBxPceg9c+CJIOjLtQ
YDr32NJ9nDNcobFZLRCJUqm2Hod6ZKvSvPcKFL5sQG1CaCnd0MZMXpksAQD5CvXDwEOnZ6yj3Wi6
zmkDFCfazm7QhHuQoBzxOQzYqaAIdYkw39/daSetkN8Loazk1Jrt0D3nLX1OVrBNt5G0/bM+QdpM
wCFTAzZJN1hF2Qh70QCKPUpBZdK9JFkkIxnSm/sRFcaSeMSJKcEEeXHJ9QLAxO3+qoQBiLnHqQrn
oDIaFpuLa+7AZfgudT6XDXdIFIeeWr7aSNoETAHEadYJJ8g0j0EtRFeIDNuAmZ35EzQ5/iLcXE0n
4x9Jf8B7hFbibWh32b4Qs6q1TJLeXt21vsfVea8nlvOIUrXg+j4mIHD7BrvKKyKu7Ag7h2i2teEh
ZJfjrTGB6tXV2n6l5uvuSHXOwdd9C5bpFFP6nY7iO0bSieg07I/AMcFdfgF/ua+FgaFk0P5RrV6Q
Or0MC/NtVLhgiUxPbSNBL3bLYXnojIRPOeaNieRy26Jsv2clldUNI+9DAMIffmRGfx5PZXft/nim
wrXM1YOlBS4U3fYk5IqOLNQimvDy4QsiEIyYL14/lZsH9lKAA63s7yYP9FcUBS6AEGmeMdtIV9+E
f4t7Qm9qMuHsXJuM78qwnxzkiIzzDlNuODLfxun1a4XepdiV+YpxBnPHLaz7Nl9NsSewlOKPxAhB
YLhjretIi46DMRmQGk+YXY63jqxxiCKu1BDY5D2ogK3PBQRWAf9Ia8YTxv8oUK9+CGlHB6RdcWIm
wNoW8acDYVKPGbj5hc4i2sAdMI8sfs1O8ueRNEciDMCv4ZLVHenY++hugOoPlghoiwFrVPZUEYFx
Kob6UVUfcxIp6fBYdBVRmM7PbOPtztJvnjEoafBgsuiTwspi+C0RX7ruyCbjO3NY0VgGTqYVfKG5
Q1XYVbyXvsa833nYb4cbGvspFzN9TMkI9KPVzEz2sGuz6AGU5VJKEzIqs/nuAyihrh61tnDhjTcB
dNcTtCpvBAc+YnsV8w1cv3yla3FMQW1K2GopLRzrRR67H/CEpUSyaK8w2f6QF4NAFR+zMyQZCwa4
86k5nwKRcyRfaemE5wmqJIO+C+7n/MrvQC/a/sQeBBVOijqnLNBdM+ybRfogYAWqUzHq52GgDKFS
rNcXeUenLwZ43My585XiTqL2MF8eRz/fGlV+IfNmSDyZdFyI1BSwCAOD8Uhx9D0cKa6/JuYoyjMt
+gx8aAvrBOxeS/rWGMbK52p5Pp4EM2jEofQlmzLoioeQJWOtfiMAbOhXWiszoyM4ZWuAXSn36Q1U
i4HI5LVkFnFJANe9ouUT0F9CTqy8FpZhDbTjGFnIAdcpdfrprRqbQS3vsstCm9CwykqM/q00gNGq
T5lkBOSRU4TG8sPYaBwMO1UqVxmP9u+XkqqS4ungBkikHMlDuydrwHpRqeyFVHEVqsioiN7Q4iTp
c0O0gtilUO8Pi8js5eAKgW+UeI+5tQyu48aBqEc8IB6mxK8rm5qLCjZpRFnN2lukOGOcAe/QFSKs
70HODDbdTQkaA+r+s0Z+Qjlo6M2AmBcr+TvQgniAooPr1p/l662uGyhdX3Wsgva5n7v26N3mK0TI
dKM18Raz1iXWvWdZcI/eFsirdHGnnHuZNFdimYo7mLPHzJtKCDLiI7jEIU80IKqXcHUwPFNAbFUY
sArKtRKSWOh6jiO8pMP6TMJoS1121N39ILVhXNO7KXwA01o8rEFE6T6StSWMNRqIBSX0zHZv8nhR
mwWPjZEwTgAwmz8f+w6UWdz+UnfumKSLYSVbTdeUlN+fxVZ4Zvm0DnXw2Er9XrRm8mR2rSswb5XF
qTMLuXbpEDrMlXjN3kcwvqfCC7nU0FzPhqGxrJhRm7ciz4A/w9Qaqj2eagHihFsKfBwVTaA90vl4
pVi2ITgX8fn12+FYNLqcGVNwRE1yzWX7fb/8I+JuW1aSQz1nxJSY5cCthYJgm1hxtufYK8asP+CT
UMKJNp7w1/SwwUhMeJ+RBlK+H4/ZsEt5z5Kd+3JtJiSptmlIgtEEX/ze5rGO1/EcczNDBeUrPgLM
h0ikaDa+9C73LmRmnBbnNdIZSkPePmsKLwri/ky9ALBKgaAcz1ekeKq5z6uiKP8Qr3n50J9ttKjP
z/pAaplogf0kwoGues7E4k4mun/gi/YsJ4bnPsFouTb6k2scK+EhkKt3SJIfEKgrclcZ2n4T0kzN
QyswwQOidBJSHtO0CuNx0/NMFbSAekZa/mBQwEu7zauyfDxjA/knJmbNqUE2WLta3taCM8d+Gojb
6xJYAMvFtxNrv+rAbyn8BTm3XIzKi260B8t4EBJrCa87cncxSXnonVHXGr+8hLD5wXBdU7DpKbXN
Gnc3fHqNQUwFxrzsnNI3bxRk7aHe1srVaR2q/A679t/JPv1TK3kpGYHWQPVgZ/MFjKY1NllPR4/b
yetaWrim8YP1c9C8DdTSpIn0oiiRUXLz7eZ2kp4Oq8olyD4toFeWBwK54ahV6VeR0gLopyxHnEq3
CLOZqNldtipQNmtDyjQvwGdR1mQI2BcUstmiVYo55MntepymHbVoOXvtNH8NmlNiFZ+wkVRFd7Xf
mdd2RSjxusNaB05tma3fVbdsO/t9F5ZoYTLsMgWdgm5V1Y1Yd3A3HFlRkUdHjlgNCu1SK1UQYA6A
Nva9b7ERpM1VP5NnLmBqwdinY3ufv0WhcGER+LGlG+xVsr2UYDszW3PrX1o2GheE4IQ/LdVSGGFo
VW5tQCKsoDTQCue6FPZzvZqa7zGt0CotlHNwKHelxNwNzyJmC+VSX3En6tmg/8+jN6nl+cZmUUrm
uobo56EapMAfMM8PoRjUq58HUxRmhWhYcbEAt71MVZIfqbwVSaLKI/OV/vsSi5PRQSdryUgMScEB
tY08umzRGJCFu1Opki9HwktuSJlL/61AyOEuhpgU8ygZFKOkXriv2N4R4qvpaxlGRTgN876FoxRx
dibMRIPhSHvAGVE+l15qBhiDhJvqw4Wltgo6hU1J1rxbnBBsqfRNvvtTMUF7G0wgbolCrHi9EjRL
6zcVPAdePY6wQIM1M4ULzkRtVsrKi5wqxr6eSB5q6LQmo10JgXXaMs3ysu/xu5HseiconbCqGZZg
FaEmqFziwG1G6kHcjSwvegLZKsNYMjfuFRaNoHXY8pn1UUPH6rxknbUkeQqUopgYvh9z02cX401Q
LQX5ib3xfVhNT+EmNmFdVrV1BUbP30ZiK8jfKl0ZqpJ51EEZOewCtecgs9Z69eM1olzJEBxv4TUu
uYuP5nDiLVZSpfpAZJ+UQJ9V2r1eksLNYO7l/Ql3nQsSH8aZj+N2E1tLwVogic0JTm4a4VTg8Dkh
Zr+tKTHRLQd+hyTt6Bbtx5mMvRXjnRf2E5sCffN+GkpojvfRwHehY1cXcl9RTgQbK4RmkY2X6UMj
2VKXR0TH5AvjEfkNdFN3PW4whIHB+9/hWhfXfz+vVzFpWo+tSKMBQzlqe6FVKDV2R85haky4iTfg
hsppKYqP5SbbsfQBFU91/9+NzmW6ty5yff7J31C45XbjftLzDlMelEbn90x5jcAn33UG5r6tsVH6
CUmCUoxSVvF7afXYifvKjZ44pH2nWBOwfaf8Tdqp4z81CzTpFLV5nScNx3+xDvZYwlIXLKAofzWX
1k3ClEiFdpsOEXp4I4kc6KiE/+4kyO+W3hIV5UO/qxuoSjK1OF13iQIZItFTZmGn2X2Q01LUnP3Y
i5cOpEaxHwneTnOQlEKrMxK0QI2EHQPr1e8QrrqAwcST+f1XsywhAaKDiYlxcNCg7MlMkbCVHxbz
VbyCyhGQYOS+rXdXnNL2AcBCeVXh3waUSL4NgPBKbv7XFr6MGXm49AKKO3pRGBfEkM7PfmIfcmGC
kNZaBYGhTHA7qCfTKWXaVt6eDUprs0XVXSclfYF5FqGmdyerQYcgkG9bHIbcElGmPH8gNT/OCieK
MtEx5YbpaRPSV6IqjcDi+pRFKL5N2FflPkUfaDwnyXNvdw394Au95A96E3+6rdKq3zAYpHhA0bJu
lfbeQ/3Cn0db/h44tBQMio+GYR6sktcdokiUMI00oaemX1Y0scmfpxYnm30D4MfQ7fyCEvXvWYeO
XS9wiiDGSiZ6rtx7Kuw7njCRKOirSK741Or/WsJMizYuOEfXXR6pP4uP9GZNOGPYLT9aTDaj9m1S
IfzA8WdYGVEg37tgKh6WP8h6kf90tTxwtdDXW25qI2uKcTs6/Cr+LNQMrZuYGXF41UlMpyxO5/Dy
58Gn2gRN9ZvmHKA7nwLmInpEIncH4n4/wXJRTrda1cHl8Zo9XJe2wi7gk2nat/qRxEvDMCK6aFIr
KyDYvd3IKH6wtDQ4KHrLy6+y0jhcISRKfWhuvwVCFeRuL1cg6F13fQfaWJVpUPcdJm/Yci5tOHJ2
dmqQg36F/k7zsFZoCuIUYRNhSwFZbZ//8u116Mp7lz7xwpjKiJU9dNHkJHWQqsqBKvGu5ySwX/TK
K4B0zrNl4HmJUlfexNa+ww8eH8ThRMIwHcYk+4x5LliEzbeBdNTFCrg0xj7g4fGOhB/NEOOa6zAl
i/uMH5l+75aaMxC5KxtvwycJVN0Djs1KZHymKFdvXHmafONgwTXmw2cbZgztLXrMLRoO8JZBYuyl
MH3YAPILh9+VcwMFagE1bNbeU6ADCo1reJW/YIRRjSVLUUOrTr8s0LsrRBASRpc2U5ysdWjk0cvd
W9ZaQTRBWcSjZM+IAaNVCELUsRqIrX/J6SL7jI7eQCOj9WZ7EW5RUCum5wE9ChVeKtjKoUDOWfo8
W1+9qqDV6Bk2M5dRAF+WOXoKvdCRyiaWHMzjYW41aKau7FoNtBOuJi9R6W4XDT1gO/MOGPiVD97R
GVITCq9y8tWSU5ZiewVidarwMe1qCYQeu/M8ra0C3l15+tx13NagunbWBFxGWQrvQi+DFBho7Wvh
rB2Sg6Y5aRmdWo2Yae6pWjPotUf/ZAjVrJvkcPxm0Dj8JIeTtqGylsMCFT8x6I+g7y/VbfsQFU9k
QL1Fyd2FDGaBdtasLiDl7TPVvGV7E//KL0CwD0a9jn/Ibt2tLLqo1HGDJTIE903b4Hlk8JOqTU7D
0w6AFNpawlJz0ADtUWbmmUMnR5CRJvoohkmGySfz9P7EXB2Q2qIQoAU1ZYGfLDkQ69BAZaQfQEuO
gv/mmMSCc6huCubTsJjs5GxVRyrNt++ANbRLgiyJj1ZSDrG9PDmHi38S0hYnBfBHk98kRnPj4Mk7
RF2V48aL75kX3l6ds6cz+1GlzR9ulTnRSkwmFJqITthHG3PfQe0fc0kNcUHigacAGSxQ3JzV+bT2
bHN+9txHJpkOwkTFbVH4VhF8Wkp5lhhuESBmLiHIBpLvTMue69DNVwQ42mAFzEJdezjbUJVzJ5h6
jT01slEmtz/Os/rf5c3CjR8B2Pn3WnGKdNawAYbyagFtWHLzXxjEHS5PdwdkoGyaTN84IQ5eOqgL
YcqO8/mYOZuiQC4b60PFJvg6oZp0nursaq0dZnhpYVgraEWCXTGajA0iSPOqV98ojd0EBRGwRjo3
T9mNL3d6igBpGey/hSIlk6KZiuenCSTFerBjtPGzzJPotsKeOm8D7lQBlsiewzLZAjRdfBwgQqT0
NeKuhFaMU8f9uiN2oTy83rBhWobohY4okpuFtGtUB5SuT/SHJQtu3cZ0hv/qksvmCmeJEz8PfrsE
Veu1E1Mn3/O1MlvwoQNjP/nBOz9yx8YpCu/LXiOJkSFezRpwJZZtQoL+jU1CXothFopZjPeysXR7
AumOIGQmz4GGYNFVyw4bRmnBf8rpNtxvjFwczyZ2Niou2YijOa62GWVhj7LVRw8KCMQvCQGhBhQC
CLd7oVlcZgfrkldtiIdcxmeFuBTiaGl7toN+wy0a9eEm9RXHK71Cqa8accfk69VibcLgCEufJH9+
xVisSQPv4J4sk/uzwYcSvjBJ2qeePjQYQ9QPQsJOVViTYPC9rknULpcTrEU5JINscRIKVBACECdV
HqRyoiEhQDc5hkMA+0a4d3XZBD7+YfJwDTwV2n8EAYsQJ4cNt7gKSBwEy6frv2Xge6GUKdwT/dBY
MQRPAExdtHd9KH/e5dARLTVWoGSSVHfD9KFpv5VdinCmjRw35XJOk+KgBoWtGhTysZtJF2+28rb6
LF+VD+sRUIWlGnkBfa2OF8JuEg3u3QBm1dEzRjbraUcUbk8g1RbiN2l3UQgG876FUI+u91qt+4js
SNOaD9GdIFCXSO0RGNz2cdG0tYYOAyk8llSIJcni/SIb4Pw1YEY9lGh4IWiy+76zmye5DRTG+ZDx
w8SH/WRHIYGsi29StI7LwHJc+jqrWUySOSq1CVDlCEog+LpyQvchUp6XTHKBVIQyK/0pJUYLT7WO
CBEuiHZ348s3v9U5ODPZtO7aABN2enNcLzBaBhLWMYulM9R2JapRG0Hu2hItYLo6nsv1emhdBP3+
+YsgcmC69sWAKMGQ3I2r0TxbsJYl6bRpelbNvtFuyXQQe1gXw32umquSn4L1W85nqHguQpmuu3W0
hSjImjcK87fPgeE1s45U5NRyh7kgznp1OUXWIr7ivEhXlAazSIYjxi+3lX1+FbHyLTP4rUV8glck
6x9+pCTdPPcawrKvG2IODVAamGVnepgboogjsE8W1q2KrYC5FcVo+m1hxKgY8xxDkhnPe1og4QW4
4IQWjBE9OyaNWbbensH8o3ZtcWM3iq7myiPIzC5MwWWcSX5lh59pIcMDI3uUWs70QgUEddhyuNMN
V0EUALGZ3BotDfKlRmTSeVNmybPditvfX5ScfXg2FKMLppmq3SjI7Rlj+I1WZ6pm+k1gyG7ndkFw
K4eWSY+QMC4XNGW3Pt74tjupKeabjE30tEV8YJKViydGIgrSogGqGl+gzGGgVMcg2bdf70J4Sj00
cZ3ZOTJHv6wThPOm3gXmvFGrE3lqpJRRqbo3g9dOa58UbGGVeNWATXuezewXi2/tA7X+P+Moe0aP
EKjQiwISiDOCuADB5WBpKurg62mE5tbjglje0ebGfRUr+KjBqeaGFNh0jxJuwf7HBeB7HlxFxWrQ
iW+5bKrtCgySJ3UcjJAqF0Cw3c/gY7P0mZf1t9hj1uH8xoCGtsgXn7qPXA30sbwcGgBxWR5MknRW
9L4JafQDHAJfxC8GDEOJY9TECuQ0i6/SwBZyh2WhF7YMe1eq+ILxyoVIfVUMt6SHNFc2H88Ewz6j
HJO5po1UE4qILhIFuRDBnrODutMx1x9jRdfwM6TKVcVB+YdKYcbwzUp544n3GyDePQfg5aUEyBX8
vZ7k33mvrYTwn19G5D6B34m06nqlAPXxjtxFxnOounQ6k5kyOn0tWOLupJQezG/M/5ELMqhEE8IO
/y1J28rb1OqMK7nFaEkvTsCvAKfGceoqRqX3JwVI+FH40/S2JGVGBsxO34Yg4Gd6Fn0X8vjY67qh
An/TA5/te7hcbpe9+0ArSfb48ptzJVF/++7KwnKlq6IGcahqycuLjVv4OhUhCzrNglmEnIOgpmL5
GTtfMHC0V1lwBbQ8yQzMiqIKoE+xlFlsJUQ60xlWsAj4XcmhVlfCaXOc5iSqsMeAZ79vGh3A4n0F
UrZmlBVOI4RlfxEql7wr1msvxAMK2mVi+Cx2oOn0AH7jUZNP2VYr/z8LXwNxqMAJqCmyfi3rvmUE
Q2t/wlYsVUfx+xFrm01BdTpCRw+rY02fIslS/dPZT2m+d+fIkwVMQ9D8CsERe0pL37JPnucVDeRO
oW18LeAaq2U9HveZiHLuAeovQjEp21azSmOIGPAoBVJBFjGeXhCO16RM9+S0JoxbtI1XyJRuFWru
pJt+5HQVuVcvU2pcXV2eWtljWoQMLP6wbFVI/zzGrgG675rQnjX4ejZWNYcuh8KgHkJd+Uqtm2vv
6kyh7N1aKuDGeZRzFfA52Q9yPG05sqjngI6AUz3AHCJ5SHMuaWA8d7ZwRCyinBbghMD0paz42olO
JUVpMWW3TDTe6CiX9JKaOjQ/IZTBJn2YtBTwl2mlpqrMhCUIYjsjF+27mWU4MxQPV3P60OWJGoK0
XUQ725Tbzo15yc+bh22Rm+auZ3WCpElOVG4dbYZaLDiX6osd75PZwqYSMiMhmjvMtBEjwfrGFqo7
BPeI2UkRGAqkK0yIGPXRCrY0t92IrJIL1ziKKS0C/3WGoVHjNGQqqCYB3qKck6vJr0+3siIiiVjv
BnfCQsTE+v6iWZghslj3ikZObrnZKRSUqfdSiCOBmFCbjhEDhQp8YptfyuoT9WA3jXHt/WGR/K6p
smIWm/jSK3oVAKxJhyOCjWP4y4ixtj7ejfDeVoFjzrJvXb3XcsIdewuIY5GOdfeZI78jKkef6lvP
vr8IozNEJF508LBpryaVZ9e/+tye7qcxBz9SDWT+TOtlw+EY8TOLv1xcsXZr2ADuIrc9efhevPvP
NnJ1L3zHj0YFR9RKdHaDf92czeN2meGs39N8EtqAMYdDbzT96Hv8cNw6aIJ/cV7qEJK/biZ9rRHU
Mb9lSxn4WDPj0CaP17KXrzY9vHkBacdW192sbN2FFnQS7lxdR4+eXZEx7G2p9jRJaM0bgWKPiTCH
/7te2biXsFzzk1C0eOni0oCu3WeV2bWR1XruECb/5Itar/3bJh63Z0efSuUBYGTcxsLrXyckQ6Wg
GSvD9xFe55pyGpei9b+91OlHRVD0vhhkMfwrz0BkmNrDGdyBEPQ5ULv7KO7212kSQ75wPzktBOVd
6oRKFXSQyPCexw5f5kxLxI7pG5uxbb/AtKPt+VpibYD6jM244CxHbIftt17Vk0WlXfvlEm9h3CPH
CDOls+vBjyINpJcF+9XsWRMpkn5WnEK+KMTJtNF6NWWpicI3pOrmt0zmkI7mo6O5EPF4xOE59kCQ
H1kFdrzqn+Mi4+MaHzGPbrtPPo72gkIM9J/+7NFfNWPckNwzrbtl1hhRK19ah3UzBP2v4YeI/WnI
ZJvNEw9EgMHQlqKTf7P75ChhllxKT5O+pxIqDBWs5tigE72U61Ds9TuGjybj0hfl7phUsP5Ai9Fr
dwJS93zBXmowGDmgHVEZ27QF9DesZhUoEw9jGaXjssDonegTAm2Rp+q1i8brWyZoGawjbUtM6Adh
Kilvm8WMZHeoP/uV5ERBi8PfCB/MScTU7cyXtgmF2n4pjBQo36m0SSQhbRQPybaPe3ybTyxfBOag
5/j8oqaY1ZCsmX6FXrdjnDXu3ZnzXbqjdS9SPRBgLiGX5R41np1jyRsHQ6EHCCNSGNNtubeRG/3/
eQLo+A/afeTi4P8Xw5vPsxmhUJc3FV2FF0nLLU6d9G+u3g/dMCmdSMkOm8fGmFTqgSdFAGjit0gQ
qedimU6mvViGAQbI9XRrwwVR8gKxHwPg2d08QPYIdwxjqW/L7Oo39iYqiEFajS4oj0PbNGv79ah0
vxZkD5eK7puFwYwanJUD50J23wPqUefh9QZFQpJdXJ+7qSXsuOlcBgVSQ3W5cGoOpKJ/wEDcp5r0
Qtk2gD+xvFAUe+spfZfTyKLdg5cauqeTS+7kP9zgd8x9+oEvDFuMkmICQFOLWy0Jg3sdym2p1FjY
wzjJWYsKadMVYkpHNYG3mo6ofa/tqFRR0WFu4uEcJreNOoO22NDwEHrisp09eKeTxqbH/7FKJG1P
GiT2DMsS/0xjk+J0T4XmfkS8Dc09Ty0bT+dMiIw9SfF89vqHT13nhraIHTRSbbPJ1qDsPMJXHwpc
MwUBoJx//IGCGa2N+Vkm8Ir47/mHkKHgGvOXsS0LWtMFwVlmx/SMWyvcWH/SJ1w1hUK0Mr6Whr+V
UtS2UVecMSoc8Ut7wZ+LSO6bfyRiWsUzPOSU+L/rk0AXy/42OAz1W92zTPWuATF2Xc4k7uKcp4rv
7+PgmP3iYfiSBMtDrZg+K97A5hfIPeXkur/v56egs3R6lgQTN6C6HFdHRKbEr2PmF7yAT6s0i7Vn
hlTmoAfrU7no5i/Z6hNZwyrzP0aVRDktpE0ExGgoSOxHL0IrdQPGTRQVjL8rLbaYlDlXnp7ZM9OQ
IS2VfH7y/ccN7nCo2UAMXqmwb0VeIhDKKo6UOKb5cSyFLXV8rb3FJGFWrgSfPwAeCRZYPKIZ9TP9
jxDo2ShLALfiq/V6FXONu8U32HmIYYgTGT/K3na9lWO7t+EhxAco0k6UfAkkdvoIPHdDsz+3MzDs
j4AIS65EQ23luzVYumAP+XnXJDDGDBmqI6Ys/U0eQ4zXcYQTBLgdEIhJaivubzBfxJwx+RpwkRj2
fXf/Q43BDnuCdgQs1YlAbytXzY4qwm6T+UAAVaScl5usy76uy8i0KBZZVGT1a9NGtEoczYhSmh7v
OWAlAnb4xssUhsxXtRMYZ0XmjNXC+Vs2t2jEXVbsOPnuBlEzajA0FxRXNVdZqJQ45y9kfDPl45/n
Rf2Vc10q1xYSXOSyEZC8Nv9Yu/mS/+5aIpCC3MhoE5mu+jg9jYnJNYl7CGsujrJ2afPMWD9kqa9K
vtstiWOPt7mczJDwsYhDLaI5V8ezfLgwfvlS/xjpnHtfvV0Bm22fd/0SAc4J9dRYS0Ildh1cAEj2
eMAaHbY5tv/8vuxhnkOKqatvlgpJlcLZvdlSD5bSPGktcbzi9zXP7yHQXhLWLKKFn8USpW+xvkXL
1IOLrDP9sPEjp0oMz1Ksee9mK1HYTtP6SwSJYzMWo5Sh6YVmBWLk5F05owLhZCZSUqzETfixgchl
4Bkf9/kOdyFmiRSOBzxFEfW7GEMJWAaOxFP80k6yOuV0X/rpOdgZ0hlVaoV+CBS3Ge4ysxcz+QNz
b5CDDFBCu0mnI/bx4sA/p2IysPB2+8lQie1sApsbFl7CDcmzAdeoZKcTL091rbwFZaGAr9iI3iAd
gYo6gUeoy7kH5givO/RMHK/NSFrQ7p5j27gMmBth/MJTKbCVBUU7iPzPfffX32GQ15j3pXIsGTfs
eylg2am+EclRoYexRngINP7ii0e8FubOkUX0WkOqrWY67wEWgnz9yLKhqfDtwTm+3j+CuxE10yzn
P8pKg3kywkxLVN1ro1LKOpUHa/I0WrkMCsk+9HQfW4Wb/sSkEDecsAFs0Rv7J7HDxurwwl4almtM
eAB8XM59CArPKexVNP71SAIawYT7vPTU8Y6fNMyNHGs9J5ou9KDxFnQ3duiev2i7QqXwIrGf9xmv
udWBjNhDDV9mqcICZ3oXo7rFlne6Vuya7ebEMnRp2ShVzztKlrljfKgRkka4hxhpQA6yKLVw50sw
rWJwZ8GlkYj7Nok82NfP4cKN3eOGYBNZxNQt2WtYv1eN3lU1Cr1tBJBUIMdnY64nqJr+rG9hgpm0
9lDpxV4SQmNZ4kbuSUEE2WAPLs4O+82Q3RbJheR8uVs44ss5k/HH4LTNM+r6oNB4NcqZ+e3gSU5w
4pOJywrkIrL9fVyP9wuJB6F4YSrx34QBZmade6phHTFIA1+m0vPtSzWjig4T/8yGEmLotPLRxezP
qzXSh4tkLnnnnlhKluqHYLvWy1Mc/jcZTW6daBNkagsgna/Ag00kUszXX8CT28y3jJ7PghOzmeQj
1tfmzpo+leK4nMmXIC7nCR8uezjw4FNFSPFyBoLhblWY6URYg9xQm/2O0fBrlPJwwPqIrBtzvuTK
uNEmZW8ObUqom/9+hy0OdaISqzsNQ84fISyROBDNQ78N99s6XuYnrXFQ4uKOzYQ20qXfk4NlhFig
Em7NEx2ULQR47DxCYyYgqpNZIfKVhYn+UNxJ7Acf3CQxgwwlh7ksx6G5/mc/MlwyhTfSohSfYTTb
KIx2+NVUB1QM45Ndfh+Cg7D5c7kDKDhLQUHD2nmHGHXa7q9thka7Nohs2w94NgRTdIBmBXM3r9Dz
30/M8rxlo9FdDRqKKSe0cVtKpq1MJtQIXFwFgJujhl8kcwnFx8XWNCDBC2sM85GMaBGUFSK1QaMM
Nk1euUeClTjVGr2EN8BrLJNYzpOZ7Zv+MGyXt3bu0HYNqcnVpqgNnHEXLzcgE245OoQP0H/Pi7oB
JfZbFUOaFkfmIh1KDsfhOic2zP+8koYW/SP7+eh7fuohhaebUax3u8Pl3a50oR5m8nezSf9cjvT+
jd6QWCq1vFhYRo0cWV0CWWClakziOx04nox2Q9h13YMyfw+EJ/Jl8MIsyvqefYfmcYXvMY6zjtEU
KFd/4g3hXzxdek3nwvNJvN6oXrrwDJCg/UbJo6HAIkKOcgTylmxuo0vq5IoGoWLLGTSvdD0TBHX9
tqlJqF56153XPtCje9ZekEbq3eBjxV0THNrvhV6+FCX+GrbnOesSfhHiNhOdPYxpqsC1BIkd7CIN
2uJTzt+tBv9XqzH9TdVf9hpda78mmNesR7G0Hr+PVrNmx436vHzDOdGDPXKMfkw1723oTyyiEK7Q
EwmcPkDyhpWCCfgpWLVSQHCstGpZY/f8SUK5Qxq1d+z17eXXjWaVJHUMXEohJ5NQghfxCSm2F0+E
GU3LtM6P1daIk8q6KYqsbSY1r83JM0mJmhwPjHPHe9jroCLyz3yEo0ILvGbQ44Pw1wnXtjjRfSTa
5D4bCDcrQbrlzjPMqGUaan4oGLb9mrtkZlpQ1NbqMsAxUm1R9J6sUEYafeENR/b3M6lJuoN8dDXI
4mNUBWFlwkQgQpIhgdw9MPiFFQr8/+ykZnBlK1gEFq1rjQ2/Wcrunw8YjhTn31itVh3glT+e3WX1
aVNfyMcspWr61c5Dohs6IKNidzd2tHRjYaSJexK4IvQJ6RjCaXAMpH93vJLPMfy6RN6qerBSCLyP
/4WiUEAKfwJtvtYT8+Nn8434pwroTWcC7dJfeOKE12/yboAfOae5ky8ZyeaVg/lNV0Fm62snzEQJ
1hcBCFAZ47tLAjiV9LUnppWCi2Y+2W3tE9DSw0+GnLf1uL5crRqHlBpFuR94wIeOlCdTwZv2MlvY
oRFITstyZAwN51f2ULU/OSUjyNG3O/zxPfs9YaC1FR76SsFsuLcuUch0ce+7b77jBhimJTgdBjcX
HBq+KiD/ipmrBnNj7JUoCc4PVAA0rTLhm4cQ9amhnmWWe52j8M1jtYwhPLc2DJqmb0B7zADjtEsK
9aJgPJ49ciQwsNYK1qsZ1Mndi7xA8lTWYxhgefRjG5GuG543In7ymnfakXQlWsIqRbNk3g1OEinO
4pS4dJd8eRtZM61233gMZSx3LtpSD1utT04hOlgDykUgH6oTRWO4s2FThCYaspWdb8AQ0/xHs7aL
yfzr8RtXLxOKyAZ4eHSMba4WZvQTdm9GWEe3NIs00q7mBmmXVC+3/g15rqAqZ7wtL7jJ+M+4SXq4
i6U41u8QxIcFdib2UWPLDbJVHUPJQMZX2Cod5yZvICsaflauI5Ftwr7LpjzjYjpXF4m/L1nyjjFS
g+Mh8ILrKt8lr7neZrDSsX7y5Ys8gQd4jN5R9VUzIfu3fgxiF9czZL82EFSTQ56jhje7KzOlLJk1
7pXczxeUp73jnB9mkPGQmNIn5/rrVkd7cGcEr96+XMsKUb3XiKgNattBH5pg1mBcOC8e2KocAffz
gHgq64GB2OOgcF49A3qHim8nbrlMllfSsXNDvnkOTvuaEiXo2cMtz7qi9u5di6zC0bP1iYihETWn
9pE0UpjSzb4AjB4b8Av6ThwKVd6ClR7IOBSPs6LH6cWYBVFpe0+hICqRJhjPU1pPngvENCtdCIHg
lWKfdqNpmTuw1LJwjeIB3p9A5cJcr95Z6a7gLEcCldifuWT3s/EeNcR3rf2fvXPWF6iYEm6Yetvp
bf03TAiAyjWJIXCDC6m96Ah6Y+NvZrV7IrQWdPGsT2GRtaNOj7GvZw42jR65zp2bKQXRROy2odTL
uZT7r4eU+s1fhtmK2tPKm7Rc5cRNn4CHsb/g0TL1htCtGd61ADwe3Ne4Wg8v2msFy3SRRdHTPLUV
aaR+pls+ZZ0/HJmvxnSqjz+bOay1Qe/3jE94TfDLhx7zZ9B0GIyUgXPgXNsx00+nqNtgOwhIr+yf
HC1WWU+FE43IUtbjKnEaOowcxu+FNiIQHzPvL+wXV4O/vgwjVPjf040seKJFgRPctqKpKfOFuDjt
Yh32vfZ7jFOwIEh3DnM56aPbmbYLSvZt7ucVSqzmYXXJfkYfbHlybWaU8+urxnRvUihQUjDSamfA
2ekWk72XdEX7cFpWso1HFJQoE81/t3FOz+m4C4lINx/38Ol88bnkuNnBPtXde5AzKOG+i6sAaIe1
79gbnEVY8ZC06QYXeeMkLlIo+7b+YARIF6wUTEpKDCC0pL7IACMrHIhJbeCLpnwKQN8342Ha3JOb
Jr4cjjpcyAn1TC1P5ZP08Kk7jq5kul4lQGg0IHYxrwLqboqzjLWq2/BiAsHLgoIxkb0W8L0RYs7j
qtHb4gS1H4BBrv1+sFU202WPm74pQfig7DZI1ywmbDjaGYaSjRh5wVAOViWFZ6QqtLGtDbcHILbB
NrsV8lMKM/kU5kZ95M5sqiLaM57S0IsH9w00BuZKblJiVPhxXMNyfY3xlqZmn925CoeL7m/7dD52
fOSpsyMC+Gn3y3cw+UWrQKP6SrJQC98O/xGjwdmozIh3IPtdWlek945Odd83YEterVkgioG2VGmA
X3a4OVjmCajGtpoRxFRlQnup0dIzxW+G4wktBl1fe2lsSarpnbzDsupOWgM3VsB42oJH/E2boI6m
JImvjy5Tpr0C1yMHJrMMcyOxqeTAYkj4us07/zOISj/Jj5XtkK9zNb9kNq+XFiz2p8WWiPkokTOC
ejxRkJpzEm4D6TmKZIXIjc8/rdhaLYuoH5chPpL6FRh8G7kQ8hD68qH5T7kEvBI/QZjSq4nyUciN
Mjxzo91vpOF+rkK87fMIdkV5cWSTk2dmej9Aheui0NRPf/3PPTfpeij/N858Fns04PxnwxM3Kl97
MpmKB4ukNsb6Z0NWnbsHXQiMuumt7xKfKvDzyyHI9Femafw6WKz5mgfk6uoY4sq/Rj41eTwxm2D/
vJ8DXJwxKYEDgotAUKg3jVMT2oj6/l0Pcn4727sA8B7DZYunf20TEaRFWbde7Pmj/+WjKm9Gs3Pa
+VQ/117qWqNssfQkXUgkDHl6ZWYwIGsrF8UHs1XC8NDVHoYU4qf9bW6cmETFVSmE+Oqb3om0zP35
BpjPL1+dI0gRoYRZ67ghNS11evFdmddtBuky7uCz3FEqGwDzfIgaauhpYMdCG04v2VK5DmF86PCv
z6nYAIWMhdTXfRASYipRjS2RiUmbdYgLorIaaDgTt06TcNdI5RMBeexwEY4ckPaw/BHxkkKu56S7
L5dI45hMy4uRcuwHJsW/qK23JQg53xVKfgu9AFlAkptTy5AVQy2EG9K+h6VwoH6NklBg0QeYhLeW
8LKJQt3XCpheHg6cRerHnoskO0hlX/eRZPni/mT7kdLXdA0FoNH2BdeuApip0b8m4e4lH2RvvxV3
Vg1wVm38dRSiMHBq3CIUKwzNOFtU2PMng5mpU5YSIvZUWsW1Lmz/EkOEY4lAQFx0vaOPiYiOUc1J
mudCLcR4sM6J7ktq6IglmdR09Sc/8cVDwpnsVP2SyuVNWMm5j9cQq+IbbxBxxi9wOWwRQEGf3g9C
4zPAZUSziX+XHU0GxsjWa1XGBgqthKpP/S4aXUkwnQXMeLU/pe+GrAt23i1zT7DCz9rQZ3ESxPsO
XlOXHzZRTvC2v4CsUhhz3vh0sel0s7wtj5b72lEgFxmyf9sFMcghV/ayW7t2Ts2fH7uHUu9x0/Hf
zbEInfEYTBCR1Jo8a3o7bIGC+h1YV5TJutirTD+PrnJJ70x+e4OH+6KRURyEloL+D/fYiWKgi84C
Cazy0J4xy/hDCkl37vs/9fOkWbE/lhpVhpaGZhTXA8m2jUytVnc1np8hpt9dRcqFEIooGik6ut/T
nf+xzWlqdM5nYQ1ngQeiOunKvybj5KWjg5Rqbu1+Im8o7XJM2Pluvp43fpdqDqSL1ty5bM2RS93G
pRuXJZvJE1WOAhjG4sE7eaFUg/gwF3838MvfabKA7QsNgLC87YVUdUjvd//MTUQNTW+6Xsl+0vIw
SGrL6qDS++428szO9XhWOid1FnObICOSAhLeP2F9gcMTtIr8X2cgqF8ym7diFp+1ofCIxLKez7Nf
F/WCFzMYrqEF/sJuMPEMUVgFIKCrt9J3EUZHPAL3ne1ZyGuyIGJFS0nUKLJ2oAIqLA+SkLYQnELP
E9C+8phFgFiHTU4lofBzF9r3/PFvs4DczMUJ5eaaA5GWe38wZWe5V3DVyUfn4ABH9061flwkEDnk
+nRzKs/k1BjyBZZVE0lbkFSG6ydvzByF0nE24NVz3Vr8HsutoBU6lX68QbfovvekmrvAOqq3l8Ei
GawUJwyJ2til9bHl7qU3T7XfJY/IuGrCyDnjSIp0kbGhyNI3w4XuzOX59NlhPGiVpTVKejWM5TSa
jgSeFF6TijE6ToIT4zpQhBrhJZFWB8yEEdGrG/T79t10w+xpr1zaJQjI5Wf5K2cUHQPyHvMAbEMo
PPotyMAlOu6EG4UTAPs8ss1vRuw5BlBQjttesQsczyoQznrnfk7aOeQepmim/LFtAONw+PVaRIJJ
07EdTE1yut7PFKonzGleKHF4svOGr0zEBwOle/B/uKhz3i9j0tPbzOCMdYfFZvFgFuxe8DDGgUdY
V00yhZ+/OU5gEviIQ8a0UyX5G2L0ru1lpSoAFuHl435IZ635M3sIoYxzLFw/u+Lx4Ieg4Cz5dB7/
KQ/rSNSslEfexwbeDMgYmmejqRlU6p31dShVPoaqesHzn9BkU+QYOW4y1eXIdI0ySaLvb2GDZ4AF
TeAr/r8CUQvG/zZGCjHEXQaFjRXUhv5OKbEh4UGzTB22eBsyxxxb/1f84FAG8MrKoDMOkLRqiGkN
KC0l8QUlsrVekWpYosP6h3V6kg6TNRCnV2zkEc2OzjYe2UhgftPYS1S0thpVka88R3A7CpZ8rRa5
SqtBddz0aGY2evwVeLbpA1yCeo2J4RLLVpySdsAEBRBqFSkVwjavUFSgjGeWC49Lakl3n2xfXgTn
05aZHVeUM6YukI2+TS7UypitEBDcEmpGTuCc7iOIZa3PtYifQdwnmFV05j2ULLC4pz6YLG+wK1ea
/IFGloTOmTUH0cpRfRalmcEmP/BGrka1Mfkj8Ysc+CQzEorNiXndKhp+wYKlZ17U7DJCNhkJ9zrc
CiI54fn9TOrAnHzMygwJgdaewXb0+tFSfvSLhWi7c2+VeCPRrbl+9uYa45FGZcNkAdvmRn3WqZlf
Bty+zdb8GbkD26HR8RWXwAO2xhzMhzTV2qgZuZwiyDZ2qSMaag5pY5BoH+7nER6ULMiYyhLPkEfZ
gGtVQACWRNHDm7OZWIDHsyiZ+bCjG/w4ZOe3VnD8v/qNxVvAx5B02gzACikryoT6j5wrIKqPGGER
OJhcFzkltc5wphsIWZURPQ+FoHbFFddGz8TQXTM8gGN4l4Bxnyqj+qHIvkLWIs5FWmjh39MjuMP/
SChJ/9OHuD5gANJTf3+T7ABiYGh/eRycu/YEEh4lPNMmaR+x5+to06oR0ooFpZyNw0250sU7HEI9
8CoTBoScOCE61eTslJkx3C2VCtuZwStvvkKWRBE17LvtzFcbnmZkh3VAtyPteJYuC9zlaVNeio9Z
iaY3ofiHg6e0ICyVY7lvsX9qliyw85nlQnsCh82fGk8QFQ0+7XlAUMsUe0ydkR1BXIoK1tdKj+kR
OPnLjdN2o3jJa0A8hmKxA+0c/vFzdPxIKRBCfReKXWPowe7wb0tov9Yjv+LRVmDQHDzFf5X7TIeI
JpD7fIv4ytSfnYB+0LNcDr0w3PSKvya71/ugan8Ybzi8aryarVUx72RhDdF6KhZtIv+8v+IS7Ym3
U9VbyGF5x/ZQ86W6HQExB1eq4dmDacw6k/4F0J+E6ph0865Jug696UQFH8FVVsdlyjyJopW7bB7a
zKfZL0i0nsvLgq0PjU61isifp88BbVoHXUu62VJMijyWzyGzxAw4ZF8QeEpYRbK9gWxRPn8D9cRQ
0k7DFKPqQZcYdhbCwlsmUIA7ze4pqSWgEICcsyxb+Z1tv0SPc0u60vzAzkaka8gmTZuXg9L8AzuM
TUKRuaGZ9VuhHpGIbvClA9aaowLsgQbgH9k7rojUy8+U2LQXBRC4zklr1jfQNAr6pQKM1VALg2vL
7ezPWIzUgqFGDuf4X4PBW5WtoHUQCM9L129NBDJlz/GnjCyO2xBnd4p0hCsk/t4HhkYRxPIfxXK0
QD73NQ2VHlg9ZpDWI5/jRWBXK5GBpINrwcoXR6bAq/LBLZBEyzCs7BMzls5IxMokJ7AK15FdAOTG
MIheaTWrZ1/LMHeDgFAzOPlLOe2DxYlJ34qfabO8F1QehooQdLxCPaO8GjD0BoNB/9KYiCN5DC9B
a5Jj0Xbq5ww7DxNscJW3YYvpgN5deIaPCv5SGObdl3e6z8l3oLYcIpyxCQzXHHx41aqFsvQfWOKx
7FquN7qp4PZFXpr0Pwne40Y9pnQpIVZEYC8V/UiONzUgZeyHm0KNCqFntQfMt5hKGlpWWge6AuZv
zFgLnYCiwc6hJR3QzibMmeY0yEsClXSXHJ1AvkMl3hmgBKETJc8j8YM6dRQw+3l8tVAZjpzqMi+D
XIcpSZplEOB+fYBUmo6BpC78QGA3Sa1RiNET1rOjydCZRuYAf6w1bApFGVYNzUAAbl4fSMvHM5Bm
Fo/D701yaR5j+H5hJw27ZBQap055KCgNKFKR46q5bDiGlKz1wMV0EUzYj9r+81oZN0wPWY5cDX1o
7eA2zg+GDGbxU4t0l/VlP4RgSB3MM37PCRm11j57Zk5Cc04rYmPUFbV68vSHy8b6OvQ+pLfDEZa0
lPHdBL+uCTxAlgLDfa9MXXvDSZ+5HPIXyf3BGtKJatBO0I9JDInNQcCLDTEAybwUY9GRqyUXu7Qz
w9oaUheVu4ewYjjvHhvLh5yfEP6ioEmMYavKCbZOG7Y2R6NV52Qo85nlASNEynBOimkkbiHTgHCN
0SXiVcAwTzJIuYNB5S7qxWtM9lLYhu4a6WDZl2RBphPiBwpUFkIncnmXIlEyx5dJXWyFHYC+xxuD
d1WUACfYmm1vl8PBQOiwmjvx2LTgeG3/z2r7s4M4t5+km57w+Uh4OwkSVqSFs9rFK8hrdSDahFzM
+svkguobb1a5wAdH0vKb7A6w3ZTgkUOxUeP/Yw+sV/cOI5hDytXwL42Vxj9T4s6C/ARRCg/irFoZ
lfsu9tISzcHsZFVmWFd2C9czbYvm+WB168kYMJr0I3QB6eY/lCCABYJ/OCZcENc+tVACAHHqT4Be
YDkhnxCwQxwglhqM9NRXu471fPO8RmP+e8cLziG8Owb/Y2MazCT+mICTc6NNYZNKydaM2ldBWQSD
u/Ai0oJgxnL17liI7thr1lJBp9pzyj2N1MpV6bdy1PzqHyU/Cvc1V/hCoHWRRxge/xEXz+74Y+hJ
jtekKGD5XovAEV92rpGCZ8ieW21cNGq9OQ0Tzys9BWj7LGHafHwhVEat7piUgApY6ByGiBnh28MP
JdHWpQRnszMFWqgb4KuFpXIyBqmfogtpfgVcSOGXHVUHbRo3ls+61TE6TaYITH0LH/x5IZhJzlF8
kBpMTYLlzBxxmps7sKSR1L90FVofDkT90sl7oHdFecsCEOzI7GPBuStKNCx2FdAWVPVPx5jra+0+
eSnAxh5HF3FPxzwdCI4XH0OFIUfxAlGpI70It1AlnutN8hrvygVplUoCm9FqqLflyKAVhDoWa7pQ
7T6QLJWn7Y0Qpy2m3tS81AAxpa3SjxyJhzT7IXjcU1LFEQ9n4cLykoAGCYGcFDvciE6MIwKIillu
4hQO9HlRMUoqbblEx0q2EYpqYiFi+PLYHD7AsxZ389EWUbep+W+yIpobb7VNgAUmB/rHXuulCya6
r0Cmo0n2+rf9wZMEEsod/PFmkBJVSvOFoEPwgY0GujQ5z+mHMDxw4GVlCpcHODPUmsUhwwQG/49d
N+uRsVtv1Z3u/nIT2K+chW7h+xt7y7PnFTeByaySzT5N261o+amSkqX/3s42SEWG7Ua7dUOEHkhV
pw03H3Mk5bT5lTtqvvu4BOlpbypRo41H9IeadsFmaSwEFEarn8+582oyMT9j5a4zXEnKBRgnhEb0
00dZSwDCef+OeuGkZOAvT2HPEydmsR2SzX0YDAio+9yXuP0mI06Rf74D32M/ZA4ezjZnARel1n5Y
64e9DMEx5X5QgKUJV3kNEBDiYmq3xl/4NwfYqPSIlNb9EC3mWp/LfXcSxhcss+Dc+dex4DflBDNr
AR6YSt2XhYEH1f6ZrWwiU38IdxvsPOup13DQe6/5iz7yrDtqE87dW8hAESCEE/7FwOsFsWE62VWG
YC8FYs940nM9euITw0cZs7hdOAG/tongh2rwNjYkM3/O4bbpVYoIYQH3oQ4GrYAdE8+cg7N6iwZS
NyB4TUoUg4Q7jUUVXA5zO+7pX6zWVW+S3EI+Y1sSO1OI3WB50NeS0nBz1WApG6dINOhIwp5lL8mL
A0GIRMy8f82kytsSmTyUSLqx7hGEL+kM9uCP2QNLqK0KsEdHI78k7xGJOWyzvz+TyX9yclnKoyBP
mlTZLHq3NuB+5egNfwPJMgy9Akbq4w149Hu0YIf0SO1hyCYesmkEcJpXrQJMcFHJjVWpJ1igF3fh
uRN9HZXfO8QLDVN/Jj3SfHUnoIARtYPdphlRL0F6eTKg4lxAG3qkW/amXGdmpDW9dTf8agX7oQa5
nTNjj1jSd8eAOv/biStGtnh2uJE58pJLSXoZ8J5sTIA2MDK11Ybr8w/yTWbc4lEzoKbnbvqRSooW
LiprY/4I2RzTwCM15RkLXHdkghGjZ2chEl94BlueE2Ejr0Dr/rdMvvcs7+jL8vN+IrrV12vffaiH
eyLerCx02xiOaVXy95S1HO3cAMxRsF2w5/QO4Wp+vPmfUNAW59VJTc3f6W00kQopE+m5hTpejh7S
dw6Ondbmt4L1IJbc/LXcP7kmlMZ1VZkSI1QMWlig+TZU57TH5HQuJlNpcn1DJmmRyw0wE9IZcB5s
95YyXJk79UjyUsTe2ZyvfKbWs5qZeKDShV4roWfhqj954aCa8S66mOeZfF2iQw/ZDyBYUs7EuhoA
wIwSshZ1hd0Kk3/LKdhJMpbJTvQRvXnPkS9VTeFIxTQ+f2dzXjlh9aRjlAgDKT2BCy3GKVS9WuET
Xl2HrQtiW7jwSgIOB0NVyJKpvpM0ZHaDkOFm3Df665P96fpxUylhz99+LXLA120kBmIq3gE72iFR
BANoRiPtKkBbkdBQVRnuOX6wvnJ7/rehQ52AqmMcIvM+rUc/tDErdKHAQjH4/ePsxXHYh/+KJcG+
EoWIsp10UiaqKfYhPC6EoU53i0uur4+46Jbd/m0KTJMZqTPEnro/cTnIsPcrPUzNGQK/jER1Vlq5
n4qaTGH/99sUlX4zn81e0qNLpr1k+OhCnMrmcmi0CIVkAj93vId6fDc/rCUng4XsWKXi01GLuv+M
3WkG7RQ0e3qBls23pGRwsMpTV481wmG4cxTIOeu1paVELiB8VGF1FB1CHDbUwhihddLcSYHKmlUC
z/214OUQtglCdxpCLAgFGqYXWyWLDVKfoQu0mxVJRXyyvmZO2pmD1IfdP8hHFrKBiUUOhiblI6JQ
SRh0jbi6oQ52uO8UVIn7O5wYwY6qxONuOfI67DLoiQCQJhd/pw8QJljEQAXXlR+UeJ6ya1YbJaTy
25jwl0+NBUyUpxw3UQpNNoZ7TVBBBaPvRRVedSLv6bmoc8DAwlivgZ2YBSOL1w/wHop1LlWXM4zL
fX6NzWgCIF0mxAM3wZQhLHJXrpgO9OOVmym9FyAQA5Fdnm5I9TjV1vMRURaL5twq55NPmH0Um3Hq
Va5RQQG2wZdFLq2ksyCa0+GkjWL5SAVNJRKgGTJRSDtudaQOUHp7CAWCfEjmkDP591YBLn4Rcv4s
riKl4CtwmjpU3fr0KsJbe+RIz+2FLw1F1fxLZ2MpYM9vAYOZ2Cj/BFMDx4SyNo56lNyZVEC/8hJ+
avdBAUjU2esv1QbtRPR5+KrqNjQCxGKPZ9Vp0lt0n5XVFq8pC7VltpngJdj5q1fsV3s0dPGwmSRV
xKmY7kcFPrbWhYBpTwjuaphM0uz6VZDBdMPsQtXgBHrMPL3+yF+CKlxAOlbS5AsI3Guj3sJCnL86
moTyRh35lpsRGkh/7agvDo7GPHQIyIa6IPDmxC3BpoTatA3CuGwXxCKVza1C6aArC9rmdw/JQxps
URpZFHmNvDqo0/A0XC2rKRRePP0go+JHOBfUhqJkW3uqX5fJE3mcyf5a0l7DqTVnhdKtLLlKrA65
fGn88WJadPNXew9xiJkUxLKyyOEOFv0FJvvPsz3zUJREFG4sac9uUfU6IdImMkcMW9P1qRx7Lhxd
C7pvzJjJzbTZ1DBJYI24DwzZiIGE3lXdE+8KIi/LCpvusJGB2ciJBISZHJpQAbqReo/8WBPswycw
PxuK+Q4udB2rpUuwmFkIcEuc4BPJYccbJ27xGq3icnXfWQOIScQqMdC9YRZNowkoywYdvyFVX1Dq
jogZ1y5V0vFfzzodPFpuVECSgqlL/Gw8oVOkPkMMF6oje+gCx6OinchH9/FBWu9V8ysT/yZKqcz0
Gu5ETGI3ziSvPaznEjeBU31ACcu58PDKoslPT/CYEP+kuRPVHhHlDC8u/4cn8oXcdS4g6bxTU+tt
NHbfYo/z4v54C826xDaM/Vg21I14WY7jhbztMYF/M/iw+uF7joFBb/+h5kNOjAXeJNsHF7fTFuJi
fMOHtx5DHy0+f4BKCg/6Kjx6GeA2a1uEl+gvoKfL8Y6ABa/DlLcquWC72VtR/PfUbyaX/2l1b6U3
iKuj9a8z32+HwmHzBME224ySRt+NFzS5pewdI7GuMk5mryrLZuIe07tdrcTcXfcYBKxaZQyMpz46
i5/aAoMGY8O5eU3hejZYmGoecz0w3pkKqEUTCnRx4ahal3luclkcW5oKB5G3a/gtFc6JlLJ16ZNY
64DUkaETcNHpiJb5kFtIU+qCE7yMYEpxfE8xtjMBD7ZZd19zhSlH7SYnNFmR9kXHBFZO2A9fW5S1
jdO/TsVR7QQXJOhSE5693pXuFNdQ1xIY5dBLwemqh30isYgq5F/5ADCgtb1kLK6LZ4NbXxiLz0Uj
2tLLvGXA+M6NMe3vg7PBFoJ1rgMuYtZUKadR2lhCNN+OrPMJXGqy5RZek15ziCa1VSNtCPnsso5/
LwSpqJ8udxZ/lsTVS395MkuYpu43hykSVbpheulk3Qh37MlvqHOdLuGW+8u+PN0c5cDMGS3WDLAf
XqxHDCIjd+u1dUVvt7AUdeWWe6ZSgrEuUlv14Sf/TGMcuPZSdxjPCQzwYD9WlIgM2FrpULUgLyB2
AohGHo9joL6l6IkQCU8wgS/+RDFAHth0pMP/c8to0uQ71Hly+yEQqt5W+zh42GwJBgxtmTR7pFBp
HXzxSkVIJh9qpu3NPqx8Le7XC8/K3V15ghhh2AMaMlOgofeZNMoqgJ5BJdgIiEOgw4iS7+l8WGx1
6Wy8WMoT0IzlVx+LXP2w4gIga72gJrznOP6cEdYYNiVgOJhQKLfagXfOwRjsvSZ9XGNaedubjIl2
PuXdtRKdJZYGwlD+IXGAfYhpjyodu1h2EE7UJxLidX7hugDIWX/E5F/Ett3S44pFVOsdUUV+eIHJ
DUiLvRr+vQv67PMiOyMxhRDy+6uDK5w1GH6THNiOjc+1BC/ZMUHlUmtsqyb+XazkRlcbQmn8jSJk
+9Ad5xRsSWbkcHlkTi+ehoT2EzIEqZLcu+KIk0iUmVUX9cnDRjwdgXlExqVZkX5l+UG+OhmPaoig
NWdqwjeMXyv0rL8pLt5PqcX9uXiaSLC7grKunWaxxrfmXbhWfGx4i457Q4jTzIwABkEVKpTucs1h
OPQ01JnPspadf4vmqLTVybYpYEwgvCNrUQeKa3BHRahZBoOOWXPQT0VydmRjYxcrUHL86JCJHmru
v2UaqgE9ODMRlxFWY7QH+Bk4IqOxAzAr4CN7/2r1CoL5x0Lb+SiWZBUjPQK9I/QowfpXi1Jol8Gl
XUIOV0H0MfkFJ6haCnkyaBCuZyHIq47FtrbTLFq3RbrNhh3YrzRNjDdod/V9PJLoicgkZwu5d9+I
rUKmnDZOWRT9rth8B6voCsWAJKtGLbmu64lfJu9vsvM7HQyRkpxGjQsBOzE0daAc8BKi5fhu+i52
ETuYDnTTlcVZ3RRc1OxNbukjGymmrkgYqGitMdOSNLeN7m4WC6LLqTvf2uo/6hkCZzAv0H/1IrzM
uEvFQ+n0hQ6IZFuNix/+aXExxZBGEwuT2VxHdXg1V3iyk1IoFvW1/4ew1MaGitc2inMK70sxZGo1
Ngx9f2Px1+3MUVBmN9oE1PtNe4ef+Rab2HSTaghgGYBMFdVIxBH20sjTUlnhCj5SuPmBODLkxPR1
OI0SUUt/OrvNCBBI+/SCvKacfkLpvk1Dak7yuA9hgDQNnw+IuL/PRR17oE7/ClgL7NaNs47/hs4S
Q+M+SxMyhWOJgPfIKEgXA/mHXA+YLwKv2zEwcUGSdTl2zF2GVxPLwNzLkwtxlaDaHFLLLTzzOjGA
qusOD4jVTYQROmA/D16YLvXkuiE6mNSOeaETU7uF6CXAPkJD0SC2I71ctIMAsDgicdZlzOtzhyT6
FejDt0A7uPT6N31h3gs6GWQuXFVUn8uG7xEUsHRMFwH/4iiSsHJCzazc4NlpwPXXacexXDzCl3D+
sdzF46FIGqowsX9CEsYjZkKt7XE3mMG9+maGG27pVQjLeYwEdomdDFQlINRgMe2ijZgfjm1A486l
WwMqGo1SM9O8JIvZi0jNZQsEKCDILPoQpxa9JCXkL95x9LEM0YZXsN38qVKyI/afOBGYzGLEB8C3
hdM/PTH01POc37x+X1P837y9DhqUmvhUJMOPuZTW2Dr1EOrW5e3Td0qHE5RzfDPQ/M3gsggZNRx5
BxJU7nt3ZKI62G4PVH8Ho6w0FKGv8hfioxgbV48+hVfOcxVSdjpErSFNMdvEYJedlGsV+XhNn2hD
5Tr5x6l17Aqzn/NNMYEbrAEyaNptXZ97le4LiO/D0EL+M3iyqDMUWFCbfpAzMXEYLDHs4DJ4S/ov
XKINRibGopvROljY6y0cOVJ8FHgWCSvUqCV/GfS1/rXoJ+cavP4OYz0WlP47sZfySRXCy1IlQBU3
LZYKK0McJ3wJgePGxpEzy8Jev7k5K9uPIccil77ZAJet4xHZlUITbMXy3A14MQo3zHgj2wnd0zAQ
0Z6Q6Xyj7nC1h+i5aJyvKcMcIKYlNnnGEXOEgIKsIMroMZFtJKFX6m7g2D/tt7OP+8Do5KzkJ//c
0GOpCah28qFG9xwgoN9Q+fiSBK+aimO9SKDzgagzNRi5AWX97w6HY1/LkmVR09K636jI1dQfrnro
Kmg1Q+JQK8LwBjq0a5okKBNnSvPqlTXqYTkwjSVDudfOet1tlQ+cayGzQjlHmyNDlRWNivUXrQkC
dHmq4z0q/5bHKupmNz3rY0Omq68Y3j+gwl6HQ4w7fsIjwscYaMFDdD0L5bQJhAqRrx9eLZAySyL1
l1Abee6UwNSW4UNi6yO2pc0jf3P2y0L0yh9Rssovx8zAta3dYmvsbdP4HCA5flt5KtlSDbRExdpM
NXEE9X4w1CDsd2w4iB2neDmeeZGZfGkJ/O3jE2BtNWv5/jCo6PRIhpm3xtfhvy0OSVsyas/ChO95
6ihBlYAdMC8savLgI69+qGcuThXxdays4ZHofla9b6+5fvBTo3zY+PR8MotVuaYi/R0TmONg630H
6cTUkhuja/Fz1mqmIIuvsH5lLGN4QXg+GD18/g+9BXyU+/GqcVXMUeruzLPQhPmtJLuK3riTL1Ud
vM36UkrgAOOeeiGTMjOXvhL7af4bcFFDZxKz/jJ36VcAcOyqVmklieA9h8sDpODw5l7Lp8HFWvRu
UMoPQF8QWnaRioUjuSBY/eHIoss7T6PmgRKymBFJNP6/J2QkPCBB9tT0loWUZLXceAeuinHAfOAb
W8sjFEDcdbMiD8yDn31w4dbcZVVRyCDL8F1VC4c2yCybkEUOCymPi5IBXH3rBIzuQrxWgX8r14eh
7ZB76g/vhjqxnST4SPYQm3e02MQ6+mtik3SwWqPb7vS2HXf0Je2GIR+SQHLeDh+wypbXlHq52as/
T+qfZ9kwqB/xry72kzzmnphrkYE8oh+s8iXf3l0857UBgPwI+W6JpNHBiAAOOvdwW9o6XLoCFKeX
k5DhIVH5ODTlGm2as5JVVLFI8Gp5tZFnlZLP9arcHNqs5VoXc+sbQy0msb79JVx0b6ptPeXRil43
Hflk6lBBnT7DJW67pUgHOwZaYTF8Zy10xOKtID0xJVMOX66kk72whZMtMtEGRz7LDVVkHC7jVSSG
6CAcmqztA44DJdxrIj8Nt+iUHn4GWt6qRzW2OahEbjLT8UuVtwjgBhFnR8ikaWdldCfoYL8udsfV
Tb2Qs9GSGLA8grHmw63CI67nX4jGJqVyo0ZP+7Tgcbp35k7ur7DNbH/4JBSJotey0DcWnNVwvjqf
QznzSzUbcBw91ehGCaR9buMWOmRBuYjpv8ag4g2gLXR4nFlhugegBIZou1NL5tq+wqLPzATg3eaV
Ye82HbmBU5JwcfuQjohfYWuvJy9wiDpPwOkc3+0pQyLARssHiJJyfYDydADP1pnCIpT3pA6Eg70K
A+38Zk+GhHzinFrd4JIT+xp7Obwjk+vb5Flrx4KKYLtNFHnQ+4UvDWI7/hfjQqjmdxIchmo+xEa2
e00ay2BYHzphqyCYRXJUsK9RCAn953CO9zCMbbIIrH4mq5WyqfcBg60PIxGD9nCCnjBSjG2yMHmO
ukf7bDqtu+Q4Dz9Ru58/REDAEZo+qddvpuph2DPjQv744ZXOly2xjujUcC89PzkLtrZUAwXU+0au
FEptmKXP8e0TNY2T9Nifhbq/kN/fSCptr8jgWs+sHY2NLazAIaKI8Q4gEHsYF97PFGMO6uSCA0QM
KKu3qX+CyOHVb9OVBM1ju8TMagt7ud62CsJ0HWtlTpbgOVKGwTY2XdkRd54t/Ue0j6zZHqYn7VXm
p/DtpD4p8oN2UE25KiDPae6dPPDm7uxcRlSTYi9EG920JUAxKdmVPJ+dlld6Ni57iG+LvtODXEwe
T2249jhsS1s2WdlqN5qR+01D60xfNJq0Kx6gcWl6QC/Om/9h2yM7lyZKCEXP0ZthsAoxdn7Dl+iy
a67r+8NeUSpYJafyi3DYuTKktuL2PdmMG/V9nHWm02/r+kLeqcV/lJzZaCDMzbqTQ+6Hm7S5teg0
jFxY8z7QL32onrRUdWF/vBVOx7T4r4LCObp5VzSiD1fAX2yQf1BVMeDbIsshj9ktcq7wbK8idZg8
7xXTUTe1HiVs1N62t2d1UqoxLLQ8Qt3+YG60Mzqa3gUzQM+knO8WvbbWMuVirFlawwvAIDp+KLEd
F+HPVap04QjTL0RBYUtrqi+LphqLzI8vd2AYRqPtpdLUMvwfs5P1Zdjnb+v00eUdqANdivFOznWt
6hjYxqzlXW7qELNVchNx0x6wY6lRz2oLottifdfKTjJTq1lRjVH5BxXgEZJjEbiQMGtzGivIKfp3
pB4fqn2jQjhJNB422mts4cC5f19c+Bb1Eqd9O4g7ePLK7/E3BU4ANKkWe3U+2ABlAeG44qSybCss
4xivW6bPjN6FAv4vJxpRZVdMIJS1G0jNczDrp+hidMDCJrRH2fTu1nMlsPj3Haa/72vULwXg6ViU
e6lPDsWICTl11VW+2mIL++271ifYSgp2rObGQ4pmxylx3TE3jf0PpwYlAPx6UGhTBy2wDGNvBMC0
qJTqKq3bDL4VFWHqyEHHcfQg+JM77xlps2NwCwcMPGLhZvHgoWz+yGLhtTlXYvmvFE4Ps1uPH4We
ZNCYqTi01s9OR/Xt0UFIZ2Ae5c9PuS6pl906eAJ2b/gpeO/+RSNgmvxqlBx9YgrOdsaJ3imk4Cnm
c33KN72Bzuteu05mcNoO0eh0UwJWZmmqGqD2swvoSM88iAiBt6q9CR1J4KGjJuLXhyf/fcqHZ3lt
pOUbweYmcUXt0VpYX4IFsza0tmOhX1ifX3freFA7MFiD0oR0Z0Ejl25ymcfAuDc+TtYcx2fknoq0
Uj+ekynmnRZmCS2hNUO2UqOVh075JWCTTqetVp/aGj9wHUnjqgTqg4qfAxrQ4UAcnb4OMWcPiVw5
7ALiLMulHPoJZMjLXsrtY6SKnzKhLFDFESOn1aNxkekKPbvK17xTIlhAkpH16//sinunNX81i1GA
UJOKdW225AEWK/wbu7pSD+Dc88SlfGt+wLkwHhACd1PjZ4Z3qa7i7q21UYfIaaLCb4g0HGUXSoaz
QB5KpSJF+3D1+7I1id65SKb1PBPsZPcnr2iwhn27hSGdxSdELwyDWhoGg0EzuiYkdhHJZGpc1DQV
XZGMh/BVsHOAmnkDt1jJZMti4YUybMk/8dl1ourKF4+iORaNKfAW5o9I0FySEpFXel3azo8WeLRZ
yWOJVdE23J3s3UXU/tSIpOtfe4Mi28X6/gUHbvqiGgR58ToxVmPcTSJ4peiildFZXEDXOedc24bo
vRboxXgDWoZ1nTD8+FYMJGC6D4MXQH+DSKaappdLKzQB2ArdPIzf+fkW7fW062CmFM2xVtQd7C2p
kYDweSJ/vrAPREA8qKoe31otyXv1ARlQh6iHu/k+sDMx0Eg0LxNUCL+0o7oXNAm74Dvsfo8SLWMl
ypSloEXJx3Ybe5E6fKZdUYxwfM940Xbt66Ho7q4NtSu8NNcX1FLphB1c6wDeJje2272OPm24tluu
ri8b0Sj8R7NZltR/F5b5W9/LMNdpyYGlcnO+e0xVlMN83VRt8sMcS9c60/V5GK5CQT54W/NmD1AL
1HZqAXND2wPl4qtjQVnIVp6JesBqdxAwEN5Oj9XNntu7Pbv/yRYBW9iUbbj7UxTHGOvUjCn6qV0S
1iPWh5MFf4Jfv003hCfBLb4oH7nRA4dXUFHGIDj9ueH3p4Uq8P/lkk8flSQD8c/xB+x83J7H7sVl
lcrS6GmTMRoh4GD0oSwjhdFiAHjnTgJTmaXVl46q9XXeh+ItGJokdXZglCoUYMguINePNyLMFVbt
2ONsO0Vz01n5Ixz0N6F4Dx1F3q6q5s8iteAppbI8vneDaSUKTIioQJPgJ8avMOM3Dp7/KIy6R5sq
x3j/dD6J5zXT0VHWvHAVQx/M0jFjiSZL/qikYNT8VavP5oQRdyNJLlZ0mT5kCMd5fXhmj8WzBMCm
o+8sy4Z1P6Qp7qOhCHT+N7FwYjAKkc9lnfmQXZswmqRi3somiC9bLlqv4A9fqHc7IdXAgaliLMOl
txB3C60LBFmATQsntP/LC86wmFxyWteiEpkOGclElfUwh5kNTU33AqVBUbZla8bnp9qCkbm/NHaC
HHAEDwPyccJxnqZyQ/sqctP2zNTTIQeYfubdtgSyC4cHc6YC6yI5pBc2s90++pKmOam+TMq0+Gs3
+z0OJ7508Au1j4fdVfLHYsJPuXeFJygis2xJv7+Y1ybbW61I56gsiQhttfH6wavBsEseeY3CP1s/
PxvzIqG2vuyPLxup1rcuR/r0gmKvtI/3QpFGiONObBS7nBvlzRReTv+bRtgCTaeGVQqfrKh4J4Oi
YUxSMvVVGGThjSzuSz+57BPeiFOHi65DTxBZIOmxr6rle9UhscMyQXBNVYnJUuVi9BzBKTHPe1hq
grYJoZTYs1vsb4rphge0P0C8Qn9AA4hLjBu3T8HVuZsuwQFJRtKeHMYB+87tmH4//+qfryvb9lAV
0i9fx6uOa9Jxg38ZK6R0kxW8Bg802DqWLnUXYqUGTazbaPd2CQSpBfAKG/t8h0BwihWckuk9Spqn
YQJzqgTtxLak4njISXzuCIWIac9/Fj10fDn3o8hCEieIho7maKbwoZrpncsv+buI0tgfBYdCAUDI
VOE86e4mHNzGNa8K3ntMaXoNuHZQotc6pgAJpFKGDEVZ+xAUBewEg8dfFFy1OVZYg34bYRZEfhXZ
Q9yu+vwDx2QG4MiZokZQB4iOFzU/oiD8DQ65SOxufAnAKNbKiQuxsArNFuFfxJW+RH7e2nhoInc2
Dvskdqlc9wyUmY0Zl2NVg00v6UFUYWnoHzeMw/+KMQ61s+8ZyjLmCUeQcsia9pSbsdMQlE2ad4ns
k2WgeF4lLJigfm3Qzy7kNQYtkIhcKFb504a0l+3vmAvvwDPzC6xnwy7ma9HvFnFKfj8xM+gc1iDp
2oIv/nni4rh69ZrFaqkbtYdTWS6rHuU0//H5GBSZu4qx0PiImh4RozhAJqsD8IGi+LUaUeYwb5nb
OIAMzcn8xapqduwqgoq7ZtBe7GJD7RvfS0MFhiDDpUBX6+JeikquhJn/m0DyWtM/M1eGR6RiTDAw
+A5sGSPb6jeUKaAdYAVUWgPhm3dFjjFYO5tqiUHHJYmYD8MzeZxAvZyPZ9Z9LVqYeQmSeyb8bDZ3
J2D0wkCD/EBHHifR8Y1PdfbmB1UiJUGIL5gnAy4veLzRMiPV8B9PYYuLroT0P162YaF1b0pM88vG
Jg03TxF76csKQV77X70WU43ka0mTmCYTixJ0norzD72jcuYEygTVeiCL6k/+yRe3VESFdi0s9JmB
Za0q5uBticlMES1HyRhYE5m1tOVEAHG0DVAOMzN5dtM52GKAUh7gQQ1QO7TU3m+1hrx5rH3ljAlz
BkM+TR4T1eH0ijO6nCdnsQ6yFz1XBOdh6YwrtbDesroccaWxuUdwqJKqmQ4i1TQTEv4QBg39Xv1v
BZ3qkQa4rAfvjiOVTywLsT5PhV4tptPwp6izoexoE1Cmt9n8hpY3HbT6PLPktsHN7sIPmHmKwFxn
BXAevLbVMpjgXUdVxQEZqJzgew4uirdcdv9cSyxLzmNLtWCcRZDvnzXre7kEPi1i4rv24AA8+i8T
v71hu7topzk+Q506PQ3+++brxOmLTggRsSzrHuQu1PCuH5DW49BVd45CqBx837LPYlGnglBN+c4j
6nEOjtlKnLw4T+WGHSyXEJfEtBKQj1MGtPJTbCLVvFq04xduk9IyA0cng2TX4/6dqXyAS/rBK4R0
R4khddVt3Ll2qHxia5dLrYDagpNw0ojfDdEL4GVgVy24JExs0OEsC+I/gxhWevS5kjVUpqXZK/z5
fq3YcWexHTt2/9BOHTXAw54t8DH3Cptj9Nv2yRhJzc1nooyNIje8D1TmFx6BdGuLju1VFjJhAi9e
ipa1IpQb9DrLic9gNtBcFEUCUdAOssbJP3SpLenQQ9vd1E6Rm1vK9zpHJv22PMxM62rIIpBS2aS/
VfCGQVDrwG7v07mDB9WNxxqRKlidZ2F7hXg48gMHbOJ3nVTpiCpnH57LkF/jeGhQd+LCfaZ2HL01
aOH+vh1Iu6TAxi2uk5evcvzhNwqElnbK5UWyO9GfYh9yf27W5ECaAIWIGYD1+RPX18s3CjIo3ayD
K0xevdCGy+f1bjGOsrcst5502jhuCeot26fSCCu4kcPPIanrX1ZeNcDQx7aTWXYM6Gr9GRx9azdK
Lz7Hp6o4t5gFTDwgEOfTYi3nv/rBoUVIPxvxUPdLMvMsHWm69kb+DFK23nTgItg2Bpw5NtU5IHLr
+NA3ecDiRklYi/YNjVT8C5rWU9TKKVUZCWfJfFcDWmaaCEQtQoYPBfoCqSSStpM0LRL4ILt+T7YA
7dzyqS8bREBaM8WW5JnhbLznlJg4tJXSVC7X28Gz8apEWRvjtfvp6gD02F710GV1fioOMBnRwgd2
HPw3Ph7S0ueWzOQgDjOP2qMlLuRowq+KbHhlokM4F1/dnlbn6jSw2YQtDx9Ejttlrtcs0mUlxXDP
wE82fn0XGOVA9j2d1SqTatLwmJ3pHJOV1NNzKfq0av1mUwNOlReH2aKH7HFIxRMeIiJLotCBFnhJ
uv7kpMBWOhWZMPYrobhhAYDXDGv4eBc+e3i07owjCmq/WQS4upty+/1/T83Sx/kD2GF9wye2kX69
2RWW1pfGK65bf/e8Ivep8YjpZ8e+vFSN7z5ztZbtkwdacie2HLzl2MY8FKcmFGsE4jDQyUKFVW2n
+jD5nT615aLcVE8fRr1PEkqsiI5zrQG5/dzuf6XCd4BU9bhkaHcgkXz2lkpfPaJiDLoReZyRqYZc
cAaGq4iV5bCXQZdIJZZEgxV8ES8OmbYD0/ty9t71x4sqfuScpEgxEEohWlAsYYP8xahM/7R4yhM/
85OKc6oObGDKhY6tOFtXb+GfFOyzrjIB0jtOCWS0h0saIXxmafo55+fyjeFU2N01u5OuGQc+RfdM
X7hrisCoyYTVOyr61Y0kUAcPCcGMvGMWfc0CQYSRGWqBWZ8BCpHNPRF8oR9QmXdqw60SX6BnjPRs
l3cJaWU5SKS2KBkTFI3eCHiNFHuL8kCC8vNes0G0JjWelL2ZZcNZlPGX3wmLSEr2fu2KdWNbKogP
pUD6IVQ9vtLf+n57sikUts65zDu4qc4/XJgFWWhw8WeiNL+jZ4D/smYV0GHDuU3KHa+WSZBf/RRy
FsdgmUSxoOaIxeJ3s2+0AjHgPJheh7IJ7OGm+CZHQU9Y7Z4WPJq2H6ii27t4ClvdE+L73fnHJbeZ
Xwo9bYyBao2ZzseZ877gtVjmMeONpA+NuNztlfIObzjrjqDwmehmf1I3iow52jpEWTeLvuOK4Emh
NoGWKpbchcrXTgUnOPfswMo+/mZlEASSfUAZmY9AFXa68ogxFtvk3VqEcd2cnXOs6NNDOEU5ip9V
LQ4aznWXzAHgl9OqkM+ZXzuBBlXavEl1BAdP9zpytZP6VlHjR38Y2OltpyLo/xz2vmdyYE/kkCvq
dLAStjxsDqVje1ip89otT7FK7jZKkohiry+puG4y1Q8MEFnuB0++MY4yN96SxLjMUV89dK0ZhtMX
p7CJMzQB2ElL+DmOM9zdbqMximmuKadMkSfWdrTdwpKnCGxEhZbEhwvWnobay535iZhc+kyhWYKg
6S7PQAssFcNkV9vrz4MMNpKt1N32echG7sllk/WsA+/MO2niUTvJ2B/z9nV/fEe/jvP7FEEloE2W
6o/haXAC9yO4wCuDghu7brQGqzIwQ2u6tKrkasRm9eCxLYUkuaQGL/ItmHQzGBpSj/yhUb2VNP75
VkQu/mVpvdqcrk818ose8cfBd2YG1H/cC2jjGL3ESD8tE8kDZG7aRWI4VFsmBzMvlPBmjLmdaYQ5
lIWM7DTlr9tpLXzVvS8F7RmzlpaHsuKxdGSFBhzvmwDoph9ONzykrU3UoBIm4c2NZgwF9uTH/Hrl
cnODfm2y5/FliNNnxye/Zzu6uqyIuvUdQWWMUpoSGBa00g/PkZkQIXmjugoIMwUP+DB7rrfkIbzY
4AOITYgASflkvOicwEdLWHrtnzuh7v0dzJPP7qn/MqIzIfzc7Z1Kb7mzLmi8+cgKKS9XIBi6sdkk
ctvnhxzNBXT95ez3mdxpeNO9xtvpHIvqosgNlSIIeiWBHlwWrIxSgyCccm1P5i93TohX78NwJyk4
pDLaOgIrGmZn+7DQsZwa8GQ9srlqOPJLhR2EGbcxQt1+DUryc0UzmVTVkKzW8fgKfe4XL/KT9WKt
9TVwe0Q1HfMVELWVvvDaGKA2tJxno8GSlHxo7W4q5ad6c33XVqSyBXe0/bTFoFj3ReeYa10hmLLW
vGoCJqUWWUKovsbbFKzhz3atN1Q5qrqMX+2l7Gs9KL4AD30YPSAzpgn5hbRm3ZEyP44rYOIZ22Pu
yDtVd5SJhxg/0Sdet5c/zFy33M9F1hXNDY5aSQo0dw/KOjmAWpXqkWmh0fxJksIuJa3sktr1mDDT
tXw5otv50a3/MEpl0jMEI00kQ0p+GflcWnYPRKBID3nf6B1Zl4KKV94pB+2FieB+0/AZ5p6TLsKp
i5tC9kYjBnWA/RcqIEEU6K/MZM/fVu9YHabuA3PmEVAgQX3pHf1HuPucvFay5PeN54r8Dniv1NBB
qac2JpkWZHrRKtktTo5yPGrZ61nFgG0BLCIjvfHiXQo2VaaRNOtEnJ9rh2wbZyXyxuVFvA5F20ma
iCaxYiJv9UjuQNBFKSZIqxnlRVgzQ1NVicSLeaAmi/o177ei2MPBBZ9na1PK2yjy7HgObVPBursN
0sUsVrkV82TCPiP2olsxeUwrTd5EJ5DcP/bQraV3LnClKSeKrC9uknil28xTsUlet5AUBxNcPndi
56IqK5OmjQ35IIGEek53KBKh11ruT9IY+PvqRLZ3lEAmaTLdu3Vc8eXAlvSd3jqKOOg/BYW+3e/W
hGrqXz2+r5Ius8G+x23U766bqFtxSNRlGqf8crZIDu0Tr5mzinRd7yBBbEyAZp5VJfpFxuVavTHk
xUOYahgksAyJQ5AorvIpWeJCKvxXELh1450HqXKEBUjO0TjcIlsSKmWdusIjQFWVCHVM1tKBBAYD
N89ovf0+Q3ugsHYUTSTOPnvG9zSrU02yGT1GtdBGe4Wp7tBF06xNlGnD8U/3wmshy9jUaTbhkm7+
UgFuiU3a4Z+xCtGUraZtCLcNr6Sa83JmIFltyvdtr4/tz89ck9peckVC0G1lOtIZ8IsuL0sBWQne
wm4hproVYX+pRPHf90EP24h17zy0NzXZrlmEcYRcxwhvlPZizh3bAfOO0inXd5cS9wCA/+hoiIJO
RSVMIQcGKqASX4mYXUXygSsuE99kZiblRFlsk4lKs3AiEhV2Xr93zEnyx4oVXjQDuV/3Rvkrib2s
TYgmAgegnlnklDq1KhxJDWSg9ExzvXEhgOvuzLW4HC6WJYY3zWj5aPfVYfYtrYB1kHHjsIV1zHgP
cbSeXVAAOMl8WJIE0kbZa1VBuFMO6FFERrmK3UZMSmGtkYV8xTQ18RPQhoNQvAaDfVBOZvNmr+vf
24c64C1pPem8Uj/NE56eGMNOSeivGV6XTN8kDvlrWJ1FDh2UFSn5gVS3/Nsi4GnLC9t0Vc1BfcMk
n9XUhHtZ6/gvWzBVQKZWs4TTpS6Ow1YopGL9+r5zlg/t63Q2LRGYMicKXQk2VMJaiJ34sSj0ilTZ
632i8VYSifFz2bkoNAbquHTBntxTnng1ZTtbsjB6IBUp8dPcOUaKdxIayJxlMf6H9oe7MJj8We5d
LiRooMRwmod69OcyWrLtLcODioU9qNN19083UlSnSprDwhgtzNemgYeoLjkPeGxiIHizWflr/3rn
7U8AIYraCDbwGHlSjM9kOHeoyJ96NpgYarQeiuhNb9f7j36AwA8ydsECcvNbI36psyUboNbWHVK8
7Cb39v/fZi8appR+yCHiL+h6zvO/tfzfOPaHffqMAADK7YmcuHwrWT1ewdr6NF537dKdondAXj5B
6qBaxmWcquRIUU4zdsErwS2VwMqCt7NpqHSKDW+z4ZCW4kRQigxZod5DoXDRVcCfX6y7EyatyeBs
CEwiQjRA6jm++oz1BrTNeVLMdBVvKuLlL7xnLcHV4ByKEcjuKMHpGk8TiOChZUXbeRO+q1IDa3mg
wHkaboEP4Tx6BWPES86pkdxjz4oeezUey1L6Tf4hvVv+ZjI/XSOmgxRqxqT0nfY/T81eUxyMjTSv
YxstxGd24sWq01pkMMY8eQftFMPwE/TRoHaYUd7D0BRdffkt/AKU0cKqtQraXSNaymRUIyZkpCH2
BNGysj70nsicIhSdvI/9fJtHmrrcmCeJdZYuXU1rsnClJYjVM3SusfMYxa3DzEhCI+xUWPID0gAL
HdZcXvAxZnsUVt4ib/ldmWIHiGacVAN0mDETVU3G+hSAV4EUMm3E+OE6bnk+/5Lnhe4FtfzJCdk3
R/mT6q4eKHwIgee2sdXQPt3L52pSoCZb2cFFRcPIrDauogeNkLPhIPOOkt4Xo+WZBTYuw58epuUv
Zrppr9fkPwQps9zSwJX7PvAauErNjFZALug3tuUgagyPf2y3mfR31NdWyxfK2mhKriyXXKyefUMw
VRPo8hvH72LwE1sCET1x15khyhPKPNq1jJe0wWYJS8OZGxK8vIEahipM8wOS2slvw84jsZo5ISDl
3VHn25c5mDboaahv8qjL5zo+9R5JDUQ0YjbYn4d1ooMt8X9B/C/dthvF+S03zz+fBUuiyluy0s7W
xlrdHpYZO16olPnmod85ArmMzPufbjQc2XswFUdEBPlnNnm7Mapnkv2zNkPeC1MlsomX/4asqf+F
q83srtXMdNyo8W95ypiBKQWGvl/VnIEcK5nrEc3XnmK6PpVtEUug+xxjbyzQlRlaTnEFimrYrHAR
1KUzrE7FEsDQIvmlvu/gpoeqvZdnLLDA2CAblXFqw7IQscJjLHOiD33k8/TKcFUehJMungvr2ji4
gTi0IMjjtr6IRR5kVWevBNZGNtFJn/TQiXdTvCyizcpRy3lo2jzHxisQIp1HtRREywwHodMlbAVE
OS0SVJfDfdrlzAjvi7s55nhLhM6P4R2GJHsFbMvp9miA5DwMVeMfhnYwInUWNpoPbynIe7X0aFcW
BsyndU94+sK48qrowouOxk+Pnu8mHgDZAqdm85M9NnBl8slo16vr//eS/zUvpk+tAHm8CBCkWPos
fsmUCDsI2G1tadWCilaic13LMiBUb7eOinVnmWagrmMh/GQHXHzytz2WOBjx1Ragr0//KqVjQPP9
Gez4dMSLhzXgAZI4VjTgrFapa6JpiB4yj6n/2O7mtVbgbn1NsShsSvo2K3EIHSVh46rfR11LP1lR
tdJ/3DaWu5kqQgdGKFFrDt7wNkYwNIC0n79E2xy5BymPULmYeqkvOjpvMntxNafEGgW1caBC0Pum
SPe9ASPoTT2K3KlnxphTp0KzPLdSA2GWrxGZf6K25io/67NRgtyzJ1LI9VuLlNkdfHCe4uoBw/6h
5oDnxDrnqhAWMRFKHJTU34KHmHRwDAXUO6t8dzHJl029qyO8zavbmuCS74q+3zkVxt+wyPAJc7MF
o747M8wSjAWmh0Efy8J++j0zdf1/1YTNFg9QKd+LAxT4dclDcHlyXmFA0of3vzGDRSSENIn5RNMl
Wcv8DArPzS32xc6GQ2proS8RRTXIbLV5dSVBApcyArn2Ga7YkUBE4a7fQIZkhAG3DLmJqGT/0LAz
01gS7RB7cLcVAoSlo1dA1JHh1zLr7wv8XNTk2w5gXWC5ihDZyMQqIk3/znZqPgSfzD3MPXSC/eri
75Lucupc2KR+gSFilguYSp16lHZda9KbMuHzXyJHJgWIq9juCWYG4Yfn+0WE10cgY9z4lFG/PxE6
+W/e9xevBAueArbn9c7T4oQuddOUvizKvRM4MXPzWbNjY0pYTALwDyd+jOsyLbcTJVIbzO3AAFpj
FTJZmJrCX2ywLEO5u1Q8DbzTHfkhVWNdvoGSG8jmlax6ZjFtqzyxWQ1mVlA9LkQRKEjGpAIIuxvS
dfvSP+RfnmPapL06LzEfG9eUg4OvVFHHCdkECJKPCUL84qlK/1iU2VSiEV1r7eSzLQH/UsbA7z6+
9/My3Z8hEg5V8VwS45pCyQ/8XPbqKVBROU234Z29GxYZnmDp6Z1QA1LF6k6gOB8pABWCgmpEJavn
27HSdGt4djY/ZthwVRXgnbg9rPJTtLSVuD2qAlAzCTNoNwUznnMmINCnIVIwWq2/gjXDTH1dr3rs
iTsXD9s3LfaN0riPIPm0aBocqgTFmlPAlI8K0tspUrsJUPtHAdUWe5IgSxV5myGJrWQhWP+92Ne9
zfy/CTVyLZFkK/hjus5ZxplxpEJr/IdJZYgNH39vn2VAarwGTRiA9pJjiNZm19qviS3BJ2vwO1/X
t2ziKR9cUF07yMqZACgyMLaFlv48AaZ1H21/ZnIyqjDEsdboOAiT2AmmBr1gJ9NHsp6EQJHo5mjI
THk15hUXP96AP7gUe4Pe12aR4PsZEuucfjrqJtj6sc90OMH29t3MjM5IJlwhgpw1nk99qKLxBmY3
vKNrtm4CAX/BVw/G/nqLy6w0YOgQXyDRWhThrIcy+ubW07lO+5DZeDSxDpc4IbT4NcHt02Lx55OH
ISSDbwtSkxCqzZfuboSbVL8J8SRRyDfSrqIhd6gpc8rMZN30Ni6WP4gS3QIsNqIVZ3i2V2YqILbz
edeSzlHC9FuXDprIBYrgHlsDs0jFUbVq/mZ2jnQ5ScM273wchQp7mcuR4BqZNHSNr8DScC//mmZR
DEDBf8q8ktibqHJkcxLCTEjtj1fU8VVUppJ6ad5aRHdOveMYT7D7wGEHnHyLWkQIoEzoN/nNGSmQ
P0uOtnvLSIkCkezVbQGMBENIezbB3Jj3D6ml9igz3ZkSdk79mgLH6TKO583dGcAae6NUhEpBNGHj
Lhs3s4PJzMPb8jDzFaUANF4sG1yZpG2Ej2NjUlNx7lfQaXIczYLtfe/0GXIiUCVMuc46shD3LPD/
TU76A+SQ/RNMmZPBpRfy9H27xHEZrtyHoFqGr6gaflbFJcaAdOhKmZcTc2VGfhnGoAec4MjEOcEN
gYCsMP1ZW57BTpSoPHwteqxZRv/iF+xote8AGMG1igvorEO0f2lLNCdlixBK64xtKR2SdU9uv3bh
Tyf8ubktg3kFG9yqiibfSPe+Ww/qzbHRvYL/VdsiygeEOqcKploqynII+s09k0tKRGYTsN8bLbdz
cEueSEuqWGXh7dG6KWbOm/EjYg2ixHqkF41/+TFYw1OidOBBml8doWNJAQnOqW3SYHGaFmlvFemX
hhpYGyY2lkUW11UddJIerQyFPM1ybZaTb9u/rFbpH9Dg0BjU837zM4E3WMzwPfNjuzHCQwAKASFA
5w2qKqhc5rHOXWIZYVJ9jADDwqTuCZ4s2qdM29DT81062Oxj3v9TGywnrUjk+iUDb9ujE1H66rIo
IPfkhNvt02qvUBPZzFgMBITaNXZgPe1TWBHWhrarajYvR2bzPgKS2YPVRcaTzxg/zFOHho14Dj30
K8VmIq/UTpwa8DUg5Py3nV2Xrx4ovHSr/YXgN9KOd10N3dt8c0EaiA8tHHLksBh0KMkybEyLe9SF
Si0SD8PLcOiIndSwSdqR/bEGQORES/DxxiXDLx3xeVtSdNzqYdq3U8tBBqNwqGSSOE0buSwg2FuI
QyycM+jdUZxSI4tLjwyWFJjAcPDcmmjyB1HgkV12lg5/0JvN7YSZ8fJGk7xlHht9wxBgi2VQeh4s
v1WgQKz0Xaa00b6ZL84ozCmOdbkNioe0ghLj92ChQp3J+fpXoSs9lxvR8sj4kdI2mgYC8euGlo+Q
lvRQ2rhI3fmZj7tmOSeZVOs5RlkBSyxv0kLqQQtnlllczFDdPXEfKOvWd2sU4zyean9B8mQ6W40c
qwSr0krmhqYCR0hBHTNyRFzmDKSgJKcJdpyaglTpXtDFUtQPbtSN1xvAGGJZ15Jn/Iz+COf+AALX
+fv8ZEeIvYcJj9crr4M0VUPMRMcFmMHBu7CSFBCGYa4O25BZtyibFp6B52AtQ7s2D6PZIZEMfOqA
eFe1Ig1ZcRMSw1tO99kwd818u4074/NjKv9TVXAt/F0GqLMQQxM3uL6mLYOuUgGLAMpdhH5oBSsB
CMbF6ZFdm9FYamdjWoJiaVe6/DiEn5uaOYmyYb9dHpup4vf683Toq1X0CXuhSkdSMWFnvXymSXQm
dou1Kr7nSPvhPXfnXWNj6KFOsFD0GSSfi/nzJ4jkRZxnGlzp3U07wBsZhFLecTwYy4h6XgaDzOQC
IzWxVLqjfgUGFu6PAa00ga5WxG1s/twiCqaTTYt3zJ+XRUpoJqq95/DZO6E9qn9KWeB4jbaYrT4W
Y+FJE+Z1lF+7Lhi0cj6eze/PSI6re1lr56Ge/NeGg3rRz4jHaweXnd4Zfa4vQ9LE+eHhko2HHAfa
dfcF+mvwtnbGQUlvuPSGi9KHaaqEnW/xcF+fg+uEZWlKvqu+9tXuA0loBpHL78uWncEFJ2lVwcfW
4yLT48hpaz0VitqwlkUbPMaHqpRkOJhBBUVh7JhbBLGxWHsOwssRPcEVfayywETD1CnUr2T7M7bx
skBiFGLsmIG+T7aYGiyAB0WTaUUxC4Wgk+XYHdxMAbxNOcfBpiZ2CPcvrsH5EERv7sMvXONlK6RK
T4+0gkfB0Q4XFapVZXTM/ViFj6EhrzgKvS0SWGV5E9SoYjBTudEZvDW/L7OIm4/Pr9R9ef+LzEzu
nCqwifSApvliFf/sJHWMa0U4bjOygPQvRrieFbHQ8nNu6YGVDOn0GBQ4RvhLusqnp5DfuySW1oOZ
eEF/Nuxfn3xIb8hjBo+z+KY2Jbilt3BkMF0cK3afYK+bqqlhPiCVlm9KNV2qx9YtRbkYIAv/NN89
eEPApUbOlFL4M5GYO7RIi5PD5ejRj+17tML/q0zYgJJVoiH5lNO2FAapXMXvJnW2NyV6v2S/zVvJ
i+BJxvfAyYl1jZmSUNiMTxigyIVMvKsoXukwBJyvMJSo3PyMgfqFgpifctdpbGbHme8H8FJCbVut
zUv5Qb4HYHydZCpGGc6b3vPCJyziL/zbwBKgckbl7KXH8TKpAuMthD40780mGuM0m2W0KJ50unqu
vURr/B0heKoDBZmOeQqCOgoO/kx1LAd7TpyxxJd4O1Ne929DshrgGLBr+eyzcvJt4zjk89vd9SNm
oP43HX7PAwNMGoYz8nDQJQFl6O+CDVOOBHlLs9b3EzBZ4cpe2DcaNMmMXHkpFIup1fWXsLcd3XKT
6MhZ8/yHo6ojjZFSe1GjfznhiSdLAthIUmEafUlHt00ybCPiFTzmkXlWYqzAx0bCUpa2LCiffhhr
a3BEh9RLUkHEkACyHS4VsxdIGUsh8zlg8FJ/tZVXghpiezumJOEszg57O8TjUxyZ5m0kjUr7+mIa
cPpDtxj1OcOBl1JDye3awafj+zreDaQcIq8Z26VbQVlMh0oWtJzrTzCyIdjt7XH5qUO2TfXopCWf
CDyd6YKL2PEfcIfASKR40NNgfcuoVlINM3nArz6WY0bCevdzXCXHZmJwPL3EZNkBZep+gY+xH1Kj
vUSuKGtbPQVXCCA9glgPUH8OQYCEUCQHK5hcokS0VgelC01vZBY+JifGNO5wm04cRFCnwzF47bNi
c/nU2OSweWTgxUImeu+2zrYxAlbRO6uYyjdQa2KMB6WZT5E3IG3CVB8Zsknj9BBgLmkSKpFDqp7q
nCOCOhihMC28ZTsHyd+4ovLJfYALbOAjecmmDg/CSSR2iva3EFDHsDiE5qsXvZ1CXzi8mL5CpXag
Pm0TT41U5CNRyMl4+EHLwspuwdWA53tgK0pQK7J8DYwbl/5wkdnzWCY+rREAYV6xT6uu7I1PYuMC
sbGfn//4x37jUQVaIHe6x2Zj8OuJZMdeBhPt97v4/dNP4DCLCNc9STh78PpccicM5Ndlnqr4B68V
kynGHMIHc5IWsTHq2DcJkW/XQA7/f0K5i12MnmPExr2HjNAXP4+9ZsWTs1+pUWevC6Aky9jBbIdU
gXMIElmuH2SS5RnJ3JKc3xy15wIw4g4ReTvcwBmvwBnmjFu+6GRVeAbzpFsrd+QsH5c7EHgc12CN
zV6JrWMHZ+AGQWU6xGIdyJ0QmfZdi5P1KaKpvCBZII2SVfPVd0ZAn6kfKxcnZM6mC5ehT7RAHbTz
1reY3hqSKraJiipeeT0B7y/4KCYSMYq4xHcwX9i1JUunS44eoRBlzmywAnID4iJ1iX/SfXcbddtB
Z2s4907+FpAkQusHf1u7y67iqd5t7AaeYlTuoHbhCwP1wxr9w2Qz5E6AFBRhecDNBPfSaQPzEhKJ
NQNnKSdplhl6HgjslNMCSxMdctvUW1Lr1go8fQYomtId3AKlTXwLYozt91CVnOlvFxHVyFXmBz0E
4CH4c/KTZUYXJJ/0CrlLlR4q+/izECghoE54YXTNWAW30CsR9hvjt3Z5USUmYWIQCZrSGu+HLqGP
eqCviwBleLccE0XBVAY1gMNKkl/PgTsEDsFGs4zrcGcZa+dGHGNXy7mRYzNMT3rq2jaGxDxDimB8
MnoajMhg1jYCV9Gg7/OrzNnsMgMM21sYopescwikPnwBEgcbWLO1q1s3Ot67B+bFvIvDajCeR68+
x5hIcP6Rusl3IZJuHQEflAvs8SBD5UZK8+fdHLo5RU3uq++1Ht6jVHvq5tz82KJUEoVnzbVsRfe7
dGBZsa0+3QSug6uJvaeSE5LX50AnNkbz6x9JBE568Ni900eApd7e2RcwQCsVPORZUnvCSRiyVowX
W11xDOoIldCfbhLzaT0a4mQFz7dWF7rNgmOYylz3WRY4tB2Jz6WFurfZGEK9XbnZ3VBDvOXzczoS
oivmapeIsChLlBqbkVtMEAX+NDCAUreOaYOclBOE7cMssF7EtH3Sa67yWi86BXEsheIIIOmz7/oE
o3cQ0hfTkeBJK5Nd4phQmU260dxzdSiNhulrywh7EAVwSVC8PmjVKCn9X+oxorC+KZwHTzP9YiQe
y3NCd6+z96z3rZpeHe6TE3UnPmLMw8UeUDs44AutRcsSfOEQaX0GpCSelbgoV6eTQydiB/5G/WZM
aYs7/5BVh+weYT+iTg03kBiDS1lVWMT7v80Ys9/K6hK9QltqC7GUZRGQ4el+BIXhem3BWzRrLx0G
fFKj3Lp7rqSgWqeOolCGzr4yRAFlBE8thSnqQFLyvlMW4GxqBuMDnhTOeq3XOHkWYwL+si/mJGYl
cFLfpsMRHOZ7/4b8jUSf68GDDZfbX/k+1osRcg+vJuWTHz/CEBjtv5SVXWvk00PAqRZDkJcm+Dif
xzse+OqWRyTwpFcGV2gJ7vFhCxgKlTeVVRM3bZy+QVsyxfNMvyeh1ecZGI2FjoubCKLnvO6/pZ+8
K97OKeTrwV3pxAnviDmZfpFrYe7IGhe4oF8WQKeXHMlUdtxkL5gx18sDIWfnA6RCBqLP35i9366p
/C3ODXNt8UrFk4lbtqG0vUlt70016hBk96MHiiG5Vjq1zov28T916qPssiUkUqPS08oXgGR7y7hX
ODZOq8ARUD5dfTujG8UniYN7gOIXQvrWPYWb6VXKybtgjxWM/86WTOSMl0Iwx0Tv/1tIUkqb13eN
mNE61JtfKB5q0qAQd2xZVe7MfMUEm/RuH1l8tMsK2LN+sQeUIbK2iWhW14Th62fqFXR0ixsTfVW3
3uf9u9P7PKz3UL061ZqgiVcOtT06I4Z31QVUxqZf+uPD+OfzXrgEofEMUOD3XtYdn+9RVuMbo7Ij
E29qEj298/EH0kWQts73c7f2trMVCnBFkKZ5bkYeCwJctBxP0i5DX8bvoba8DbeM1y9D7yautQWz
yLMWMjQpzfOP7QhxVe/zwzIxyH7sU4m3x/Ien6C5hKBf+H4T+Hszh442fK6+sJhlEG2dJOlDqXAO
CdIMIRw5bwy1KBUVHumhR8y/nEAumwJbRlvisOTRorcEU6MJAKCe4Cu09e6GYtV2gWxmjguJVnPA
i7cbM4q6rmIb8iIxwlci/3+sWR4EMyJu6tUW+BwYQkBQScZx8AzRJkO6X4sHoxk5ZfZObDZiooGZ
320rTLJMlwEBTnkBgT8JgAx52OLL0SATMcSXaSZWUCvPhRVpY7xKSxudm2grUTH/pXhr4LoZB+gE
jNJS1+4wKtds7VmDOmPSexMZGOVjg83EhiCf1U/dV6lPrJ9GKUJJmioeyHG70/2/usNax85rbbUu
ulP9TUl3eYjoLw+HNqWF0G3tBHIBANbqqbX5q/kGGdDeALtLzbfWYQ2tFFKeP2v1BGjNeEZtyiNL
bc8K+m9vAcIExImpf5DyhclPuqp9JMClo7Ui0EL0Ny6kRuWtyTDwcgYVTmVUMefdkTS9oqATuQex
Z1ps0/8PCb8lI5FPDIiM6FhM5ldRUyMvwiYwQlJOQNKUQwz45fHTjY/P8yfaG38hS8wIkQy3RiYJ
7gEnJ7YOhLHiYvmz3RJbt5g4mO5tNtrgTEzv/ToMon6abDOh2Alqt6ClwGrpmVCaWfYl8q75RuoO
q1xYU0RmwgcMLQ0PMFMkPOAQ8dHOh6A86HmkoCphLsjUS/81slszbzvyQVsJgVLERpNZWXrCs0CH
+JkLahrHlhFRzZQ86pJDIYzcvK2mI0jdT1RiYdGKPR5V54G1Wi9NBpgCbRkiLLc+JLcTQg5bqLlv
Z4gRdUvvx83oRm7w+99BrQJnouFphXmBEtBAJKBX92M3hCQZhYofETcDwsus6HvrdEudMFkDOBj+
kwGhdzbO9hw5wZwEQ8X1toE2P9ppV8TLVZU4Bn5LJtqy+hcaie3aq4sUGqzBAT8VldFACE1SxDft
r6aVdDI32v9zrRO4Dcqi6JEJtyLWDCqN72Qb9KBSnE6Sie3NAADPENmzTOXl6puKiTa/87JWWCKc
4voYzWhLR2xlJszrLovj7mDC/Zh5M77GBsN+aW5T5uDunf4cqQ9TVG91V496mKv+liHO/PZypJMX
h5VfY5SwdYDGZcchOahYgJfLSfrl3ObstPiSEIQ3jPcaaftgkwWMZthEVAiZYaaXy0Ar5gxGu31s
Tct/QvF65eT05fhBHhQQmdlS5DY9kl31FUj1T6ZyjiW75ISLFrxLk99mWuR8TNWzw9cAvLSCdpRx
6S5hyt52LjSNWRpR5jVpXBQnvz1UUp6BegjfLP0SpJBoaXeVQP3aAuZjqvq0aXuh8VEUWQzpbWgB
EROqV6fNgSsYJ/ugNOx24gYlhrFu1qE0qg4sZy2C72o74CdO24Hqo37MeXzrdi+npAn6hjJSa2ep
NpdIl9cbh0JpB/jBUqlEwjfAbWx0PHoAf+mKAQnaMdU7n9LdyYtU6ATTz92Ap2fe/O5FFKJ6qFYg
qVvyH202zivX+mp+QtqhiUWodOumgX3hlyGSOPPvuSYh2E8u/0+akR4tcfuKA1+b3X7DsdphwuXl
wlspPDGXBoqtm+iDgb7rafkjhGcVzdlHPmwAs5VetXBakAJLKD4I8n4Ne25VJ3VXHz9i3EHT1uYK
1xxssxLAmDxjdEcRcihLrZ2rBo2/I5SO7WWcJKfT+tqOjzLJUd3CFn7Mg0r1j08i4VKHwqX4XKEb
sZFhPguj5SkwtleClqOKQ08Fz2joz4MiQ49M0IGSZuLUS3E36aD5mj+/02iMuLMAXfxFhhuOjBG1
2+DL1WoSAROj5+eIaLfYiqH/qt98HFWwXzE2q5R9d7uhT1amBepSmOvyLHVylPRTK0SRUmQzdRM9
vcJp/7+GzaxOKBUmas5qdsvWAHdKKLQQarAkH6tobrk9VgQK3VaRsU+7RctQoJ6YpyYWSvMZ0mhu
8+alAfKtTxXwPzMMTsIEMfAT16z0UQ1dF+TztgoSaTPJsOgzdl417dQzvGPVh0XK5voCTEAfLwSm
RE2MZg52yFWJrP3t7dWt721QNj8SZ6SOsdoF/US+ZuGEQVjbLbQfJd0gP5cex7Ik84eSA5pE9WpI
oBS5pK2yrkaY9+ckfhLk+ZXtyZiynKImH4bvFizCIyNzK1zjb6ecYAJk/Uh1Z42X77XVW94oA+RC
wbe92PgnzuydGh8l4nzIQE6zLe+4ACovdZgi9XZWTZbyLgfyJ3odxjTigEI5PavZ/D5CUPTx8nh2
3nNsXcolmSfRRUcAIlenkkpihQxQ25JXlZ7ZBNIuJ5Acy5YT7zkMLuZv+DfsHVh7IZA381Ev5iR5
XbEpFkujIT4G0EOqqwlBLjovoIlLPD9JdsssWFEEDTe4S6J7h1baTGAWvsc+shBFhXg/aWzEo74N
/ZGE8B11qJ2iUZBA5Z5cb9Kq40Sp/BUNq/6lT+uoBXFoYBQOkCPsLeWdZArSLJ/jo4rSf7/gacuu
g//GtvCrCwiMXwOscfN6pgQtmQy9TBreeCsumvJCUjHAzvUjxfBJxguEO0Qm1tVh/QaWT+oZduhT
QKiEET3DtBHJYRw17Sx98+dI6sj6ZhEGCyyw8ywu2oEVrm0lTDVIUpKYd8tWF2q/gsWCnsEEUSKw
sfuytURK1sfNBpkB0nls7hOWM+hQUXTcBogceIkNpbfQ28BglR00qJxZ+DilVP5Rw3e28woH0GIA
sEaxP6FltR89snx8CUkrg53GRosjMfIai8PFTiBVACgFzTp+FsBtk1/maMSikGM5gMVaXOpDD/Ig
2oJYfvWj3lEuOyD5mnjDs6El6BqWU0x3NK2NExLngxFMfWXX9v9lNs6GCqDZ53zV4m2nEOkVHra5
DIsv+VBcsWw2pmecfJ2Oga5bmxC8hnKOsizpANv3/zeoiWSa/PPhS25iVUK+kyQAb6FLyI6oVuyd
LnkEEPhm/YWo/S3gtYhEJscXObfqh8hvjIeMDNhE0Cj2Y3nWl/8cSF2663hRj558tTULlNuuWilO
uIMRIZVafc7kWi0Y95+zUGyVUZqoouM2AQsX95RrZUb0507eCWRDFrA+kdIw2BmBQIpqh01mDrt1
4j9me975s0PQU0+JEHVgnQQipSCtmoyO6j/Z4fCbdxdwrz02IT11y6IUxSC2vr7sLKHUyXkcquhk
0fmgNxbsOgfeCag47PNM+MzoR3RqnXbABsEkjaKeJbcsR1genMCScHW54pAAh0Y/SsGnz7SPBV/w
zfQSofevvxgCK/TsvN+4cp4vNVAVUMJLasyj91qjX5Fm9ASC9Z0llFsPMEXKs6W5+r3DEf5EKK/N
Zm0xTCIA7k9KR8AsuKGSzb8XHocKhC0vhcztQCsONkZgTDE80lcLyMliYnsaAJ9r/nCS5+SXcNOG
E1gsJEVbENKxFJjtsCn+CKzOhgYuFMK5k+j6Gy2bGUfGs9Fj9YCYJSeEDUdkbGr7mVWV53aSjJm0
ktTdN2YU8x85tTkzb4JZF0Swhs+X0jlZ9JPdzlSR9enLsPC8ZsJ5gHz8vY2oOLRrhu/H5NNKJNDS
ZRc5jhKp06jP5Y2bM8iF6SV/sij7owvg1/Rfo/074fZbDt0TS4mkQtmPBebK5t4+aon2jT+kDqJI
yV86LFMGzA920cUIL/55X6PUyT51i6IKkpgtGl+Pk1o3PYQeXyH2Nia2r2bZYo/+6Lyj0ChRN/If
B5F+LAwKf7djvrhVMoS4uNjjMC8jXp8Xfm//aTx4U9tWfrKrhDEH0aV+uJVwI5dyJhR/XBpzQqmC
999qGAgbWVmaGK3N1BVCPyyHY80cnCXSqO5REmr8nq826+4fGlpXCDqREfa6K0ETSCMZwoYYOl7h
aoezWuCdcF1wqHoKEr5f/3CUlhZJtBlAzRPnS2foExGbrgYoBwWrIixyVSvrbS0ag/Y1eNOnu3ph
BZmWLYKTJWIN0za88e28hLOB64q0bNAroHTZR4H7uVUrK11gc865GDVIFUVSMXnkhf19QOYslsBJ
h5kpFbxS6YPjVYzE1AadU56gkKw3sImIx7wgdqy7R+ezD4VJzTTHT56HOaubveuEWPd9w8bm4rXe
Fc+CtDNgAkLc3EYcY8nDdZom2poMDvT13N6w7Yd+SGO9+4kZzDAftDgdv3Dkcp3XhVzY/h105hhX
VzJScnB5doL0zU/CyausbPuZOgzywp23JMik0zIpYMl2kT/jQP6Ih/VgN6FIF+3uYP5tUPbvVBGB
k29zg41rTUrjVtjOszt+qEZ1RuLUA9I0pD40z3xKMJed1y7iyF9yVl9HYhs0cesoR/JtEyjwB/q8
+1JH+lww6uQxI643E6FnwEN7RsLVGhXXPNk8+sIEIlT8uqKfZxDgSechf0ZTzTf7Wu1qcudW8xT7
mClniJ+7MvVl8MzxQWoj1sb4g0I95HNSy7akCbwni9Xr0MLTV3oEg4o/Qd6fv1E+aYy6S41EGxZd
bcH2GCbFKfgAHv7bp/23cnBsuZrNwZhiDNY5jv4OSLQp0vfpslWEWGW+/Vjns2dYhZT+1Frd1cQF
p6c+G1Otyuxz2J+q4KYKPCrtgqX+Q4PqAhkGxePJOXvmQzHacygXVC1k86twGZ/5WqwZwcLMtozx
kE8BEZs5EwY/vZnQg8ER22AP0SBxkNKUkKHUNcZAKx5g0MmStX3U74lKvC3SRitq2uXbZiTbxrMh
ODMLct6JvKrzTeT71loaQDKEFLLHVzLl+EdyHy6JsUiXJyP3W55FdosnJivI5M4f2TgI6/c3uwDt
LbpaoR5fiFkgaZAZjgrJO7SLq9g7OlAn3ub1FXXofoNGTHC6Y/k4TDCB8mkmJBh2+v7ImSAQRu4+
IlZQkQTtPfiIk0jVbJ+P5C7y/TV0Eooymo5e8JIG8UYhYKVdRR8ajGF3X2C1bFYeLqb6FNt1d3u4
beUcY7hckPnSS23sAJRpYzSpUvsRYaUmkcqXB7uFr29tqNmlqGdZwM/9cJBMKjU00rl7qmleB8sG
8O0DeFz/lsGWns9MHoGbJsydbwqvuCajeO2uiT6pumjZ0qgFqGQV4nogxgY0WrDnVvGvO+FrE/eB
p2UimxkE2bP2md5xo7QL9Fh4Q9fIJYg/Ye1hmgLCtJSLCxyC1Bk+V87TdxyBEg+ZuJqAE9pEL5Wu
lgHouccnKjDeU2FvouInR5HD06wg/gW9jXnz6E4RFQKoyuQ5yaJnv+37QuFuZjYg/obok29qEsDy
CKVYwYpoq9ZDLWw1XF1cAn9tfA1Gj8YNBk5kdA9R+Hav7h3GDL1CHaRoH+3PUmFVUSikQjIvllOc
ZVL7WF8KiLvMj1fibJQOKCoSclaADnRQFrPL2xcAUKXWiqHn3amFSolu0qolO1GGii0/55cCXVwh
TvpqQ+WdJEA9kRUwjtMYuqszB5glO8Aei1o7vwGtgttz6yJp0nTl9/6bzna2wza+iR3aMx7qX3VN
ypjos24EGvxgZT9rakeoOKf3fxUtTvhklD9h2OVXpP/GzrQ2DlZiNYJcPKYnju2SmE1viPj4jfIa
+ZOdD1pWlel2kSDOQJPzrG/41/CiVGwoS4A7ffE1rWpuaZm+Fo3iYyoD8FXIxrnWbhd0gIxFwqpA
i6U3pE4dDI7rWO/Jox4CWmeEe7X4grAVMiPKDvGyU1h1NgJeLfLfbYBhlvAlZWJv6ol1FEIKAZCJ
CO+zkEVyosYoLaBjFjsGHyJltzPOY54VPeoYvAR6sLxuFxmqBVYHgH/x8f5iXJdBSAc+xHmxpAJb
v8STO1JZhEOJfiEX2/d45NxPZOlLPG97AUMg709N3WPta5j83sR9miOG7LUvmCVFf0rW1Ozv/T4T
Dy4Ygh0g6UgGcEbEnd9LxL2Jmsw4jQkR3Zqi+G0EIrJSQIfliWRA5ylBJ+aLdVQfCYMCZ4A51xi+
bLBFsMdqSC+nK1nK3l4GShMbqnSQ6Z1p5kEYtnBZ0ySAJlJC8qFlxCwihsQOvz4bSNdNhbxC5D0B
E1ovS/g3Nyn8L14I6c1XugvdscjLhyxoYtXom+yh4j9FfKEH2k5eJnhxHl0JCuolLiDKRvJHk8lu
25DxpM2KgunZfWNgHRTxh0/29/vjDSQmTxe+V8DQOUb16iPOgiAzCTPp+gMNUZWrHMmSeNbSZugt
nDUQGFtVnbyx4ye2aD92HKH5HOA/THs3MzlejhacTs+UdupP6Fud5irhWtfiNlQT3zdDdnmldoXd
nP83Cj5oPVtDm4FgBvXFQE8iNiyIZe08EhwkukhEDgb8DCjcjo+ZJxkmyEUZhMe6GQ/RCD1yd2Zp
J5arCAV+Pfb4H80dS55s4unQDWeOzx8W4mfAzcVg/4OcPRg2P59twohZuffZ04HpPYTVdTrJVCAT
dxrGe0KO8FSiQ+kXH+xgnEQynLxbw1+JNmOUmbtlImBlEgQoc0JgZNKQAb/PP7lRWcdINjnqR9Io
ukIuJ19Skfm3Sc2aNoZ7jrxoCySXk0mL+vpyvViWO3j5SPhFj7Y+YICPv/t1+Lb5JBI/ZNQz90jA
Yvea/qL1DvjstJjomgasZkJwPfMg/my1hzRSg7EaVDhsOq0AZ/H2pIpm9WXNRNdUcHoNdZx1Wdfr
4CeTqeK3uV6x3GDDe5z8dR7MUpYgBmx7OZmkpCk/RHtqRY5biXPiqFTyVU5ucVboxY0XgnD0ppUu
dEG+SPcMEkeloqK+duHiukyZOTlhS+zQLCPAkNn1IXDS0MFHR4M/OtYxEEgaXdYhnCzMyeRpTih1
VVesj3ucl5yO9WttMVW8nh269y2F7DV3Prr5rwQ44uDT9sQi3CGQeakeUxypshrnHsf7h/2G8dyA
GjN4BbL3+NDeAC/wG/mtOP/oN+n9IJfmQdj8BdTViv1gpEt43YuEQay/x1sfT3iOBjjn6keOFLIQ
Ae1cSgl8c321i/nG+wZtnV0VK0dvIlieDa7CZ/wUzAQVs3EMkoiAyIJ1S+x5iAkf2mNmyy54iKIc
BOy6UmkRFMdHRTJ86/coXop8nI3qapd09KNWsV2nrElXVnH6/djBYJG9dBDpC9poeDrBDhjS0g4Q
yYgYgqAnrpZt9XjbxcLiY42UiN3CuHUmPKo6uQgS/nlmssGMxwY2BexXoth1LxZTzzpujuLxoM2N
egWPlLCblqjvRD0YHkj3FH8m5P3oIQR5NGPsYgmX9gQkkE+0Ca7PqBluPCUlWmPvTNXMkFC7hpso
PqACXu/ZydRLQycudDFvhbe09ucCMIJRHOwE0dUOtENYh8tO4heNs5s4+uRWEfbDXGWCqNBlffK4
kuDFx7vTTLZaACgs2EGSkezpIrVBLFrM1/yr0IwbSJ6xEqFKEBpJlela/w1twkZycG7cD078UqXr
daZQIwddsIOE73yMXJF3pEA4FAg2uLD92lnO66aHTuqlcDcFZN2z/DoTQYZfiRLxEtjN3BCTllBF
TMLm7zd3UAYvja0SKQ6LNdtMSA5jcoOJqJ/lcxi7AKXNgCCEPGpqPhphmEWCL5OjXuh6EoqDQOrO
ZCInv4+WP2mJof+Pz6BBMa8ol/mKUQwjBAlg1eHW2m/iGqb5522r3gpZOUqnw1HIexvDfLMnegP9
QOT76WoXda+fRPfvbid2hg48KjWOYzHmMdn22uGBlQuXPpbt6mGwO+OBgFy8zGJb6ajpqiJXSiYu
+8sQ1PYQ8EDyHlT5ZegZB9LyNNydxprGCNrXM2gyB94LuAPUj75xCw3fzGA31HcuhyQgslq85hWY
8NDJRyxcVpKyRV5fFWCm1wn4IaDBRmCOL7HVPZsBk8BehN6Tu+oTWDL23PO19JbHv5l6Km72bvRP
S2H7WWX7VaTwVwq3gaiXiOmpJ9AGP/NU5mEEmdEMv9UPWiAFMexnTTiVgw143c/X9lz6BYNWTKdH
cSv0uJvJmfnILdLo3neEo3FAgeYSvxOg2McJqbhyAGVD2Tv7YOC56iN+sTQ1KEV6NVXtjeYxqgKs
kYdpPOUobFy2JnlPG9D+/WPnSGxvFxBe0+Cq4LMX0zGi4gOTSKaaPjZObyBRvGZ7jJkQX2PD5JTU
rBWnET3NpMq6q0pUkt6aaSlRSay0r68pnE8BX9oTuZCSkETogPEm6YMV4B7rY8JpFpqSXaDGIR9w
vQzJgghFXwX7XHNp3UzP3EY4g9h6CL5q0iad0PLC2/8PAg7AekKFaP5fpoARL5TjHQKouY/7+e8P
ZqLfqYP1uOjoMnaDaXMkYS6X/G7mUJOhdriHOBr7Vef+w48ZvAhLaqcI3jU0ifmrprbQFkEZ2nQG
B7WV125O6iMb1xlPyfROZOcaNyjoGyzTIOU06h9S0iyVm824qilXtwpB6p0Zif/5jzr5PpzLl7Sf
IIrFbVbBcD6RNdpEkYP+jPlwa612aLyD3zqO9PclKCeA0Lre88gjT1Pv3my2aLNlrwJW5bJoaBkM
2oN64XtcA4NHkE3JauyH8lefgPffEieqq2hcrSpVgKqqZlT9M6djTFof2Nod4XoG8ium+lWMcPy8
aHvLeJUwgo+geME/6MeVajtAos60eFhaqh61u5DSKbAHKCvUnIPV86emGV/60xpPEDpvXbtrQqZ+
0CsiNuWDW/IO1WpNSU4kNwWoyaegusbXne61snzgf/CCFeEArg0Gf7iIJIBYArg3qVOT3/7wwPXb
kT6kiiy89iim2PQ0yBN9leIq7r4JJKCmdRCttPEbT+m2lt+LDyLe0PEvccFnQ8soXEgjNZ1DEn2U
3EedxSr8iPSsFAoSZSPuaBZXd113mO0ZpY1r+wBZ2WGzclzDBGhW6FZTNVtzQfqoreDt1ztZsiIN
tOAus+drxfXXZwiEygw5dyuG/dgEGzu5/JJSt5KEsGevMyrT0BQosarYS+4SGI3bf2ue4laMyO2F
RKQUvrNiMaR5IOD1AaZOR8NzQuOMSeA8Wl+5WJPOb3+1CsYTzgdx+KGE+n/2CB8x3J5+Q3wSJb5D
GSOyNhX/lfy1EfFiuzDEZSV09K/kjyzWy++R0qOGs27DgDWiO0hfp4l+2Hichz/ilLAp+xZ0LcDS
upjSNu3mXxSLrSvWF9x8/0IhiHDgzZiSLYkjappJj6JelVYJC6aDos3Fc13OdSLfbIjQazwDS81z
IM9dJUcns0RRnmzw/i/wMCKF0HakVmB4Khj+yeHq1AsT1+QNyfsCfKYk/ypSFHPRu0lv14SC5eGZ
0BEFw/pUwLkfBmA+JoWtJB0iIAzU1Nzvya3qDkkln06rM+ZDCY4uk4gmytDyK6h3bOt3w68KablI
FBjX5e+GKJEkd4hcejWP+8h3vzCHONJRDIdAP3eBU89UeuC38gWsT3MaJWTL3hGDfiVrkDGc2V3F
eZKJVFGlrFgqpVdSJbnvhZrDHtDBR4OxTAq7IWYwR0pJHayDqPa+dVD2CcCpXq61O1LNUXTON9sr
f7SsjT+LbMB0w6Hulk3rEv3xSCzWJKQPyX2FarmbiXCtMPe3cpoaBlYXKJ57tM9FfTawC6Sb38SQ
TFfb9fy73YNQhOHgGTpFzSqNaMpYGojN9OB+EIYOIHEEbJ/PFS/ZSFzo6/mBKUWMy+qb32/URqKU
B4OWOcXFiWaDfs+Fi2L8ocERqV953ENfg/0BRzxOFqCthvK3nTH8C4/KGFuT24fHDy8KNdXDaE2H
2xgTMyOAvAGGxuSO1IjduKRoiDXICXDsXr0pGbXvDAFH4MFr2gYNnWgNqU4PQTQz5l6/gQpnathU
A4LTuy0t8geHnE8e3jr4mot+XAXqHe1Qhn1046EeqvT6fO4dgkvNFtP4dDQ5hypsuDF1hY8RUxUe
zpcxZApmCdUtOqaT1ln41b2jQoqdF2hdTqDoHxEaJY/+wGLaLD9u6yax5Pq6BRRobZ41IXjCH6tN
GHQT1RlY4iwOsIcnTjoWk9ZdNsjM6CRuMD9sFxVbwqU3/4aYaYHe2PvvOmlRZldq/gCD14XibYAC
+ehHf14g6bpjDRQ3uH/SAh9bssHmLABjvXZBz+suYCVSvoPCs18ZzR2s/KxX00EDstJVuVL+UyDb
QGIxWlnGDhGfdhr4+08KVPvF1lgcZCoqwopW9lWVhvql9jdWIi3Zxz22EnnudBJlTJKq+FiVdwh0
yIBUL4akjBA+rVcP3YeBvwoWte0fXdEHXf4OyPXKfVNMVhKQ5Thckn2Lw93pkaanvIs2aWJBkTSn
TQYTHOyiSdVTznd+7eydw6uYlLxImHxlppIMKTlIQa/R+cLkTJmZKv2UAzAqsCxkR0jmbxrFGkTd
CAGBOwE5vxIM2w9RrTBUglxszOvI+fGRJw4Be5RJi0lXLsH1ThtXyRTQLoO1sNpAH4+lfbn809ix
zbiuB5Bz/ZZc2c1WDGNU+TqFmXgUR6wpgvkmE7ZHGz/LzcY07WB3goHNallybmmM5swAu8vFWihz
HxMG+Leainb/sNCpnZ8rejklhlfYqzddERas5DHEZ9tFOlZls4N4Cv/tub79IqggftwMB5gwn2h7
uMtCunXpDTixSWb+xGLQfowDoQbxxlxzgcrCYhNoLcBQBDXMjKMLrw/IlqpJVtAO2bKRKq7c5gN7
r4hQgjHLFeZfdQ9zaB42AJAab983ZZ6LOOY5cX8N/BGCWAaacGyFhBZZjn5ae+Z/hFTZs7mE2TRR
uNcySzWQLPkFSPKdDcbWzElpG2jZYK7JbWBNML6Jzt+gcgT4eDsmMAmVRl0J8vxxbWy0ofxTaHok
yAg5ARG+EVZIgH/mD3T+quCbERHI+IXP0FnVJotTtRNF5SN5ioPQAMOgfMyKFnE9+DIIJQPb1THr
25J/wPtMo1vaXD0EaSm03jToyUYhVklPMAISH0EKYpKR8wJjH5wi6tA/DfoKOwQ6SE+YT6oQxH8A
ThP9rKMxJxmxgzrYhKZIX9pjqcP1UJpXaFGhBLBWsHJPX1lOqMAQ77l+KsjzINlslDmFzD6UbDMQ
n+qOkKmLSxGrt15mbWTYR+UE6HlHShtmAdQStZnQsoG5ROh3ewyNb1L7fCyRUUv0ldsGxMCweQVL
ixQZH5VDEdElUYe54mOPIq+LkUksM0Y73sMoNAbAshk34UtI1psaJSpzCTFUpTtCKCqFAEr/pIIS
E0z9qZ7iRPgs5dyAI41EyqVmpLVYtYKcLYrNA7ClUTyXqtnOaHnpEMqjt6HmjC1uRgGzoqPhSfuc
B5bPSNoGSUiKYvrmUBAwXjca/UDQxoQ8uk7nOrj5BXt6CTGM7OwUXrSRIAGr87P6tR8t2To4GZa6
CpCUZdENEh90MHV4zJaFUv9BTnheXu/BHtmU6+koUz7ZM5p64Vvf/XF/tEZJGcaEmQEB5hfNX6bK
zdfkkB+nhUq/SfpTnyk4UJy5a9CAGfyBNKoZ0FfYpHugxfVuTVaLE6ErF2j9NaJ0B3qQH0QeIMQj
t0QpTdTT61FQMLIxv1evuVNa7Ro1ghtP7bQFgnaZi0PyQvwJU1aHdmfmRPfiTBYMoCDf7e96MvtL
76KPs6jKkhcE2T+E90wTPuh7/+ZHiGF+L7X8H7CoWRawTOOzn3mcB1ecgoKCM7pLnE0l6fbirGaq
pMV2rgVvfGJt1isAl/AtezuOSaBd+8Pj14ogrUpfRvxD11IgE/GeMxRWuHe0eqmshngDzsgNichM
/7cV/lA0ydMj1mSLm3s72LGmNurGs9UN1rw5gqYmZuz+4Xi99envzn/yIK8psOK4BYsbN/gcwM/2
FFgCQrSks13vvJUPJi6MnHV+ebOvDrBS+Q/h3w1XJOX71TQQAicxdRCjxWv3EWaK3ukEHrwz04Z2
1VhyG8GtphZkvmfIMAMn+JL1XXTnKp1XRzAtfOcbxlWh05gqSGfk7FmXrowxKfAY/7EJ85+fkBjj
7Ak46FAVPnw032WuhP/vuuagrETzAwMaRSpRxFiGjAiwAoywKQJvpI3Am7alepJf+V4JpHgXZ8vv
7dneJgMyhWmo67bZqPYleyp1HCR8GgkQRa5oHnvwBwELMQwVHvbMipjT40iPFhIDuXJk/pCeYoMG
ojGWKN61Ix9o2ytEPP1hp2zaoDrNXwqr3VjbvVRoVgfkKGGQB1gZfug0VcurMpgCU0axF96kuasx
vSCDEYPWQV/ogso8AH/CGowr02h3aABNQNp0yPtCb7NOSTZCamInhIgmwC3viu0ZJcTLMuTwMlJh
v3dNeo8JdqpRjwX4zYv3159oN6hEY0tOCUQRMscINsuJnw7F2JQ9iL5N5XFLZNhuJBhKRioRa6Ch
5Ng4SQy7PTfERgU3VNBOq4AsROAV+9SK17aEDiEQ5DeK1kF8njD1VhPOFAlL4m1c/YcFhK4LaRCR
oVAAHdIAdzdjATzVL8T0NdO3WGYf26FRrQdNmaqxSCOwQqKizsPyew7UJM2WpCKkMqY0GEkHrAQA
EDHuNs7n07+mxQ6XrQ+r5XfV2zbulGKUCCahrdBhTHH0Rjlyqq2yyB1an2SQXbmcc2NxusMer6s8
KosESykViUgdsP2J1e2iQcxOrPZb06nFlPLZJRNpJqcKIrVFsRbdZlysBvtNzIakBA+RpnlqpCPP
Ruu6hFRdkXKLE49N2HQGtgje4FfMKV5Fcveh3efUFGMYi+YlTx4RlwS0UEVrz1JBp6WniankmJyD
JTeTXhUx+XH6QnjsaqKJjIkHcrKeAedpLGLcix++SBbL7ey+qq0i/Wrx0BvBBq4vD5yy0P161l4x
ILsmyMnP9R0E0Zd3+V20QmM4rp2qTKies6cNa0Dwo7jpE6JH7glOfBGTPjDoHq4juX+GvM7UiZ+J
tLr9MskKSWfWZBn5saFmvHylc7/qru7qiGbPaYonT2Cry4ELcNV1BGxmPmLDQL+MJDaDwbunP8P5
emQZjv1/Fm2GISFKEf+fOjXVuHmNKwMDWA/o7nfZ1TnoZUIUjOHGdFIDJ7zfjW/jtyQTl0kMndYm
oo36inkQ7+Up5v6alU2h7EKd8v7cJsGIhElv63gSL5qJZaBx+2LeXoEHhmkVCQ8ZOcctChIY+Ex/
r7v8C8+zyubF5euqKA5Iz2AO/YGERDlvJ5JAZgIjpE7qGcZ0t9e7Xtv0FqraPL4JuBKDo0jJU6D+
d6gu1JpPmeJnjJmte8IeezgLnzNYi4fFpWtgSe9EEAp4XUPZayY3vPpJ0WAOq8tBFKeDB1fLBtE1
Du2ONWCXeUQeuLYSyEOlEE/zqVWnRlAjfDg4LTrunNrMFiW0KCIkszd4ld14oWJRF/HsQkITUpj+
DGyndOdY06nqfYz6uR6aLz8iPradlC62tlS8R8aoj6VBHPQ8K8H6xETZPmI7o8ua42USn33HWCO4
fOcZCVRZt/TFFfvLgTd5xHw+C+og3F2WOeb8E2tyLm33Oy84kMqd0puU3cm8lOf8YT7NIViW1R0T
nosq4FWakODbnoO9kkKmxLidQ/KSV9ACJOU/0D5kUsD3YeK2xCzMTGZLLk0uM1NZaMf14YmV3z8r
kz3/azXLKyChoM+8S/MN0x01EHpTXDI+HfjRV/0KRCgaMoOLSu+vPOXmRLyr2qStkc0Jq6Hf3Mzw
gJ8V4ZlHbh5e7PvbMVGi7wiNW6+SMYHDFHef9Pnc8OIMQp2TqbnccjokZf/nBgAEThZ05xFYZgac
tIWtNEk+5drWWaD4YeHV77Hgl+1QMhPZG0k7ELc5V/tBwvux84OMyfJBTEeTdcdgAqUeW8L574og
ZRqLM3SBf3duaQ57b2f8xgUSquGVzhYo/B2T4HtGlxrVkzwLiMNg8nveeMJCnjOorLevYfQKOg2G
bE0tXbPF6bnreqe9wKNDwe33H/114+aB4HinVPrM2XS86AF05MGUno7vmLvbtjdhCyOZG/r3KHy7
y+iwIN8xstqQmlhIitEbzG6/ZF7/2U9K7SpUBi62cTjNuDuS4CtQOJERpFPoM1S9KbfGdxy1sE3B
wok3GXKR/e1fp0mbQ/8QAx/ZzYnx7bn3lL7S2dxsPkpAYrrx6gMEYTFB2hKZI0GIAikDrbTiuDGd
NfH36Uv/uSUuh6TFa/jl5kzYdzTvLAHX1uob3usYkL/htwSzaCZUNAmgw/P94GU6DLkYmSEiQ6xI
ccricL34BL4fhtycQZxJz9ZfFKQskMt69vodpdC6AQ5rRv/ddeqz1VvFAlvU/PpG6ta3fw8AiP9+
VgOcw5MWU+AQPgFYPTPFN3VppBV4rAZqZPujh+Fo/hUP5j8PcPQNO5/undKZErITdJ8jbTvEjjmA
sDiQvnKlRUkKV0zxz/U9eeNCQwHOXn9Yp1Py0joArDVVIE8sSujHq71YSo7eTKoy9KhrKc9+/4Pr
OteJyUzXt8/wewaKTiIJzepdEdP1Hq+TSpu/5CxyRhN4uYfNlQ2SgVz1Ah2gsY3j6EcrPfVhK38D
z+XpJ9znz8JwBvVIgnwXAqrB7ryi0AfCKWgXQgls2Z9mAi3wHx4tqcEJJ0vbF4wl8Yjhd1UeJDgl
deqBIj0Xaa8GkV+2gLCW9wnWm1CpTqWCeF4xP+a5gM/8+gu8R+HISJHvls8JtndWSQDQ+sdPmkB0
RyDS/vWAxV8wlrymfVs5cVNbO34PbbdZCTbu3PJ+347vJWP3CIxTCYQgyclwdlk/4iI47RVsc0Ui
h/tofNEGTKQNX0Hso6DwLa/goOQPsCBIzclE39pdYZ7YPkebMyTxddk2M56BHX7+7SAPlK9bI5vJ
ZxAJqcLuiOPFATjghCBMVA1Eg+ioh1fs2bHQPLqlCojWrqRbmReaGBQHye3slgIgbLg65DvY0qG5
4gKPbAqIfo/uZmjxMJ+QkXMEVe/OTUvH9pRklL+VOfJDb5SyN52UgHW22gp8ZeuY2xkA6DcX3SKW
feLGWGtAkn7sXBmSFIT+4/MM2LsAcIYU3E+vdFDsnkoZztHivtNsd/PmyuinRG9VbDL8OSsACMCk
8c8GGzunQp0lzTElWkDUoBZ7OMnbk2Y9E5iNS7f7VGeoQiZ15Ngv1AlJepOPZT1nIeN/t3gVDYdL
idzQbuuoV1/i9v4YJynZa5GnX0UVEmxXgtIAb4zcH7w6wGz7i4Q+XdTdx0Q7DPXDMrvU0KQzjSp6
AYtZwqPMHTu+ke5zflvyHT9HB7KWdF6ylS+rZY59sUrxdk4ymIcMv8uS7WOUGwl2YLIZhI1NdsY8
r3JMCBvle8PW0unb0shcInU/2lEr4ZMH88Dfem15KfgcS7EBvnrZeXMJi6FUVealINpGDc7ft1Hq
k0i/8EkNYCTRbEsPItmKJKVCWRpHSL8dQPfCX0ldpO7fvmrvdsl8tD9LQnx+cR5UI5s5qNOz1WaP
XSolse5IkVz/zbId6A0hQKHdJIj/gZScRL0npyOYFEEU/brC0up+yryE1hbZ2VQ9pfNyyuoAg7r3
R9c7nvv+EptX4xBhrDggKJwlg4xjUzLV6WUDv/0hLTlSgiucoP7nJmIqnDN5I7t5dxTNknwZmgyD
tnkTS68yvTORQiRWRqs/i5jz+YiGaLUZU4Rh13cgMS1x26dtZoa9v/xH5DgyRUAkXlpb8vBHZK6M
e8JpwUbrVkNUPIBQi8WsfKGgNFhVCAl8nPUWKQVX1oSpH3gtbmHpljDf/NV3TeK0s+QFhp7l4bcC
VnZ7eJNI7ihI7oYojSZCk+oqjIlXH2cDUCHPbjSYtOEn5gjCOS83+Mm3LUV4jptbm5urC1xw/fOg
D/XYnpCjGhvYDO4XmtUAPnlKtBqwordxpvtvpWJ9ojT8YNRdyLLCfLXIzbUMK12N+EDBjWnvG+tQ
dys/hooHNQOS7/uKjgGOcREdRmL8iNYzCwJhED54c33hQqACyo5d0G3KBVm5fCM3S60rzW5eqCcm
kuj73W4urqNHjIpzKRQhfdRz0Ct3dNdLXcfKYj9KeMPQ+l/60qAHgx4qW7Tfm1ySZH86g2hvC9DB
9Dtku7YZoqoCbxrmp+H9h7Sc0kzIZg9DAtzcsH42a5PrVNPznkicr9kCq77BzLFI09IZSCbKshmk
smczao1ejVNTcr7CC1mLV5krA/PPbfIsq8V36MXA2AauNlQnMFuMMgJKQcqRom4Sa5OCpmaTeEWH
aNdhcJdjuSlsDjew/UZfAneEEScTRtYlFuN417vYE5ieH4DRope5WPY6Wd94RS8M3GFc/T4llbUa
fkHAHEiNhGn7aehkWBcsgxIk3BO7NY/U0s01nlSnVUWPbJscLOZPKZqy+VId0YVD2ew5ZkpIPA4e
qRJzsjG8Y4Bvuu0xc8cnJSuSX0GEIe+5Ehol8oJJsiC+Lji3xcWAeYehRbbnVZPhiT86tyblioow
16cKqIPMliMY/Q+UJcrw8Em40KjwIx8XFtphdsG67vDWeG3eymYwDl0f89ZiBJzc1n/zXHcekJGo
G8rIpHP3sEci6piHN8/NmLUOkHN8ZOaQafDk+nbqtpPHXxueqkSUybaBtSpiM25k6VQnfN5hCJvm
y/YB1Zm9HASbgTtMX2ezB4Pb+haNxNW0AMAmEv+PnKWwSPCVV/OWhqcgfrL+MGvD8wrnyVPbbCDE
+Rr6pXFDNHUWiSYqQrP8s7GxbdZgXQ1bLOqravSwmZO1a9g5oS6vMPwd1Ssb1ZnvstUGd7BVLu8/
EnU35Tq0gjZsD/2JaIeMI0hapxZYp9hjpwvNajb0kXhTe+xzeQHWU5oD1uuqXnw3Y6l7zTULCEkY
uDa41hjePGG2MTA97wDIOljdUyxJ5y+Joui/NI2YNnxpTtEU4ItT/QoQFZJyWxMrV6Kib8Ah8WnS
+3ETdGdmPzu9qSf7nl5co5St2Kw0KrVDOWQTONf2d28EryJ/moYLmPgeQq+CAe8FnoymepiTe3SG
a37mvzKJccSPUVuFEe+8U8JD814DpMDkLky2Ef2KFjYQyBNShV9i+N3+X0sHkWsCgbHW2d2SCbr6
wHMwiwPcIZrc2LoSVPWhgAWaLBxnlLDCxIgPP9J9sMNW7JxE9NeXzEAc2SCXSGNOcTZ1ltPPa2Bg
ltx7LmqfgXchRt2vZWJTVb926Mvd60vhNwkr70u2OaXb9C66qmgLjVwiR9rWM/uB5ynI7SmR2A8E
/mXIBC8LyB1kGnEozxWVlAIWLbd2PoMKQFd6PyTquJ3sc5fCfNAZO/zGrfwPk/EcLlRL7wWeg7Vh
hxbwYK3LLWsyIohSPqYv+gV56gzUW3WYW2E8PGUTrdKhSSuks80yeWYYwiQS903E0vm86yfx8yPX
FMA3Wb7FcLyTKZEdc+5h1BZDH2LSZoXNcz+72plBdjPv7sV37zyXnxOZMnESrpd1AOk960xT//mQ
FalomiSz3Zv49NzTE158khRedOzWqTneHoGtW9GJaZEE7iManE65E5m1X1LtMYvRzMseOJAdac90
7+69oLLLBPk6oR3AeLu+K8QA7DCwZa3tPQsPbkP+SkX7u8kuXm0M0QCYcztFzrsQfxiiqZsvZV3l
dOWSy2/itFyEBsIXAmnx+FigLVh2f5uZsLs6YnWBmVm6kFMM63UDXd3UAjVfS7AaaqnsgWvFSMar
U386jud1BuUqD0cf1k4bT5r+8V/edgIOGXR0uxmf4qmYGCt819hh+51KWLwa6rr+Ef4l6BHuafx6
q2b/wP6KmNXR0Bvf1lE/Ut6dgWFHcMtnAI80gkUjhuQqok1NbVkgZJP+9okX4pTqC3hyYnA15nDe
owXIPfQR+A/XpOX3mdZR4AK3Ct0rNJtgl1m2uP3lAF/+VsD00EDVhgiQEfyaiyXgYqUruXd2z6mp
u+n8WZnLqbeH/kZQUZn5hSVA5jOZ/TX7+DXZ89e4RkPQN3ABA4Opwub1Z2lchVGIJa5ajcZLrTD7
GNnOiS5KEUprM/gC+GqbbUCU4g45ac240j5ll27kO3MqFeSaUlLWy2lSeG91xD8hRBmCPdoF2QPN
NNzu+THZzUUj0C6V5RufOimlhxk3yUxlTLBEsGuXlcRa7nepbdFhPnRG2RrTRuQpR9it5R34uoxU
gXWlTNVwwmBpindLO0L9JM3aK++Snb8QsyPm0CXIfXLgwKKCuSTThv5X0DcXoKdPCUC+FAwHnlNv
Om1xoZucVWj0HN1wIux1DPXW4BW6E/aqitatlecKjv0LXeDTCkoOhdJ/UcPp6zy6wXYTB/gJBHJj
SAbgEe/s/9FTKoVM5z+XZnlNNjUOIc4CBQTw8u5SeZZ4DGwP7+NLLp1HgNtdHab3iHx/stoeGwII
ibVpVBAIti1NRuoG/6QKjPMyfjwAMxz0738843rPDfRHmaBm/p2WENTFH9ocgYSIPey0uMj8/mon
4foQbVSU7s6sLclj245oVgUSRNHtzKw65ImcGzvBFGrjm3Mh/59YDE77tFlC1BtPDbwI+gteAlCj
4tkkPziKcpJ3ZT3Y6MerjVXEOEy3yLSyrjaVHXbXWjHWNITUT3HYuaCkw/J11/e4FZ5MBc/0N7xI
e3fAak4gUp3rtn1gSr2aVmuq/LKG5rZ2FrUmFaUaDiLhgpjGhDOiXRHGW9LUfVmNs+0xgiNrWVWP
ma2LNCevVEChoJs3yjvqeUFHxebcitSP0LcHbJTeoQW5Cm+JY77BlkukWFr2lxAIdpZi9TCG3yRp
/6cdllx1SHOz4PSJGgs1dQQN6lN+ftEgjs90WGYa4GLSVZYiIeUxhrKJEetiIxQaGmWEAQGKD+7S
ecdqLyBLu7a5CJ1BoOrYa2DGEEjT9Gn5bhKdQjASKupyyC8eTYFAHOtvDI6lzS8fjUIGDpc/Ypfo
GhlmSX6nHIG4aH9gU9INiKHu9H0bzHYRjCtLVMomBmfAL+KOmKV91t1ZUALg2/J7xBq+thbR5hh/
3yGGVgPq4iSuuh/luLmSzGX8eaY5D2QdIKdWxDkZ/t7rNGYtBWDsf/8ChZNQZpLY2PFuVtR4vW8p
dxBssN7e5Ols7Uxw6NThLmBaTiEHPtaAx6+XBFsHPbcnV1Nk6TDF7Nkpp14tEvRb4kCTLf0HiHDS
adZ7RBSblGSQINoK34vjE9TJdgjeKaZgsNL0C/dI4iFEm6j332bEN13ph/hv/47x/DeQ8tpAGcQA
ORdgpe+ew4iDFIBEEVdM8/JlGMbRxax/Kfd3tE4G23JoL8CQLX7g4lDGREigi0inyQXOg5SqEEaK
Tl8sXph5zEPeE43q0a4So9BQlffrEodlFMpup40+LE1MSieClXu1phzbI7G5ZGxWSIz5W/it4itq
50cv+110cOAjWbXJsQx2QMR//mpKdIRLkHDZNesP9VbiKxdg+ltaS34djSjXEK3Fz3XOx6DmOgNr
YkzC2mniMzUEg6GpoZ7nJKI/i8B7lz9TjcEBCHK+uo04WRbGyDoY57O8v0aqmm3QQ3hIW+9JLg++
UJVn/L8ZLrFpmMH+8gKjZxdgiTEhWVXiQ1C+PvyV0Yuzg5YUp52+C3LQJPxG1qzO77Wsx4NnkGw5
aSR2ycJ1ViKG7NTgyKUVl5hHiWcrj87weUC/m/qaCGwnfyqgiuK6NGTsBVwfF8yGjSbAD7369JAP
qmyx4Jmt4UGRhg1j2AZ8FxxP0wctv68uLsKuudt1Yt7511MxJ5cwKtKZgYR4CGg7GRRdSx4PpbYk
7aT8hy4J0H+c7Ipec09dgF+M+TBMJjORESKc+6JVbkl5jMr+F8qHPp35ozOkmbtWsW1aVo6ofTgh
o1gE6HgyzcSTXnkqk12I8VnPtHaLDPiHZg7UJrsykMaEMOdy+f7rx07SVffr1WhM1/KyQPqEgtex
nlwZ/wLZ9jhoiB/6Ej7mPsXAp9//kqMSzPV71aS7iOTx7zueFN3/m6GrHqwt+CsepGEpf1ak455k
VFOi8uJboZkJbshbG8YcYCpecfCb8F5gOf1wHEs9jyFkEzNwZZIg6XhnN+1U3FHV+pPa1ygRFIBI
NAPf5lUnh1+wqSIusIPhzZKS9bP5QIhMaUC9alW6JiAQxp1YqautIvITLxkG4rldldbP+y2HrIth
nONInxwAXAFva9Y4X7Z7DMwLSz3ERTiJevv/l4VH6qbf+bv8Oy+dvpC173Bj4y48OBgAbB1dvDYs
KNjUqlJ3JKdui5LHse+WpV+ZbbGPo2QjBroSU3KXbqJPrOFtOLXyfMh0kIMTQ173QlSI8WGtBY92
mvwIXJM3pI1ce724Dfw1xaPxLFQe9etqARy7yCtA/NY00S/yLs5n9TCTcH/eBJxKucy1wTqXXWeh
FV+I/PEl3vZEW2AixxBF1p/SLEDVfL58wOodM1Bk2WE/+dcq4v6o4+fv3ntbJfVvcOMSFmR4AFXy
qsSlZWz0iRo07bEW6GYX/Buny91qAEmZlkb7pGxJlhvewTZSjHwMcBy5zwRQQzigr/ky57h+IjIW
uj5hElneVLyD9p2tgXTjUclrpS/cVFAPUczE9QD4ogSe/0Emd0GA5z2asLw3MtMI5oqPcQsWssht
x1twQ5oflHIhnbBlAmLuyqb4+auSU6T2UVblNum4KQ1+RJCJ2FTJtfEz7ujpcYzRe776y+YIo1r3
v0tNM49Jml6RGqxF7K6etNOcm80mpMIELgArswxT3lv8DTQA43mQl4i6l+BchzRHCMsvh/owvp1q
a0nZHyXOH+/YVMs5fmGggb6GVYszLmX/QxtjfYGYK9QLB+h7yyfv0ntFZ/rCROhI7jM4BBV6c+90
QmWLh/SuqUwUdXmHs1m99PcWaeOOBxUFzwL+jyDpdsGlraFrvmHfo7JgYZGaV05buqFOiiqwD7Sy
jbTJNcLZUbUGxZFuYtNbnAVYr6o5w8/Mw+FOQc8V4i4Rf4MA52lNsvKyaXFshSk8PPpPqJ8IDCKV
l8eQuML8R8CUSCBA8iCnizbEOuOXGyevqiWF6QR2eoYhzGlLfSUnqPOqE5J7SNeu51BWutmGbRsi
HXBMCy3QVJKYvtGUUqPewcbhfq4MD8F75Kwgps9M+LPmgrqFRgzHQQv9mEpDrch2eJBlII9UBHwH
EWY2Z78eIQhLIPbmCe5DAyMnJvMuQ3wb5SLHsBh9ubGb4mKwVy30QAVOURk56pqQfQJ2yGJhXk0e
c5boGahqR8BkVGOQnG33dzHDexzoOlJGmp2IorbEmck8VBy187q/i0oBPJC+sDFxGhPalCEkjJjp
Euxvv4wzC9oPCi7Q8E4KTZbfPI6Ko1pwAfdy1gTmW5Ycj95deU5Oo1KSKnLWpfjmQ403azSUoDzh
fFL7MZt+1rrq9/X3p5LNOYKxY884bfCgRX7d2oRUQxbxxlFPDnOIzxfzv6x3S7NEzVrVVB99/hP4
5jc4wD20cBtB6OEwRvF2u0wd/TcFZ3zaMgpB42Epg3v9YA8vzm3s6+dGuLyjC597V/tE5RNvNMj4
+k29al3YVe3F30Vvp6MEPUSp3zcc1yDyTAxNDxYytVqiHoCCiihJuVejtIYKbgXSA5xhjx0bJCAQ
m8IfbPmkY5D1Zo4uOBdD0m8vpMWmd0XvD7fJqVcz3q4uYvWeCWkOYP4jJL9Cv9khEsaQnkO/H2SY
iyFz+1f5cQaN3gxC2fu7W3pBHf1R1ovHLtLZ7/Br3n6gbWfGdOHw8Pwxs7imlBqha3a5x8rMTLZa
pYr6f0MoJ8ytQT1T84g9cFbOZo31garsYEmKpuXXsKdVVskKK8ujNPs3ecRaGX8hi8KONRyg8XH+
Lys2NUH7uiDscpVrw74Zs1REdupyN2D8HyZAghufKgafinN5Eln0opTvmPy4MOoyL6Ccm8vlXWSb
KQK9nnG1R2JNIGkK4F6lyRRBQ5TzErYPv7wsAWVAPgalMIljOP5JSE7YEO50miRCDe7tFa2nPIZb
YBU17YBWqxU7AWSlu5NwJjVfkpJx5fXNEhbixDXdwM01P8y8PkyUcsu1V4zSYpHPjTp+xD5DO4yX
3nR3yEFc32m7AY/weGryOQVyRJTLjFHThi+w9P8nfY6jS7ZBkrro/WJILOhJwUkACeGbT7wzzDlt
wY36SpvHQ1SnnVvB2bN8J6V/KtlkcIzoORjziJXB70kOga7MWh4fu/8uff5EM5Evn5x2lS3FTxZg
zttOWGKWhhBfOZzxKMppd8ayFfWCvpkJZV0UBUmlEac75lrEC4C5yPU4gPa4DGz63RJbljy0wqAr
hEE85i8/kR7j9SbtPFe2uKAibrO7SuPBd/HkYAdmV1efwHbsSmzbkfMgiWqXzG/9M+YFPTOMVugp
K9ym/G+XPZULCjZGEjxzb3rjt6CkWlDPDLl5+27qICKEHAA5A4yPp9UvqBEVe/jOT9CDjvA73Fdv
AmipCbrMhb9NI61Wygk7dakOon0fagFRatmVgvht9YtQsNIoRLMsRfkprW+NoQ9djfv1DU3VAPB5
xVatWIxa8sdkSAyvcIgTxznwpo9pqC5FvranxiZsWQnUSEgukegcsXzODMVMEhOJlOqDquMZR/At
LKxSjQfdKPujsmciZeIakaq3GQ+PiS8zONk1g0M8tNkrWQTS9S7jwXl5tFVqBb0Fw8uyD4RyjHHn
aJ6G9Elb3yPOYRlVmDJwCBXxWA28G9k7v/6YCMB14vW6wGUB5Hgp7npGj7aOC2jWnFd252cqMjeW
Hn9lbrH+bnC7izO5/D+2mzD6ydT2gB/TJfezZmP8xhQRFY3Zcbwc7kylf24BX3zFj6DSsIUs1sJr
8lX34yNYaiyZjfN9fxEM09lddTV2dxifWYM7nvj35doiG+PMntClGyKdXBYxfQcYeZVNNEaX1czv
o98NMNXDoZ7mengmFHjKGsHfG18tfYzGPY8o3kIykXuc8Y8pYKqOn39HOUJzi0caxgKjXh2YO7N3
9s+6vR+kd0NRlbZQLor8qzP7HyWCD2nEEEYeyBbNkRPgKjQVdLZaz6+jbjR3W19iYrzBGi+OEu5M
wLuYjdAavN/Sbf2uy+QlKDsFFSPU1hGJ5EsJnEo6SpaaRf9NWdW+pa1kOydeB0CAnzhkGAloFwWr
k3tavIRYgf7mMV4ur2nKeRYd7utcjNtw919l2t/0QXfrNgv2FYRTKf1YTtU4/UihAEw/VzYj05qJ
0gIdAHPchnXBBziPVrFg/Bsdnz9hYgVmd2cAFYCnB1Lznq+qQZ9v1LFBfpxtCGWB4Od00+ixKMCT
5IK0yea3swJ2boFaMiYJZpA7Jzhp7ki/GbO9G7FoAjHxcttEMWWj0WXzlR9VFh0O0ng1/iymHDNU
5MmNgaTQqJIWah1V/S3SXcFkp9iADAHwNRvRdrYgaLNUIPmqxxc626DJaNsXJenOD4b2ExsLdsAA
QIkm4k2MF/dAd6e9By7ojD82/gie3MPY+AX1VTi58bBNPomm26jPQUozaP++RFPHqoGkjU2j2sAb
DtVuHw5tNi+5H1PMYeDxywH0jiYxaGeXkOUsFSVBOf3VekfbFYKvqkm86kYgnSh6HV2JBCMQPp1t
Koq3FhvQaq5/ZZMbD7pW2bHuiB5oSEAv3HKaskFBDkClgj6ic6YRqnC0D7oUWUVoeWbHmV7C9qAy
QJQABBCBpjEcN/uaVDjHtrF93I4kuRHMvCSHMWCYRiiqnI2gIjaXP5NViDZ/AK91Dx4keJW2KKLN
iwdc1t+xlnRAIqiGmAU7NH+V5tmahIrqIzSGcsYCEQJMzcJ1P/LlHp7T4MdEeFt61uQeO3GDA96Z
sFnqSj4rvcsYFHF4fqG2EcS7s3ySuT6DdCqGQj7nrO74fWANjM3INOe0Sh4XkvDySp++9zoB2fCn
eQRfYrBWygDd9TK4Gtb/hIftHfCi+rsgmDoSCa7DvKRKmBVTkth5udFzTUqOraZeGrsfHciNW98T
T8BGhgPxXCLUpTMPnrPd3hJUHv7Ge6RvBeJbFZNwlosrESed2mNOxZao/mL4yQW/rNQkQtzSE+Kz
xw6QzcTv6QAnuhnQrYYYjjTn7jE1/Dagoj5/PoINB5FOgbBREtus79W/YaJ0IvmrNX8Bd55epSdV
TRKTfvcIR0ToVFsAUx9DCmXutlZSGezybqKASihGxBsKjO24VE1aL+4SEUPshtBqz4qdK4jNEeIN
PflNwBybuom4LGK8gziE+56kvaANCy+quvqnGYasffDr1Aev/KnqChYpCatdo0MDOCAKynAMx3Vn
1xs9M/g+tEbI4J+3ezTKNip3LgWG1gnbtDT0zc+yI+Ot32PDk42TZLkGHyQ5LNaWnBdG1nW36oHp
7LZKWbMvjMqlVliZqEJUrPDQ21kLldqoBF+UyUEddVynXEIuoslMOWu6JqniO0lJw/Fh87YnDSrv
YGH9+fhmRPoYaXyjocyQxKjeJJ2EUhvzzvdRdm+mLMUv6UdKkFzpXE515wPrqElWD6JgnJ5k/NCT
aJ4lIiY9DGKBRh8RNNNqq32J0R8JzaG4e+0z5xDd2gsTwoY70VpRw/CEM2uXabax6pMHyhgG5U+/
HZfb9lSGELezd3aL1Ym4QCg2nm/k/Dl6e33nu0/zSQEi0rYVkqtKv++yOUpeuwxKgEhDHoHPskA0
6Gf1YtPgZwMsP6pvD8lDyEtZbG/Jrj4RRSfQTdhHM2lRM7o3OpQ5WLgTlO4nv5KbPcDig5HwsX3g
sDvG61iTQTxHn0gtzBJVMha/lr/wxky4YcU3y1Hz+r9SrJ3hSPYjz7HSsMwIUglxpOVkmvoKtXqT
Bh5Yu7jZsZbEg2xYy/YluK3SfOuN7QcxSOBKyzC2mNGi5Gc6m32I8ppeV2tB7ZoYTwNLFmtoRoQP
zK/t0+BGXh9+yy4kj12aEJEtbzuvT7Pm6wFYj8O5BRmHEZOlzAdct6ikmgE1OqI8ohol79G6ErJo
AAMaEiIXMXN5DcqDe3yhKQntNgPKsqzT8WnsL01aCnNu4JYq7ZLdEaq7CpZgWLffrWE+RkwcVrzZ
zTQcM3Eugc5G7mCA6BFy02wQyrKriJ/SMlHEFl2rhlPZBNpxgHIxFqNQxhIPTOr2glcPtZJe3N8d
VXD671YAfzWNRQ2caZvGAFNLytygwAbkxBlibmNyi4R8olYRf/V3CxFI460Twn3DXInTeZTdJfER
aKKSK8X1sC5JEuNln7qbyMJasMHfYMXLO494JtMfiEZHzp73zujOJfIdY10bG9BEuADvPKEPgZBN
5gWW+PpXkrK3pwfAWAf0ccI6op/ruGlLWd3bDmfmUINXgueuif9YJ09Ap3H4Jragww4BXAp6+vIK
sJP/L+mWFis6FgjHlwLgBwwARwzKB7PnL2vC4xwJblVsesAXLFj/16lyKswjuIeE0u9snJkls06z
FJA/vunhLFpXG0I4sZz8KiEDXckdqbKQqz4a93XY/vqDbNP1dYoygLS3DxXuVElYfZXPzbPnyNZq
UWM+dCy6tlPPgP9Quo9v8qyk7xhLA9XxIO1EzyWC+3vIByM85cF7rPXN8XDcO0SwlXZ+Ra6GovtE
j3gjZ9waKw5Cs8qWdszSRPAvwea+AuGDpLMzo594ALlf47wI0KQtY3tZWtZXpxvcW79eKmxMF6BA
+Blc5J7MOZcUp2V5iPeqNCdcW66rsdji8j9U8qAitXFkkRPsbZN5pjVft7J/2djmxa65GJuJ+OzY
I4yCd2vTt1DPA2bjAjEArmvUzQud6qgcLPLztUZHU320p5mpuZGgHL5kOZojnh5WaxXDn7BQ0b5c
s4P8gccr/u3O2FPBnYMckSfrcDYvyyysJUwW+b2VC1U0afPbCMlijqkXCDdVzEOyL0/IbHgqo/EW
2G6oLBs7+dhNrJc9EdfTbw1YsmtjI0we9Dz00dD/fl0+OjW5Wf+lblbEa8WiYxVoZqCTjBBpDEHk
z4yN5t+8tWljhq8zByzmLW2QNDek39noG4Ji/t3sxfMw0DO35fSt6y3UM8QBnvpV4eNVnVW77ARn
FrVIAJ8i/5ubzqK8vnzPs/S9DXfk1guRPjrIVGSLWsj5ceFOA5l4BeUNXBfEGwlsiBtWfZJ6qhxl
yDkruKbSOaRP1pYNGP5gWHKkA6ktH1rbKseCTjRagS3veIJpXm+2J+63ky3Tftf/UMA+1sC5Lgr+
VSHdLXsnZ6xhnjgosR5ipvhIoetpU3cowX5XD+Tjy16K9NM/4dDrl97miNMAyhfEPFFCXnXvAX85
ij0gkT8K6W0CxTMo0GlPghczPNaLt3+NIQntWkPxY8wWoEPgKSBW2NLES7v/KVstkw/R1u0ume7C
cTk/V6xdCOxKzN0K6QDSlcvcAFA4YXc15Csi6bUz6yhg6UZWdkhOlLPN64o+zxd2d/ErdT7a3Rjj
p58PnFg9dwS+DBiMZIMIChm70Uqcwn6yGYA04gb6Xtyzw5TGg/K9a6zZxWftZoTfnIsKv1K9nDV4
S6COlVANUGuogt0MjCqUEoBTn+0RAjH5oM6IZFUgOVtbcvTV7/qSiy1m3bk7ucXNsH50Wlr9VYsc
mdvm+Mp7+AmWrSixzZdWi2MOH8OWqs8ts6sIZNNT+F1CL43DwpOCloyvJuauSCE2t8y3+DD26q3p
bfBQMwGHrXv7rWzuDXjmeLlubt5GMIe1ODZ6Q8GZCwgP7tSB31FXjvwKFjPGO6mayb/6sOyUUz/f
cMN6B4hxXKmFTZ78BoZ4WD1HQ+QjKb5Jx5R17fcnspbvFVbSQcmzxNVxlJpJicMXmfGwMXCL2j92
oaVp8GfmHeggjLkvTNPCTwwgXZ+AOrcBRVYw8GNmAOu4FsiTBuhDvnAtUaRepmMxB9NdDEK5iV4z
I2t9hHZbiXv8ni8vyK+e8KZIcCQRQeV4Ft2/4IDuhgOmV38nhHlTc6vvBGKPxm1ekzHpErDb4aqM
GtsJB9jtkAhhixioYHjGYxFwkxcut/DkiWviFSE4fVuzRRtKrMN6UZQf9ek+KN/Z31wLURbb+j6s
LcqhAetTULKbiS8FxvDR834hkdDw9QIelErWy3ICX0AtUCvfQb4tg08+Vw1Ajl32VJb0WAgelYYx
W6Bwc4u65ZwM/oFzh5fBEGGKrnqEt657zQiIG/l8EAHtjEFbW3Jguyc3AOHRgcZyRJehzCbTexhu
1rvRSuuwo6XAR6PLolxFFh3XaO9cf/3mqPFBoN6G/4+ubbMHNaf41n6kzitDbxjXO76L9aXfFj1y
dhMutjUzTZTnkEodSaU0LIKW6oAl4iAXKVGsLBNvgt0pKyYHxZSAUBaJOT3s3l1jw9OI/rxAEHHN
w33Bzdwc7iD/OwcZhJCFh+1BE86CR+nmCFEvgzfT7n+XC6Sf3NP5/TWGVZgjAABWIqMsZ/Tyhhvs
Zk8HuOBR8MGma8IsIUNva5SRZ5ElKWHHaNjPJgGLvu026u8hpv2e3DgdVofAXNqAM3FFftmbu3Zv
RMG/pHQYH4FOdY3DvMVoeanAyVJvEXxAq/0LQTFaP38I/8vfF82z3SCWhHbZLt1NwTtVszjrqA5q
2GjmtkUK8MD1UgnVaHVwZE89tH3iA7KjidjrQPAqpWmtxdbd0bX3YbBsNVjnqupVDh+VGZDYJd9O
D3AFxxl88ibgsu4htyVAZqaPnnyLwOKAsq5Tgh5eGGb9MbMojjEYNpC1k9kxbd62kRbuCWWyisUY
fVL4ZDTd9EwtcxK95KyVjcOcbAWCMwnSRbjZ74GuB0On+k4uzzzgkP7XStYEJlG1xUJcNq5Tdha4
WSJ8HmPaM/xhbISoTHUmr1nepb69/Y5YRFe6sZ8484A2uoKebOuBR6PdmslJIA2zaoctxo2z0Qa5
c6Jn20zhmkjaCOTbB2BibFbyjy6thFh0SxkHWSUIDDulEOBQLpKteo07B1oaBfQdQr4vQdh1fgOe
TUKm8wSVJotXgC+hVgjWXb0PzGXIEs+KfgbBMdhJBGxrpTh8FSant45PoaSzVOnME+x0W3R2psYp
y+SxepCaHXL+AdH6WxCv0VFYc97p+vdXGp2cMyUcKHxhVGTLJyX/EAJG1AhTWmDmwcPPIIKiM0+A
JtqsOhmxOtO071cHWWYfXEm364jYUSMLY9vwbbvy1SNmndqRkGldD9ApAPs3463v2N+7Hth1JSGk
1DGUqS5qYijNCI4zlNuTzhxcYthkAgzQkhPKSzfJaFkdEPVcuEKota7lN4F4O0rBRjo/LGG4Vs2O
TQamcTPww/SOF9hn8m5P3i1/mo9ooaiBsJ6RT/fpP/wNRRZZkFMHHO2X2gcRoprzoIMXFfzvrMK7
9Vh/NF7YiA7i31pXUsDYFDKGZYD//M1jfcrnG9HoFWTl2cu4hgzdrWzo3H78bRzWaJyko9nXZYAR
J4X9EXO+Jjq6+0noYllMnbgdHEBuJyCSE4iIvpNvnbjAxwaw6SrUKp9029mAbmLcZvku7BCUC24D
MEyV6MspCnIgs3K+34IgO1/u+KlxpFclfWWxJ0WUXWBNfQ63wkIEQVxtTBbBrXkZN/A5/ex5aJSZ
/nfVSx0WuTUj92aSl2cg4kfxgK2+BrcQ3Y2scIjjrhob+RZZ2FqB0tNBdc4u7mQKeX0MeMNksW7x
sxkAHnlehy8C0tEDexad7E6AJ/RiXXbU2VpmxWSAfRpEquMLbsDgAQ8/SLopttLHvano6dpDZENq
U9dOB/hSKJG918pbxKFVzTy0uweRY9Ifmf/dehWWL40SIIrtnnfgw3hJ7pP1otJXdsXp4Vaem0ez
1yNIsycYCyVeTgNrTZND0L8wTwQGyA7r8ysgABiYqtHLWNcwCPaldi29Xr8J/1yddAOu1s8/TdgM
v/41CxFmSiyM3587dTmuIHsd6taygBI3kab07kLnYifuYG4QCDdw5w2sQHkzIAhXpZ9MX2T3W7pQ
WiENmgoc+fWslZW5XRVFfc8eCBntkzFJ95ATq8DJ90BQ+VNzU3URfxiTEQcHIWsW8PIcS6ORkdaB
vAWmQJp74lHNaSzpHVVmVwmczYQsKgtwViiUYKyaUxbUzJITO44D28lOnROTa3tfwKFbBPsbFnwg
w+c8rdt2qPiKhzFcshRR3jje257PUvZJksSjsVpzGYjok9mKVLNXWnt1+d9aMf0TcCRcWl03QM97
Pu9ibS/gcy0HyYUS5J5ZWXvWo5W1Du7eXqeZrSPIsYq719GAp7f4QNEy9tqYol+gyKu2bNVmcckZ
VMSywa7krAGpqZQKiPruapi9uECS6cqFXht3/57cdJPKzwrNfzHVtUOZ0Bq5qFcuSfc4SrEh2tJs
4MtAcNJynL5Bnic9zz5ZogzOdmHwun+YupzzTX9v62YS13Op4MJ+rBrnBaEuhr2mBwvYtDc0HqUE
+zodPc+zN2MqycY0AfnXLgfaTd2lLlr5VDb/0wa41djaWw1ZcM5QUzvm6WEwXxX70rgj7jxFdDcT
/0QC5W3egwMjBrFK4h4ycZTocQ2DmszFWLNAZ1dXR47sdl5y/saLSnOZm/Kjxt3Y6n0y1sspASal
MhGVr09gX97wxoSE+qtkyFbWORDc8CLqnLSTgNGUjCnH91Fehyh3En5J8wHMw2iv486KDgzoMvTt
g6ngdYPacoz+HJHDQEsLO19aR7dXl39OdeO7VJVpsIMjRBL6+avRPF56y6VQ1Nmjus9xun9RTX3Q
i2N8bLaNs5NIzoDwZp5S+WEzoFUkDsIa2/owNlCcnq8ostxxhaIaHr5hnzom4PedVZlheNS5oLgl
UW3MZy9hZ2wMa88CGKF/2IBGxWjmWxsLSmfspzXD92xtkX9sOCUudJKFm7aVdRxvY0npJP4tV/N6
Ef3QNLiBkT7f/pM8f5lcR1YqNsd57lJpO5vpLTbW6BAxgcwL8gY5lzIOotRND3NLbcznAjEStDVR
P7/xGeI8rwvUMuk7HjQSniYsEMcPsUU90shwVknXYtsvVtb7+2A7dymCTyyNkSd1PjMi7Wl3n3ay
NYwKbHVqtfJUxcH0CIQfB+fFdd6561xva9seuDvBxksRvWz2ti4AS3tNZ6P3AEflFqFixybYx2uk
aq2wBNGO3XsPYVSEP2hZlwrhad46NQ+Drc0pOyNl2c9oobhah0b/qs0B+7yIFEoRGMR7DKiN01Ke
C1vMRT2oxjDnN5Xu4VAdJsDS72TwBmN07e/oHytustX8ylPo9PW6fWeYSCMp8Txri75oevglFLhM
r1xxbX3q7e7+liD4WmJmH0/11K/SwUuQWaSUkENbDiJRTCQlPpby9tBSAxer9V9TOPPsOiZo44aP
ln/Rbrn9JvNy3WZ0AwESwxKTCeyOi8BbYdozB+VGB77Gwpu+bfL0cMlKX0dcaZVhHTXnYkGrdNNh
nTQoOwj6ifoO3DHqV1kc82uHsN5X74lSO7z/N2KBqUqMuLVhFknKUJv+Q0CknBFYNCttJ1dd16IJ
dsQmqvEqk+TBgxChyOmlPs493MgJA1cjCpTP+294uJ6hOUTd4Yw7dgNrD7VOwLePAAHO+5z7RnAE
EUx5Dq60XOaKwUolGxqSbjr1ElfLvv17W4kt/JeTrKD3HggidMxmgk/JmzD7brKQvLtAD4VxEQeL
XW3RpWXZ7TLvMzg02gQ6vd3/ZZ0Q9zWW1dYcqTxWf5za+LmDKRDVjTn8pOfMtnBevIsMJ7nSvMdT
gDDZBGrp0nT117E6qElE2IbL38SB3wztmiW5jw2YYwNguOg5A9sZaWHy57UwQyaHcGt5RQp4MtZq
tTYP9ylNvjpmhHYevPwcH5WROIkrYA49up2Q/2mtEWEmxlwbeE5ReyME6uw4Eqkyfozi8AzMIL6N
/fuXrK4znEovO/Q7AyIRWoqbjJoydKoQ0+gwcGPOlLc7t4luSrIGUFhQ0BLaaa9MV1ZuTc8HKkt3
zfzg0l4yvk7fAmvj+ASLA6x+5AVHs1NKKGaXni27gKkCsTgz3vqWYzNqJGbHv/pEOKXckd7RUjbl
GQ87HOWR3DUXm0VL9d8NuNRVrLXX8lwdSZE0ZgvdBtQGgDgpxhyfUCrS1eQnFLTSWQSytvYEnlAX
2wFZ+uBrA+JmwVE2YJJpjisHaR5iDwVHxVizZLT9jT2PyaXL8qKRVrJ6U2ES61W6qQGLYgxomwjL
H8/zSXjJ8/Hp9WQURaZq27ZshpR9V9+vaNy1uXG6/v0u7WlqPeCrkzGB9o5+fj2g23mfsmrJnunU
eAc1cqZ5PuXhSHuzXpOJ7zZ8ENkh8McY0ew2I6QoyTJ9K/8EZRhM28shI3JNXazS+HZOiegaSu/F
n03yoiUODwAJF0L7YkOikDTVnIP0JwNDY78YYYuwtVvaQYjZxCpi88IGqmAWfODHOUf50RuI2BDD
n3d4/5Db5L1pCu+wr7pP6OsO9N5i2ZGCmw1cm+f/wIjshX2rT/Apk+MuqSUZM7eJkCPyhfi5RxhB
Kcm8v+B4VqgyG1KSXqDSGEDmwOgV69W8kJ5IIK+Xcgt4MExo+jnYKFB317cf0Kj4G5wU64ja9QEG
wKH8jQ2jHsxVhOGCghK9Onm0K64CO0XXUJChZnFORJ1KPzKV9/6fJKXGUZzztq7XIHp5dGGlbtI2
cLmET2Py/3e5/+d/NbpDcpaBW2Vap9ttMDlz2VdO3gqF9lbE7Q1GH1sCSSqnqVxZ6A4Xu7fJ9gdR
ztM1SWGsEWN8xGKFL4Ucwlc2unRoZpdcyfcbnLQFd2aSpXtkPV5Strwe3jOHrMSjzZGm5nY8XN1Z
SM1n5nOygI87nW8rmVZf4lqTrMH5nFwdlAEPJVueAi5plJAedxKUiGl/AXevDemJZY8xJdRQMK89
38iF5HfTnpnj+doNeUhPH6/NkVxBpS0DzJc7qYYarR7Z/2kL3deeUJfjrnEKBr64Uv3t+QL6QsLU
KHzHBqGE2C4PrIAurSSFqAHt7aZD8y/QN0rW1iHNnvI+CLSAKtudqFgfZCo5+OTQX/svyiIWszwp
wgz+jVEwidBzhmk0U0MicZ4gCjEnjcw3aQquWgFFg4BTuT6t4bnvg5ct0Hwm8eSKsebS7Y9HCDIV
aBD67mwTTHHDewILY4cUt3AsxD8F2eWvzlY5EfcMGZPUYPmwnbCc2HUPL3jbnSYhJGxQ2kMmowHE
m8gsLFfgZb0R4Wg9tVSw9vSOoKbtXkGoTzJW5Tw89aTDIzqe6Keqon5xCXq1e7poL+hEr1TUWC5N
3n1Qh6toYL61oD3x4axHAX9nrr2/m7MTgxyZPi9Tx6d1IjGIv2CjKk3sgQzoRLrUJpx6U0Ik0gJ9
gebLO8mBthzNnClr7TqMLcbrKnfkYEDYcCnjNLbaBX6eEBMtA//KjQr9V7ZXySq+625cXX9U+ghN
J4cAdLy/G5mKJPbEeRLB/wWRVDfxZZEqXL+GvHUYPPhAVHLAb20bSjb0G5lJumZdVrVyheQoTdPK
mKC31/7uUmpbRB6FYxn5/JhMp/QVutu6PdObKXCH063tqTsW75+92/MTH7E047vUrbIDFp8SrF+H
vqpk9SJYqgZtLsEO1UX77RcTXlYf1JHWxgW9w0foW0na0NlWc1EKZjXQIRAJJj3r3GAqa5xKwX9x
PESOTbgnzAXJMTLOUjF9/ItdMV8z5ayydiVxpsWhDM54Py4VR9I8xbi+gC4ZIGrG7ilyxaIELJTx
XZdnh/XqI1VXMrbFahBFELB8Pdj4CEi9fOOHkBLcno0uukG6iLLoJnif5Rz40KwaR3b/GnB6F+Ku
psDjBTT6fs2T5TYSdNZnkd6wYJNTKcx5d1r0UgeOYABQWvhB4y8A+QMlujkBjnNGoEVW+LAmNgWm
2UQl/th6991ZmrJe8oRjkRSTzcMnSF4SVRaf3f5rYrE6u7HeZuKp4kIngVYv5A8UYU6MUlrYGDY4
U5Pf3PuX4loO4IpxajAQ4xPX0kIcnqfblBWB9syoQ2eaGzO7k+EXbhSeFgKy6op5SlHICGqY2ZBm
Z02MuHIw6geYYrwy9jivq/gtPNlmgsB+flE8/J9wqajVIgS3gIMdwejG73obUiFYpHjEsvJ0r1ig
7aTXglU//hlR6aC5TOtuj3iBlQ1PunBT+WW7ZrhOk/ALGvubWZA1AEPyBn5Y0NTVwAsn+rCOmqRt
Nricd7zpTggYlIhG2VZAyZmX9h95TA5cgmVGZeAn9qG/IUrdtCyL9hY/nY9h1Fn7LYp5soYxugti
+R0JDo6fAeLiHdAthMwjq+N+gPnfesg69t2Za12mjWVKyUu508qYIOQE0fSNBEB6vJbNnE6lpCQx
2cuWI3rYWtSrqFhT9r15O6Y/gKLExg1yCC9L0G13Cl6xCUT+9J2DCq3QVoDghmf/pdq0Oc5+ZzUW
URsjyne/3t6YSd//16mKS9KhnVsDbp/ykP4Dgx+iZ0ta1PsNFrdMU3yJIjqE4GCmyIEahTt8w+WW
9UdNHayyVt+bWTa1h5DtLdjPqNY1tyGe2Mo0rjDYfQpl8hsDOYdshb1aqzh8XU8YziQTSwjsUx/f
i/bQNoLqf1uDykP+lW5BrlKK5qRfzma/9c6/kuWjEHXJCu6xfokgmVnQkjhfXdv7U+V5AzwhiQdM
lnjzRCi4FAXaGV0+IdYaf1J2iH1CGcnN2+DVB7AnHuHt8L+yx+UXQOAqbHFLh7tkVVTW0cDdr6d8
CbxNVKnkpxRN1wkVrNqC9FYmhfCpVz+QPAdjm4r9YGYq3KB9zwQTjNwL+b/s66U+ZOdAoNy+Qu88
woxjdYLa2QoI1MdI3Wjmt2DO2hJhEOmg2DmwSpfv3jvz87y8HzWgQqvFO4ikrKjG2EQoz6XGI6AK
6Kl24EmC1eUIKl38dD6VvoVwa55CPokPeh1fs3gvxL8vRrEhEIv/BEwUkoRyCaRGQIgJ6VPk2Fqs
Y0q6tIgMT1aG/nNnWskpJA++UgwsexhptD/Ro3o+/XSzxfNHtqkPsz7WvWEArWf+fSW49B7dxDEm
3pgkInXI7rZ758wNRUjxCGwczZY1wnxqOZV7qxqQFgkWExAHyi6FPiqRD7RfG6fbIKXSd/AORHxQ
qbPKe1nHezEvEn1SVDCwspzAKYDhX/SKkY+yvuOAqzgfiK46P/3ZPNVFOoaAj0+0AXkpwMtIa++W
sd2HJ0Czz8eeAnAozRgGD7DztDp7JaqV+mVcWfuVCjc6dT4Bchc+VI9GIoKPURfDkp1O41naOySy
CjSbsNx5D7HmMX2qZWDrPBxVhjQHvCnaNRqi1MK9B4gYHfqTvR2zZuQ7QPsD+BgqeUT91eS5S9++
raezbmuA5lTjsfvwjyW1ziSOnCDO9uVE2zg/AsjwZVzkouxZf3iOwI7PCfkgk+ZFaCU1C6Z3ecz+
Z8UGfpg0pIRRT7g3Tv7avCGhUl1yfr5jxWoyNfRatRiriZwEctp3AeMEi2t7P02MuSaMO0LNXASw
dKaDC7EijHNuJAo7L+cGtawD8x6z1bVTfjVXcMuzEYOVMZ7QyyJeLyUY86i3cb5UTgFpr59+RH3X
KhvMN14XLuKM7/37jVefIPz6siMXjsIxEg9GIdEduSXbNjs4yj9rB9cR2eQP3hv+4VDOrLEXPUHu
9EPGjIHp0Djuh52yFSG39kJhYzcrsggDDlZYAmta1h/RSYB0gvzEpcjJjcgSt26kpYVIvYbLWFld
B4oqViiUF7Ij5J/a2fYZZ8c4EsHqVrSh3M6TOdvCh1VaCceaO2Nf+EwiPQdzq6cmIHHpMiLJWBUO
tOa0TxX1TFgEUZQvvCRchC6wxvYOG2j5KnCeT8LosJ39eFzeSL724QKAPXedrQKccaPRDfPpxcsf
VT07/FNO+Y6K94Xw5LuvO2OqKN2ZULObKKLz+bgQ8ausFZtPCuC565hw1/dgRTC4I7XfknHbVtLK
Aa2N0Qb/XTC3xMf5J2XR9XXGmuJ34PssgPuizuh34k8xmMk2t9unYUsDaie0hDPnIzcGy7ae7hZO
VUDsRuMJUaNQyiVMlJe6Qwa+JR4qKXBzXk5yDQLoP+lOSOsp/PSojqP14xj6rZgDdf0xcZOdoSvJ
6x8cZIOVQ/0sbDnYQX6mSq4LAvBYSx6w+ia7xWZji+uHcQcXhM7UVUo/2Vd0GgoTUbARc9xRQ7nz
Roj9unEl/mdwt1RWg/nHaFtK5/BIOW3WvMvUw7LDs34SLRRHF31k/WSb5ne4nWL4Sf/ootWgjIP2
9zrJg/GgKMWH4Ui35wa8H+cH4DLtj0kWF/cmBdu47xm9IT3vV320lNnrWV0Te/FioBiNX5y/b+Uh
ROWHr1l33fcMI/zbEnPDBy1TIR2jXZNc540g+MocGjDtlseK9x0yE10NhDN6vtS1IabjrN0/JvKR
neNr358YoG3b0H9EPbJ2s/8qfPMSw6Hd4/LSLIaTyKYH3RcwwDgqO5r4yubIJrVFoBGzG4zmXpn7
0cogmTwcmf1aYO/Z4YtcM+qnjDiMats9/8pOR4m4TTrnoaRI++BuLkDNfZ8ENzbo9Z/pCgD9oc1v
dxQq1AGEuuwJhHVUXlrTAaX3ZmGb7PELplS+eOwktWDdNTe6w+nt8LXc6vdLsKcgBJqXpXkgIBCH
UqgLPO0h+z+f8GxAw1LXnpzr9horsae7GwDeMl2Tz93PM//UFKMpbUqYyxk6Uw3c/vJVuyFZXwou
3GycmJT8WmPOe8As4xvmXtrhqhDjKCZvl0MUBCvBLoZH31ErJtjnkiUAVufQfM1RQCz6JmfhoMS6
WuZ6Hqu44kwUeYQrs/U4KTXS9xYghnXEI/MrJyIxCfYt9AgvATu9ddcEvka26KfSn+spHXVXgKh2
J2gEKEqKyspVBH4xfNv4Qpe1y+ZBZLW0y0BCnchzhfzo69PscdaFKiiCgxPWR5FPhZJZd3MqzJYR
Di4dyxIeO8YQ/LNx05YmqmSePyIK+fxrKh/AGl0yZ/vwhhtbOpwECJJ7kTxn6zPfYVkH0v21hpT9
eprXfuw2Z7D/UHPuPSTxsg7QlUyOBOlhmYv+2ptxdxHTAzOmG+NTieGeLc7sAZoKzL0/r+5K1gn/
d9W/w4oJoTDxoBtsBv6QoP/MvIWIch6D7zV2qZSO7w8DQqD8spnPJrGPK/RlNEwkCFyjOR3WArlg
O75FnIF29SqSSO1Sa1at6CUzUc9RVEG7bql6MnbhqRwhQxOef4LhyQH6faC0GmqXYm4kaESarupP
HooOBtfL6UzbDd2gvluNWv4L2jmECFu4AkZB1lcrDzOmffuF5TqmGffq6TL+0HMGs2OyDomf154F
gTivLs5XUsRlnqvYZhkWVpMsk6U7c1Em3qqLlPB8Ek6K2HT/bF2PMYL4b2wV7hmQXbvIsuMTE8pH
U9hTJfRvQ4BV/ZfHXYAZLcxtaO0G/r5yFZB7W7Rq9WMPuE2y+4yysI/vUBGGU9QSqVS8mY0aTq9p
F8Gh60K+hVYPwqzoRvGMrhXJtLJC6fNLhtqm28XgUF3BFSWUULLNL6weRXAuAf36DL6/R2Fbt2pf
UKPapsaHV82Ni32n2gRkjuqpo4zxOUhFBGuBZGpRXf3VV8fL5opwgk4QU5jJEcHw/z7WZWBYHrHQ
P66Vx8r+n7lV17VGxFceO6ey0ufnA+EuR3gXzJTr6+3WQG1X/xRf10AOItFKjC8p9hpACv74Ueh4
7MiCNKEjOcXGpArezVXDqg9asQtQSUgjoyBPD7ITnu2wT/lnZS+ux4nJULCA7/dCzCCTQFgfYThA
ro+bAJNKdXkoApw+B4ZaeueKbeQFQn120z1/tI+n3lfsMUm1HVGJRngevN8TgCW3kB5PeJNhMAHX
9ZkMDdv7YLbmnUMQRrV8gjvc9y8nP7GBosAUnhUaCuPdugBmxtQk9QOse28hRph8q4VCRiYnntbY
LTWRtn4ueE7ZVImjWsu2MVdDNiDVY6EYnhUCz8ZEa/Ak8/ZrGQUxMBE1hQLwhg8TBdZ3qNsEEW/U
7ReXiKBISJlM4lDFBOYgQS3p8k3AK/pVcase3u3xm5AWJ7qC1mO0Td5cTkKIN0TTBcZ4cbSwGpAF
GJr0wyIIGAAaFIv9Fz6x1ROpT3lyUach+IcyQ7l1+gdpiZL9AqWAEeG0Vvz1a0TZl9bOjkD8cGpO
YghYbV9wn92IkzREsbjHfI/p8EP47arxRPVWqvkoaYzVIn5Vv7B6vzWt6uNOhoQhLpbCLadk5XxN
sqmkyiB3YaIqh3xkCHYp0kNtxZTlyqHfrYvTgnQ6NW4u8jNEZB+gSRfiFW5JSwAEBkjClcqQubVu
6Qa1TcfZ0W8yT6UQftTiCwA6AV+4OqIM3lQef7jh3EXUzMFFyXxGgri2EUKtPL5Apm5ktbYy83XP
1Yn5meCL+UV5JuwCtDatHqw2IrREqnV5YnZTuXDss+Dpfu/c/xBF9abF9hXfz3o3+maaMpngMeDp
jxh8r5F3cQr5wtWg5I4og886f7kxv+NZn4ck0wSAf7oozARqIUNwEv7geL77z+bKhw/tv6mWxGiF
Pd0OyEfw5/YRGPkeUeHaVW/0To1P5a7RJryBH2XKObt9WflgMhr9AfReoL8KFAZjxR0C33EOZ33n
iVoIht+hEE4Cv7lsQiGaHSrHKULIRCOCGp9HbZ+xooELTr7Q3LSGJGYqTp77Btff3UCEHFzcwrcA
InLwO091l4nn1WXSNwov/6S0Zru7n+u2Py8qtoDO0jwgooBFF+JMTISBltjOM0ivFkePdHFrDDVV
pPEJTDbEdqFkbVBQ/3/KK1/VVpEqpwDrLq4FkriYVeyYRiaX4x/VEu9HWqlSldLQJIJPzSNElMQl
7zLHEE5dfs4uHqspOcPLj7QefHtKWCv0U2QKd9YgXhj6DCMrhj+oR0mEZhwTb7fGxWfABvDNiXPZ
6VR8WhYC7JbfjnT8fX7Tz1ev4zyM/lXGQRGwNr6scz603i39TDvrD1or8m/Rhh9V6PmlPArm4nzw
vj87/zIjMA07Gha2aQVmvXUGsCafU2dBffh/C6PmWODFA92CJNibdUq5xaZfiDYhueXe5YqXOKwM
3goHx0quhNO++OY90XNrfRcYCn5eU0syyA0HUghqf1yR+PGuVD6mAeR/NGlFZQAlkK+cktnZK6nX
swoK+P2j/cqrLuUvIFjFudDR+rgbUS31bDtnSvExB82G9kuxxUR80p4dwiCm0L7EkhyhqyIMODQd
RNEFFu9dPmnKhD1D4JijdlChMisXf0ebDqxK5wo9P4FUR/FFIdba/PtsJ2NAaq5mlc7hq1SYdZIr
R+I4oECgLZ2rSfHSF05IkOF1Gx4LkSlHC0jRyWGlTKorPuUR4TynRYWz0twricCqpOlRo7ohRMiE
Cn+IobwctR5WBI69lb10Eq9loAxU21RqLe1P3rRP0jZv3lYyN2Ie9mvj6g3SkVNfv9kJkyRhmZEH
zbyaRSJjusA7q0Elbt7XqwUyRrMEx8rfqOrNQCXiFoGP1w4iV2EBsTpDL/r+G3P/wg5NHGLEXb7m
w7t79aDUbmgKC7rJvetKYyWjuGHqD1SuYW/o660T9eLYR/D80ewcdaUWPYv09/BB5YF2W62nGrE3
9L9TQfzCqUe79YflCnuIxTDodUSDT2YgLeNPlcXJ4mxQW2Vr9GlHkB0QqgW1K8RkJ/4rUqr1qENL
41c05vMUQhKz86mOOZQz/X+0U/t/dnqH2ZzJuuXjjU6/KU24p5nnvspdv+kHaisv4ya2kC/nkW5d
RazLjg4vQFHUukceSGsndus9u81bK+L4Q58LGaUUnIvdyId98vor+6/xCLeyKH8yy4XDm9Krmv1V
mgUfHmpBGkSQQ1ltVEX7eS5Z5VovBTUl222zon/0S1nPJgv0dMUDlJS/6849ZGQqOLrnuy1QTxuZ
WNeMaExY7WyGvuq2Mbi8937F/6WR0nX7jUrZbMuimnwpwr+cTvJeTSr5dD64C4ZYfF3rj5ZDmDkg
Z3KFbSu/mg/j7jEBbe8lsSol/pBsBz6k5aaRC46aiHYNRs4CSuA4e8737ho3EIJqb7XqEYzMVLot
fjeUmZE7CkiQfridjPm8yKsy1md6QSsmOF2fiROIrD58fqZFaPeY92ERdNoyoLtgAinxV03KZ0Z+
ddnePt3b97Du4MPyJU3bNpjo3WlwFBP3FqWc4drjUeL7mLNOgzstEuj9mn+RDGUfnD+RtR5fuXHi
EuAqTNDxUDOn8hfW0aYhNArusgIbcM+J/21FQ8u65qezHNQdjX+JQokJXNLqjhI9hghOytrhGtTj
xbn14f4SVf0tDIzb3Vbrnp0u2N/ITmJ29pm4+qczEwnTzqx+n4SaAi95XPLbq/q+bK5JSX1Sj0A2
X2k+O1jCff0Qstku0rrimErFSzego9P7eTVycROnGwM/BwSz+XkCn9oGsuEzM1c5ecphLhrlgRBP
gLjUXjkYMp+Q+11GfeHKSJ4cFp2i71FOrFYX6+Zy9Cr027iv66cDKyndlJu4uzjSiBNActJ+7OdK
sMKm57CvSAhj8EFqfoZwpErOd053BkKK8MyTkxDXBbRIfkoF8rWy1e9x2zhLA+INyWHSf4QsLj2P
NEieHsvpwaNAldnXrF0O8wZpukIbRFrhbDhS5U9XD8ucmqRM0RPVquJT0bPt1PPNW7j31KswVhlP
kBUcukINQ050vahd6cRt2N6cVfkUu9r98ue0r7Q0YQdn7OQy4Sg8guU8Zzq9gNIC00FjD/RBpNPo
iG41nqIVuSpSjrhxCFinCc9LKEMeKn98qh3kPCqeUCSS70pOeEZHT7CfoXLgr68yFWmM4+CQSyt5
XA0nIDfCLKhvkYvHC5U7e16x6BC48QS2efnEftZes4QkIFY3/DyD0atjSy0kERwNDj9+daQqFbem
uC1kkUY2DAY1Kp1Pscfi0+aFnnDRk3Inv/IXOrdlPUGZps7fqCdJgTZB+bSiiRbrPn2AJfASFdJQ
JtxB5ZOBlCA4WMWY60eaTjfJZt7UTWDMzYbqOHwS6Mu9WkpQbkH8pU1kQWXryMq+FHaj6GuRuMCU
blizbY+Im3B0HjH4RAbp/g0CzDePT5tng5BNuKCs6Az6otFAPTOb5xDqKCWrnCVAKp3QpelfvR5o
zE8UKihahureHZ5rMw9aEH5KEt+C9V8MV2XoCeVnkDjxJI2z6t51+VzokKV4SXLhczWQj+k5EHFb
KM0If4pXl2RurP34WHB1T2HA6WEt3tFC9FcDpoQNaIvEZlNvJDSapY9Qo8SVlaYIdPxgehzdHDp+
r/UaZGtwI6xYKX3iwPr9v+wUYusJLihX6Tj9gbONHFZJwP0ynJidYY2DucHyAZDBLp+G3ohS/WnF
zTrtDTCWCnf0KaEuTBf8ZA5TMWvMRRSV3PnnAeRvyjZwyKjG9Ot6ddFqfY8tZMV162u0Aim2z5+X
4tAsMTz2FYZLgq34AlRejwXquHkQ4eOw5nKmwKixdAqZbc2nXu0DkeLUxnEPG3ighTx/8g9Cw1q7
CbyqsPDtpZClnrtXnpebvP3X9xGs6uBiAgSqcFIk5ROWN+JSnyzqd6NTLG2Q7LZN9luiHEb8veKe
sxM5oyg68Xo6y65AEMLCiNIgtvBu+wqd9bmRdnjWv2yiIx25KfFJxu/DV0vG1tL1GZHHXy/oQ1ym
+INn1kg+0QDd+Lx9dWfMq6rOO1F+MbLE86UE2RpV6Lp0c47j0+Zm2x6eCJRMoFhzlcFb732uenyK
TrBDrC+0K3Liz5bLQ+bP5VTNmNy81qwjkt/0p8aGcHxWksmqWoab8Zq2JA+CcOan4vRNrJ2XBgAc
io0GyGWms+/hpynF4Io5Sk++Y9ff0SRErzm2hPuX+5UpF9i4XTePOgQou4uohlZEwqE/r8xotEsS
CrKYKWyr1Nj4jgKMLl21kj1SdikN2Z/UEIAqSz9FqtvLt8U6m39jXIaQLaZga4Zobn8cbkcs2Zrm
qygn8yq9wzRqWcvpvgGRCLesV5s0fE2lQgjilePKnyjhG1IRFXISNJiqlA7tuP9rhGLC2lYV10+2
2Uu/EgnDDdcrTQlzVuqUBsufMt7gqiKvPhSA79OAA7wN/Oy3Z7rcUUR0WbEnoHDoWQKLSOHQKXqc
u7CWlCMbLsM7QSY7YTuTjzjp4jErlr94J7F/p5sIVygdskJbTYJdOduvbkxnHbmBynY6eK/OgQFw
5f1gTU/D7v7RL3vMJh6SV7QaM6rZJSPO+Jl8Xk8Iw+oeagSfbnec7+sVau67ONOM8K8MMxPmKLSS
Qz6NLiExKCmLPmq6z6vYqbH0mp3BmuAuRTNaNTuf4Vop8AYYTFAkipkHQlkeNeLcHl6HZquh+xm6
uBJCKLCShQ1M5FdpS66+vZlTC2VmXUrCY53ohMNTyqibfvweoI7dJnW8AYN664PF3c0PNfYhRq/g
ptO/VjPIM2nSJONAuPQJCqRjVtjaudf9E7Zl1034S9cLHBJ53t1vEiy0sZGR5b0Ii9qFmuLRwLYS
TtLtwmIopxbZkiwVd536Ufpe0Cj7NPUWvbmnVc4jSjE+YyBj06NUGQfCiia4LvnNLLiNxoeHHSoU
jtwrBRo5UPNyIGm/MFPDTm94f5mk4K+puMgcRPj8zOawp9va7wgQSTNDbCAW6eAHYHk7xphWEgv4
357KrQ2OsV8iJcw3yFsvrhWHDdxgQFaKm/8dYA0wJW/OKswlqYekgXPCAOW9a31C6kKR7+xb8RzL
BO/mNuDnjr7xYc7kAmsOJm7u9hiFxhOhQDKkR37K3vw3mRjmuWsCuCkU+wbSE+fDNPBWXEap7vuT
6qj3uto78DRxCFZU+CD8ddnFSg62dPe55Cu4PLasBh7vtthco55w3lIsT+Q8weEA6fMJC1BWQ+5C
iBtbk8J+NMHyHz6kqEE391mFZrWy5EDxIQAVckYMvvawH7QYys+fxUJ/pyC6Ivj5S4/BL61FAwHm
XyujZE7h37b3avlW2xzbJ3aZtKHJQXvooNCuT9cPclAfqdnil9VEMyqmJH3Fnmgp7FLtXyIL5GOO
i5R5WeSIty/ct7/16RuLKMMDF7k5a/UfpIaKwQLW6ulTOS5xZt8PKW/GmnwkS8wsPvs2Ux6SMtXK
HTl10opcx0PTIvdKNYEOag4x7SXX+vF4vV5JWc+tdk267spYmxh8IZNtzXgTqN2xj3s8HrDvPsPn
5zrv/mJn/sWg2EsNtaYZdAPFT7hXwN7EO+ZU3wllU8IovW1hzpB6o7/pXQFDHvBpmZOg2dfkST02
55byLv8JIuTruv2OiXw76JrfbT7pzEVgozY6ILi77q3ETYOryTrxQ1CgQEozxQZWS5prn8FLb0pI
RhRu46gOinR0ZL3qZfOFq98p76/TVM55yBrhEOY2wTWxcv6FVjESih07l57afztX5Cy9qHT74Rge
DF8VJgCKDvCRrJqsraXVDPIe41kJjhdf/Av6ngXvAPT8HbPlbuho2im+Laz32pn30TmB+OFWWopO
WjOUEtMtMFxOKtUaXKcnJaOITRoRu2bTaOc0quYtishG/lnB7u7ndhAgNPos26clvPSFkJwCRbOz
IK3wxC0oxL8Kc5IPa2viYfUfXqthx8O9ar8yWOJHz65XA4zT2aW6I8iEFB0ircfoKVvLtgsWIgYH
/agYD5HNXvz71sJi9N8AnrWnuPcjrTcsR5oQU+uhmYetAQ8GhNhwHrdZaVZglmjlcApfosc32hc/
BOBQUq1hqhYKmjTiMhGYYGEqmuVnhCGwQ3wHJGZiT7D9ECCGqbg3oVeF4dnZ8WI/xhmw/2ZzDf+w
1o/bW0DffS7vnWGUtaL/0OmHZfo/pDTAuZkULe+LFXtWJRY0KllZjUYbub9jR7G7KyfFCGwrKcPh
cZ/I9LZY0ValsKN7C0FF5s9ARC/6TPm+VSd6Ahhl9XDWUkW+994Wto/atxvK2nEzDw7ZnXVVW++a
Rve4J22tk4tGHtxZpX0gbSt8YE8AwX+hjsqdIi8EeFfQJD4b3ET80wK+wl3sC3aMD6v811NJxDe8
ldSeGnTom+RYlDWdLqOEKgvnzPBwyNV5i6LB2Qe4YqmU8BbqtKLu/uAhGtJaJ1TNCsDL1C8joHfP
Hp6hWmWslzD55FT4wx19rtklmuCgGrc2ejjgNsGNr/i9vfo8PzbcnRf1e4YIPr7+KRTONTBl+Xka
EsMq71izBwIU25HT7lv6ovVq6spkNb9m9lvcs/jsW66oob6U94S0EYZQ+NHLc7c0qaVkdPIgWTHH
/zSWokWj4wtxY2i3Y+CRrAoH8XpOx4fkswXxQTIKuvtH0E+e4W794tBqVnwxoFW7j8J+ps3cc501
44+E4qCGPZw5/JdROZlqbQr1R04Az6TdcZdKXpkW4/1uYlRI7s65ZAAWuJoxW4GO0PIZkRUTgmue
4gQcBPNgUvkw+oVTjFUBTbSq35p9gUK+MfKm40xUlhB71rm9R54LYZKFPsymyBcmnaxc2w4kqGXn
TNf6lzrqxJ/Ix+ELl1DezUs8v53TFTqZ8+ezac+8AuLLoXnusTQJVxo5SHotDm2LIoQUIMd3Fqio
VH+vAOcaNWtATR9h37xap7/hQ6D9e8DQXmRGFn1QW2W969swN5TSZNegdlCKFBabTR0pDMZBeto0
sAsN/1e/EiXanmjGKv4Jvtc7sUmV6Kz2BjQNXIRfZ5GoNyRZDZJ1CQFfotOKK2ag7VmXiEsswr6W
m5j2t+A8WgDOYEEc1gAnTLy81YSnTS6CXJ222ZS8n7pvOCQeQPQwAZdpGvG1d+g9ktntx7o8l/6g
tCaYkXjMi9oNsmIeMgv0/lXMyOchMlmcm2hUAFGm3QxSoSJmzvqNOtSSajjkQfh2l1lElB7i76LY
Fk+c1jQybL7BqcQx4eCfRQeBUM6DWXE/OsxV3Ndzt+9tPlwXqMN48Y3Q7LuZr3wMwDNgbsEJ8ddZ
1nkpFthJXjchJSOQuz9jI7VxxQG9P0idfwNiMqSqWxu7jYUXCkgXdfNrzTaHbCxZYpxOhRKVSZ1e
kH4ASKhkwRm3nykb7nOwhmHii7WaPQY+jHTFdiYGEv+LgDmK7MSrmFwInZufhPF1v+g4mJuqHLB6
HVzftAp0pO80uc35vvfaO4RkkBjg2mDU69yf8rLA9xeIi9nBOoZoO10HVoC+ZaYJn3ayB9ImPxhh
dCwScu7F1Djzt4hn6mB5D0BEfqUYg/4FrJde5UGNR8eobJuz6C7PBAltNzOqhipLNcAKZ+ui48yc
fVFJXjV/yo/+NbEZHYG75fXXO/1tIzFf2WTNANCDvrpP5cR7qJXhrJI5rxIP4LC9EC4iHoV+ecjY
4aJ6F2fkAugAOyitBmD5o5qXQWr1tDuKHgPUOsBao8RldC1RKTmjnNzIGyPC4iuRuFeVd73Chd/G
IIp0PFLLw7KV/YEWuugLa/Ylm1BHCKBIQxGxiU42I2lAvHjCVJVS+KAjhmBzRv3HnuqiP3PrrKlX
/1EZ8Ov8pODTKJZGG3P0FokUaxwmEy6qxKV9rdtl/koMX4bPoMznllBO8BNjBDGiS22S8G1PLrIo
MC3Ow/gU6CfduL3t7q4NtOdDBh0DeWyNZOdAkk+tO2WjEmiwyOHk7tIYtHPC0PMowispaYVg9ZFp
kptZcXBFPYpwq+VbUeeWtt27nMa0MWPmEo7KO6yGQzvIq8/DwEIso5Z6BXYTWmzSn/r3cJHrLN0L
pFzScif9hOr5WzyeobyXIPyex3HcXixpPP6WN3XHQe7t5n8Os79x8U5TiuF4pw7PLDlHp3AbbdSV
fU1FkF7e3JJi7pQXFUJJ3lfre/vhGBJdrcEbbw9Ygkqa2KoU7N9Z2u38IALzo5wv4gHdcIw08GbL
tn6CghYQT0PDcBFz5nm+wT0Vw9hgBJmV0YN4/pqT5zIAp7BTGNcFIaIuZRTH7rfl8wUyAa4oelUn
NIWNuYIPPBdU2SjppGCNWj/YmgdsaUE35LkiGhiaJhRuw5inchryrCxV9rMr0mMKymB6BBf2gjYB
67ecD+kDkOP6uEz52eFkSPOsGcwiAAlWbkxFlyCDbrjQbeLgSZKwJPgNvxpS4bGxKmPcVzeubgdg
49JVrX0NuJRoOvg2yJjxF41uWjx/gqAK0OP4tW9s2vkVazywBbXUReWgcoMVllMXR7P7dmRgxu34
xg5ERm9AFZhaxuvThafTg8YH2zM2pCfgJ7IE7ZotvQNf6f5bqu6cG5+KNL1E7qPnnffC7nggvrlY
+4jQ38STlQ79s5vCC9SCKYbx4T244GujWZPTnUYkwFv/s0z1pEKRxEoldLH7hWLFeM1o8Q8tn6Tm
rfnl69ObKG+Ke10BfL1kwByWnGwXEVtOiQfIL0e6REtkPmMrOy9zyUDYaaxjYdVDI8vpIgptFh06
KYi1XVc9lFYUA53RRsoOd/6kyMMYLe0rX3YbNzxxKkkg+vGROb3Y3Zdu+wcwL4DhsJ88TF3hn4ze
02VOf8dLLORwmeUaPKpg2X24tHqfCIFHsZPWbobKPIq9A4OU0ZgjjENaRlPTt2mA7gQEAxq7Emfc
uDGIElFe4XGIrwnRR8x+5jYJbDj0dJ9VGJYo0m1s3MpBrEF6nFl7QAmBKa0WYICEZBnrwLeMB578
aEfQd9/fLQzyfXbVoAHhjSJZlackMc6FyPjbN7kO2OzGioSZDW1FIDTT9N3FOXWesae6EfVwcqki
HX5llPnaV5w1h9TMTfOHfb0MivjDJFuodQZfu4bwAx76ZJfHr2GgckRbWBf0pE+DvztjYCUX6bhn
1vIE0paB2tR9EuLwqV6cwuHfsigQJKeT2t8JEmdksKJxoGNzpZuqHl6jDG9m8TYqWj3Q2jDIWkNX
+YWRsw8H5U76uxDsaGSvHaXS+K810yCHLFlJlUmieQhpN5xO8CdVp3Z4Z1mC8Fb1Tx56ORcgt+V9
8i8OmMBUyhny8TQIh6/RqwNLMygYb5wO3aC0byf02KY1VOFY1DgWbx4m2tkMP2VXou5msihEmMLB
nYV3sJvXka57VNqdGM6NeLXZzyZ1u4a6KQJ5hgDu1wDRXyS0MNS09mt07QFXZLf5eA+2FrndoOlZ
mDUJs9k0+0SNHNsBA7Gtu6mjzq1FQFwJSE0znQJmgG5W45IpFfwXMBSobLcQ1pCN5TIv0gUy8jLw
qN+VxOthvaVWUS9AX/Jd5UrDqAYF2awPEwQck3UcDInWwzczj8QoQZyTMXEY8tz/LY5nbV5uZUKd
72Zjp54Mi9mBm8TkgI/Pvvmf2zlhazOfHip9FSvkSxHyv62RZYWG9QilJLAo/9LWz83rVOwM0/Uc
Yxou3mKMIg8HsjTyqoVlYwYPGoYLH+fZmHpuGJQE4VJSBjEHFFc6ncDa6BryB0fkEZ8USqg595gV
mdr46ERVQKuS30RMTemxmeEnkaIdMz9b8y6YnrS+eo2TPvtWVC8XmqmpRn7dcblnUWU9xGAb+NHv
P906U25/TzApcTnn4aCbCHxwnsNf43oIOtZy5HpQ9WDr83/Pgc1BklUInBgGAP614cDzpII6n30P
8869nLturBCZLVDEGw00s2LLxc8eeV4bq2ps+VJE4InKhDAPzlOKO3nQWtufPw5DlBX6QtFdXmpu
ushrrbmin8jr1lhatv5ccZ5xmPg9C0cne8tMSSFGnRan0qeL3N/Q+g7NuJ5oRdC+5SRJoGTPlXac
y+UY4iYW86SM/etp/AbjCqo+juPIEgxVrMb8voudwPcHzuAqZwkIf8PJJi0UjnwVIcpIKtsb5BFx
LF4zAPi3mzx4WOsLzQ7sxo337AFNvDfyYyhW05PSypSOe2o2f/aiu/CH5Vd9NG/gwa98Vt7CbCl/
VxD9hqIUubvM93AQcjUbc2+5mxDEY9uUJ+vTx3Wd30xU8OjWZIgG+rHHmGwDYSkvxH5o+TKRuv5M
hgO6sAIafV744+OMZDn1Y7S55X51B4MNoKr9hcE382JpbnXrkkSEUXVnUWvLsd9hqa1MgTBo3hu6
AxOiBokzXEQKburlIQ5tgqmfG38/ZCj4oLVO+CKXmv778l8kbuq682kW52MRDo+kW1HSWkZC7ou6
7QRoA71r0jRBb4GQD2iHBOBwgM92VXPJkFrhYHPafAzD9Ohl/r+CSEzRGmEFpmV+3jrwrnT8cla/
ic4xfaq30gVW9+Mt27K+8xmqJWTa5gMi0v3LIDQDMIDbBP8uBxIBwIPFiX6LqtGpjHANL9jyhV+0
R3jDh0tZ06idMko+FniXqi22t/vs/ijCbewOFBUZm6sxxTo1+o55OO5bCSV813TRPN//BUkL6tXL
ntd/yBVT1eZXCTKHB/NxMlAZYYY/4V3DQDLoMjIGKEUUtyfZywaelZJYm9Fdht+EWhi8kUkmQBEk
Q7+BtUPgWDRuz/zC6eBeCxx6kMw4Dt5F6kQJneLkBQXwN6wGoLJd5JR0cY8HxbUk4xH+4ffzG18D
EBXjxv+P5YO10moUiProwXkWQmochVFy90ltB3Hv+5Z5AGT9ycV9BU8hmnwa0aatSvGG+lm0lzlG
L+AG3XiW+0vIiYBcc6N5E4ZIkTfGPUDTM76Q3OFbmU4xXXn2IHXhHXICVxdRG08ggcT0bRs115RK
t4Ar+VdRVTQJqG4E1NF427b0LfVyhNxGerPLuZPBGsd4syzA6EULgeexzlv/882l6lFcsvVDcbHR
RdH4zawtlQKliaUFbuohdO70oxvsH7e/NP4qJCAoAoWFoy2Si+6PlYKFGVkQVbu8qKeJjU8BFBPF
vc7msDwTAjCdVEwzpQkFhYm8Y5OeNRYsi5Qq2irG0wNmPXIb18T14lUsZdaI3JNREeZSvuzYnzPS
J6TVRK3eIHXSfOpjP+jIZwIvkGMmobNLRhFvj1B+VKFPCLaak1uhjG6i1yGvjMYCLobsh2/JfqS2
Ryv3jQw6iRTBQxSN54l3Gy9j9Bz0F251l+dDjPmwLuoWbxPXLatGMxgavZzr9nCJNhfm75P68OsS
79jLOGI1NVvqLMD3SMwsekEtDXMZ+18bJHBnHD64PuhMgdh37jIkIYduThrY+sDNDIDfW4itOf1c
55HNDGlPdOVIskuwhqHMyCgndFpbvCxDjOGn5ffoT+bixqQg3rCWCeUxzN2YBxwKqx3Sok008xtS
EfsV+rH+dOJBQOSH4UWHGYwecm5deXFtoqDJyfRmWhskENCCFb2XZGq2ky+EuUttUgHR0+EbPsvm
oY6q/VAqDtvW9RrjcaP8csiY3D+a7HPTwFoLMCaeojRMeRPoegitSXyOogGAy/2EHzFVqEyzjDli
kIxx6NsCQKOfpeANrrSQOAZuOQ/B5dBZ1P+yzppw7H25WU0e34RCsa+505BY415/Ax/hUSzygQhB
O0nAElZdnxAkv3bNm/usB2aH6IJQdw35TqoUuK0fn1PJanTWXkHDBHvNtF91OjMXMbxfItv2GZok
NBa76chsvpa5aRqsd3P/Fe8QFZP+pVOpDKn+/Ilx+4hppkNIAtevlukLiUFs3SfJKUREW7zygEEo
LxowyigH3jl3gxDxC+Ae/zvSHC4nQSMYGJyVqO/UlKYCkd3lu4B5DlEQG6talw2ZuGG/LsDFB95s
solJhxxxfyc8pZFIx/lJiuGK1kZYNkFBl39fbGLCWAoKQhy5bKAPNoVi8pmoWhc5QMkXIyvuwT42
4TIzPrSgn7oFrnddvmO6fY6OVfyCRGH2MfKPLpFbc2/wb5mWIdY7P9C+cIhuf8pI5Q4q/vikvWKx
0RgHhPOAy8HXShr656oRsTTe3rugTJtr/3/EWmX4AHlba4BlfiBNRPoy+vdGXLSLZDFSMKDke07v
xEI5yHnlx/KT4y9tL7Uo2KlgxLvH2SqidFAyP5khIgTDNVVtJ0NuP4vl2YwvQlfWpVUFXz+PLt+w
uvOHaEOd3gcS3KAY0Pe9mMpUe9dDeONhlLB+KA07XVm+XW4S2h9+Ne7o4khNR3LVDAU6ZVdopKzy
UfQcIMi9KdnTIKIceDsCngiXDg3IoTiL10SJMA+x1TUheHFcIBjEXcjTzz1mJ/jcjE5C/G7MotuG
S/M3PlcraMJY8ExuQSlsGMFTWbzpANFjUAPFLaURe9SkZMj0SXmSm3N5iJDvSfqWjRnwQ1/tREqc
umvcDk2gpUN3HnNHHR24osg5j3Vb3ZoXWM0c9Aqd+ef6g+C0NFqXyjrCfuOFAxtHm/tq/7Uky61u
RDf6RVoXbxqmlMK1j6k3gBqrEefcWjVccsI5IDWnNCUSQ592ivUbflxKrXDu4KMEI7wQZFcWFmMh
W5MkrfHwU9OuzU09I8+xtbvLciEkDQ0GbSL7rdWvDUI5aJ86n5zCVx7uvW15nSlNBj8Z8dLc3xcY
gmNEirBpJmLq/G/E2GWb/r1kkuUuhG9ZdjdRcJDWk4qBizl9CvVHnZg33ZiHmnVJcuJTpJWRT2tW
oXTRN4LHwLwra4Uqff5JCqYqZ+Ddfovp+XITWuWWk3eCo83PdzMvBwc4xzYvAVhMmUJCeZ23jeq+
GBzQIvKASmvqgAylXAUZy8VaS4Qo4SfNqdMqr0k+ZWFj63yxX4IR3tE07IWTkDthCQosk75d+RZm
fs5BV2Ae+fyGEIJO7VruLcMAdjsvG6iTGGQ82b8o83NMPdKVQWLdp5wIgyrUBD2j/Cgq0tHMTJ42
PY6vsijsoGh6VWJKni5xw2RrOcr6bTMM6ASQXZuOpwblAZCsd49gTwfkWXMhvjVzZyzjMZvWjvKB
i+bUCa5b5qz9e4jqv+laiF9ljaBMSeC0BZB9gLzn9fORXvqJkpbKPEbNTD9ZYtgo87ULu4HDJROM
4lXz/YYeHr6A2VRcmOaknXpWyfqDSeu3og43OOzbQjcaXmzc27mU12AHiLVB29hImzS26Ne+yIFq
5nyN5N0lHvxJ/wSmp9ZWLNKiZ4SlBGiDSHotPlgtAr6XxYpVKOGYHFlMEiZ1UH5WF6fW/3dvp5mw
+ScXJvYY+FFCYe3lJclx8akZWn+bcJZ7uu4cQy7bfYt5ysXaOcDJl5BjK7fSlifV88P/sdgzAfFo
hw3Fuc7Zv2UNgMkUSB/sl7XkYLHN2UJ89R6VzBLPd8Ivgs9JClR5e5bZEiZyK3B0vPBLKhMq8TsL
XDCLYJQR7ljQS5at7+AsDjOd7HjE3m6akHYgXQaDB0Qts+HvguAeznqkYgGXpVtSIIjpwbT6HasY
jV0PutufQvbWNoUJmqPVXXKjXhRzJKJnatCs9Kn3zZiJzBAwdAOA3vHZ4yxv5yqCVAWcr+nvDLTj
lFcXgDWH1BtrXoIrFahPCd1KCJLRpTuat+C408z0G2qvlyHBtd55qZf3dYmRyUtEpBC8Zptsw0tL
AIFVwYgl1yDFVZ0g4uu8EQ4mhS30piucpRvP3dxzYr8F1DU3FJ/3Ba/0mdkHDsJ/0mso0JOI8GiJ
RoFQOMFj6/CQS2UfSrRuJVLVGyihiWWS2kBQjJiQ5+7WFLJnqMZ+syMLax310soUaOMypsE6d4Pj
H/Im5xxUW3DIVW/5QpBwXqqPVJW7fCrnm2sJ8yL+kcXImCHGcwzQAvP7iIlzB0KtFqJn2BPKjcND
1OFsx/p9J81uLJN+1GuYU3MFc2mdF+ULAJ10mTrc3hy0I2YBoQz/GT1Wvr7bzZ6YnGKgcd1GJdi5
EePkG25t0G2m0ZB7SHy7TiBDZ1T9VR1+fwnPeIa1mtHYV/Gfe3odVR2oq4dmWkR8b3htPUiVfcYj
fofiuxjBstEl/uGdZX0N4Ae0xH7rxqOQUEXgjUuh0j8DGaHbAkIn6Fd14rFijBbnTi426r19fsTb
0c+WgVDFO8zVPvu/AZutjCpkNXqjYRoxNe8MYTQeQYFBnjPRX6akfrLwSfjJCQ2cU1Vxxhoh6y8k
tkg7LWvnJVCW6/kt4PLvcIWsE4dNP5edlryU+MaF2Z/XbqTqYiV9Q+D8gmKEeuRMlniFAD/16T7H
tpr0vTbmm7syYUEx7dPS8dERSxpfyTc3ZgFIeZm7joqDL/PqeVyjAyImATptS+Qwa2+cYWtK6XKP
Scz5f0mO0+V6hq3bca58BpvslqdVu0kY9UskMACM8c1M8jagTMI6Z/INSmRgy4b98sGDE98IawG2
o1EDSjin1afTVcHL6T81SO1c3QGugJ+qA6lsAInYGGeOx3F0d/t7nXv+GsAx6ogyFK1jgidB6AlH
O3wsQr3NIoZeb4lBX4kuY6CwqZsod/amGiAt39Zpn3CI1vQ2/O2iEopErYeo9d6ZBwueHzugdruj
wP8BuLJ66uux57EiBe1o/Ace/49lR2ejalSddLIM86OnZSStOAQx7vaVtx37ipPhn67ZtPJboCVN
iEkqQqGhvHHkoxhjxDgpqWZQ5CpVl9LcEkYEVEwxMR0yQ7hjgi0UYu+LvVYsdcGjs3ImTQnsSmuY
1cMwS4YwvXhsJiTbAvIbxsmFm8zHqW1GzNp0jyhbQPeU/Jn9ddPqX3O3LtjwJS1yU9qDo53a5kKe
vt42bCIvRmZTjTi6+4kNH0gwWrqCrYWGcd5EqqceraddyI4zDeNJlwdmCCuus0VFP3Amkcy1O/1w
qHgLMn3SQ4knpSP4aB39IUf0Hi0Gjd8kdTCK13r9LeCxFqTO8t5ql7mzMjl6fb9+M7fBwOhMTlXT
Gl+VOkcCvKrCF0qwoZplR2y0Y/c9uBUZxGwr5EKGUsfnXjTqx8B0nskxfHrIz6WGnNg+jg/Albsv
injmeN419kYRLSC1o2SPBHaAt2LHmbQ7aTqGy/i5Oa8b9FxpdSWusn3FQh5OnQtwZh/8a3ep4qP9
ocAn8Ki/xDoaF6U6MxNbYe07GYDha4ruIjaDN4lYr0L0p9SR3Is2hw+v/IsNpgrEchmmAnH07XWY
Ai/GH+2Aj9ortC12ZMLM5AAJlQl6l8zw8ANMzVD6FeIBoj75YVVadKQ8kr3LCAg8GKwxE+yPJ9+x
ho6NFe8bVEBVyR09HyvwUEnij4NBziYOCMD++8E6vVN7zh1bI/+5x95RwGRHLFHtKaS5rnB1/mRv
TB7E2j6MiDjgNLZmBtbX+gNLSVjwMbbrxDD4dyjKK+IIo43pJCZ11pLdbxm37jQVaLz3l4x9IDuB
pSp3wTHX22lTb6wye1O4DQIWbp8VfqaolRURHrN5ZVhDuBu1tDXfnlfsyBuYrTYuYj7jnqVz2IMH
NgwclHfuR3vxqrmHaqicjNcel+c/T+DZFRjZDjWNSqk9fQaicgDwCRIbeOcSvBQKkID+kCGN/aPM
7Ffvojl74/PUVvnDUsHbR3otrEsqktTBDKBMXSZZujcC+8gYy4qZGd9jlrRGcJ41tMEKEDhlCB+K
vuwru6Bz4xg01niSFmZ8J9zo3m6gBahmBTHs/Y9uIGI8lmXz3FdoMzcrZ9LiDt0p1b9Uqcy5Ykjl
JX4D46df5x2WshYN5IaiXT0FKkiDLDUNwJBEE0qXuL5XMfyK/GTkDfBgoQxB7YjeBQZUwYQCOp1B
bDjdyaugQwzox6EnC3G41NEPNCeVIRNP0Ei4nGLlrIF39H9WYmG0Xc/OLT51qezQjLPeaUmX8ERl
5b68Rddawe8/ZhDn6KQgfRyR8S2iKKiOM86ykREO7zdqbKSl5dXMuFcxY7Hi54osmX4wf7jx+S9E
D3hzoBmovEF2MH6F5Q6y0ZpktOZTZyMGpKl7xfLMJrLZdhiwkreh9Db/B1fSZvMqfx51iUVJSzbV
qytWuiE7CLps+feo6ldKASrQh/lPnUgoHs7/Sl148C1/y4YUCaMprgGiPBVEK8hcQsZb7jxluEfv
4d57cNBbTFARowLf6ZrGAiQO7ionpY20Sq7uzbP+53ngAwBqtvxO3apZSyFokF24xNFXNg6wCP1n
EYcgORwmzi71XBbuXJ1EzLgFdToqRbHsl+1VeUaKUlr7Yr2E3m/pR7Ik4N+cHB2zkySX3xJ93j+q
Mijm5qRdhdY4WSNR2Rr5XhhB6LLJfBX+YXiJ4FmNa7ArAkhvbq8GuHL2X5bY7J86N5V7t+hIR2F+
CHmkXzVVJj+l+tVXv1WLeLgN0ys2Nyr9/prn4SgquoOl/A/reGjv2VVIV/J5z3hwkVj2K1HuDM0p
l3CkAGdKqg51cV4GueYs0lyNp9e0q5itACSjf04ZfgdTkr6gudU+G6DHjBLIbbA2TWjpnISeU0fh
Vki0pi41N1pCpOGvS75Xxyw37xW2twOI70gxaDEIolCGiiXAKjkEh5jtt3T5uq1aJYEgpAhVfzC1
fH4SCgnTMQ2msyW8l7hiRmdpcq2Vqe0oAhKgxQvahn70dzw36z3SNji8CVnwKXhtBHJ7ByGNfaJF
NQnU7VjyQS/kdfV+TFDuEzfEiMoIzGnIk+IxRzx0W2lWc4HH/z880ZPgMJyxLrjo4Zdj8IxPbrVM
rqXtVsIg73lHtnKMt2gbqhg/Q1XHZEsWBLiHcg1y5TcYq93XtjIZx9Oz/jSgNk8/lKPv6Pf7dy7k
yI3NfvxgnMUuFS2/WTkyWh/fnFUuKOl7PZzzmXrBIAu81Vm46qL8Xi7364mWjjLUsGoZipeXyeJj
j7cOsy6LLm58Jknz9P/e5lsj/KhiRe6IKNIFTaM8Eg+2RlH4zSgiH6CLlhaIwtoxeAV60lZvc3tA
3/ZPl2U/YLzbYGYS+Lf47zXKnJtUfJyOujSBnAFghPuZH8I7IytD+RVZVqfXN8whxKmKNqUvtfW+
wO18r8aH7QFSvoYW4+fCQLuBwpeLjh/TjFROgRJ9K0tlHnbx0Ji+6WAHGvFj/51RtisnwMRD7sYN
VAs7pOGNKcN6Qj19KIkL7GfWt48Bad/wqIiHcLhoKHakZ2/GV1g/pSvt3H400TZ54CJHHBToaXH7
NYGdaiiloFTFk0WzQ2/XMep1rSVW2gXvOeCnTarp2V8pB4CeyZLIeBlkkHnTbnE5v90ysIxBltzK
FQgYHnavBIyKCJ7Gsi0zlbjgyQpJh5VB3EOoaeKnU8Q5dFs5NRySDGhPtI7tqbxMIUAYscFVMDaf
H2OGqP34W+x+isLGZ+uS4GnAj2/OVg9qxeh/+dSAhqQbby0kYi3NIjm/gFE/6WwARSWtbeVzcKb/
J8i1WfaV7DRos1XIED5AlkHFovo+7BbirhxrfzY6+Bzs5hfmI/jd7xAUixU6XYYI6oDqb8MCzBTJ
DJFVvwpj1is42mqjrvGNeiPPx6OtG7ViSIlAjVhWRsumCMHRpzCb7X8PRG+K+aDnEc2uIf53b8ZU
lbkjS9aU/Pnbl875EXHe/QqZBFQpt4KrPyRsx7ikRszs2bTD+qTPpTng1tm3dkObqEnrTH4FMNWP
O64ie+7FUneWva/q2IjjT9spBZGA77WyM+2GoDAEsZguY90mt9uvzMvJnh7tl8bquv3aWn3lNNtK
Mx6QiQYL3NX/mSBjORboN+nbwXqGyiw/uBJWlBj/dx2ldzU9DYYjORC3+EeDyluQgNQ+89YFk1dR
lAH6EVzkUm/5g9OpImLSaScgpf1k1h1MNbGXrfYCwz9Xa9HNgg9g5XidgxpCEv5vUg4RTKTJvn9d
Z73+V3YEf6CXl7jERMCmU333+tDuczsiAJeDqpvx2p36KgYRKXPxIG4KKluJgkmDdH5BEcZ8H6Z2
Tj5+t3JQncjwaHApXNWTlIZxeJmvX/ZU66TIsu54szitd0Yc9O2jcIYbHcQjgK7od05zN5FOcB31
WOr/xHtNZhz5Ul+HQOa4U0INvwT01Fa2ENdQFJoeXINTAPo/7wr50ELRFxxrL3+TGQfSM1iorgVx
+dC5SMIussOZ9auW9iO7ycfHpIJ+G9frpAYjvdXbljYqR3ptKBW1+N02Kc2ziteDxGfQQI3vbMPv
ebU1SSFuoxLVxj9Hj9tSxaPH8HZhdPwTni3WnYkTJjGuYy2Jc8Tl4VWLr2HPw+qdnweo1vX2JgR2
B+3GhqQp13p68WtuG4eQ8Cxv5/DQEhiRVN2ixQYch2LfwOD2lVIJwJArEQqwDG9AbM1btFN5eR7z
oHWAJc06hu1TOhsRpPCqeygu0XWBm+PDDi//8dfuulzwnB4vYziE3dsD8wYc9sjBuFGd05zMqXKj
5Uy9lxxsadYSZCTQ5L3w/K7Rfi4Ii4lZTE/F8Zi2vGdZWQc3wQpbQ8/UJ3sPr3dqDqHw1QNt3ThA
UuE03F69CBhvOL4JcvxW9O0u/vuNYx54mGobucmSbciMaIzgPMlIoqzje8I7VmEGs200XkpT4ffQ
3sIJhVcawi8iWenYwiiOp+CDexKc4oj9J1shIRp80zPzLuDRvOWvigZ0iiiinlPWtOlWgQl9cE9q
M20h4nC/Cr2BQfXmkL3phzyVol+puSGNmsC5rRY4KnP15VH7OJmtZYqQC8aouwrZ2Q74C7CoDhOG
o3Br7GgjF/OznBPVx7nTaEoJDlyyobVphBB3anityDVE62kHOXpI8KfHgd5WZFv5egRGoKU44pyT
j1Be0VkootjIwbucwB2OQBEctwD2WpyiHZciT5UC0atmDwmFqa3P8qrUho79ZZrUAZi4GjO5zaLf
PhgOTvL7MzaS5PKAzUwKWnkCP7tQEPXBrT65npngKKv12srN8Rfgcsyaz2bVE9zWKH/iORJLf6f9
QLopFaN4cIabpnRqt+fE3xIxwvmxreI5SP4sjj43wuzn0Qzk/g2VCGa0z3BYLbu7K+A0TDLdxIp9
iivfFfpGJAlQ12WfZ9/o6tLKLV0ZZ+AsjPlFZCCD8R3uw8r3yuDpu8aXEse2kJeDJCsacCshJMlN
Lop9rjUJVdbOnb7CjZHW1rGOPVkthFV1IYebb38mhJn94LpKYnLGLtmdw6t1wOGXjsryXvg+oN24
n9YLRVhJWJN1u5dc9rXrTWIOEJ9tTErnwBRM7/t3hozwC5Zu76kUxbuOhEqV5YgqmeHPoFeeHc7a
j3osUrUhmIXTZXhpQpECj7KwDAo8dQznFBhUUcSijnlfNxAMBgkqjKSy1dNw4YL/+gLZ8GH1Nlum
JzquZqLx9ql6Zsby2lRP/alNHE/T/N9+nmsuHTpajWeatH3UxA2wC0Zij3CtkjsqqIrng83htKjA
DvzXo8+8o2sdLrmfVONI6/MqVC8EDMkRDRav4JQe8Cet6wLO5otXgHVCX584EQVSfpc3wkLx2qoR
eAKPLVOPdF8HumV3mcK5WXFWZ8Y5jo/okIrn830fTruHeMdhqu6L4Er5w5e6tp/+723OtRfXy6qG
x29AuijehnQCEIGw87FsgFe+6TqyH7zanmQQVc+pr8ckRBWSytFMeQFDlcyoHcqDjptoDcBKQzhX
zlJzDA34nAbZB06zdewxavZ2EKUntQyIz5UXHhptWvFeIdBLzZ8ryISyWR/C3YPcSdYgLN9GyBge
pYoOy6YEEOjq3ZROg//Qy/miKLDBQ8K5RuMQAUQzFdzjV+nwtWpvP/hjrp+fyK8wWbVuGJP7btDL
bzQwfDmHyYGhs3eWgyFxVMABDazAyeG26FntYYErBZ/MZfKIB6hUzqxSs5RrqhSGgrsl1NX1kX1h
Azn1OOSCQirEIoRDlExv2+4azSCopJOJpXoPNFB9L8UC1n1wj0ifkwTjpT1qgRZSDokMsmOOiqlt
rq8eOaM5kfPXkjfbpwv7ju37dclpT+tLHdvciGM0IPUbb7ppqKFdWCZf84cQqYM5J6aKfKZvLkN3
s0JEyFLBb9g4wK39ZGGCCHdkjNlI6OF9eRCJgZyXqidjv61GbdyXvClAmLEdCoywJZOblRgfQByK
h3to74DB8COVsKnk6FzfSyawFFZAiWZ4AqxWZgYKsV3HoN9a4Zj4VwQ5jzqI5rMNtHEvR2odFkGe
HeWYVIkucc9tv+MQKEkzGXW49jeTMxbrnFGkHhngXnMSqod9E2l4nKLV529d4/NNZCC2MYS/az7e
oqJ4ZR375IP5WIGB5wf0xXn8/QaQisf3QFRag2w/8w3X90u3F202zjbiq2QH1dh0AsOdCDiPYuvz
ik/pSGezKLmHjGKnJALs/R2PjKs1nILotngZqpUDg1PF/p4Ht1qg3gGM9pT5txnICQp/c921vfbT
5iHBK2uKEf7vunMizEI/Z3TrCFbhvtDzTWl/Mhh6ljbaShRtT/5PFhuhnmAoTFc3eonmRYKy2hqc
nJex/vRlERcEgOm05nwk8NTniGzvqHsGprvXOYIL0sHmx/evNptiaunDkbXSsNovSzx49ainDbK7
ZzcOFltGafprSR8YKZbvrOAI5dXinb9VEb4UWp5c7DPjhQRI2Fx18TC/UqmEGhh9T78wNJ0d3WpS
dEa0yzuALYSg/1DlfUcukAr/kKvJi/FBbcAbZkLCxx5RQu/kQEsuM3yj8Ctpz7CIEuOfvoWFQWQp
Zt3F3mI6yuXBqTtW3ea1PqlyuAfLj6pIEeLIXw75ssBUECro72tqXiB+NLyZQYz/uWyDtiuqxstR
YLaRUWxQaeBDxpk4j77PktGDmxRpStV/U6XTaeFVj9UwyaMLeJhwE6EdRQ2VM/zBD8BQFRF7rT4j
X0s/t2DVW03QQzXH6b7SuLW2l1cTJ8i9LYtb0YhLGZynB60pMHWRgjjK1a29tEFUCSKRPz8alUlM
t9iADSXe5noW0jBzbwB1DNKbTNGJd2ZgdhVm4Fs3BgqLp5glMpY8PCh5ZmDwMJNzWJJB5HDXGJsG
DH1XW8MEhsCDaw++bVKtMmPyalNAczTVEQFynCuUXGdBDUbnilMdSzDbMjdL48j+G0G7cWUSo6bs
Slq58toeKkVDz9JXRBOZAAbCdE9zPkm16HchoSAr8YLuaIIVQE7nO0XkiiPMVUuS0U+UWqV9gA0e
QI5CdjZjpDXDB2mEx4ieyWXvgk+DWwkPQbuIR5CgAHtL8nUqU2c5iLLluSBw02LO/c/t2VUHYtP5
T88KpO9lHMPHD1hG5OmnvAe46eqJ7Ij0wWVHTii38NS2eRtigw4VjbANbAJmR2BsBlVcCFMu68iB
AWygho2iIgY/VeJAMFT4P2WRFtG0Rly3Q3GB9hEc1MEJh6dAZcgfUZPyMU2P2kG8GijLfeVYHxWL
cfUljStOttvWXNeJ7CqGLqlOcsG0LGOa210Z29vSFumtllp+84u8VpLl5EHB3Iuyn5K7FZpNrOXL
oV+d2SJ67T0QF2BFGwgROoc08MiNDGwT8G2uDQbWr7ObYbd1DdKyG6xaSK52Jucokgye91jS9wji
G6PsXZj06cwECKyQ1NFBY75jmdehIxxRLeITWoh+kSC44TFqmngY2UIZdlilDcDqJv9MQYqLc9PG
gA57sRgoLzGVkgxy25T+AQOXJ9cl5qPh7gObym80Na7Kzsn7Ra9siWfODWkNbtCk/t/LM/6OdTxf
foLh5AJ9xUQ/qADSQ4bRFidNZw02gPxVdnJTXFxZ5CIDwpPQTg8WuJvyeUQ7tMn1mEBDEPZGKnPK
JXSOwAxRJJSsTrXmiAuKX3oNWvirxRQQDrwoesvbuvXyNqzZczrDxMA0/nLK1SSMvnY2t6ugNtXT
X36X/iCP8HA6qwMAFNSqlnqZBLb22FpLBKyDuWWKVo79f60oZFtQQKcpbBjBFVbvjwdeDvGCknxm
lZ//K/wd0NJ/a+JGqgNEZ0zHSyJsB2/xCHuckO9wnQsVzzhHBD3xob3liNs6NYxF+le49l7n0oK3
j1HF+hOWat+ERTqA0tZZMOIG5GGM+UX4TzSa4z/dYKutEuej7WjsISP6ldMpWFc2E6/O5Zz2rGXg
QBasweuXyXZUxSVpT+MHO7Kn/0zGHfJFCdiVacOkzwVHEiNGsjfTMgB+ReltNTz4OzLhO5TwsvJB
Xed/SxANkwv/a4ZdRT/r6H3WcRc/TDRLa+pDQO9YHum88a43HO9tDQT6qy/zQXFG4Kull41nnh/x
zgMwY/o7GZi0pMRvMi+q5lm8/xj+efPGeXjDZFQI1uq+DOyR9CmSr33WHMYjnrl4tnO5WSVv7L+z
+jVuPe9siPaFMk8vaFBjHnzPKEcKWTS3V5DTtt90dIhMM3N6VViFXhTq5VdG5urlqq1YRFipeWUB
zhuMTigQcMt84hN4E+KLlPWrMzkccj3TjNhybJ5agFrZwzf1q731W+wENshyVwGJjHn+kBnYuKXS
nA5d3i4U8PI8VH6L1ZNimPxAkI9Y8/vzgDYAeml/dF8rboD5saaEHmFjyFVbpfvQ9tJLbMBnv8tE
heCzkAST0KkDofbEOAnTPfKpnI6g9TjCDYrojQ3eViu7u3biWvGZY/sjI/MW5UnWkqsfhCESLFw7
nSAmUQBYOKMEAC6OTWltdeh3DGZOmJI0lv2Ep56M55x6j5KcJ0L3g5x/BKKcW8CoRfuFSvGS/ccv
smnMgz44bu/7+0E7FXXzPkqgwLwB8qC1PVcqAEYbn6hdqAfUmaKf3pSMDn+Bw2e4/WnRbsHE+v3k
FN/ID5LiSPm2L+f+HjMfLsU3MvR11xJzxokUmLoXdh4dmAwUk+EBdfmUtNHuvJ1CeeDorRinzIi3
Z79a4OYLzx5ErEb/VEdpmocIDEbqWldO9dZQucbB113I1GHIwnB9EgPH/oE3dTbyG2vRurVYXY1a
9Y0NTYCjtZIgfcYuaOCoVBDVVp7rqMQK68UOxc225NFsYt51hqhs/DjN3fy+9o2Cbvnz2eoVQUed
vI6X77BYFND6pIGETbMmoFiTQUKSsRUAfc7CHGKoJ5aqGbRySkGu7HO+wJe3VVBek/JF6MfpZ4T8
9KomGCu9Xb/FbVqK1l/y0e+3hOIPN6a46vjl+Zb5GWGThyvSTMM/LYu4TmadU2yLeoQFvAF3Idj5
h3NXW7q07nPeHc3HYbMMLuheCYg7h+UuB7h98X/4S23c7gP3iQ3ddkpbd+5ImXmEeTSm+9uu5l7t
Z8U/UTwC/DnspnsmHvOs5bOZOgEdcdLvsezRrXI7ixjpNeOmD7G1pM211f5oFBQC6q68yoTxyKg9
EMkv+jB3HjkLNKV24hV26YpHqANs3gO56VZIEsbxNDfmAnauga3xZ4fpCPMNetdC5+e35746h036
Dhm5dzyW8rUTsl/xhPjuqufiiELtyiAUgv/Az4boyRyc5JQjMnZ8m6YgV3YTVPD0PdwbsmSylBwI
L6fZmFJeH1Yc3s92uXJgRwgT8MedFhhHs/3Om8eBiWLGNIZ9dRJlc+NI3D3lZRSim56MnZ/2IQqY
7jXQqX/k8mxOXgANZAX5j85OSWQ8X47nz/wKF+rM1X/QpMrfqb0iWEw39HycUfTGwW3HGDH3Xyob
/4VJEZirwQfrX5TN/gJMEmsNae2itrLY7KPGVWrXYVz59kjQvfBe2x/m3W1cOXgk+c0R1QWcUtW6
hb/7AJG5pTVNpgqFqsiLL4HPEHTdVdTCzlGa/JRUF+8lczA91yjaETKJJZqlcVt7hqnvC1XwL2pO
5jtkJuYLQqu6Nmb0Vne+ZkXSWDd4DN7ng8g41fH7+0CAfFYHvBSMqjn5pjKl7A/TU+T276Ha7Wv8
jVSE6Z+pGeOOgznhPoetQpLB364hHQsywl7DWYh+OgT2QByB2v76JCSxf762EF0RzGLBIT18zB2A
Oi5E4+npM6BumypZctkp2/+t72GRR0k0jF4QD5Wdc6SFmeWhUIRhzDGdC481QhGpa835dtkiiLD6
IefkMzoxLgU5E/MSYJlFHdnXmZEk/6xvMDoszClw5JiRIlymeHeq0tFdIftDfCPrPTje4lrt/kIs
C3+Eye9+lZ+o6PEVX7UOtxK/2Z2s8Rml+X93puUKAFAFJgAR8JhySyDkGies3qhmkrhuZmDKqawh
3foLaGr5LLDhS60Q6GJykxvGyAqKb1j3n4dTfdObh8DHnOvel89i/QsuI5iWqN33NxsJ4V+43hBH
+2hOAfmhUgZ+1FB2VyZmTE87lWb69Un9hbefTpiWFhPnNBAPBwoe5JflwV9uCB153aXxOY/N2RnF
L0EhakRdhcSwxgO5x6u5E9+pSOaiNQLx+lZlhYhnWYqs7Ca3MRpMW03GhCSDzRX0AiSKgNmInTnJ
PuBXJovGzAS89EozEJUkVJ7Aap3NZECOJ7F3Uz0jnkqHT5wkip18P1ydK/Bn/iRZdbIiHf/X5Nve
Szd0u8V5+zScBLWSz4g6Yv88prKSL2ysesRRh+PBDWlBDLWgOFTML2z38UcJz61eMEBgAWw8djCQ
SuoE2jn8CQh81FqJMkqZntvtOftegvq4PGeNRunFgsYmVhHF8gK6YkGGA0oshD9ccn5EdaQyCQUG
Ya8r1FyaIiIVihzzPqiLtlHWykhfdjEGBpXQIjw14taj3RgoCD+WCBj71YLaw/GTdSnsOV6OKJn5
p+EDrJid0jG+9kXSgd7CDuj47+NiPE0bieo3eoh+rW2l1iiOkm/0sW6jSKi4ErqYkwdl0OR1EyNP
G+1vtCI5E6U21QvDKPgm0ayPdNtmUqArreHoYGksu9UQpErAjg8+g7FfXN6nblJR9xHxaPn21CCa
7lGHg3GoaNQUrzXOpQjYkY0OsaagOXd94ymiTESCyakHxiuTUinJAVY87Gc+aPiJIqwtutfm8UZd
jzNjuDL/W6PIg/S/mMXC6F+QFDO/Nqu0Hqp2NXmSwTSCYm4XGOY3z16wyiSsVW3dfkin7nqaVUOo
C3Vr78AMoPraOLewi4a6AALbqwEQKAXBWTmw48XHAIjVmg1wZucocbSG34RgmZ76C9+igK3eWWYQ
eHGgBEIqI1IxQCCt/9xwaoRzhdKABlbRXLymVEGq3CoWXioMvF0jQuymATuLbSvKVit13E/D/KJ9
F/RuDJCpOZnX4fpO/z5MxYNDAmGKqahQOf92muZntTT2qwQz3E0dBiyU+5eAyq7hAbyPq4xahb6O
TxuWBZf1c0BqYvm863PU7Aqy2zSSpA4ydtpxJAvA8d+LXPx4dudYyVt5dakSnRqK1NE/zCm1djRp
iuPURBEwJpXmlOXtaJmoRdFRpVLhlHEZZtOAqlokIg1Aa1FekwNdWQJFo9RzVCGcSNk2DBNknGMp
VjdMT1qZeN9np7n6m5Okz+4ySEMXXOaJoY8mdb9CTC+dFjPw8IQfP2O2ubYJYROo+9gTt2vgvo5o
7zYnkxmMNGHOuDFebFIDkBGQmQVJB3X1mxRnA6i174H76UZVDNlFAR3yXKbmI4S5dwdUkS0e/wfH
+FGMikBqyymRlbJWGYvWcj40a9AQa2k4sizbfono/7t2J3/dhjEee6oSLLMioBkBOjlTzAe/DfoJ
cY8BJIZnKuo84jbZcaG+afRlExQidEW8O9GBkasb6kfvXimOkp5sUssLqETpvfVvzwFL30/fSxet
TlqtpI500Ly0x4SQce9W0q4VA+fHOzyKAbJEXoIrotXXpTGBEHXhE8hQZA2QKH5mcfZbAr8hhNWO
LoC3vevrxJhZlsaQVmZz9UH7KNZ2Vdwx0TjpMPuoCmO2vhtTOAlXNxMMOcoU+HNfOoiD6UTXFzlz
zx6MAxpAT/AfMockY6qPJmsE29B3Y+CVR2xlg4wi5h5V4ja/gHQWM5LI7+Cxd5Cir8Dcu78GfF3K
jqzz2QMe1g5Iv/vi+vyJols1n2sHGghblRueh4fv7kxVjnnUqID8flN4SQ9LV343zUFtOxSar8Fq
fQsB3Wm1KhwH050TOfr82DlqNBoXL5PFKA3tfPN8YPD2gvOohsHKiZpsKTdELHhYHm8Fw21XQ6cc
t9xbX0wMBaBTK+KBj1fw0GgCBVIMSitpXjJbsK5MvHM/kSBH0EsFF5w2xLDVpZ4XFDrsrZ3X+lQH
bFAhuMhy6Qawp03H1hUvaySkEEPvj/6qOGH0Z7BS7xh6YZLruiyf/gg7eG+2qUYQZx3o0CXnqBXL
wihsUPZ8tDTYet7fzAMkl7Mj+mkG2jHdrFujFPhVsmKxwV270RIgeXQtPd8QGg5aZrdn8Kp9n9x/
5/tN0dfnwC5Bh3KvFXN/heG6kd47Ms1eeAJBwFreZTP/82HdGQcUXQ9SSSRkoPauzPOPAALoGWLF
oIInmZ6WJDpfKx708lj3JRfeN5+igU0OH+8eWV4yvWzB/4nj6KLI5NzJdWjniA1uvjIHXMSgfSiW
xwJ8Sj0c8cH641qX0gPlC89iET+AJmPuFxuCUu3D5kqNHMhwflNRpPGinm4ZzLhWvNiauFh85UTE
8E1O5BOhJ5norGD+LE8uaoiYUnxcY4mhd4WamkQY7e22fUErETk+T9bhiEEvkgwzn/CCZF4+urih
ojpimBMMAri1HzUAKyEH0mELvMXXOAr54tog2MrJORfoRLPWjl+cwHuLUcSzH4EOGOATDm9BjJly
YoVBRH/b+RkU4UfIHSJ72LrUvQDR+BDMhLrYN+mHmiEDQNvVFjmV97MOUE9np7hwAlqjjtpsPXtO
sCW5C9X5YOa7e2nwR360dtQPD+QQ9x2tsRFaM8OG/9nk2HnPIT7stC0T1MHrkJ91R2aEpnYqpJkQ
dpKcs13ERVDp/XAJJExwzWR++9+sJZkHB/NcqGQkmdJxSF7BHpmGlwxOzekuIZccfsQJOTBVJ+Nk
242ZF7AKTpOH/5qPnTRqmP4ABMH8wG7XHRkPFP3I4i7mLSSPall6AqMdSaZuG5DdlwpsQT+clrFZ
LJkeDthi6Vz2u9xnyjEnNt5HXD3dOdWXQOAorozc+74lM0/m+VhI1hDKhotuB0vgFSF54yaQvsOk
Mr4n1ZhyEYfV+vytwU5XQFzQOMn6Mo4youRg2MKqHplGjE+Lk7QlxkOxSbV3eu/J7ITZSlJMQF55
++cm8LH+c9l9hXdn8+tASSGyk25s8KLr27+fAUVceiEi5uZ4i4uOMRY+YK9EkHEBP6rJx2Ua5Uhi
2a0WYNDPslFfvxg+JEBNktrOsi5KnjyvcL8mXUFEPOxrZrQSjQeD6xn3BoeoGbR5enMGMbBDZaDD
PfeGuyrZgJHVoefgOZ23ZWGmhxTqG5OG3OwnhtrtTqVPNsnZcyKf/TOzc+FxeXGyoDGYHd3Ztke7
JfyRqnL4uSmwBZM9lmECZ5d4s+Ss42cIXWbTU6X8rJHV0NEQHMspCwd2CFSiJDQRj4l/owsEjFHL
+gthvSRsD+udZvWsCE4srS8ooOzXe/BVVyg/vEfaJrGw51zWD64UrDGSwrEAfson0zBdxgmXbc2y
ioy9alYJ+H24lvRqIzXvyS03P4VS7XoabQ/dRcIxK6jlHPQmXGYtYokVKHK6Ar/FBHlYHxToZhzl
nqgGLygFaH9yLpEL6zf8emlmOtF6xot5IF4QT/RoLbAbD8g9gEFpW4xQIoz8brScAla+6M79V0MO
99VP3DCtTl6mpY3XaIrQ3UBMSOG8zfyz3UoQxKQOmv5AtIk3/6hes81tIRFi8OdGt6YTaMQRIsGX
nnbhbOYptSwMCxdmtBCqgAKr+D7BSj6BR9zIu7fSjZs25HX/Q7C4tUrgNX16DgwUZdY6ASWiK6+H
asC9VIXMvymBn10YMugmMhGltRIUrPx01tu1hnMKpzsFvZAYWgUSyitxqft6R9huQD1cvQ4aNqKz
e/7odBABwydOZvoXZ94S/rpt1aMmheRCrHrI3cJwsijOZzMxAFeAQCYX0a4NqxFyhjgI901F/DmB
sj3tVcgDTCpn0YXAC7dfgaJQ+6bEWYP2DMmRVE7vUQirH8CxDHZuqso5RqWL6mqTjrCATdZZnlHc
6FnV+O2ie3zUkZaSzFK3jkPsWv19LciAILOBEJi4UKkHVqUUHuWL1X+iT8n65rQg3e7wBf5biVIc
L7qsONn2pea7W6XQAfGHeR/l5V5iSZox4355peZUGtlU5aI7GvZLROn5vM+hQY/MfS6Zqhtn77MS
qNz2ENOpHzUJuvCuChlXgyXBrH9kCt8DTWgktJ/OBdDhGxeZnMk3jnTn+MAiY97hl7jB69MNCtGk
h5S6CDLt7OSWF4Z5DOWlmr5zXmYG88Zb/1X9PwuK/vBtrc4KrVGvEACAjQYR9zmPuHCaR1c+3OBE
2Z5ANoP92IwsevnfpWhbG0LmXKEfeOFwycuCdZEk2M9+MFxuWjCGK7wRDvfwOKAYMNdA3P+31o+o
zw74U6/vP5xJlEeBT3Rdiw1IXoeNDDt3HW1L+66OytRqFc7g2TqLEuGVuTl/zjLULifFiJ0tfaGo
x1+vxQm6uAbFyMid0ydKg66UR9QKKBVYl0BZeTvHrOyJCOzzV5doTcPPoIYFwEVqorel55/EJQFr
1M8TT7molZRW3ahuX/+mI5kqWmkx99c5Z2BK/LV+MW6RudaTpKeuZKWCbHeKrQYCL/ZxvMuumuwm
Pk+vzeSAvELG2z/tpa5oKrEdnu7t/4eK10gAqYdr7GLFpCxQo6VYCuIpTtY3ovxlWClyInHgAr3Q
prj6rZtu/RmoEcv7/0l4k0v5jpt+nO5JMkyJZKrcv0r2YIawx/3fMZhrIYRSUMIypWaO7PIR0nsO
81XEIvojXf7uRzyzklGpdTxPbD7o4W25lHq455qSaxT7+KWF2HjiEobahomrEsyUdb07AB/WJ3KS
EdsW1HotwiAWjuvUu1WKffNwLEyUgLOs0liNcoI076CiszehnbrR7saBF28qFoMV0Skfez+gTpn0
XkuqfuAZD3mmwoHk+f1EuEtvDbxUN3xr3debMVHljDHAGq0QKPQfL7SWelyFsEXiUxM5z5LioQS4
uvtinNO8hNc8I5f05n1KiWq0WPNpZzgR6UONs60DB+7oWaBC0dXld0wnfex/aaFD6TeSVsaxo3ub
fdwTS9M2HVZbh86iPxnvnPGyoBQOuN7XOKVFiukD3WgqfwwlDvTSiHSnuBosII5GTxoYMN4CEvfQ
X7aHWbr6KKSRDqsJhs/lLird9Q0+RuSIR5WloaDjAI0WDQsK6pe2SQ0nuaLPT0jjRA31rbxzdrVJ
OBMmgHPkajcqtGC487nfwMT5vWd9xdS6jhXrTY1qBYuqzifb3kaOo0wmcZMPs22wYNUV5rgMgSPw
qMKBfCg9Na8L1zFGaNf76dV6VCRrm9wwvgvlm9Y1CfQYdqB0BaeJuW71tpFoPx8MHVY1dEeKjA2T
1YMZHLcyC57h81tYV2Cj4PMOe2XEXlnQa8GRJvjBkr03Up4OEfFA8COD4rB1Hq2sjZCPp6nsmdcH
Up+XsXsoCy9pLf0BPF+PcYCQbFAQNwQVrS36R99w1qZzdFb48C7DPq57tQPONinoUfVhki/d9LyW
k1gQktC/uxR/THRvkSZrkJlWOXqTVNdsJrDpAMoyXGwmiJ+NloFfm7NF9qv8kydMf3W/xJl8VGac
ejvStZanJDCjqopAkLMTLJ1gzrsHx/X877u/FNaHeuUjUPG4I5wHL16z8azdtTiG0fn/gMz8tF4Y
lJ+m+1eK8vhbcMpVTzp2JZcTffv//9yVpBkpEYbH2ZRvBWxucy0t2143bunO7efoR5rneQuRQuGQ
WXOwr32T9gWdmwEM8a8oF201oGPjNjqcFA7ov4imxEFBfbwKc4LYoGrtem3DQKFHbH7PNwRfX+y3
EMKBtifim17t/Z8gGNyNKFr2XILngq09pBqnWfi/wMLKLD3SXUFkZt/Y3zahLME7XgopYUVPGaRB
evLun0N0NNZJ4iR7A/KBd2HKmLwB3O9nGJePqMfcg3qlwFqvP3DMADxohZAXrdGme2Uu/prCpjV+
hLH2lcvpWPHnaHnps9Mf4pyJ//adiZk2vfalFhuD/rHdDbFE7IWcbht82zBI2klVn7+9eovOw9Cg
eSHX1VJaVi/APCyJ/obRbZq3CcosaBnyTtJG63RkAwaI0udIZ5m68vv5HO/iaEda39J2c5sm2wON
r2dImXvZC4S5YztnnztF+qnwlUJObQx4jGFIbeayDU7THblcIK/sxTjBwYI26dASSFc8EsH6eRJK
jXWxqTiat9XCbGRaE5VO6vlOm0Pd+BhpLYADsIprmdHFVM8TD1xwxTAqpXeZGhQJJBxVXQvuMaTW
OhWNR9L5huvy84x2rLb8VwcIAR5PI4yu4iXS8VhNo3gPj9Mn7sWz4WEbmzYazrTpHK2H/Ubrrv4N
PGB6yrAOluix9MjtoStgxpP7Zmk5LmH9qywGWC8qJwt8kfLMPd8TkLPcEcV14jF3/dPm2wlQVQIb
z2yEJE+6N9xd94wbyNH3evhHdfV+D/G10Vs6fM2bBRtBjifE1fcVppENoMBxQ0w+EV5N2E9VPrLy
Wr4hdQ+LclHFv/2c4BjkDtYiBgwHmQ6mQRcT6eNYufQTL3VvUWcOIb+R/qWOdwgV0gmaH5+6ZJFv
Jg5oeDy71GWx+BGROyvy2ivo3n5fO+aGUOmXP+7Y6DJQEy4f4lkJXjnBjRsIp2nAmkGtS8gZ2EWs
o+ik8dDCcMK+OccfsSnrPg70mYEgfwi58OXWYyIEs5Alwv7dXWxK9AmuWbPd8okyUCdxBlLamh2W
7sxLukMd9LodNfguyLLfWuhplk5R6j02MtUrZEkfrhTroWIdTH3l7VwjK/tqdqsFmX3vONelqJkm
bh9sCDw1U8Z/R0SVOlk/dvP3HhFsEVj7FspUPjTwjrjzq5tJ/730ohQEyLUO0Zgy4fzHt0678plQ
BV/l/2ZcN3cBh7lduoUcaK0ezLe6Vlz/L+C6Tn6xBYaVGCy0m/yziX/YTxF7qab7p646gdJZy+e3
2HpIDRfH6Kid2gEzqyTbOqDdHHQtgG6XVUi1KsDwODI7vyRmZS8eotxc0azHmWYhZl+CBf3BTmLL
SH9440UuBG6+LbetDKoVFaR9upKLjliox1QUFHZCjHHFPwocxD2Dpj+cxHyP7lTfBnVIdPMNOuOQ
KKS0oKvyRK4I3P28wqNgLd/mguXX2QPDoJG0DG4UoxforLB74hox+JJnutnmqpsRnl2XUgYy+LES
erSk8AqO6jlA8+XIQyGBcNQWLUlina7oQGbf7mNTnL8c5R/Wq87RAjCSHl+liZe6zvbg5j3LdKDQ
EbEXWn+DsaQNkmLWW229FdfMN+XikLRB/Ke8ym4aMdMuFL6xeQZlt6HjRGVZMK2mskn1Xq1zfqiS
lGVrbC9hR8YCxShpsodSQCVfb88P6djAJaglRvIxl7xBAP4GWOZsN8nuWykhwb6He0etTmMntMWV
Gb0a6HHtlpfSDoksnQ+EwtNVyqk+K5r8d029AJopMmJyIW+yExHW+ygeqRghZLiK9Wn9dfaIxpIJ
OMRHdOrrkk6bDMZisDvqtCA/dfda8Rl8/6bsNHwrmB5CyfKmWYaAShLrhMaRa/A64T3PRCZXi/I9
QQZ0xHKbPs+gLSLSrQo0fUEgg/LnqwZTlilUo9GzNDBOrmD/kL876YhI5aBU9CjJoKWqkR+Oe6Ao
MEQGQmiRVvYbFLD+V+DQTAkF9uXA2XlL/C8eZ3uvppmE0evWdYTh6gZzPdxMQmC/HQuS/Yj4U1Ey
YM4SgY4LQaOrnLmj2KgmNytDJrMAJ9YDdwCqNGDxv12OakJoRcZ+AAYXnuunCCG7bMKi4eVk0+/i
uBGvnwbpR4sWFmvymK1TLHtPZ5Tc820WkQGSiKS3XbkdCyJRHl3CCrNl3D/+TIvClOZHZtCP0Y58
f8rLQAByVXSwLWqqWe38C0M7p4cCFzClTSCVXvoL4EKJlREtNJ+/N8K5VmwSmCYAh4Hq3f6RT/7f
cxti4+rKdkyb/IZOuaZwAoRG0v/0+XI2lnw9OQE5zlSOGQnQd9VZX+7sgDBXI/yyP84lkAdvNMM/
rCQ8a08KScZnQl4CzBzu4TGbL8/dAyRig/VvRUJTXfJ2PudfzxOk2doLqdwpI+UeK2vPMQPHKkU5
NwaAzItuCXUxwSX2Q/qqgxgcQrxEWu6u0Vo8/6nD19iLE/3eSx++iICNuW5EC88bcdR5nojB2Lxc
0Fo8GLRfR45iDDZNILueLrLQfa6/nMGI1lwmR5/6wns2i2rre93SwzCxU7sNNsGzq6ruyGbGPs0w
jcTHkovL7vosZvZjF1uHytsGh6xu9PvHS9XW0uXEoa5GtMTRr29xes6yHt8ZTmGwY7AT1mwEkN6q
aCXpplj6NfVNNfu4VZodiuRghwS5Rxq/OdXBJ02hnO08SKjVefEr1FCHZfWgZBBMSCj0e2DeJV1W
9N9jK6A2sG1BXn84HJEJ9KPgtNpUVZ3UZ4Xhi3focYEsL6u11GAULD5pWK611b3csYvsiIkVpIkW
IBcMav3vpU3tf8ydsLdsPLflbiEGOWa2szDEtnPG9ftk5cy0bhO5IGGSZXRxfn/QSuwyWvV2c+/Q
C4wIprKjtlWC8Ke9cWaeoei1VktXwniNowjxwUSlQV0L1dYO/Tculy2c4D2LJ6mpSwaM5uGnWgWH
muX4aTAmPOsRa1+nLIT8MF0ymvZpNA++dUlywdEays3zK0HhgrGizfCVyF2m2FYz8LWd/wwMUvTZ
ABAQur4HGIXY25r3oBENErBVUHOKGpskhF+/SPewEczfzNFrJX5q+nMODwI08VEevbfyfdxc3OOj
6uBH9RkR8WZ49H0TtZU3HH5qAzgXQrshiKZMniDKsV906lSntlr1gFJndnnA66ThDdzCP+N7Zwfa
DGCae/eqqC1YFSquYRc8z+OQpL/VSwLlnOqsWGpXdQcFpNpz6wAGcJhibr45t/O/c960wbAsw27K
8B1miKIXoZa3ho5E7eblFCyk1Gsma6hanCngoVGCQWalc8qM7Zgmr/g2R2RKiocLMPn4t6nLwr0W
Ih32OR97YUISnAZ27VIrj6JYNM1xQVCeZqyerXmcAjXkDM7Whzq+/L/nRPEvkXl3kTQdY/tf3bcE
3Ic1i3YyXqIiJGnspcQer5XZhAZpNwabRttGxUjpowf6o4sKrIzamG5LguJSZDKYWABaSlk/D0K+
EsAdU4JHow7VeN33JNDU2AcDMYujECg2tmFFzvISv1pDCfthMgXbs5EutUgFF2ytKoXlf+qGhY1F
oCPG/bTfBk1foEKzHCktjuk3XPKeescn9UpD7O80LbC9+n27hpKwZixXMtqGh0n3TxSuo1y6fUQb
/wnqR7yBRSpkSq8KxTnuou5SM/eAJks3pE8ItxQWriMIzA3sQ3pvidMwPYS4/u+fmLqPovcUaWvB
X9UzM4zxC+uFucrKrKgZP7oHda2HyLbBlGirAACLSD9UcGTjlnHgkdU3n/Iv7PqGvuUwMXyL9WgS
PVTkRAwjIM4eC15tsjH7Ef8YqmnTpU7ojNLdyIVU/lbYljGdGMQ9EMWi/TMUDlzcqnWXhm+KOTcx
5v0zJYbpX/10BbhPwF0OTicl9hBQCp3v0eKT1zrmBW6ohUhOBMx4d7o+IIZC9Ce/PZDX6nvgNcFi
jH5ump1jyiLRdQ4fIIKvHh0evo1WH12XIqvBber04EkDhjzXzwtJYU/D0d0q1NfnK1zhYvsshQEV
3/zY+Hr411YyO1bECjU1IKpOz11xs9AbGEzVxnIc+Em9Xt39rOvuiMPmStWZl7QwRo/CltB5Qy4/
aGxQJI6Lbz/oCw842xvSwFk/cwOpJEMyrSN3Vifj1yJse7//JNaN3nY8diKWRaXdQ2ruSH7QQD3E
/pXn65HJVuAwhve+KvFws/Ig+OivDJht/aD2p4WMWapDjWVMSmxvVEW5mI5GKe+BFqSINp6eReBc
bkAZO7ybJKil8ntHSathrnvKCcXk0eUGUPz8+HN3GvgEX132cGDxMysIStTk7TuayVVL5vaqxVBJ
jKOj0E8PvqjzBSS+sssOuyG5O7pVFzgW595GiO49Z+f5YZOCkIAFp4DeyCNiyz42Biid21N+Ae06
QtucH2fucODQrzY35ZaibYbGgHzZugj13wEhCLDIqkX6dUJ4e59Ari6Yy9zjtrbMWUFM4p6FqW7u
iNXcqJ9QGd3Nm7XXyfWd2GiIOV4LnZDZbGk5Wj++YC/HjbcL7qomR8wjrx2hnjA0mSW7WE5FH0FK
+AJqi/yHRD0YjH92it20GdeHQI0ubYZeugQ2oF4iv9NmjIauNYAhfIkg8nG0M+6wSnaf8zteF91x
M+1YYjR/KKUHnFouRZqP3z0DeruehMYJt3SgKXdlLx6hDNgfU2DD/BNZ/xnD5s79AE+mVVN1p238
j8g6ERNaueuIlU8bpFcSFFLpOW0szmdC64IPeyJ2wgi8JkVoHIIBGEyR+1JReXne0NaZQhSrT8jH
tUdC3uUvzlSTEppq/xCZpyJUZ9Df1QCXeOltY+TuO3v310GbYmu23tru7D35+x7GazkeQSmqgVet
tU41D53Cb2ge+kaLvbLrw6W8qAY4z1LuqPxITIUUwSmvQlkKe+vIFot9j7MhJWSZTgTbKbvROJcW
+0+cwh4FjD2b+jC6/0oZe+vnQuuDmB7G3gjwUR5RmQU0WVDI7vcF4Zbf+ZMcui+UKWJVIR1lEB7+
nis0SZzDDSqwkz1RLLPWpArNy5tzoUFNosZd1dlFU1k0TqBBhoFQcqRzeHPXD4LQ0q75ZQsAF1IU
DYG2MucKEkZF47DVvHGdlfatHbIMz9HcM8hXTH6Xm/ApbOekpZo5uHwlpL/+jTtlcPPzMylwMoze
VhGmipKLakwiZ30UoeB0EdxsOKSMYtU0LyrV/JNZJtfT344ofl0TVpATUlO808kes5iNLrggGOef
uJbKOdrncYZJsJFhKgSmPpb1sg09GnG5NyijXZ7Ocf6PVO5zglqhLDirFzd8K/rYZXXG99jtP8by
1bE+291yJxzDuFZPNiWP4ObOL6jWJvpMN6z3n6Y/AvnyRwfMcRU5XgGQoTju9bgA5C88Y1O3tT+q
diXT884scSb6XqTTSzYArc+ZPPdPEINQFJKU9zM/RYt9z9ymDBzN4AunU+V+Pq2JfjoxQxS+oWpz
2p6735ksJJoZrsGEQk356FXwaB4czNy/3x9GKNzuaAb8s9GZTW+Fj4WbLKr1Q0VX07Sz8ZU11ssu
1SM8Rqhc1Gyt0kC+ZHF7fFVasL4/dUmiWgcijRmVXXL0AFVquQ38kc+W4Uj6zRAs3Rvx0mUXtQjn
CG+UPeueo+D+ca+tdfGLncs0G+X0Y14iw4VFMnkGGG+X5WRlvtZg/wBDBuZuoSBQNDy21o1jIo1P
4ezo8L79o3UMTL6SLaetFMX36NQTpdHP/irLy6DJaw/1w1YrlVakmOfwi04XCXl18H6Sh3/+QMJK
1JveAfo85WdfMnL4sM3Gi1+HVOuVugan8hCva+SrpVb9b70acfto3I7L5SyvSAPVG4xfIrSDREuh
5b+Yea84gLIqDOgJ1t+1GtsfPNGXyym39wDBSzCkzsre4Y5k8tACmRWOVs5GOMAWdukzoXtAnrs3
3OCH75FiDd8fZuk+DR4JqR54fM1HvGtsgyOKeqq6GaMTRr/1tgJTQXpiqqphWe0MyYF7VOg0ydUr
8kKWLfNLm8GUjIGknjlgFyfKr/l91pBb2Q2yD1LzfLyUkHrDvifDThc/h9Z0I7+KpuK55r2CmKsW
+z60fek/IS4QGCLlafbmVtrRoqSuTyUMbBGcDR0kRMHFuCUlDyxq/CX1mK9uFQSMyKb6Ht6zy6sA
/ojbiW9TjNav1OiEWWlBuCuo73lMgmULz+BLs/s6bMr58uUXOea9iIt/d5nd/y/dYJSro20R0RBl
xkDdSs47ku1JwUrIsvYS0Mp8DHygqOBhhDa/N9UKR8QpLorcp+tZxGOmtme01aC/wiqyVgMqbLxf
B0IMriHzzmbwzGqWNZpuYqkQK+BV3O1gd8LXc2H76etJZG9qR47OfppsDyxOOYpOJLusw+ufBkKl
x9RHfAUGT5WoGWnrRUcdPKJve52AlCSlMLzuOVGvsPnXEt24LsEoL/ZTskSliuC8mmsCrqR6LILa
Qs0FTLI5Ye7fA/GKoLRaryS/UeNCaPuARhWoAzox/iyig4A3XwcOptDbJjCuFGftsYOc/pNkKDYS
sC5hJv1klgtQ6ZyLTfGrFK8g1CeNaDx/03MuOaC58k0uuksBobZ+BGqucfSy18n5q43Uu1UiRm9O
/EsE/KS8V9WXUhCjG1NE4NWnNzGS6FriN1zberKILp/3/EhZ8g89AwA9lFPqtBxuXnNbCAXVhEff
TvlzzfhTnADhhmTClCewzfnkE6VkP8J/1N8wlMK5/QshpLNeQjJwfM3/QM6PslG1tf7+bgmbPkP+
ocGbkEs9v0b40c/RjTdqi079o2b8dO3I1yq0IZ8uxOrjcEd8s6aB8oePqF5oyy0IpwclvxCAYu5w
/f6+HzIHQOvnvZKzTUHqeXDGfr3TwQ6DLckwihx73P+mZUMw49LFdC2mFHViTVieRbwfKo9FIVXt
Fc9gf32CRDX+Ii6RqE4+eaF3hZDajLdKqCY5VPGcJpZfY0aJ5aL+6dXWPaA8cGiZC8hsCZtGJhY8
vXrvVgzIL5F8ev59MGXPJLAXZ0jsXlcKACy/hCLoQP9nknwQiBHbZKmbJCqU34VMRLAErEPYQPK9
vD3EFmYzbG60i1otH/StyNTVoQoZd759bcWs+uIYxknIt3LTl9Iot6dCFtttwcO4QWfzjgdYNZas
/yZq3RIQFOnSZYKSYm279bK7X56VYK0SvDECGfQG5vr+m1UQ1m6/uFOsAlIOWdE8XML7CC0nFBQw
qQV7yfvrYbJCRTAl0KI/MjcBND7TrHCIwUybrC4EnbWox00ItruE0X621aD9hnaqPLWx1NDLJ0mY
2AJfi4EvN7//NyZXyI17S9AHGgeamdW/bvMUciwSaZ2NSNveQ4Y+xcMCzE12sB2PlJkMSWfWLoXz
ZDZRj2vSvXukxm6t7YrvRW3SBDRQuQBa5EKW1IieSAaG7FHXpQqKBp0hMGHE3X9bwWD0L8tO+zqH
B/zL0beB+vkegMpr3kZrFIhwZUiie2Fd/pUbnpUE7zK/wCq2FxmU/eKIhvkchv1dU6r4+KWZnhKZ
2F4mn8uUGfXcILWSkZcZBk8yUPCR9IvQQXdRk9vO+HHVI+Syh9b0fK11E+/G5JM298OelAG+8H3U
M1pFF0w1VP+w5Cj0gOAWp1yfcmQhT2XzSas2d7d8mtxZnIdK+yqYARuAUZ8TsZQYO0djffjr2sRq
iXPqgI80sJPq/HVzsYdzzgcEwZYPJtCd5/MFoL7yP78B2tWQyQgTuw5QkzN+YbZs5xz8uwJ8f+cn
fW1gRKZc1cAkS1aXMiEt+8WGupIwjhKatdC220BstUOgBJfuEj1/0CP5h5weqcKkSar4HdMX/X1v
SrAZE1yX01Ta9NZW3wmDvya7sHT+XXIGwudaoi4Z25i1A+cWbraZR4vcdOjHF5+dSFgqRTlT7Od1
TJpr8G94zkWlUm/QpMKQ8l2nCLLzupSzWY1Njo9boInBiX4IONeGhCQ25mpyUbhCrwDD+nwnpNqj
KA6M0FwYLA5SturKpQqVgi58qPN6s5pblyt5iTk5v8/t86t8ysoo/n9qYZrotkoPCBIWiMLlj+W9
Cr82ZNxsj0c8bKitWaYtNHba7jYZN9CWSejISJAGB/MQFkHTNRIxgtFNqwrmSf2ZAGK/0a6B4bno
uVtMXSatNYitNRXAL4WEe8/FvHtDt5WY6mxq0Nlt4+Q36/1Blv7V728nzD7KXGIR0ay5fz3ma+OV
bZCDIW1e+VS9aRY5HTF+ICCf56080GhiHZFrf5V2mGuCRqylJUAOChYy0A0vHzz9NTc1kjyuDfG7
AYMRmgElBVt6Uhw3JwGG0jGm9ub+A1OSp+BWPuT3YI/NLFK1rolJtYY3HBIC11RmvzemhUr/yGs4
CamvBr7MIAtGtX1jl7qwJVmzzt999kW183ELsFJZO2AP7pVOPRnmMYINXE6pTtv8ow6261f/8YYz
xHY9slw5UyiRIGY5ka63zM+HpjI4i1BtcYCEwjzFBBNu03orMredRdx+zOxwzgJlyV3jynh/naRi
mB2ekTEbKiy5aUMHoyhv4hYOz5x466PXjK5RjBcGG/ce+0M+nQXHSje+gKwH+QIp31pFZ+rqL28Q
3h+jLPPTBFEVjpI+9TPdTOD4CfE5UYR75JgWvVI+FPbiqEx23tnEJ7kVtRQqSMENoGbFlO0z1Enr
YvgMT9kdmTkc0UQXlzP8iAV72eG7lrHrIokR2OVXt4rClLaRLkM9fRIa93bc2KHK5gfdJxAdc6iN
CYapfZi5Fv/2L6njBUcuCuR3Lpgn5V7s8Cw+3TrGSeER25mG8mCdSuKds7sw8OhtSzF/XgHW6FKf
CgQy31/6fGjshbBa51Mc4AjccLJm94GcXIPzFjFo3SsyfpQSsa/VFi3LIA6eudZJwY+aLR7F3m1a
4F9YgYYbsE9pKwn7X/ujgq5DowWvYbsjfYYweCoeuTuZvncjechV2+6VGs4r+cGF1hoHuaq170b6
rsLFbDXtq6bHMEFea2iq5u7eu2bj5OfE4oxBO73GCl53Ic+Rzre7cisnSYJrq8j1/jD69lE/5ums
ss7jbcdYqGVX6e1YbwCwZNQchKQ9FrvhyWX5c2/mqx6MW7f/pVpoMwQ5EB/DVXDX0P5GGmkIQYuA
4g0qhNySiZFp2xhSEYF+wnnIrV9YYU4+oAkh2DEJwMiau5/LwRZWuRIrX+NDAvP7QKfGHK98hgvC
tchKVucVfftt0QfegJEXEwZBFKewHZWSMXZAx5+IPKfLFTx3azKdZt00pZdK/4e+2hcLGDjki93F
8ktMk99mgwUJGvUEUlDjvX03UM3lstmUQ1eH8ov9RntLAAI6R70AahYW1weT08SNMyhzzBDNlWWw
m3CQq9qM7gtHwieqQeFNoVlPM5jg+XRLiZ1lnAAqnbOcjtwIfrtdhyjfJqJBazmnDVO4eRknlJ6A
RYsi4DV7Ka1XsXCSKykWZZ7BQAjJ2fXpARvfKHDVX6nRCXlZBhzQOqJzqyf+RtyqxsVb88mHOv2m
cJ9szbbpLKzQhlaaS6lQSjoNRgVAGklGnFQYb4+mIBiIdAbfayII520hgzUXZo0wXkl1iELt8m/+
FR92B+V9SS2mcoyZdAQ+DG7Pg32c6ecI6GLdfbMSR2Q1nHNznBmbDmPruG0DTuu4M3doJOge5CPm
xiVLS7DWPlSG4h72kfM4nUcmKHfLlKsOfljFrHUGCHbu7mV1TJEiQmM77wP7SlATwfe/Cr4Dh4qQ
t8QRIMI/Y/bsPPgw4trMcpx5cXTX6+i/m9WocWlRBuH6WJvAf+P2xArDC/YGmu3xjAAZ7y7GFTvY
5XwvaFUn3AFPiiqu8f1Pr3O7Fqr0K7Mugqzyi2Va0yC+qXn05PkSqQbD3SjCEXZN5xpCLq+Ry5GN
es2WTZFJPs9x2Ij9IAW7WS/eqEWpi+SvE0UGTenDL4+9lfXFsEnzs8iCObp78R2WQiVBWj8oVvGy
/Xi4+qjwXwUSq9IDEMBJ3DXOJ3stRD5H0bH1ZwkW7d7ivUb/UfQOspNHsjv/13nEd5OxPgV5U0LN
x+cLt/6gKgwB5032mpHuIF5CoBorlug9Ru6TFGnaShxvVCT4jEqzZ3d5biTjGSFav/+Q9fWXRyrh
y9aq/AJycEJ9n4gwiFjU2OOc1aRTqDT66VYRQsCugYdFhSym0VTSmTvpKEEm9H+Cwap9u7/gkx52
SXrji9dieN0pHEqv226Fl3tZnDK/WFuKz0tIaSHj93msyShpop4NHBfQELKn4Bu2D7JtMTrcG5Vb
+EGx96ktN9sEUu8M+DnO1+rGHeOX+T1kXg0ImPYIkCcpMXkV4Ld7zJyjSBEITf/Zr/oYhBVeVJb6
YwKVs+Q7aSdNPPNxi8zB8g3pbK2tG/Q2duH2U3KqBQUmBaLsOSc/AXZnSHaEuF2aiSChzst3VMTL
RC3i4vQuQHYVzu1HCInWJM+XSloDkkZwGEm3BVtLvV6LwUnG09DrsV0FXutGlxN9XbnxnfekCY+C
21Nq6u73RzxwS6iWIHoTXVbMWNb7ckn4b+NPR+5OTsRjg1TPWY1S05JsA++SMpzwGwxvMc82d37k
LFifXSc9LgnR5DAiD6ZBih5UGuUfZyh5OoAsuJt/xbxqy41Y84qSJLh5YXDj2C3kkG3IMK5Gdqr6
J81GwuazScBsAeiem5q4dym9aaoow+rhRyiB3n2N7yLjtmRF13d+T3OBdHDUC3VyJm21bjQ6vzq2
bQmibwIVMZ9M6MvmFnziRjN2zVLP1lEIksdhrtWQsP86S0nN+xczWjGkq41zK33LSUX/KbWT+Zqt
VbxkKl6QDVJD20yTH/bnUUvwCmMQA2DfWMNkT3+kmlEMqlA+X5K1cQXsk/6Qtu49lkznKneXHVsz
/GKcAUero3Et98M5uD9+s8g8Kv+YCoKQgCxLNN8OBGXorRSpVd3OpJPM6wuPvdlbUDmgqKppJmZ/
By8WYS6MZK06byzZGwdzI0T5HZkK91SkQUh7BZ7XblfeGj4pd6EexPw4QhogSIK0PGqB5Z6fE4KV
If3MipeFKZY2exRTGYqU0d3RiiEUvQu9jnIIkcivPvngm+wrxaHpkCphQn3LDL0cZKA+2KOmjohz
lRUT4TcEZI0POEJtVp7qR79fe5hgzOPTVFvIKpM50NeZa6YrAMU3+giFa4krgPGF/rkNo7bybWro
YBi2j0A5di/3oVkj3f7P0Edxh5otG5y5SZ8v38j74pVcPmV5Ok0FYlHxrBLitFF4K1B0ifUrol8o
eGrop/iGtF1XBk+H/UlNw1DQyznYVKsz5zukG+zcYBtDWsV4ubXntBnUZwgtTnZLBn3Ryci/Nq7S
rTd7Hv3u2sg9XyA7QF6b79uAM4j5FP9SxV8gTf3szN0ZxZKjpE0+mAyBrFLBnqUBz8wyWoVoUmIY
t18huRqOce5YpkxXEtCsQisG1kvrrar+8DigoOX85h/jE0DloJs2Mz2b7gMMGsQESYRNuUYySPb6
6VO9nc1RmboeoZzq98BUVP6lNDV9IFwYkOfkJUhKiqd0phyKBgjHDTszMuCxIBtOk0BQizUiqn0X
9qBnEkgYg+9yvtsBBUmT+JG3eBuQYE1Nd6/g+smLtXBwVW447BUuEBxAftaCv+N6iCv8W8sQrwTF
9sV0N90Sa9X8EHxnuDrECo0/s5mZJNsXcR/J/GfRQkQ0h0w2OcvPfXlE5rfa7g6uOzoogQ9OBKwd
cq2tAt1SnHAvySh9DW+CdR8ZwOiaa7j4wa115efkih2O5IKRgGGIPDGA98LfygPtJkxKTQ5zoNAS
LX+yvphWgkrfzZ3G8D+ClKMwbwz5KtJrl5inD/MegrmgSZ/Y3JCOPxOdi7Muq6onlYK7zKee9KVX
9oBAHs61ob/spqa+sXp+CGaPs0cImCttQHxW44L7GgN68uukUgEcjmzjSE4k7S6kNSoPOqcNFj8c
vJaTZFHgFO9UfUyBOro8QAuWgYfP+E2e1BCbqDnLExKS92MoXFCkvrLrt0wlKPROY2ycyg7+IX5p
snqfjUSVK8nQXkJr69pTs9ChJs76hkZPMcxXwSQkixzn7q1XbA0mCO1tCcEKjOtUK2c/3W09ajmk
NhIILI32NdaQUT9Wgq0A0/ZCYmMBtIjuLd2GHj5i/KnKIco/0Lk0N0Qh+TfZuNJR6fdoY/IzKAKQ
hpfvht5liHBbtApDgNz6s1SM66Q65GNmATnZAfprTOZNTb/k4CbwtTvin7Aq17/f5JA7yIVZZjbe
l0zq5+tBn7uUEWqAR4g/r+K+WoYQ2YQAgOC0Vd6NtzKm1BQwlOzKF6c5/rkoKtezYwdKfo3xZ4H7
84OfhPY2EqJSuT3/Ud0kcFfL5yuf5lfQD8o/Eh2XbeQm4CzowB3vFYGcRzgYKVUq/5IVeg4mgWHA
+eKCP0wnQJbbmfBLsW3PhkCkPUyIrp+KLHDzP23DUJs/OrBeY/D7WaVLfuRH/8AOAoTMbJXp4gTj
HeWTTX1H31M1HVJYykQI/P+a+5r82wE1ck3z4irNeiR8MrLzo9kBGUUjSyYvDgU05faQa7olCRx3
q+H9clvBnLuFYgtw7nZcQ8qyU419xEna3/qe6jQlPwZGhjFUbkwXXbaShT8d/T6GotkkOl8s7KIm
6JfEGnHynttmZKFcu2DZGAn3nHWWOwj8KBurBTVCIRQEy5JUEyJsgtGyxaC/p1qLjyuwMsggqFNE
NkgFkYgzaFUDuij8seEuS6vbmoSKaD4DvD2p/+sq50b+mBeXn+IS+rQUw5IHh/CZwEv72gE+O+Cc
4xVoM0MPENhIZs05qUszUHSXwr5wjl5N7NXlMpYRxpWmL4vk6F1Nx7+zOgBvHjVFocGFtRlVrXpJ
I07QgQGkLETBKCXUvw04+u0yHgZN+ShmjjGd28ZXg/rf5yXh6X6LcyKM3Z2rhCbKz9X6Ucl5sQML
K6kq+5ffIU+g7rAPATsRj4yJPa5Oj5A8h62UogNcX4eFK6R27y2KTFTzskMxcwKEg/E4phrMKTRw
thU8+33limCnZUYJDjCR0vKQ5iVlYFEEmaPlHT/Js8+b+oyRqsnfGsz/0e7Ernum+VOqR5BZf+hY
uLizXneMiJzSrtbZbPOK+o0IwUdlE754MJEyyp0BxS4W3sIqeZm3szlW9UoIG9nEP7rIeUgGLAnk
rg6eAvsa1znceipIFoDxdTXqcFdhaih52nAKOvoGNdkyZYzueFlmmQIfRjEfc5k0SSJG/gthi2pK
VTmLuyh0ISs50Dc+8fXw6R902TM0QxoMd4JUBFPTCPlXPBPbBnusAb6tsrDjkQ/opBU/2/0aANnH
VPNq2YjMVHiIp7L6g32qIxJRdtLRuumjzqt3+fIZFfpr4DLSEr5LkWAiA+wxMzghvtI/KfZEDpWF
loqDoj8t0GysmQsZc4YEIanei7PR6+joE1ep2fc0I3RXFOLjWthmE6JQtkNENdFjFxDnkN4hZqYF
k3lQcgSbYHZviBz2HWGR/Jbz4f+x2MYtEUWA4U4r4DhEnbnfOROGetNOdpEaN7fcv7wseZMqSm1f
iYCu+CYMNtwkwmx7vgXEfqbLvMDuk2YvWZthT9TJIbJyETNXmOhfhL3S3He9lnK9l8q0bukp3OEx
cskejLFbgfsWwitHcld+j67rtIOUfU6c7mZaqiXysk+npCamtehDZwpfdfPIRBFz3uV5iBnoDSyc
GBavK9nxjPNun9Y7cP8lEd4GKFmiPj/WtaoZ44BexUwpHMA7Tfc6Pp7bRuibI4lUTwX4NmsjPTKU
uvhw4ApdMKLS4SS9GOGkGl03T8FDEBM9VxrY4uxNeMKDEAbJ83azYr5LZMX8lDEf0DrNV0AVL9KJ
cHP06oKkl35NtYZ/xkbfKMEBZNDtfRDQqQ8POgn1ny0aV/CwywOTWGh7C0qULXKLnhTDpAwiiTRK
JmjcMAUwCmz6A6oTT7PoOVP13USDysYoUkDwB3qhvE6ZXYAfugmhl+RmA0rEU6YRSd/HAmoq994P
pOTsFfbeKKsRb063x4QJMD0S60GQfrQVLV+AjX2mtRP7PlPh4PNyw/XXhEOSZXzWVyMYhDwV5Uwv
QPGZY1vtwTQBWUbUqyMT+j+WFI4DV2sUbvQYyOWZUyB+rPV7N3FNOLZHSMBMNVx5uk8ZuwURmdJ5
HWVMErHo+F8e+/4jvDrzNQ+yzZYsArr/vqL+jA65M8duqvcT+luNj4scYsRxIPlM378untEVxM3b
TLj6/8CIT2PslQ9LXN/42zG0kxo8Q1qc0QYSxNxvVE5igmDpE1SJyxiajZJCz8048o1NwZS2J3pq
LYjXkU4Tk9Gg6Mcl1CdRAVFv1MIx5Zdpr9YsiJBFSgiq0+ws8ho7dCFZTpOXYF5P+6qdCzOgaebN
K+Mw0pJYC949okuvWK+5fq8/mAP5JuIePO5Ezokxcqnt7g3kDB6pH+d6yGnRznUGn3wssll6qnun
7eu8riU8V297x6Kam6t+GHQZ4VoG2LgWg4XBTby+dOfBXJlVn0Xx1lIq+nbpVecFJPulLftZayia
aVMuyXEba/uw69Yo2wRZTSYJGgSZYZY2VGERomAQQBWCNu8KHx9VrufPleuEhZCJeb3bVDTUWzKN
VJDaDiRPHjbnwniAdaxUNifKjq49eLBCqiDJy0b13BLTS/TWL3vM4Oh721AV1pEug357dHHtLfkT
aCrE30ACLbRzQPEQwPe3YtrcPI/6JddTVa1/EvlmbL0zSNH2TZWmUDl5ptSDklesbDDBP5TMzQzk
FJ92zucONfZuO9qK+NnKwJp5nMiBD1ZZTbtdFpoVLR/yFgd445w/rvGgiTwO6G4rlBr7ihfml+IG
D+xPltL41+9QjZG3hMWi/Hj4zUNlLFm5ib2cqIrgIbSwS3Og4kqAQ+yPGcJUGgTJQSygoDE/woq2
V7BfZEEA+IvHnnUkgvSXBIjrjUzDtuekqTq3OrUqVgP+V2vH0JU/eZWu7xhWWU7lXf4MHVuu0btk
lOoqgnrGzgXH9kqmQKsFqn8CPqZLp/O8+4adfeoZScN7Kt9MsENvuJVLtPU3iOZEWuyy/FYL0u3g
+sJUmzHPWSEE3oL7QFX2dFjcczLS44vopKNEs8tI2vXEAmfDh1kzwG69OmzewZeYehHhFFDIx3+3
B8c9+twh+71jLIUWAapZAz6dh75wsSz6rAPKy1mJCZajzoYRuaPyyPTx4tFvKr+HeDfPZlN3RP0r
natclKFrFZkFDNbvSq/HhhL9TMFva4MM+7jdr6rKyfFBrpW4R00K0cXUMqbtthDGyNbIiHeCTLtz
hnSWIEmiwcARtP+BOy3o3GgGZ3PtuTqbuCdY/4o8QY5nH82wS2yE9J1fl3jzZXv1Hg357KS5WPlZ
SLTk+NjxiPgwq+vm7sEPOPY0pCudf3guaNzv82pSBnM/2xasWN4Yoi7Qg6if94leiPNnlA4Q8mS9
iCUcRCpxenZe+9cBoMfYecaLl0fLOTC2iC54DWxk6fIITP6UV0Tt4113UJQrNe4Y7Ls1wDUi6N6k
L0CnvR5+X5PvYev/CU/gO6A+b8TIwZpcNmWF3HgDHdfZ7I1bs0prHXzk98sFqV3/8BxvC8e5kgU1
i7FHLsSA6DnT31/f2bcZb2eYqy621hfPtYZjwolG9jyh5hokr0XXX8EIXfnROzmP9aYfnQSDouhA
WAaSqAwljzE9op7eiSTB2MQVzIg1UATeEt7AhhrrglQ+AJwYmV7pLLH9q7JkO+7FZ3xtCcRgLNvo
lN8DmxU4HNBwtRbJEg0pvSMLSEZLt93BKzQAxytxUOM3YzST8TrhCyG27vNL2oIdj9hRKCnu/pkO
egS2flAkRfHNBg7uwKcCuGHtsATbLc0v7FRa5nXqjUAvBX8nAyPx9mgkazQen8YdhZdod2XP562E
0AEf61Pz75JNNjWnYsGD6KoWFuNP42djsOn76Pw7preE5fNSkAMF8vNvPYITD3vJLyJ4QQYatnsB
2pftMMI/YPxIOBIo1IAsqSRTJ3D0rRxhykp6SzfKR4El5a+OXCanjX+NRbimWXVjjo+zpehhtaqH
vjcA6a/F1h8r6S7rhbkJxcHpWj0eNffwYa45Z3/irZ93SdgsB4S7ZdBExpAHIswbuvcxgVEo4nkp
rKERN3uYDPmCO9eZrHwGf6mFy4tFpyKnt4I4UvKph635YVwGBv8MVWFLS/iZz0qGgV4Xq6vlR0Dw
S7Lbn2afxEq71crqbCbfv82mnU7uqv0zzTvb2tL5w8BwXtHrSzgJo0o2IEOdo3j5hfstXYRK1Sue
ZffZRhsNev9cB00b6Pm/nvxDjYxSlxAMt8qYFAu9qNrruAMxa2FOhaHICEUHS+n1HV/NKQduYgap
13zbQo+5fufONsGAuarGF8ybSMgbjh4xvTUk71AfuYocGzs0lPMZ/rioITAspMlUYztG7Qj/ptas
Irf+WgJEBhVNVElrr896xPhFvUIpuFHWqyV5zMJkXoCTCN5aBReWsFQZMW4QVhujz7HzpucsBxCV
J44ejIpe7RiDr0gI8UIBa4BlTy72QqmraNt+WY90a51ZXWzWJqbEhLk2wea4kqth05o/oFFLY5xz
MvcsGyLuZkFltOVow1lyth8IVlw1m7fMIHYf9RxwjZbH/0HqAFi/gWu1dEOdPRzhZELPtidWpmCk
+q6vEq8JXE/5yqunWaDfYsC+OqFK8d/i4aLmarw40JTFMjV56bylyjLLp+gN/BDo/heOUKj9W2IX
Av8WOE7AeGcFi562Dk92xmwSzYbje5o3UmFI7mM1Fxp7ei4OYmYQfcEriNZcKKr/TuVQeLNjOBcq
idW52VS0vlL1dpy15VFB6tZ3IGB9V5gVkzyh6eBwaYv5ct0YZ7buypkCMntlZBtG65YRGJWkH6Du
dbq3UeHASEicdKdCl5vC+rnjaJGrPTezMmQCL/rThCkfebTFH0ATgzIBbOOwWrxnyunccIcyeCOY
5ku68/JV0Pmi1am7MPoy/akcbS9XyxVvSbRDjZMA0sNXpdJvCNRIc+nDejysFs15JFXmM9OHkLU1
sRHfok7fxdFmlQLPBk0OrrMS5U9paa15GW8tfX4b2gNAkuLKMy1YTp7dj9U9xG84b5ZMBIStsPCq
e199uwuYZ9aFVv0O1G+r6FdZiKr2OsiDBxC4CWz6CjRV4xiElkjJ42wGRHRsy+XNoaaaIr5QbQ64
zlL65B5KNJ34Qdf5dcsNWrvfdNLlAlQ4PkatgeM7PZqyqVhHJ0zCJ40KPm/WSWn33tdytylErb0d
lLxFfSzTPoKf3/bTpNdFMWshL5cNKdRd/VRXHqOVzBZgtAekIDevxZbJVqSh0QYRVOEJDs9OjzOU
FB2B4AdCQZRBe8ylPAC0pR4m0NlHEyKKfpuumJAVmuloeyzrkuQzd+/5UMoz3UpZGxnpaMjXp85c
exwHjl8MxJkoUCWaSg3/1pGNnIfA/vB6unnDS94IyeQ9JlChLSz5+XbdkmfnmkQTwFw3/7jDAtnV
bpajurVJoDC5Dexn5SBTDzJXNBTmRVICB615d6Z6gpqMDS6gvAtP6jo4fmn/xr5E//RwcZPUfBWZ
L7F1N9J2PQkciLm5MZ5Ny4wb52tWz2v4Iz6WBYpaG9sJsTEwdcGTF+c7KsHCVB6RriOZKTMRAg45
GFvWuGplFLWOZjUGOcy2uC2LEvRcRe2NDBeFFmOEjuOcuGfdWkgr1its1a5SotIv/lS5zvjvxRzu
Eqh0uULwcPGlBmm2u11+7a5E9TfbFTG2pFeDb/MN9JHyexEAWs4Zqj5B0kWtv4UbATOyP0qcTZSN
dOoqsRpI0bQ7qL3TjGReGFf7nN8scHfRoqB0YMvP0bdDXsS1U8o+CYWPzF9zeJi8VnFaRIBCHe/h
VMIHJslhMNVPLTeIbC/4fzducTDkYMLlKlHu//NupyKgupFR46HNuZpU4bUiZb7B3cs2Ww+4xqGh
NWpN3teOdfUZb//ftw6deNNdc8zk2LLihbm4wy0jgOngGqWTGTWSQhnUsDDV8egzw8v5l+y5cZnU
iCMzbB70ad9iIBPYZRY6t1shM5CLIGK+tWjOgv3k/tnSbo6F2aF4km77JZJYZ+cWC35tldVjWj5A
c6CEp9B+kU7pwBC430rPetGC0/BZCCRYctNnwLREiYxKcJYrTlSVYHKIUlVt0JLHB4B7l5EC5RzS
oa7aGuzVs9rSqlopxfBk1pSesMruXaOj8gdy9JV5ljkTfMm5I0IVZeAyh5yLep3xIRXJoX514k/t
qCtuwMP3PXiqP20h/Z2p8XlABAL2Lqs4TN9RxGLfdLN8zejO2S1Z2B3o+KVcOXQ+ZJdxnrZzc1ef
zLszyKIBNt/dMulGh5011E7f6Mdbo2GB+2PJUcZXT4SuqgOzUSKwQww+L1Xw76nZKaXp7RmKzA+Q
iUAJlrq5g2wgxRQNESjaY9YwuvmMRe4z2lsT5h0PZGIbPYUYOIz0riIxfB1uOCs0M3T2yxxFRkCS
Pjum0mILV4w7LciSfvsgku9Wvi05v3TDQnxOPfrHSU/EKNWGyzjy135luxcI6FSOGxGb+zoOUgwv
PxGNVzOz4OOanpo2E0OD8rgkynY29sczRlevC99Ghqs0YBpsPMLSnniH07iQUPf/e4wLHYGD36Ab
OT97Wjkl0rTXl8wdbnroKxuaWAt20VmKAGWCRQI96NZNP3tM8l5FF4In4S1TjdcA6vJTkwFWinF0
aHb6XGeDw3DmgBlIpOaFXpie1ER0O9izTW4BhPAgZ/54jdiD72pacgkxrJbFzEc6Wt854eetT9CL
6z67GAegliSP8JvHdEwVN0/YGEr03AHwg8QyDNYwqoatdgEkcbR9NULsv/Qg4olnPN4I9qkaC+nh
8HPNtl4SdejzpyQ0u336fWb/XQbV8BUuubrj2WsnPEWkhsrMyCF3TfqUJ1FYRA5Mq3sWr4jpJuWt
z3xBCBE5DViwEV89NOyNP5pmRp+/wPGRQ7NOikSiVun9dSdU8lx57/QlX9AalzclrHRW28ZcrAmJ
OXoSJuQms3sCdI5Kq++ncyymgumjD4ZMfcnMKT6kqWNBln5nGYAIgm8tW/1PxL6aju2LUh5tZYZQ
vqyX9YwU0iRMpvqOgYOa05Pa2VVGm+IDcWEybqOTNeNbQy5wZunTLFO+9yX/bdjudA407RPuawoh
thuroQJbz12U1fD5tqgoGvHmwSO5+hDHT7w6ydPo+SODzpviswwI0aQ/kkuErxYjDRqfYOsHJ/Bn
mxtbC+OWMV+kvhpnAQAk9TexW9tGIqIEz85Iio6AudRlDKBqwK4br4AygCY5X890+vpmkQMlol75
VYXG1hjvUJUwrEFbjV/Kg84EWpTmYjJSkq3DBGGsSnYAPovrpPDLBRK0iJjwfY/nmAk9Q2COx2sI
f/WAtmnwCYFdckjhoWvvALdiU5xSA7PF+Z3Rca+vW7swJHf0deP/XVu1xhb/KTuZbqThQus3gAA3
HfgNmxBVpxuUCOWgB1Xi2Xi3v8m+J6F3N9Fmax7fsbKuH1wgFx+yYXsxzMC3bYWacX7mZOXtfleb
n8SzsIi/X246ukraIBzcLKa9kWp7Z794hWFUlwoIt7tnjVyilTPoePEOlQyNwrn82Yxks2xoDu3U
lfAtNTLTSbfWvjciKp7Pf43372R5nhPJfmMlQXYNktUe+8DtmI1Ktql/vNscNIuy02SRliTyenxb
thrAXj/vEVBz2fwuQSDmRDxnQ8bpfQOF31CaCD3inueS+sEyugVQIjnAgW2fH+294rm6s0tgs0hR
lkDh5f9C0RjSr/m+oF1kp9Ng7XI1OO2pfMnD6X9MoX12k0M2kd/EzrR//YaBKNNv2QR9qr1ojtZO
wi0DfWSK9bJ+/OEeH7FSKQj8tXavh/Ff3jNXGwSJgFCzgqWujVU/11+/7E7+JG/pVFNqJ5R6yE3F
Au8gMel56DVX3vf1fb4mEjrPdU0T8fRah1p37sIPPufF5RBAq0ON94lPyI+SQits68/HCa5JV7Tt
tXQa9IDkxN+34Dopatkias9ycPkQf03zbzqVNuCWGjMb27i3p3WtTfn30JMyVRsnPKo6m6QADVdV
XMEiSPjRcqjPWanPIH/EjnXfugOoKleb2PcWrzoIT+2aVO8WTfTFejBCdxLTjPBAg/8VHoR2M9ws
BtUsDddFoHqgzqP55MnidZa8PMNUyYowiNmrhTrEsC2bw65cODIiCsp8D2SWVphHjn2GuKbSUifO
Jf0K8c8tP7xHN+lUvcyCH1QPhsMgbCs+tgbGlBkLFN4vgZ0VrA1oxDayibGWWJIblTahQPmlujVq
Kwx6UyNzzPtJk9KmN9CP4+xh0wxjKIFUU91W7eescwo2hdeFFtztAwzQ3rT0UojxRJzbKvLz/jgg
DgMOIkYJaACDTaipW7b5xKn5/rA7wSeuzmSjsS96pCBXg5aLIwiAPM25b/DyPi+E1kcgAbkn+i36
kOzYlYeczgMNUSqHNMJAAZbOIcKdEbPjzRjVNoAXsK112+sm3bjxf9hrcsKoZh892Q0RCBRWDN0X
jVSuWGB+QaUTVjvDaU6MgcqR5mrU/7Qae5BfrgtiL7MKY4F2naNZvwuXS/1nsOLYvvajqh8FeyNn
+H5qlKTG+OiUYf4Ydsx/I6cre9KEK1aAWbWK6Br+30OvMJg+ioZywm0+Qwf2s1xoMW0RN7iTk2gd
9tphGuJhVHhpiqdac+3BOXAsIYXNiB7GSAv03miU0Q1O/mo6Oi0EoeHe4kkzwkJFxUj8sVrYiNYh
KCihZf/0Tv34tBvG24TlfZG2rn/tB/ZW7g7jhml+R6XDyjxcteurxk3Tf1QyRJbhhsALAu2oftPZ
Fm7tU3e29jCRBxzrQWmb38TA2XDmZBa0zNX/FGcPS7Wv1MCIG9W50ZgZAIX/amTwDBUjm4mgEOcO
XJaXw92eD3F97qHjgvkjWOwyQySs+GDEwzmFgcOdYXLOpopgEShH62wIPb/UQb5WWokpAwFPfuef
1ueccAmkLBpkPu3a/qYoBVkTcjBqkqCkxE+XxHbgAJIskJGsq8i0YD6vH4S9dDbypIOMNuM0kslu
AaczG2HzYdwESzd9slmciqMlZYJOCIrkfPITqAGS+XhZOdv1tYO1l9lTg2bfdTEyzQRMJc7tGPA8
z27h1rno4fU5hTnu3rUQ5c7aezkZoqHJqxfSc23nCO3fb7F8qkDPKaVxM4a80l+ynFj6uVraS9aG
HxYpUAdk3MdIX+FxGTzSMJAw38bR8Yt6S+qj1R4zjIUgDVe7pcR/y9UujhtGEiQahdqXs1ojlOY2
5/t5+9xbWgfDRu2xqORV/V2W1Gzi3DBJk+Iz1nzY7P06LWjOkw5sHdKih67R6I620nriOsPf7r1T
foWcIptFvNWeJNjqcLSiGZMCfLR+4a+Fv4r07h857NQCeTMXTUnO+MJR9xscdbMqspP+TUDrCAvU
MsKsRZ3338SDNfJMCIRuDdXGaXPiF6uibuHsdkJcuuPdnQkBhZjh8Kl/S4AcAtrOYkGe2/EJKq1A
SvsXNCX/c3awElu0eQikFlhz68D76glMv/Gt9z0Wm9yr2+1ftTfXhJDzUo5ECDIz+qVA14Rq/R0j
XsSHLRutx9aA4IYCkP0tHHOdHsut9Ibk947WPFLVouTbI/iWlcCC7+31LC+QajC64Dc73KaMXgWM
B6bu7vsoU5THUgyOP4KaoSlKKXBVlrzFqxxODOiWr/Gm/1EI2z55um2eZFWl/QEUBNVGRAbbmOQT
5fn2L8D97xmfiZzQXs0T70aZ8nDudxwkeTF7hhwKlW/qYoZGnj7UD1bOZPset4uIg5dPZCRRv7sB
XICBftMuwpVdJf9zKdXtuKL+Fm7DB0v9EK85L416hfULWQpaF6w1errYgO3WY+HyOf8rs6w+wrA9
TmMlwNDCgEYtcphkIzlEFGSgCvYzeVo9+zm/BxXVmJONAszhllkBNcKTIDA2bYYSagDLJWukeP+8
E9pG+DUyiA4q4GNPJ74476ReQAtWv6g2s3wy1pknyO4deIGGj2fiPHm4irLB2l7Wz/TEV9Q56qWX
8RRZ9RmSNaYdv4GVOXCkySy6m7OlCBzyXGUKtwZu/1ANGs0iwqk6Ced/QMpx30alZTaMvcP5pFKb
GqrpULceq+VRqruXgWJg+Rh4YKAmneFK+jPnaV3a8uhrcxMC2TrcP7gwgTL7MfNncIMmLQze7efv
ANYZxFw1xGDSKM661uh9Na1qZ0mgzRGLT6IzDKAgmk+4okY4pMKim9pN8ItDYrU4XCwVfWGkQ1RT
YedeBoIMD4KNWPq9HaGdQZTzyVmdgQJ5vxTqpP/iSeFD7MzwArwWlHnR68ahpUVEDycntnxwR3Xb
KP9+xca2ExppbQvoZRNSmwNEDWMAByflIbtmfavltlRkPz/xIWiwIG6FjLPNJ+HNbfdoS8BrDxNO
iNyYEyaiiGqKBE9TUdlLKNZSaFMJsjnQBSUFRD0LtZJtxZzjnzzVEiN0iWZ3jHf3J7tCmdFZavkY
d0xIBS6fChoif+w8/xRxaefJfRkJJgO7heU6RvLnX5l0hVF36SCUkkF84++O61T4UNJ/IxgmV5px
3m3Ug83U5HSv9+qnIMQy//NRO4AOZY/d8RAGRcNM3p3+1fZbNvmZ7l7UClaBRtSJWqgAYo0xjOYb
ycLKDSzGRHieh2IhcXUtJy2DQdsjLfLFKgl8foNcq9AX23/uJwvzvXlTWdCcvJGXw4vzugTH0Sg8
rD6PEO9yLOTLKU9GeyP7+G4lYPEM3eV8wPgmCOot/JX03NnZT9gznIha5BKaEmQDpOXFt3F1zWVv
lkyXS6fIcJ80eHfrVevOu8sv5JUg2ysh7s/2f7HgFcG6r0GWwts/04BkFDahBvl7uAefJcEa6jaS
gn1xsdZRWuW4ObQNiA544K6XrIZuiQo10D9M3xB4TJl0k9Ftd/Iu2ZljJkaCkoqJfXVNOGAfZglW
AmnNiompPlpA8ciCS9TSg6aeMekHn9cs5Hk+YKwe2vzpOOgBHevDkR/YszsbFS0yDt3INorkg7OA
tQ2+mS4F++eQC4gIj8tD0ve580T4J5j+k0Qi4sjDDCtDH/kzZ36d/4bTlOvtEazMgWFI/7TIk5Ix
KmtRtl4/mjpNHPL7/otwmdxah7Rd2gDXasT5ckjoYkxJqtBj5L16kZwS1NO4+4dS14yqM37NMh89
HSddL5GDC39b+wMCO9O92mUlZZRgdkmulykzaWs/L/TwIDzjJstPnc7SSfXv0xsGwTyVTA3ziRv3
FzKFOGlQXltUSc04sRE/yQgotY6UGf7i2UPqoBKwYCTXaKGBOiQ1BdZGoA5jCXZRnP6iGv2IURSj
0+OCkIXAv5YJr5eTHfFbAXxT0NduCgdRJAGXpv933oetuoEhdJ83iKBSAujYujdEFK3Tw7Zt/Hz6
TwSGMw1fMQcLnQk6e40OUq3cru+9s5aag/HacT9uI1DQXEETNi1Yh4hO4szHM+aYMtwH996WJvJp
0U2EJQ1sXzQduvwHxsN1fSQrUd83wAlE5DD+AiwjDtchlnXD43/tKbudX16XJB0uwLjyer6hsO1d
9DmYzvyGgdyeR4lhE6owe0Dn8PL5C4Y0nMw6tK36j4kegTHQbpN3cOeDgmLBuYqCWfheVqlkI7Fs
tlrhI19XoYWjM2RtI5zpFlqD7KQl72TFgqXY2eRoK/yD7npJGBbQ7SMRR0Cyek48HfKiG+GGljgv
Dm6dOxovcYDcm36XykqDgMU3Vf+50WfqEwaiKAiOO+0FxNGNwXYXgmhJgO4khO33uvBCBuubL6it
UlnBPVECKFfQ2e6khC6tEJd3gF761BLy7WtZRdYbziprjc05mG+KaVyZqJYOO39/1ngNWRhihw5y
5m/WXCE3gl+KplOBiIue+ba5v+3JTiTK13N2dsnmWJCEiG0exHSneOqfD3pkwmZFYBF4wxDIWpFm
tBpKknQFVl6n8I/LSTRhZ58CoPAVA2CLoLv/sYO1s/ShGqNnW8y/dmEfyTO459AaCeBLvlCD6C7f
axLDUu9e9fn+caMDePuMJvEnRPcYrUpssLT5NbZuuCn1qZZ2E9zmbJ6+UmdD4wx5b/xD1//shQcW
v6Cs0LZAVwbeUSgjp57sVOdFoqRMGRn2v0sMThsU3LBZAkzY9FqTMx4prfKaZ27Crn7C2xXPvnes
M2QL4FhMOwi04e7JqBF1rELc0WfA7O7GKsKob/iQ0z+juweJW0y7PZTnXOsdvoCMHsEniDIfa/C2
zs51YNkOsKxWEt/gSepmubKkcEVDOjwnW11MUG/FWrhJqw4uPFjljq1jZbXXp2d/frBacWuwkjiq
ZvxxTV/m2Bz99Bz5BvvGEWkLSFFFSHrhBGWIr1LYdfW7iQ2aRfwhGVThhwOxy39N/RLqkpAtD+VH
4XbAHIR9HlOzXJyyKtqxhnlttqJ5a0Nuc3d2rGpisguuqEB2K2WZaqgM4oNOX6+Tp174JIKPhOq3
yYKss4vq4bHmUM/g8KNewZ/SEwu9xWXEB0UYzeXKj1qX4sDRgXBiYMAzthI60Ip/GE+JoVmg5hB9
dSIABRsKSSS2kYEZHj5OVohNUFpEmQNVYGz3jEfHsFFtxz3PPQ33F8FGd6eGQ8isFFBtA6rZQUgV
oz7a4uxQFY/JbnXiE2j5lFYOXYZo2UqPI8p8xlia9HTS7rdisEwc1Ek9yGg9D9ENNKB66iAGfft8
JYSPgEdr6nDSakHh65JP6wxwx1iATutvSEplN9yTy5kBlhSpbb++znJ5HKxDU8GlJwQsTSyHIDOi
OFQm0bXhc3uVavFKagNTi+Xt1NJQV6LqeZRy+N549l01eu+lY3sRPWEYPh97ktj7rVVQck9jtyuq
40vod/2IEuo0Vq3RWIq0OefPBt7hEdGzRMFpmzPwGdc611mw8IMKquQdKeKc5g9ftzN1eQsXX8xc
J3gyLMIAFzBvBYS4Q0IJVmDvSATmwnGuNS6t3pe6lSYVd+gJqwK+uDefdhVj2ckzp/2yb8FoFlHZ
QLfEoqaDkIefjeKoruRyWYAApMgarp3JhJzrmVB2M+p73M5/HHtiXRCnGAYqMiW3oGP2kl0ZxYyh
OvWsNcUQDNjzUQQNwWpXecTz/9RsCLhDQ9C0NMnFhunx8qbCw7zWqAjI1W1CXZlbH6Ehq+kYKioC
yoGdwQ1JWZ4xDLqmxdRY/ITxR8BYhZi+23Q9B7w2ZRuGBrds9Vh9H97uItkcJHgKs+Dzb8zuvzJI
GvpsEd9Nu5qScibDKcZaMBj+sAivsX/r33zKLjH7jQBSKjrtPpbeWT6D+LtOxWuj8/PD60CGUw3W
H9w4wgfvkcgwCDR4wxBU+RPLWAhVSQ4Rdpl29uZ2dbaXQy3jLAJzXeKX54wETR197ZzMf88k4OMR
0NEplotavjMT32vwrzeMvVSf6ngIyk+eokWOzGC04PugIozIbVW96B8i8picPHKaJIzlD2X3RR+K
CMO4KF2j/XQpmEtWwfnsFIW6+qyjswRI7pT35pTsh8vaWBNXiScCZJRRzfjwPGnM43D6nATOlSrU
AHhmq1dFJ/7mEMZ6FkllUwzauiL8fDvsIxVJeIWHsVpmyuq66xgZb71FuO72bRv1F0/jph/eTgiM
Cp7XF0X0ZSjz4h7opNjn2LMsmoFF6b4DzMr2uwCcaUkQL3WrZrUTlyvcb8XoX6B0qpETs9YqayBV
10t+Z2gZCrstVg7eP10Z/KyCHTo88KQbqHCEYNjjod15dvRwdw5AAxRgtxNRT1uSLdozvxIUesp7
mcoDtG9aYqcBYJi9Gmqrz76mbja7KPpsN7MLpv5s3yk+wBSc8OQNi57Grbk7tB5+uFKFRVFb/kLy
NzWE+KlB38dXKREPX8qz8u0/YVq9a1XZACuFCBGNGcyC6vOz38uh1a4hvV36wj554uL9+qvm5mu6
G39UsyjPOtINMyRpBJkpqfSHsReXr16th5WVZri6h8jB//2vq60t/3rqd6QDutsWc+cUboO/pxS6
Zm75Z9sY977eWn8Ew3ZeJ7e1gMDccuxjKip+fpHevSEWk0dK6QHb0Hhe4wBCTpSLZmLrjcNilv5g
vOhBrxRMbGachNHGpdvTho/0fIxMdVUlG/CxJOGgt8wsfZS5T3YdN0urPunj4OsYg8HI2gkrKZs+
COy2ZcbwH+xJR0x1B+th9K9oL3Q8Bf7b22pT/PMdhceK78PeaUaOFQ4VO7EuZz8bVjoXJHK6xg87
otF0l3ucY9KtwgO8yCTh2JntWUQd7JlOfmCq/+SabAHOud0icfLh5y6wSjbCpen6R9PobCHCVpic
qGOgQ99lvsCGoXfPTt1Rj9a7J0VDhhAjtJLdo1YAfTzG4//GC8ys86pZf9eZSSEo57ECsedLtBLC
3rwTI9dX0B2LcfZdiI18s3m/dabwiLa+XNOCEcFFKsR4E+AVO1FjvOO8RSkj2sGMvdYIFufd8BOR
dAHZPzci/gN4Q6XcXODtsn0/2Z7+3CdT8yAiU/2MOC9/HcceQVI0twpF/Rbcbu6vCiaxUSc9ts31
EoneGDfyf3cv/CStOCbbu/pNYkdcPaFk7mPdpMa4UPCDP1JtbXGXR0c7lhfNvAhUcxnfvjQbm+MZ
JR7OChzpoUlA0t0AKNNVz9z14+QxT9VNgtsmGJ9QM5Vkx87kvmORmJsrHJryIU8xGJfz2OeozZgP
+zwC26uyhU3T/W0bVwJayFdvz4dHCrAts9lALs4pv/4XeEin4Rnw+AANmS38JZ03c3JPXLy59QGc
65FZp1MdX8QKvZ8tVSxi6Z3RXbXjhEwFPCmFGqZ8+MFH7VD94OSzRoOLDqm+445sX7RIPaeQw+yU
rkjm/r+e91vyts8ppuo1f+EJrEEg9OeCAUt7HXi8ZmHyd8Yo1nPRFLZJ9eY2VnRvmv1ABoXfOZWX
0893IGsfrP/P34xs04u6rsVbpu2veMQS0zMrUqYl/Sy8D0glL+mj8S/wHdGcWvYctTLabSF+oq2P
EqJPQ+iPTlSvl5l4lmG0yub8eGjDJQJgOFPHZcZOHqxNv5zMbyswBIaF60YOZpq2cHe+I8mymB18
0ff+tFz5+EKocCLRUNGQUHZPy9VKfXtiQMzvNl2HlOT8ZlHzVHuWZ31EaxKVCcB5IiT89/rLwHrt
CyHAiIgwdOOLJ6dpdMO0vif+L31fBPdpZ4fkVTEejguuJty56hPTS5Uargb9CRH0QN/2axBI4Chb
UFe07tHBRuVv3oSWOJoMHFqSs/a9dgH2PrXAdoRWmiNCiPD60TbxDzapIp7TBs5e506a+0D2KTzS
4Phl6gC0kTQqoku/TTdlOMuym1Lq8qj4pCcY0Lfryav1D8YSgDOSV4qiwUvpQBnwmO29Z79A/krR
43JNSwmX9DPmbzWuTalp05YhxkCoDHBVUld57w1EaR7bEPCWcxrvOPJkaXWEdl5fC2ot1q2rbA2B
qQZS8aVmEzSlAn4eEiwVLUySH8jDRy3//qY2XO2yZgAElc1tCJdd5LBEa4/EbFSs8EtbbdhNFnVh
pHoAN4b5Wj0Da1fY9PiENyXqQ0X1AZGVWxzni77tt02cxz14e4mKtT2qs9XWze22eQ9G3X43tRD+
j9LpnTuV/w+KkpRs5Rh+0mF86qs5Y/N7NyVWKYx+wRy+uXj730MlAKSFwLJOtOlhHJlWM8C7Et8p
mvyit8n5pfNPPJT74TewqekfOlE4/SG4GDjhsGvspeXUtHlG6vgnJbPcEFUjCZHtIICOwlOWlrSK
GgXjM2HIluSviwHg1iYowIyB7A+Fg6BPWSZdu5zrQf2kXUPFCL98fsme6550Y+B5T2N5+tc+OqCK
pOgMWMgcew1hi/MjDZ+iua+sxu0LhsYVULVpj9TLCTocBFAuN3pGL1vnvOG0ldTqefezl26HmF8K
53vyUH6IqNEUznjiOur/yBDCbYxdbQHJhzshZgINbCet844nbifQbrthYx782m5KlYKrMFh7s5Iq
AOMzERjz76qs0zZ037WxdYPw4w3VYYdJX/U6TSQMb3taEScZnpZ7Y5Pkbh7CiRgFWEk6MBUWuz1Q
6dTm+bacu029e8MYHgL6cwIJeeRaNrUKS1/SG3K0pmFbj4IWMqP3vpR5gRnvwFbO5rL3M3CEKtos
2l7HdsCjXxN0ccGxsyMaLo6WcqTEM8R2JLabNhmhajSqYqT1751wJBjXY74flx/YRyqiyoWcxfK4
rYehV/1yY+6VPN6MKB1oAMdesekIa+qKRvleSbBx8RqRgTkYhH3sOTwL2b2c4EmvLHFT3AT7nEmn
ePAdDsRh7TNTIVClIEgf4IauJO/1MK2dhee37uYUdIvv3vuTRPIWfSwKO93WxHOERycKHzOYD+ed
XCdYHo80X/UZARRPjiBbl/u9jQCmJ96d1x99nOYeM5FhYa33HwgCl7s1RqqjBDHhWWg8UhPihICS
B82OiD+AsAzKUxd2tJdMiXbiBGhBEB90hqCoLt+pNZeDSktMP9h0ZWPhSvyAhLsiSnpXRWIxVRHT
3N8a9ds+GwlXfgrH/4ePRRJv4I/UCmdjYdmsd3Vp7ZpCwhWxrOsL3AhiwcVe5yifoU7JqphXhUbT
BUWe5lZxOeCA9JHIu3QKkzlFVAm5heXgN2uj4um2RC7YgajJY9fbMbodsM97aJFQ5TC5+rol6lRq
0cbK6//oz1cXwNojc/5zUHwCRmM+BBgWs2j+uTycqx0uAGn0ec3OTxDwiZJVOAmLLKiHuQTY7Uh1
r0LmLL0LdGuUYwk5coD75h/LhQh/fqeEo0Rf0B0ZZklwk860G3+NhqC6/Kg84lJujiaUq/f2BVL2
3RecNfxBoU/Kdhe7TQe7ODgDcciRmqP96G3bX3c/ZSAg48uAttOfjiwZtnNyCu0S9p90W66iqqWo
UV9JMqkARiY8/gkeP4T/jaftcybfpjfLAFfUbIgrD448E8fqyV0S+pKHeQzOj6DYrdZaS5p9qH/d
qqWFF2PF1hPuUyAYK2f3FJ16RYtcrs3X9BrKXHixiUj0a2pO2tXIsgeZzpGOJ5eHhPwP9YqXl6xX
v0y4nyKIozsKJ4OMJAs+nsRIS7s+y/T7AR+J1aGaChh76VU/Z9ZFCX4uTIqcwtpv6NAHNEeqJPt0
WokGczzBIPYrmCT7llPiF5leakTAWr1rAEFpUO1NwLd+3ICdgMnT/oRToGrNs0WW1iFX15bfO8tq
WawJ9c1BaB/lSxDocMbadQDBxfOypwkBMDgZknFLD6Y+JoVZR3C0Kqi9Fgsh0oEK+od8SryoHKy3
GT/z52IV14rCYk9vuB4UszJT9ZKjZ83/nwwVpNdd+jpD1uUjN3U7wjLtk3VKpxODRT/Tp4QGQceA
rMSuhJ42PaH2Y1OqZZAV3Tj2UdM1kMgTFMeY6tt/SxHhI5XF831hGeiF/cbV9fD/MLIWl/v56igP
NRVKqO/z3ydl8WWIrtCSkTNk9BiS5/GsREF5JU1umYFRTv9mgVLrmP/N0AkOLslhM4lDt9ckJwdO
MtEZMffZ1BOXlzV36/M8QnMWgA+lmchQLs7O8hIr9+MnCJxPRqzN6ykJqn0W2v1CI7+0YIk6WwDE
Hc8xfSfMQUE8axwJTcnW+5OHWXyDyqjHulaBluNPkgxeyCJtswQniiUNdOyAe2AGdiZqEWznqKZD
i23x3gjMbjD2LUa+pLmpVwLrgoBvg3ViIoV5T4LX9o7w5VpWp9+ElPVEwmT2unu3yAOxgXPU9INf
BlYigUNAStREdcIB3aljo0gX4r8+yrFffN4SPY08S9tVPGGpPQD8rjkUEcVyRy/GA3l4PmX3sj8E
eGvFYcH08yp7RzrPqcMuFXbBFXrsFzsYLsrlOjrLLYtP4tDI+/rHUvo5pOsJNONNSdwpscd7Sqx2
JSrnIGcizSUXn/kv1Wi2qT9I+TUnu5/6gOSNbNk6/eu5KdqDcT8Q3mhCnKwXoVtNKKuiC4GwkiSz
8k2k+cY6gwgUWIKr9K/w7bhu/we7HCx5bshmX4S3brPytegaKzxUPnI9+RMd9C+7H0y/KSj09P/J
7sBinWGvEEHNSTBOTOo+1lz/I1ASeLzBjCXbrBudm79vZ9EAxP7NggPDTFtfH/7Mo9E4aMn73t/4
I98iOEehaKtQ6evTdOVRV7Z8mg+4QE7EgITRuhJ4hsoUk/0dDooQrg3XZAHlrj4lWK6/y4pstsvv
h/Iz4N1JHPub4TmX25mErenibJVxFO3GGuZXsAG3qfKxben7Iw+QzYxTs3yTh4zEYRFGp8WYGjhE
LhQ+zQmpip82xgQ3AZiqxxBvwI03AdOzaqt8tXX8okbDVK/uE4kiZEfn25FWZl3x/dunf+N05BHK
+DxA3VKoXGzfhTPDfNevJljtRVqYvB2AVIJnST/QbjQO2fV1oPN3VXUhAK6ZjVQ1xIiMLBdIoSYe
WEJNpJd39wFg0VHAgGjlc/RRCHlEsa/yXSIrTDruvHPFhFAFUXTfqtrBDUSULxHrAi2U3Xdf5srG
21rGzre+pIB/e6KaQBEd47p9VytrA46OLDtLSxC0gRyM+hpz2yzqPNiu1dbEUb8ucYgj/AjHrAhh
X7p/hUXdBwyPG2idzMvcgk3768i+whznueUUkiXZecvFFINBEbYFUBxorp+HbIed9lVXVeqyoSvD
5wUeqAfAd+Hdy5uLQ0phUIkik+Fu5zSPthUCLU1i/s5v16lTJomv8KT9kRB6SOCmiP8WlEpQSOM3
jqjSwkrHn1Qbuei358epvjdnpka5dtwUBVgVmND6KuOSDMU4bsYZy9pi83xpbBa6AeL2sDZ9DsWH
33+kOZssuxLR+wPgKSwyQh74YwdtH9bGJ4qA6dbCeNoIWeTKU7SRKBMQ8D3zW7XOYNRbb9sSTxba
emp6YuOVzKxm4v5TSNBowrU+NAdy0v4ReIDLgLAJZZGzpqt3MEpBLCrs5YaCZoGPfAXa9KhQJZOj
L/G5bLvHj3z8MGRxQAHUQt+Hp3coj1Vz00J54Xz0Shuou8Cd40dUIs+DkYykdox3Zk2Sccoy++HU
i8grnATYc/c7MdX9BDizkGc9VjqOqrzU7GzYPzbmD6N0T4kwUe1/vTr0cVza2oRYZiEA3Ymt4RCe
/zupsHgZvgDKfl+r3PdZXkMMv+A3udHDzD/9MrO5wE7GvJpX/LPQjt64kjXiPsoeEFM8v9TrAK3e
hadyn906ASPP4bwJDlBqd8tqPv2wrlTPEux0XuG+Q2dhFE2yYzKZeinaCXEWJs2IZ7b5VBV0HCxd
+uLINRXOXCUHDFgtrKFNTC2gphey9AguXWgRoTEm1A1uQKCg4aGVKvZ8mCnmWr2iNAIP8M5mw4SF
/gqptXtngTr2hdk5cSQUDtUn4r35cpO2R2PokfUIQQDbwGkRmPyaA9NFwBGEGKfy7bhBssKTUrEF
bZpefjwyRzaYTmjMp0XHGDyGu2L6xUx+7g3A1LMAQQa6Bk7ydksbVIO2x1OB8Bfm7F6CIVgd3T7X
uUllFXMbMO7X/ZOVNAcqnR2AKEnqdlDl3nyq2eT6NjqE8znD937J9SZ/k+ZcDaZl5MdkOg7reOgT
xSTuA44LvL+nDoNemgVHfE8UZa9zwjQ1gMrWRUhxOjXjOv/pT6fSGpuevx91U6cWZVemfHTRHN/V
zc4vxdxMc2KUmEPtHf4jIWMOlZG0ZSScdeedW4S4Jz+IQBBVW1L5VVonIvOF/ZQEwlmkYqwx2t9f
qG8ZAVgo6jvJ3YHPvDRkjWUc1ebpy/5V2aKIxxMk7UpIxU1WKtaE0HCNqHlA2lx6qNqvxoOjZye6
UHwXmQrdNiQ6YhYFY3hEab9syZTYv2svV2gSspr14nGgo0vZgCx5KQrRcm2eJ8Mls/+fLu1fRhkE
oTa8a0TBTCqtLOeNctT5Vn731mjxqNIqd76uk1ZjnD/dUJc5he/ou/d12NSd7IuAkghZinGF8YC7
2QBVvQ8B+agN2PIoZ7nwk7tiXgIcaxDQlGCnGphN9riypm1yb7JiuXUmbM8YH8Joc2cZ6Kg1lfwS
uBrlrUS4a/1trUsFnL7UBNuUOd3ev+n/BVyOeQZpI2730t6lM98wXRJvRi9VFITyhiB0FAnNLLqv
ypJcYvM/qSGkwbCDdO1/8wtr5bVlHBrCo50vsx0JbuzZgtuOvfHk9g+uXj0KPKH1ya/xGOznB8bX
FYpo3zrBX1zOtlST0n4DjlKIbso82rIeJiTigXJo+UDp9BXT74VKbJYXc0eni95OwdgNkA3ED1ke
yMB+SpmUhwfydlazafJ4rU394CI11Pj9ThpP3j+gUVvLwoHakhhXY08GI8CVRemjxyasGwVi793g
aLOak5DVBC+cYKqdhWDKXEnW1X4rKVniiBwfQ+9mumSUhe2+EsH/ndNKuW1xbEhBx/8o/mNtwD9B
taXEpSi4V/UgXpdvXT4OcQ1RtCzTpjmZ54qiYJVLw+B/tEwuqe/fpfcyXR98QakVjrhMmy8T1uSr
MO4BsbkaMnr1SN5teMcxMbkuysBrfWxpP89n56U8/ESeLrG8LHBn2XqTE85PIW2yxzxEsqnxEVkE
2wALGvqT5cHQO0qqGqezANSP1c+CQ35iuL3nj6lZSZSIRrfKj+4LCRQo++xjEb9mwpnZAwew8I82
osZMyUk9F49aiIYeTEi8OSCubSUuRoB4xXubV+M4eqAt5KKAzW3BPi1DArvVUbiXZxDkXgKTJPtF
fhk/gUPHLDBomLdDJqdq143wO6Nl/1tieu6H5TW0f5yGi+QMcu6WsTOM73fqsEjfjKjWFo7G3GCw
DJzSC95AYlEfJS0iKpcERMVsS2z10WqseNMMRAhPoJqt/A6bEB79ylB1eBOXGkzmy2MIqjiMZKIy
kL4TIuJDQnRFZr1seBn3+rnSvxaD+AW6SR2tTe9XiFb3sEohzZ7mfKz0URoa26+3FvQ5HpSMnhob
nfcvYngQoAfjVuTLJ/sfu4sinpf6AoQSHH3P8DbQpLLRi59Dbc4FErQlmJkthqr6+f3UkrglOxFf
5Lg8J0wcDatqrRj02UDS3m6tSslWXjxJxgdsl/Rq/mxWAacw0sddK5EEvSmGmbnSGe40OhzvM1Yl
u0rPtDHffwl3O7Kboa4sYhOdqE2CHF0Rhh4Oa3L7OYSRmUt6VVOdmb0+y9Tb2Dex/yBYEM1SNRtD
SYHrksTy21rbNPWSgtbNnlGTGJhTn4VUl9YStpU0o+yhGx+Qd/BZDNqf0ec9XIJC/IjIEb4TG+bA
QC+4UN2ZTvehs7zhwB4BioyfRYt5fR0Dg6xzjJ2gRH3VE+0okfVrrLYrOosPJVUAsgdSq/EzY7bD
ian5HQlcPe4iTsnGZCaaPRqbt0UwxP0dbJqYMKMaOyo/X4BYVa2ULTCDDzc/iq2cVfd6ijO1IyWl
tSj2gBQcG6tmcggH9xD3m4rdMwRXtaOUyuI8G5MBE5f3z/POqMXAhmAGU438IrcKvjfaROl6ua1N
qSmS5nplbeqSReLlXrida1YNl7j8XaHXFmH4nB13y/y1/nMp8of2G2T+jb0BmtFDjxyR7D5hf+ao
bK6JGeGzkCjFCKIsjxWQYEGMuSN8R2lZgIqdAjVsdQo3UDWCI1539SxXVMV573Ug1c0TdrDsW+Ix
dOQKXGrcfPKiMzexLjvwLmb+1yY8XRx6rojDyvZL86OFZb//8JLoJtJwGvgKdvLqKER2ppYgbsA3
HR5KuC+/TRVzfCeLPnuI7P0wR8+zasbEaVAEoWzgs3IBXAqKLIPCNV3ofv89CGAF3ETAkIpg7yGX
j+7cZNbIuTtFfEe0hEYzgLQvwLF50g2UJyKj4mtYidGraq85nDPvfbTzNywlnZOtbT7NAgbV2lqi
vdFSdp7nYwu1/55akzSY4qkhvN4UwFFikHQrejNDtSAk6XB9R2C+WYRjhzzEMInTgUR7YU0IhHpQ
QDajvpUN3PhnxvymVVKcl4ZMpDihgmViIvOa32wJ+VRR6jAoViACcBRBN53+oPBNWL3YvgUGEyFR
voDbl+JOkUxwATk7LjC9yrAVHcUZrra8l1f3zQ9i2/bDC8Uq2IXe2LdSaLDhqopy0BXJ0MXAGgO3
Z15LHG9fVChwrTQHgYCtwA62B1FiGJk3/0SvhRGfx7gJjoS/9fZcGQRXZWhd4OqmEJzxAVuyuuPz
ShTqfW5bvi/hmyTNFFP25DrmOB+MzLa1ONZ6edWg9DV7kSQl1WH/QowfRw/EYOYFU/dajkjZECda
s84Zo/MRkfB4gp2hVxhqQCIihYhEpnVlnu1J7E1zKzb5fsBQqJcsJVFs8XCirvXb9fYQNaVN0kS1
GxmxY9HDO55VnOVzPjI6GTuHotRWEzkq8VjNi3aLEoY1KPbo4R6Xyrl7SkHFwyQ44U6fTFLL9StN
+A7rTDDENykjw1rUXmfmMF8fZ9mOuFDV6IknEWW43pAp0vYj6eJgvPPKMF0Dxz3605DEigSjgduA
ykVDL//UP2dIjaHlVEggb6JeqPOd0i1RgkIybTCZf6qtsaZ9cHayHQRwj+ZUp+yeK60MerCsQR0Y
EcltV9mqHMcQR+7nT+ygEatoZBYH58ScpS37gcYDLz5dDY90NNNie4UFp5C07XmxwohizpyteMf9
EaLYTa5U60t+j87e9PTVidBMHRyXXzIwu+vRYl4yNKjojrolppLHvxPUXQ83zkizq28SckLkYdPW
E2v5CcZksRikwpGZaCxeZF/5o8O5IF0OXBaKTPKtdvxZjvxxZcWv0WLW9LSY4CdyIyGAjgNo/gyq
9riqjCicy51uEqAFK3qnjCRvuF9NA10zFoWgAUrHHH88D/wgMGxJsuN+dVaMQC5+lNFiS5ec+RP7
lAPxov7/kGrxXFhuwpDniSi5z40+oftAij7USHjntflNMyrM2LH35tLzYiY7zq7JC8XdszrXGHy+
iO9l1oRw55jhqevE5okP5j2vC2C+IoA6deUYru1rAc99mUhwA21TVu5w29f5/SsIPldVTsOnMbh2
lXp/YxILjmQ/rypTmmHMLL3eWwiY60F5ZrmDoS+1RkptZCTxhbRs3eEaJKwp5yH8oaMqFmqGGHhD
NCYSqyy9SllAp9x6GfkQ6MtMQdK876ddvKjc5lRug0ffFgr+g2xbJlYe4Pv4pDWTAYLXiOjTfLN+
S+9MUB5/FA06vG1XVMNpEw9fVV4AlRnaLcZwluTuPlV5wB98bNMLBYPnNnI/7GYvajTJOuNavkLl
u1s3BYuMaWPiu1pOFCo4Kgi+XaC1RE8O3ooS241sfA3JOHjTwSgphy6qonLdlIw4fqSECHopzEOq
p1u8iEW3s5hRPTewJFA88SXf+jnMtT3pwNW2UcFoD/vG7bSEMqLGLLtUMgoCNRmz8OqxO9LYLM+w
JPUp80SK/y7PBG9ct7Vq5vBlRyDHv0MqCOvEJCq5UOPMqexlHFMIL/B+55AEI4zPNcnjTEye3lrU
tRjQklyzuzOPplxXoNS4nORCcLilgP53Ex5PlBPow9dH0zkC15Z6ZWqJPs66/kKHinG3omnPgBje
RZGcFfN2sYWq0lRkribtkuNd8G4gt/t+699r0Oa5XtJUci7tVxHKEmin06I8bcjv/4aQ5RNK1baX
RzrA7n6sQ/Rd4CnezOFtNx3uHgnhbhjfeuNrnflRRMZakaaJXvAR+7XEaUEX2SdaMppau9JLx9T7
ulYHeKacrDOPXiwaEwP3FC4GeuqJKZz0gavFj1f9MtxsqndrHeHQQ9JlrYGLd8eDsb+IJcSYozCE
vif18M8XGfo/F6IT9GGxvozsVJDi6vCOK7DJ0MHhyUVULM2C1lJjyrp3cpBWMpwaKr1MjziNfz8S
xwETzCOqevFi9Ny3qSxiFmTS0unieYqWY3gP1W7otqm4W18c1AfFtA/0K5LMdRig96Rhwjzy5grC
+OwrW2IxwyBZRqGKjbgr2gXilGpLH/M7lfWyTYDXGG8i08+wQzBq6XUMQv+3Qj2cbbsw5qqHDzbO
MdayWUktXFUuC4Le1N7qv3aYHkxpIHccXsLPuGj9rljV04yKg8aPTzUcyG8ASpaTPgoLy36MfrI9
nbOT1yYRroOO0wA+WZOEXctUnk93/T1vRpR4XUVz+Z82+YQgcwKVRbO3tujA45u6/DvP0As+BS0G
yoeM0RuG27Nt/Aa8NzTE2kTkf9FQxXmQ/2U6qV9EQLwHKG4VmhPPjUzU/lLNt9/X5/OksP/SNQsg
jZm6laKg4d+sT4Iwp8ECouULY4r3vGfx6AvcQM6nXA4yS+JjAAYEXO3+O4yi5SnwwDKWjPVcNR+W
+RSSx3I2ALVkpQhUdy+mltzq4p/5jE9fCBe+gLrG91bNmLx3Ty04om9ttcXbYjZHVeS/ItgTkICj
BbUrn5wNXVp6aPKYrqkVZjf4E6/lGB6F3gjOuuJVFsyG57Zvw2ojzdEUJK1FEIG4TV3IM9dxrweH
4zOCGyH9cFvZx3OsGZMuVUhRT9G1jAVDG3S5NlZKYKrIsVw31lGtRBSG9IWlsZ3xk66Yf2DHmnBn
VVqN/Vv2bi85h+yabppJVczogPNvprQs1J0YIUqP9VDqeX7WvzIE0RXsFelNUdNhqE+mRb/k687L
1thxI0l2S1BT1eOaHXo/mzw5g3aCeZ+IeCrjFykUqpaX5MBRreUKcYbG6hEUC9dGyh3zoQyl503g
lXYCBztJAXEv0ONwa/H/hpgUf3Zf7GS2MNgE16eo+vQzRfesSdimS6LqhZJcFbJqmYFOhChPtBxL
od7YJWz5VxsS/P9x1VvN7Z5K39eyGEDjftc5LphdryrEJg0LvYW1T7EXcoxNcLKQcuROObWQzepA
PAJZ+e1jZseuW6Io77hmcGaSqRcgg8HfxIooDQO9qwvVAZejoTcVg1evwU4BSz62xJmB17+mKiOV
JUsb4K4Yd8FfBbQtW/4yydN2pCDiQjO9dghVj4yRooOID3xqjB11LVkliV8ivybSz1HClFMYnSbk
+q4tr2UVii3qo2/lmNSWkh5wd2mbTSqP9jezDqzXmnSH2TdlzOD5rGHZkhCJyGE2OQCE6enJnzTR
AftRnGezO6kW7h6GVI4EB9xuEdnFC8IOpmXPCzvqvrFHAnRK3xYNUDq7mMqDWkPf6t76HeWazOq6
ZbU+dhG3NZSe8lvtJksO9i/i5Cx3+eTLg02851cHMyQGszJOfgwmojpAwm2loBXKyyu4ucQhEi4n
LpVmVLrNBhF7situhR3amddfl5405ZBATuwhEnQsmmxltm9SbXDGwDjUtndCFoFVcczB0DwJskoS
F51DWR/0QyU5trfjecG0nK8Ol6TmU5p4Fvint5ehrfnD11WHFge1awsjlZdDFptTDsEJr46y5yKD
Z1AJiRit/gPPgqCetyEAyOHPozj/GYESBiO/cwzOh6IFPMyaaTDV/RiZ+7HiuQkbbnklMADngVOE
m1NIc3+i9GcKYyDVPOh4EfnqxSU0LXnBmw/U/Uafdnitr/9aVeKlkxRZLmFUVGy4MruuRc6YxAVV
pyTWILGEvjH6FnHoyvzMiiRm7lSy+9YksQGcUVUrNnHNiqOI5ZxK0bTFHbF8QewrvSBcAPnd6fEX
3VT+rzXmIwlaphK+xReVwmyaIEicPkJqBPgWgnkI4VUfJy4Fl296qjvdrnwuREHBaGHENGNdSvvt
csQlMtmnoP8PeWYsL5Czj+rG9y6OFHcQHD6KkVtRjkOhW8zfqsdJ70JL1c/jmfJS+WluoYrtyE0+
dvABJ3CFswkXWhmS+DYstAP7jPcQ42JaKmrmk6Dms09OxfL2ONWk1XlD1SE1stxRASkFzipgqxhi
/ziW4tB0yJfGhWVMB+YCH9wVPBl78lEW60Vfez7rKWvls4Z0ZfHDbsrlUR+ABKPEuo5nDglsCElP
tCpwhGwNLm+pmQk4J2VZDccXiDdEILUUyxXBPH+hr5XvDfULHufMyFlu0Z4gwOBAU59hhgPnUwZH
2WOr3Wa2Cakhv9Izr25cfnbaNRJz369UOhId+VNuBQne7o+SrrrVEDfFJLqhlOLI/PkA7M++/nJ3
tlnH5I99DaNB7N0EEUorn/Z9uAUhRXXE564eDBPGcM2o5c1Rf0ZLdSKUXu7vvBZIeQJvtI/UUutE
BCChouj6ux+mZONp+aaZcWAKsJFPy2VDO9TsKliAj7xcaaiAuNlHbs4BX09gJZLL9l3oLM/bZxLd
jXFG8hBLcxEKxzWdUszHP4UFa4QDG2CGy3OHgE7WpOq8XxGN+E3KpFxlXWgA96l1o1FLwvtSA+k0
mkrR4pAwB9p0GEJkHMS3Sxo7V7JcaLFdrWdTRauRjDMqjeJkU0zS3aG2FPI+sqmoNzbD21X4sW5B
sINfZWGFFWwVE6o5gDaCy6/V17hipklNueJbx5j4daW6D6ZlGaR9Eg8DjtuChthtJdwgsayP8Cyi
5ENXoeOueJVhxqlBdpq3IRhvW/Exvazl6NpGKqn6KiMnXOWL4INDn8K17+HMaRmWgjf/NdxqQHWl
m21CNXg0WjG9PSPmkN3pqZZNK8y6zSRXKp4GLL/rJBZIFcHRCxwfv/dgRpVGAf7L/+A2Xr3BcFIa
omv5lorHQqfMSUgpBPiGUuRcTVTochq97ARwXv/iBu/6+GvZ0xJ/PE0FDqlirSGH6MkiEpXRfnJt
QTwwj500CCNt+7GdLwxV1hbci/20+JlI8BdH+Li3JZOt/Cz05LSf5QsDcnsGWt/j5qbYRrdBsWQl
RlYOG9VuwxXZHMvW/Jtcj1//zEdvK8HF/LMDM6XHvcj7HOYpoydnoeH4JWElxq2SstUCGtwT9Iuw
cQDkY+F30OBwgGUZbQ0ge88kdz7LoADiebh2EZKoebWELKlNEM9/PuYY6GRkjr1Fk6S9cRc3gIWm
AZsoxP8lw7lHe5f3p/md3vMC24WGCLGPUXG9pMZte6GIqcmICyxeDuF0vQn4Qm9QotPLIX4SJ8tC
SFLLHLvS2VHvpuOWlePG9TqxPN+AcRQokYUXk1lNpqyN8+TFjcKK5RPSLoBQVNhJ381ZRZaA+0aJ
qeh9QBJ2NNXs9N3F9VKtEyRrKIHP16JZGhobQLfIu53PvcpFgPvFeNTSIe46NIcbmk0+JyW2J+B7
f592nfBLk3BipUl7g4XdL+xhfqmMtQB9tfNBTDZqx93eDbSE0KqkhiuMLpcaq6EFwBrUBgBI87Ev
bB3RGdc2CiqzehQ7gjKkpPLoxAIDPUeSnddQS4cCnpTDOsgEIK/62Vn4jcO8/RdVpmvCPtY5G4bM
cx3xIwmIxlGyoDyLPCkysE9UiqYqBRvVYrbgbNN/aS5ESG1Df7yR8ZMlT9fGVzMKpTicT1CwSkaO
d9G+hAOYrUUmA1osJ3D01c/KtZIFYIARbpZtvqCzLuZHo4o4Jh7AQzHsmB7uWOd/KXqjfc3UhnWa
EfqnAVzmOsgBrsSwBwuEDsjDcVCu09B1GUD48ltMCN6TNAS5+ltZc2SxNVlurOapNRFXVzJ9XynP
TmQPZ0hNbLfX0Z9M26lVUs29i22KbAyv322aCf6/VyC4Xw28NGNXMCeV0s5FdXkyRw+7JJOZPHxW
e4sL/DJju6Xrk33fqHag7HgwetZpPTEshg6xB8JhPHTEWa1+ISfeX4E4DelLeX5vNBSicOckWI/E
tg1w4zctkeE2VPFLzBypwfv/0Rrb0inDyRe3Fds61LDL0UJoWkRqzjfgih+wxT0wnXYdvhl170mC
4OmxVluKHLnU9qIA0jR7kgow/bj/sqX+g7UN7qcvJYHEVI5tV1ZZ98fZSx4mHOcpZASERrn8bLni
DF+w5dxhRkhlEFZzJpTUrnbhCS0M/pW2E+H4LgeUprIQRPGMmzE2UZyVjE6eoGMJaqTRCy3w6qH9
Oq0FNmTLjE85wJCqyQMkQbntU2mBhQ54+OOWTL5zNw6t+I97lvJ8KJj11y2X1WCBnTRwldNCSElE
ZWGJvnYrciJcNwz9uC+QLe1ypsfj3vhoUaCxUUBeFU9xhipGpeonJirl1WDUWhMZNlAIcEIh9OPV
OPjs2ngH5Bid/ujjveR6GPzU+MC2vc5GVKIgd6bdSAeZ93cCYvawjugtsk8UJhPpeprIujCnbRsu
dWVdiC9YtTJ/fyVwz8NiwgjXHwmNmwLh8SkPDU9hpgRW2SDI8mbfdh/zz9ywFLG649merRGkc5wP
rF2s5EPjRU/KWWEgJbF1z28rstHX6ocCFCZiApmyh004gxUxHmyedgPyrkbsEt5J/Zpdl3KgeQUG
aWlpr+xUSYOowMfQl8oQV+VwIePaF90hUBC290vr+KOhXbKfMHI8xbQnCE1sqAfnV7we7NxlFv1H
FKVT7x5V8WwFA0d697GYpwqwlaJwQ1h432zywPd7ytbJ3xo2AXxr37XorBoYRpjwZ9ue7l1uWFmh
1epLeORbsXSCO4dAHri6Dffu1pKLA+luAxFSwt3bkbw1TbgD14e8ummfMWvy6mOWPtJOQd0ZzvXP
REo8IUyM1urUqICekNdsatW2p0GqpKONIoE5pEPYSjVbOHotx/QYGph0NSpfhCnukyIT9YCn5SFX
a3v5i8hL1L2oIwVgmppH5BPmx0/2gdulZFSHidBvVdmWReAiXJYPGqwNssroVxcH5TexNsSXIGHz
Cj8sz7QwXMV9aqa/dr59HISA4JXxlARuim6oiJBs3+XuS5fTyyz6eAALlpQ8biSe3A3aE7s4AAOV
KrkVS2JAT38g1oNhxvtfsCyfBu4gwoOTfCIth/qL/0QnR5ODxZd78dCVjOB8zMiP0nZt6R+zDE6a
khfwqDFDkLY0w6YFKIbIS+L6fBjp2Vsnx7y4tImu9STkQIWpg9zmnhnOMxsWUmlMCfSd937r2/V/
0LhJSBAyy54bt1h+R8ewnecSeSjqi6wyg/wKZRarWzcujMunsBdPV0+zHuyy37FkrkFnIZUreYIK
GAOaZjfUfDOc5EU7dQPTlYZdkXf88lZGDIEA7c4SEM4UuChh1C5NOF6eXit1Ep+kSBWFGBdAxnOl
XPBqFum0ZpPgO4Fa1Wv3IV0WkMVx38Qaw3VVXDIfzIivEoMioL9fDLxvpBo5RJwwalsXxuvyclNZ
LCnQZHRKR5VrBmSYp7xSA++Y0xR88R/gxkd7LCKvntwXEshxf/DD1As68/WgZ3xBu/GnTl5aGgqI
cvqBDAsuYBGCx6DDifOMQUsR7q3Wokio0qhvZQknNNdQji3dokdHy1E5alZ6FYLt4wiZcPooar8i
S+TS0Hs9k7IDTmfuKxWohyZYn/LsalmJ/orT8Kmh/RGrDEN95e1q4Ezq+a6nMrHSy6XnfcZVNXr7
xcpqkX2OCBuWocXKwlmUDoqx7B6ISTyl+ZOS3Wd6ulvmdsd2IFqRV582lwOwUWD2/eVWbkFR+nsV
nW003fvwWfXKaH8TQzZO98dBCMqdKgSyoIISnffIj5wJHiY1+hAxlsy+z75cYotlmsm9DCf0ILn/
EeBM2YWGi3JV3//1VHjlVhuN5RueY/E088MBNRd/x0VV3/3ZSx6MDej4trFHPekaXJaCkD1OSvYZ
+M2L3i53AF6Bgr6055ocVkIJSpPLAoYtru8qP8me0/pbdDr5/qfa9wCAlrFoBvdpQxEJvtrgIejt
XShoz3AklB5ikwnJo0ZUVFCNOMu03tKYpYWGUsoX58AogXGgz9qaKLu8+/x/0hVQFA9svIY+HAUW
9qAN5/JlXOSC3i5/tShhAYOPg8aEy5hkKKVYzw0OIkM4f68sHhXWauI3NjY8nRgHlgdcIkLgReeU
APwm+Nmi/J29ZeYDq8A22HLKwY8PB4jzAklRS0iQvp0Ifhtf3ISyeppnP4wvEE5niNdR68otOAQE
tGoe/+Nv+B01hFj6H5ZuUnD9B+YEX0X3V79NQiyLsvnXiQDnDFhlObiC6/lt13/zH7I2a6X8OCzh
JJfHLdQHGxUp74cMmSeuXFdTidgPQ0IV7v5zWwQq+G+FXVMUgB9yLS4zknJFF5f6CdgWBRpcHU8y
WU+53HksmRuO0BwlH28MA15io0Oc1ME4WiBiocszh9lT7yZYUkUrs8UKqNDUBG6VAVXFHGGTY8ng
cEr++VXcTpa9sDB6io8m7bJwy1MGzQZm3yzxYVKGBDUT54fBiggNjgmcMYdREaOhX+smskKR48Q6
uI7B8gPJBZQBHzR6pG/jJkuEpMxiRimOlsYnkeh4KRL00rC+iyYDM/VgqBMlJp7SyT9L9KCXiXnp
XYkjTevobR38WHXWY6DXkfE9yfp8qjDkWUjIGNTycXz7pVG/8oxW2V3PCECl+0y0KvJOlp7vRtU0
TH7O6Dgqe+oJVAh/TXELI3+/byAiftdB3tl5fLHrfWqXc3+KXGiS8qsCx6DAhlrQTuH3iQffwOIK
lh4NTOYqpUa7gX/SQksJrcmi/U31Ax/QdFF5Rx9Zso5CEpnJ32BBeiPPhAzMJljtE2yH7AufX2js
27zRf9oPKQhz7dy1ENHzf8fEvT0SQ6quMR2os49DZH/H7ZeJHclYOaUGFWQcecjNuT5sGFKPHrDG
Efx+lenfZUE7vGeuyf7aVmRYmZRAhVNKVQnuUxMO+16AhPRI+AePpSsg55RnNfnFqVQ29byJFQ3J
rpkKmXXDImR8J+EwquqYZbSAmQUDcncmUQK+p2Z4Ec4NgHXwbOVJXURFhA6DG1hAe7SJrQdWil+v
vXDK45mga58mSaX1YHqL8pxYOusxzVHX1RMAtHOHAfjnxh4MTH+prcxCmIB3fOyMcogGRYIVClBN
SHJ3B8cRcuNeuBw2qcgCWfwRSmsaqdz6OqnoOaxZhOFfuhjxAtAIvWLBFWtE4nJj63Wb5dJDtdck
Q+sGGC6cGiLZHwfulTB8GeLrUBYs8eQbdvp1DcDv+Ne2GmF/1fh9br1APbm+Z72oqmePwgzYKZ9k
Z5WL1UzBPh/DfQ8SbwQ6b/7aBGOtJyPsWKM7V8gTX4SgSWwxpU5hiIpQWcqZ1VOWQGf6Q31bFDBp
Gg73AQ4YAe8eRhrzUbRgQ2/NnNSm7ztKvY3wuNNS3ptxS2ri8vi/GbocMmfFXqFBYuydjMLWtcPw
OVExSsFLqbMsl7odWTKCWY503eqZGL4s9OInqpGk+1p/KHdqnLDm7OT8iu12MGv/TJjI6RJRVVJk
OpJtufBVgc6wi4H55Dx5bdC0FMB29Mkl2kvz148U1gE4ZofZrdVlGEQP9X0//cKS2F2xWGZz9Ooq
T0ibODsUPV4ZEJqPgx954iuLSGWcpEc5SKzd7B4XCxzCDLhM0gXiopluhXdIIPXlfdcMuo9ddG3t
aJi5/kNhMFIAaSnJbo/9ooJoIvvn0zjn9lhl4NF/HDEHl8roYwTpwsmcaSzCS5ITzlidwGKcDpr3
kcy12ePDhVQU83o6KNCq+MBx+pZQlMyoVwkSijHGsFXin3gxG8VkSp0oeiurwm+okQ/wS0F8FqFv
kJQMiwVBTrkRcmSXZeR9+8ljg/qmWdq/r+DD5IPvsh49AkT8RcdDZiYSOqniMlJ7igLd0dsckYwU
BqRRl8gQ4TWM8Y4I6Z/7G6qhmVYO7STkH+fuhqfnVisg8nkN+Qmm/lqLvOIug/PCUr8NOWYrerfZ
Q0awceOX8PDGrub/0RxZEYIcMHFJKQe2+hfmWGuF3LSu/hV6dVn3RblIPUq0LyRZXod1fx2IhAsV
EaqlJvW9XZZpd2987C1UU2oncIHpzXi+VH/d/SqZ6SHNWOpt09BY0/HTXE4XN6UjgFYuyExc8Nde
ycXryfmpEJRX6zndyE+ZizAKVCDj285yxBMti/ycos3a8/mpCGgouzcaUXx5eyEgPscfoqrj/ma7
sJuXWTJ4D/6KG1PdTPk1kS05GR0WpWRgfXnp7jL2Z+4td24Ar8glA3C+k4Eg3WqPSdnYvDzPDCC9
yq/CWSosYZAn465d6tXkIHngsMNm7OsWYCNooalCmahQnhxbH79ww/WqEICyyHKJ23acYYYgh/XO
1wjaU6WUeuG0NnBKs1bNamqwP1o77M6B9e9Gzeg3RxGzlgYkp5YxQb0fhcO+1fwK80167GGcT/I/
jj8yq+EAKtF8GVOmY4/9W7LJWPYZ5W7GocYbn325TEWqas2+qQ0E3rY/rHXDSOhvn88PfdWkYz7g
u9+KA9PaNr4+3LqNuSjQ8oqavDIAvK6YUNm1ovHTFr6I1Ro4lkILheO5rBjPsaRalk93FdhSA4Oh
li/fRgDpOMIb+DK9fY3/1ostWp6TlGhjimNTunGmQkes3wM/XStMrz6duQINLkYM3rQhAdppa1Kf
BoK2Ew64V/QvOTKmrfu3qNX08zSwLn3vAH+YHI8AfKUmO7GZaUQyZsj6Xd7Ct4UsbijVO6JeJrSD
e2lobAjtcdNix/tRAhCqPsdrHLwPW0o+kdyl9BO12GbrKLRkwvmLUZsII09ffbp2tIxEmLn103zM
GcgnG+ar7n+FbiLBzcFK7CyLy2gQcQaRRtDwk8hGEF05LuPIFyon76UMJ9CTnh1eFXwVRsqO8lGK
plRCprmVd2vIwaldqQGFbidH5s2JBh/uTHt+Mx2bg5t6ir3Fwzc94cDvm+uA/c/1Gcj+FrX7qAEU
OpM2iLO/wMf86F9jJEKDSXDtIvK6m9iW0dJspb+dHR18gCS8otoEItqmWZrCSY3nDGS4JQNbwmEq
Xhln1jUmRIRhz4ddw43xi/ydY24yYDu7fLSXrN1/WAym7vEUHBIIFUCZOY8fenSCn1j8w+E/3AP5
vBB0yGESM7AzCxQlx+oZJkqkLbDA2p9Q/9DKQbiOP7ue9AvSGg9FGQuzG4LlDJXBj/7jbfffMrnD
9bIba268NrQ8iBrQhzJBlHadre06QUztwyPjyMhWnB0xk8YLc5d6DMw/AoklAvdfASROsOSfLMzh
C6lRT0QZ+He7ylbdTnqb+vo1tF6b2l0dFuQFLDiPf8gIzdo2w6XZYEWq34j4E0veOhSHESLU6jbY
zvWqeFY7QmGeeHoVlo4F0jfxNZaztjacA+/H+cDnR20qpSCDXNzzu6ksDGcCEQzJr2yU/aIo5jTU
EThm3ZbJQsQwpTQ8zqp4uB7K53t+L4Z+lGspUQv+980KMFWeFFqegCAWjprhKHGnRuuk8Q3bns3w
MNKoDWDmtKFRIXA8Wif6z2ox1ZyCaGPlt1YRyfXsiruSJgkhOvKZramBgFRHC0SWiawRx5anXDKe
iQOR6WbLyI6xWeJVFQt9NFo+DwITGtHBKLVyoxfBasLj/kvlTT2vKjUv86CzcQrMygTGN9L+xrur
g2DzlturBhRV0kiWPj8M/ld2inUb/OpO+7HBa3UGZM1UsHOGl3yHv+JiOuYvtRXaQ7E4W6wYp5/M
p32dfbfUzBfbn+cQ+bqUcii3rl2UkZYBCSURZJwM0gl1SggWa7uOekQZmFwhxkew393MFrEUEi94
0wDMylnH/OKI4Kgqs1wjWd7Zkb1GIJshDEDdhkrKLTLF1DdQYaCsc2JPtecGHjckJ28OYn26nwvS
WwS17/hWYYviSfhN8JGe9pNPw1RB2B3dqqucUZE44MUwZGUw1s0XtWySgSwdxt2B/flIc6EynYIJ
YEf086U306t0SyWBF8l7bl3gO3SU1fvdDnVo0eVY0hOeEshTYMhILu+cbe/oHj3IypbT2ER1d9hD
ToqbHYD2BZQhHUpvihrgWctfpDhAibw7pPQ04NV1HpvrM7Uq//g7Ue2Jpo3Ctp2cgfhkNZ4UMA29
uum9rPIAqq1PfZkNM5g87sg2WfiKlkO6qLj4n4UbokWNkDVEaBXIY5NIAq0D6lS+pYYjXgczYjij
GRcIyEkQ/brbW1AzPkWV4BeZhQ7rGfN3g0PUXV1v8mZZgo+1OpdLu0oSHePKkCnQH9QY2jhmfPFS
R6KCAtYG3OtqjiOHuCq3Az2nw9Cg0Jc97nWlQvHa8lXVZ2pVqEtRxOtkXRR1T6d7hmrI8R0BH6oD
S2veGbEZR/ipFw4EbxA6/rrSyLnpSELs5zTz7R85BmlYVBFmv8NlxnA9UkXoZjxYCsePJ4C2bb/4
KpjkftekMGjJv9bVSlAYRvyaUIh6aEiGYcxKAmDpziiRbKi2NEizj+WgNx8qWuypRJ4/Nr1VGT/M
fsz4j9iFexB5iAF5lwiCyJwGGzEHneL1izMUH3c3sG2yvfRcjVhyGvZOqmdYrcQXPktUIf/nFgzT
AzjrpTgQHNTEG9K1Ui7qj5r1bHX4MXZ3sKgvy//Ms9zNHIyjrjgMgN181kvJ+Bkls+oLTz0Rh4tJ
sdYO26lh0cFP1uBxc746Ma+daklM0KN1H9EK2Z82v5O3lMq5Tl6t5WcsYTpHB2R8zXNnUtcd7Z4B
2+39AY9XoeLNXpy4gRyVc2BakBVQf3BQ5zXBAgWQRFnBmv6SAHKV+rSeninsMs+tOJeQek1YfgZJ
MZllY9TatJ0rGbjOJfhdmJWwfZqi6AzTTeoIq/+zeKVxId6s+nCnXGLTVtDHaFMbBdtSrQkMhv56
X16H3EcBhhKRkgJxtyAtoqn8BVyVIidrvHybeyEuWsGRxlfysnUZvtY6P8JlpPJWk8rQjYzGpprI
Sri3aLC5oU6vczMQsG8JxhwX0ViqGQdyq04I9MBEyncHSp/AF4pAez3ssgGFMfFZnvPRXfm4Fcz4
hG411+BPZLShB2AH+LkF8LxC6FeZrnl7qIjhrYdgymPXdvpe3XCOHUQ+LwszoKuP3az8jN5Q+QiD
Fx5FmN+fiZuDrlb7kw9FjNmcgCWuPrnlcPO3fz6r7DDdC1TAfDAfYJiKYvT4+nmMDtO/Zc2lV9+c
e3z7+LyOQPeEQExzLiH5iXiqBVpjmpYMYmfNKhJpQvctJ+mccRvaqHhYpyJwHHYDnaV2kiCR/PWy
FtkPddNyBfUQVgeOyVcs12FAElNtHhgrp1LJROxh2UhY8ggFglh9oC9YAPybVVoDnRvj0+QPvB1D
XjSCB3434c2805i5XZRixEe4v+6XqInVwO1R4FqQaO9FZy8Fzra3/sJ/DdFP31Z0dp/nqCeNoekF
tC+h+F4KdIpJS+jIpgXl2tXbKlLCHRKKFpKdIrR/1PUTvpUww8WvpPpQzG3SL4tu8d543MVc93a/
SqzSEsIS/jUWP4JpZC/AUpbkH7ATvn837nOGx3zFnmBEn3aWQ8FD2tzBdOAUqxaBN9QmPHo91MoU
KoMA3IvuG5nrYB3mMgG6ZYvnPiRikWHzXa0YzzsfAWcGwASsy6M8DZQHosr1B50DeJ1hvs9Ssprt
Yo7YnO0IEfXFYXbybjHpE0lukEE8+EuKVOJwkA8MvkoVAvcHG8fvEc1FCPZCy4zsT8W+GYh6thZh
iOjDTrvHDNp0iGv34Y4SHclEdJ0ltZN8bfUo0TLi6hPoIyI48Kq20BfKVGgmeTnPtALWdxKlLCNG
7ABIkkz+4vcC5vBlN8ZyKSzZQ/KxY1uLGcd7OmrACKe4F/xmhz8ACvh095cZIfCw0n6nl/KftQ9C
BGpJJ0i5ZVbg5c5iBcNq5OeboYZefIoXofeRi/4uQsg8tdNem+sxCDJhSfY2z5zQr7MOMfx0uG1E
pjJqGKtfVF0F8JMWjgBRiqNzJKr3gZpEn02fbOwEVWgS3mKaNkUn5e+UFsJ/oWry9kegIpLKRd/g
hSHp4ExZ+kJ3BTyrAz0MxVxRmwLE4uoapau6qeAmP+/GZtuW6CAWY7Xkac4P7bubalTmID/I8lBi
itipXyjJY7lmnGgpPhcUzmOEDBGl+A+vJz8yPU3o9KkWoDih5rSEnZ3990YLQRhR7ceXEzu0DwiB
JqllkCq4gcvS0wCvBgPT9bGfAqLVUxYkFFUkStW3UMMJ578g2e30MTnpFEQXdKK96cLHKQ+P3+Oh
sgqa0hrc/DApN9ZnXmdfmhPDSCsFHaZ16nApGuF6vtIodJSImkHmJFh5oUg6kBmSnBoJCFK3n7bA
U/GeSMYKNOVhDChpxItoatLHrwtHOoqhtPDpuqCa8kcXqXB6FtrybBaNLUBDCeJnNu3BbWwgnooF
WuWaaNMF5PGuPqTyBCsaWSHG0qkh6E5hiyg+1cdwmk4i27ICWEjLeahe5Sg6aGsoLAdew/uY6vqm
thmkAq6raR0T6jnxkEwUjHykpBrRIRF0aMj1+hjNo7ZYniwPY2DyieCIqApQqWodkF5V3UFnZzsk
S5bOcir62rZqf8odJBpqgSAEcxEoCk+fpxPCFt8tKbh+fgCL5M0VuCwyd8KDetn5+CMnGruIosLQ
6BSipt0JKyxwfNAS2qQa54SdWBFlhwmQTlPX8uUIofCaaJJbSUWwG1lGPTwA/GuaRM06Q+bXEYbd
MUJZCLLJBLm84cH53rfOQaAl+795kczkK3sx3zMpnOgxkJc7dFzVu9hbrSzxy8ND38vaO+yYOx/9
lxbofTYFvAqUsSmHUreDNFeNQLG0CQ9lnjUwnPlTljO1met+sk6T+W65LmOQjNP03saQf8V0HW/6
YCgc1Kc+dsAtvBoHH2ysNbKsbbv0X8d7J7hUub9g/oAd3bYor42224jdOJq+ioVBcw/gJyicbIsM
5VpFSnZYX7Jiw73isAncdyMb7FrgUlkXcW5z3nO4I2X/atR35GCHDVUysLcseBYxtGtJbwZptZqa
p8bacxyd+2NzhiaRXD7asV1aTholtb2BcUlW1+28sbyfQwP9ICWOUvFj8Y44a1fr5bWvXd5KrQPw
EHSCGhUXYxsuGKl9l/deqoBsp1kPBS/PTGBifs+5hB04mIpjgHkyCp6osedwcofwJ5rNTcFGD2+u
Z8f3q2JYNLqPpSwLv04bHhJjFKjsDmKimEknjSJcyEU6APOk5os+tbsUupQxB3d35GlceEBN+S9Y
9JKni1fK4Wt4jfnQ5KTBbn3oXiJ4T17CKs14d/iiAPIKoz5hxRC62JyNZIYOKiwwhvuzCA4tdkuQ
VglDjcxee4pYp0JdQ3jRezSvMzUb0iOe0mfabOUHoQLFVpzbb/lFkXO0W6AbPrhnARbTnWnqlsH/
j4TG9cd+azjFkadRXvOlrujOOXyp03b2s5WFmoe1hBPbxW0nPdz84l0NO+O/rXCYpm7iX6AgPUa5
jdf28wE9DvT1rPy9GjD816S0bjpVnzQzDsFJ6wzWXEwhk8ZrXuO4aaPap7DhW0yQ0vb+bU9k0LWj
t2mKFPOHt9yeUoHt75S2QuTUOP/++mo6asAiaA0oSHwUGqDl6qV3MvVFJaZ0GgQbtPGBHMx1wq/S
XpMku7X/LNVrhprhYbKZNaRuLY6oZ1xpiu4bwGqoXTyxZaHxppDAfke4KbvW41hQOiZTyGOoAD0+
bAdFPCMBIcqbVo6Btp37YfIt2kgFbj4fHVY3xJYPIwXvsIEan/1bdIcR0EBZ3xcN1IZsynLdGG1w
nVBCcFl6+ljTiHe3Jj6z0ZaVocuqmyJTAIM4olzicMnhFr7JQQ9TQRtzlg2x2hlyxMOFu9Mj902T
0zOB6NauMoLog7Ki5vvkRYUDjxG1c+YGKuBiW5i9kB/SJfjkzCDw9pAy5gSxb/JdsM7DKlSQMvE9
BoLDIGF1OZs0DYX5LMkMqDtqAE1B/+rS2AobY8PI0P7Rin/12P8fffBK7WP49IEUYti2Kph/Aoaj
6MEJeZEJn2dkZFWBnQuy8H826F22aig7jrupVW7J4O2XG9dqHnBAqeKun0iq4LHzuWd79jUXX3a5
OMzEYzwUj4He0bYWZuQf5NCavftMKsrfeE44Qv57d6nBBV7279ggFzqWImMmqUwuEseaXIrDlz1E
omim6C11RAfb1KPFklGHLRXF14zZDXHV5+n7Irvy5Dn0LLgU80rpa/h1m8zKdNs/gu4pfrDnTkVV
AMxka1SEddqu7yVWwLbCQQv2Z1tIlzPzcpaaDT0IbSObLh6mfYUFulDAsJSytqYKrAtaYZ0vgAt3
uhHW88MHC/2wSs2oCoT1wSVD46GVLqi0wVLuo4KUJwkstr7r1RSCjLD04f1Zb93wNj/w6NvwE6y1
ly8N7RnxPDQUIjb2h+5P69Tt1yKmvLHAM1O9roWVo1akQRQ+PFNC9Ac82wa5bxuvEAbhy8wgo72S
VfLudooADwiZ+hcJZkZ3C8P+5GMCplXorFBQ7oFvsHWj28Wn9kX5/FV8DmITa9iEJ6uQz3x5RxSJ
YNJLk4EojrMexmMnc5+3w+bKRYGoHhWqtPgnhCot931iplx2CM1H315/cheHEhuDts+Rtj/foBMG
TCMGpBnuRc428nPF217GlcxXH7fAQSi4sx2dH/ur+jX1mC4LtxAYDHAK1NzT1uv6I6WiqHaT/gk6
njd/LGwVgP7bXJIGdZXBDfBFYhzUIV2PhT/N5whjGj3g+mPiVdT/3bMI1daRKNxIdG92QE/7ST9y
OqcxAZgHApGO/C877frpCBggezCWhF+VCiDelNA2Ww/QZ16O5XONsGohcgoAQNheQozfq2CpfWTO
nNSXPULX+ZKdEdWfbI8F1WMnmwL00CWIMgmFpy6oEKh6COaLVwGZy576nHs/BWmwgcfPPIvhqFzi
7on65Vp398yiOPjibv+iDr/405LVRLDjeXva4ZOP37CgGiyURIM49IMXmjrGiTC42vvY71ZqmXPe
EvWsOV+8qZp3qOPHfVLO98fpFkJhroC99r1jLcL+v5w0+MRSBUS3luR+jWtv/6csZv55Ixb5dIpa
imbbFflQlxnX3FI07t18CsTusYShM7SbiHlXRc5FkuCVCMkDL6TsNghgQhXXhlqaG4FL/KMCVaWY
Q42tUr3Xz5pK2FKMsX692ldpP5IOMpPRx/l0A2Ld5Q506a3n/US5JC/r0YfV+U1Fp41GKEC2PgXA
DXbQtb8osRmtRXvy2GWFlLjRd3XnIwGxJTUtM9Zbyf2Njxsq7FENlf7wLf4sPnQdvv0DezjN+2yz
wYK3X99uSXq1BzjfLYxmO/CEBetvr3IFRrliCl6l0UBKJx6DYJjqoZfUsp25IBv2mPExUz6JryX3
OVhman13z9RGptYdBo8ZukYPPvFLpMFOkFGdqwPyDXyyqwo29q3lhyHsrUIl1424bO+HomVALaXW
BCckSsIP0MQhz8G8NFFKTA2Rd2u3I20z07hgAziQfPsMBpLyeuCg/V5tY2YqCA/DA3i2LQbEgGNR
HjVZdbeK02J2ku8mcwYmfvJeJ05G3qnifwMB0/eL30HkAiKvilclsXUdt9AXa5BQ1GkX7Un7km9P
mhZdrofedhmCpHQmxmPfKqr9NT2JXtji5SlGxEQTm3w9dilW8U7xTZcPrS/hMf9y4djfi1YkGF41
W5buE2T27pE0BxKC32nIg6RYRaWIUV1fOuAOwMrhnlAgXivmtLrnWvomRD6b/F9ztwDcyiUBLHfF
JFfHm353/C9lD568EShmgmSi688DLm6UF22XPqgY3sk4D71XbXsJcoeV6OSiKSmTa0C8j49mSwNc
K8j1bCNGTIooj6gXjK5JxAQCuKO0SjcLNvSWSdjIZKon5Rgpfzzs+cPTSmGQFoCY1c/xw0p5obUD
pIz1vM4zqQpKItfLq+X0tzpY0x7XG1C7+VjZXMcTEVOFmHsFItG4tsHRRThwEh5PXyiQMHvzF3yM
SAf+bp8TGz5EpGUpkPxV+sNrSAKUgOzb/UfWvYw+4H+2oWfkr2qxTR+mFU77lyeF5/bj/IFi4lqt
5F6UkwiOQIhwijCLg2F2fmY2uU2/MI+boieeZMiVc11LV0Ch+dUitjecwcCerBdy4bBi9KbX4YoU
qQO6Oe1Hjn2ZLk+KQUXA4j9Axcg9PXqOSms/MF44JmdY9jrc68ftBd4lNJ6o7K9cqyNz1v4cnJoO
TgLVGYYfho+IQ17TA5fNZ0HJh3mzd/08M9rKTj+rNGHegjaz20b9KPyMt7nO27xQGak08xzIbMl3
lU3SxofIeM6WIr4OeNkIEMKfd9NLIgZFSYYqF31YtwA9uFP0lSwil5omdzF5M7+bC7MPaau2JCaN
QQHtVL8YgupxQCURyyb1fHcsc7k0JgdYI5GaBhFFqTk+tPdvMZIhHOZA0xeuKiSr24VkhIn2uQOt
x8umKXSc+ZAt/8DrUfqnYZPW6hB6FXqYfiWASqGDtwLouzcKk6BOpRHzBGfdNGOy7xl76SiSqzxA
sKsNlZBRRYizohPmrrHDCPq3JuBNarelhWUtIQUX3ZSygJ0O5Edr30By53rVyLypM7N9lzlCTHly
PZ/vJ52kU7yrAu/AB/LGmvwlqXKxUKkpj19JNRogcAw6IbfVFBcQtDXWrewOQwtwD2ZtO+D//plO
YD5qZ8G52csMiRa0HJaZkOoNIxTQYdPqIx9VpkiQMLY1XVjo4QGZFPsgdpq4oIuaYsmTBX2hY0Sd
MFZmF/kqvzY0amLCFt09npWTCX0xOjPspw5nr/IYSfVCLRhZe6ewuQkJ6wy4vD7zi0Dxf1SlWkJr
Fwapy/YQWqYzbNaz81lJq+Sv0BwXPE7j7l99iSaXkXx/tbZKueGI1Kc04LtzBKYDv1hB5qiDUUKH
F2zg988gkEKbmmlRcCcXd/MQhXlj0VVRtig6tPlw2OV7WM1O3gIDKXOHM0oxJW3Lu1r9nlFFDVDw
5+qh5+KNO5Y+AHWAdcUzYSlxBdnPRyeh2MNI5O+dJ2sfXf+24oLWojzfeAQ3CbH+BW77EHoSrcAL
ZI98cnyLsrDqlCW6j21/Z+Aup54yEx+PznLYEoBAqrxqM2llwoKiBtclWy+OCQmV+hMYa/uT+Bfv
N54BcTHe0w0dxAdcPJrBvy90OuXc9BTsEPPKzHWfmYIiEbGX6XPKOiIhYYtyqoG9epb/VOcVHPg4
wXuljvGNjC0QOmME0UQQ/wXGuYPVRtl3hLLw40OK6XlutJdDiYzMbjb/Lakikl0Q3mLGSJY7DShQ
EKnZZCQN+LP2Es57AqySW/cRpWvmvFG20ldrnOrKScjwJxhqUf2tgUsXt2ZdG7yit9Gf57UvJpY7
w4cQVbC9t/iF3pTPxM2+p7mhAeKEh9kJdMcEMdPZrobrtfTELHKieCDM9akljklS0AVGakiUTYiZ
ghqaxFQb/ukoxCVEoyavJyJnvFDbWtXulD5ZFB6EwxOc2yvXOHtBhkC4gjWi/EUKQyfcuX6iBmHe
2ChfuEQK4K5UKOTGvzflkofkOTReUfJ72PakDJ7dAQheCWQ3D/w9vkw9Z1BsliRppypOpDcnP3Gg
YQCjpp4EqjPhkUZxAi5exYpUeF8A7a2wuUyxtG7nXGxVj2h4Q/fpoPAjEhUkCG9b1itX8wj7PJfR
Vwn189Momo1Vd4c+doC7/0zI4zljRqLNOAOzbdDpkkSlYMfAXntzMzNw/W8whZBWjk7Fg5j9tOaz
m0zofGfpy2gDXF4cKqiSBxDG90IzLSonWyTf7fsLQuXx9CNWocxNdCKLKC5IcffUfH8SlFgFqpsY
xOxH0O61/wsRjs2aefNWQjxmWWuRjIkapefmzh0zJWJ8PvJQVHs7QhlCwUs1oaCdwtRitu96/PXu
2O1Owzf0dh44qBxxmG7HWAN5mGxIN/3gWdbI/1w6ipY0UUeIzaYy8oodZmKKRlbchYChKQl13DMm
zVcT/9SIqAae8YrugOsgjnb4AgfkeywTzwlQJhp6sfaZNFiDBzCSNXMETyiUehja0W6kWBAVHP4e
b2DGnJJsYHhgTkcen1ds5pysOC8+dwWT8Q8Y6EonsfNfWwDyKxt1nSELa81PzxgHemU2finELoIO
hNORRBgNeSM+h1sqfBW3UsSAqst1cTKbjqk034EZxaC2FFzsRLcTybGrwoRBInklI9zOvtDq7BYy
5OuiKgVU5hGx84TdDZYWFBN26aXlDu/KaqryiYgZ4BuCFLI9PeMvkTmU/D0lBkLlaQXWgEQf8cWn
iqmTFjY548+3k8zxQFT/rerA18d8AWM5ysI98zvis3aN3VfYgt62rhB9LQ3GLXT9NfJTVsMmzq1z
jZrpC33y+HaMxMcAJfP3TlCmWJYDQ9cfj9LFu9iEkiERIpg50SI7ynZOucYM7G47itLqesvimky9
lka2nsThCBdVQ5/wic8shvNYKlhCClNI54p3NpiIPbM1fu53v11Ivn2WkITBcOKh0X1VTKLctsN5
+kqCMn1hDjjmGIfisE+KIUoxi1H+YzZoFRrzVcYfn+FhoweESx3yiawfBeYkMmtdAQFjP9S7Ddb9
JxMnFA6mCQH5DSayTj41FVPY3wVpMVT4OpSZ8vZU7IR04x4P+MIAC1Lfnz0SWRvq57gste5n+TI7
7ZPAQeezyhRaB5QAFtSgXo5Lp/xISUNfRAglPlUoPz8jwZlMojyYAQC9FCzWbr0zWyJz99bDHmlQ
gD/K8r/a2nizULIK+h8JASuKcb/H6tO2hBZqEYfRC3V60u4aXv/D4cERG7VzCs5CkU6mdmGMLfDi
tQehy4VjGv2TRkA34fg49fToxW8fbNddLEo4Kb07LjunvQHK4ZusVNQ5dKH+hbmWUdwcJhS3xSjj
NWACkjZaU/6+2gRVr96GZ6ldulJsOxsYdHhOB62xwExo4rg/kumFTbmLQZJszVwp80ryR61XsWN2
rF56mxwVO4woI/xfHY6hu0Hq+Q0q1qjGl9MXyWC0yBoZ0+cnl/4y7HNFGC9khxcKNVdYIhg/Gs9M
XkTKMQsvEXc5z6SYTvudbsfy9UdnMRYzX6ZaeJwL/jM5rR6tqaVFQqeigKPXICMovoyDG0dBnnk+
JSKAr7MZXOzo/vYi5Wyr5d6H5geWpo6efjUvEfzOV0Yb43P17lE5gkkj+vvYJXKn4WQrwpO0SW8t
98PG6NIlLhNIrMCHGw5cjsv2evtsJXIlA9AHgH+Eel3pwwdCE0kTgucX/RCBWzoFAIbFvAw/lymp
IOyOx0tqNsOcpc3zo8z41/+v3H4ORaXoT25c3+VhUNRYrPrNGsMUt7Y3gkyNvX6ZM4KUeHWCINj2
3q5oMQovl3UGGv3dB2BMT0KgWgqztoUG7VIIBXFmxOE84PXAi7UwJMQdsM5QzFj694SflyFAYy7B
CcXyR7RF8ylbnBSlN5W9YL3ujkmyycZlGF5BPRKCiotSvc0Ew+MYOXpLKcQn2Uqs45j4QjAZ24R9
EcPapx45HF4BDnUZrCrxXaoDozaI/wGAx6r6lL5VhuHVf+bCitGOIxemvku0rpM50JM2FCjSJRrs
pv/EoHruw5WyP1mk4QXGc3UT3uQiXDz+AS7vB0y5lePIS01yJdTmIuWyb/wOARZoWgStKZdBSU9/
JJeO46uUU9RGIg1ikoILw5A5rYeztAdzqHQ+V3AnbuijbgpMqlDF6ppqYt94QwS4c9zK5/hJnMJ6
CNyKyFy5Vmt1IjICCDWZOocx5OCgpJjJIGFWt62Em5tRt+G0e20JL54bc1yWDk956fpwwZisDL5f
njQHL/8JCT+kP9Nm+U7va0L0bVnw7yrotXOXA2ZIBQ0MZCB9ouJC/MRcdxhTcGMa8YsGhq+y7Xui
I5/mdcj/mIuUy0EjXFwqLr5gGxMT4KUIEmAXyiCQWteg6+kw4tE790zChVwh7ET+WpNfq+uzWPVa
uqFn4UjdbmgTTsgM1m8hZwm4djLbYIgSwXsSvVmLGZ+M3df/vFgbu8kwhDeW6ZuOYr71KX76yqYJ
XeoyKOBc//PqYdF0K1RQgwBxCecagepijv9ipEv8pzWhJYTKjq7UKKKzpUjZyd7xaI2H2qP3Ln7f
tFpjEYpbWyQnxxw/+66knCRU7CjMrtDcxrk3m5oJJcIfC/fMSW7i4fgr0RYT0IQZqHGBX/Fteeo0
YE0NjHIdjUOhplI2iEmYkeXuWWYCfVp/r8J4qzDiEaPP7ODwU+I7ZzLQTgK9bW8q+Rg2C8LCE5Ni
65YzXfSmQCzVwdCS/JgAVEp0gMjcEc97KDV8yI6ky+hrOgETPOB8nAMeRomngivfdkDe/Wsc0x66
xF6cTlEv+wuFWFeBvviP4qmig3OMjOujly6Rvl8sP3H7TVCYZVWnAvqGtSRec3wdZYntTFKQDwMk
e3I5uaZ/2PGjug5g6Yl9aEPZ2Lg2iJNj+oKo9+l6M1gPmZxVuUZ87cRO6vrpyyjNi1BvgPc7hx1c
6NWRP9O+OQl+JyhU/4FhcSStHCvm/szdg+Vfp/6kN9pZl4QSoRnwi0ij0+0td5LLR3giX8qCwqI+
HdkAUkBhjBgqdfmZ4VRDoUc5+m437SzfG92G+3LMujD/0GGnJ86xdwGKVssTumJ+QoZ1FZdtBkmJ
oFR2799lf9ctYAVWkqD32o+URWodVPlvIRF/1s7i6WOjZxpJx6P9u/ptssJQXgP07HffubYUEQSO
bsYOzCCvfMnaf3CRUCnjuHPyIwrFNFpuNb41+FmM0NFoYLN0x85bdkgY3n65nXB26x4vpjv/Nr8N
pZX1SgpzQY5vpPKiNYdXlFjFQ3HDW0qULfKH4NlBwxdw1JOl3sy6M96lyCdvB/hu+JIKaPG2Eiem
c7SCw1aDNkAbzKuYSoiqolsWGS1qwmN9LK7B2JhbLLGy+K9KN0INWrjSd+8+Z3d7N5Wtnmc/XB3s
Y8sYxZuKMwF1rzbDEF3UCrNELmzcJrAzBeQKNivqyVCCqrrA4ieuISf6mThyxFEXoNXS+bKtEHGM
s7DaLNw/XwRhnMG7Af1fcvwEcrqa1UGn0XY2iHrL2o7WV4uOSJ+dzfFRzUXAzg61V/ZfMjIdqsV8
k7QWtoH+PjkexgcxZzDZooHBT2RCgAcG06gwy9XJoO07TjJg2P0DzGe7FAPX0Yien/J/TUrd60le
SwyWTfqfrImABXdY5AGkqxu6YSBQYmXiStYcglyyLNR1xI4mUC0/gOI2pgAyOL4plLt6DKZ/EGDJ
QR8jaQoiW/It7svgitPGFzKsj25jSxpjdEtVt+3RfqRKczZNeFG12ifmtrFdzPxy+on8mCQcK/sF
AnRhzpwPOG6EREGDX/pEC8lj0Uniot4P9ny+yc6bc4T0/BbBD28KNVOSzGuRWt5VDgHnu9nCK/oF
mH0+gX68S7HyYvMtG9QWb71ENtSEYFkEYp6bXYdgOfb8UMVSTm0s8GiDTYMzM3TX7CqAbmSY9X+k
gYMdMTGXBq0e8KBTrHrHOo/x14EU9nxN7GFfuDOoqC5hFiCBr+Dn9zsUhZl70yu+VMbh1rDT4G8n
I6Fl65fcd+OpmvYHpEffYMMXONHljKAV65f8xcws9JP1Hb9ymVjZRo49DyBSNOVB5YTT7MgMGYIP
yfTV8yXgPRKWA+Q9HhQKgaaNcfLi/xJ+pCNRQ7JxamM7lUFf5bqSdOWdO8TWAhJexLghYJ/8wave
aZV/OsJCR54BKECXlHa1ekTJBK91Cm/7P0O8SjsUzLEEd/rvrj2GwTwuEmEPSCVWbgq1O9tqiljP
h4YeMqo/FQF+Pzv8LsVf/+xlMVk3BTWb/jFsJsqKDHERAAKigCv4ectx5chLQD06apbMznJFzzn3
7y3+22YVh7Z2qDqs+SmLgtKoPqAMqPYVDjCDH4mV9AynCxpzUEqyxPtvbwgGVYxL60M0xOBDke2U
iNtL5bcNAFxMbWQVr/ooD+5jabNL6QK93BCo4PTPdQGcRWUK/325VeOad6erJFS6BQZSTbrQkv0h
ejWzTEj9yLfXNBKGLX5AA8nQE1QtEHbXanet+D/2Pfk6JQaVlz3f/DTdBSoLhZLdvJvl2E+Z2BWm
9RDmTehFEiaAqXBjXG8uf7tntTb8E83Ezys40qxWb0WuHKmNQwBq44gNB+DGQ8/nFnxe43BsWDai
blBc+rc1YiDbf12sNJNSjeqHuHDECxIPZZkq8xkOljVPjepSw5KKnVNoz17Wltd5LFb8F+A3Ur7U
asXvTmWV/mOu4opH6sYqoDonLVaJh7kEEQar9lkZzGSprqGbgU4M2hOXaeCZifeOdrYdUdGLADdt
OBYWiFkvTfvoM+/J7gHR2kqlfLWumf1ulH772ZCFaM+2j2rq8Nc3LGYWaFCpxc80IxTGtXBDiL3M
3CVTi3wku9OcYBG+Iyiy2UKU49oDGjiji058bxI38rtgSTHCK+dd1OKQ571Hml7RbUNB9++V0eho
bfegX1y/yApTXTNvrKBQKL/9rtwxlqeXc64pXB6NwKmSiuZuCG6nY2KZHUzQeKxVVzxg8S5tj4uH
tU2m2hlfLFGWPcsL8V3dufDlisA4qCKcY0C0/5pm+I8JhQOnwhyRtWUo1DMAhQ6seA4tkcHp1QQ6
3NPs/ze6muE03zEXik1v/2PwOAZamxaIqrtqq2RvfmGkkwXsO81RMz44hLsRa++wKfO9ZL1QyLKe
wD3mSdJBYU/rCdgRqXpgLmKLUwovPpmsPiQyBlWOhBbXcwZfuS9uox/WMGPRCSCTr17mwxQbowQK
fGzKTRggj+GtKL8ht1ur4De9B0d7SBp5m0GcdIHDky5iEgtpAs5rALS8erMuN4J/gibNm5Rx25FQ
0rlNyIQiRDtUsJQAoi27NCHeDhLSVTpdNdhPL26T7vkObET+OHTKPVaVplhblsmQ56GlOhm5evcZ
RUue2KvB2nZyRgvJKDY6JzqacE9QB8Oy/7b1hp57fCsuJbH4xkLxzrMhF6mDhqIKxsNcgNraMB6G
5Npz6aMrqWkzgQBhYc70LpwtWuNHHQb2BCpAsXBuXtlscWzU0TNlu3ZTdQX5rFYg1E5PhSsUrDyr
xYxkCU/JFC6bxVNn5YTUH6x3+J05KJ1Ex/+Ims5VNe42FjDf1C6Km8bQ9N8QWXpbNayVcm6FHBBi
XdboDZeTyCP14PwvvD/68VtWqXFcsG4pkA2CarlT2VcSmVPwroYDdOdwEo+WIu0+Oq9RdS49bGSK
V/th8T1m9W5v8OoLiZY47F4bYgT8b+mBj451U/3ps16LSvUNB5mK6Ji1IwyCkO5soHEpbi66Z2BU
zgNKowuhNE/y/fgm5O6BNJ6Dq6+jP/qG7AeP89mXBeGgOjD8WcRNytTsFGBIZrI4We9pC+NvSfZi
K+RTyjTCOlQflg+fNx3Sm8OpFslwkF5gheMtJcXC0j66CFO7B2BT3cvXZ3Il2OndczD3VRVHIWDS
TkAiHdDc/J/2JvhSRaVOK8IFfzU+UWiy2OEHIXzdVortLqFUCMx7xDim8qjJz5xFRES4lWjbb0RJ
lAtwD10KynEM5cwMFntP0WldvwsL6NPErr7zQ1gyAzmgQJUNcGEN5YuD0pqhOyfvxX19Ioh0eSwz
WINB865cx8mhxcezOt9783ymtW6x+YSp6lfpimMCwvpmQAwLyfgTNIGUuDsVr/1wwtLFIbCh+lPF
1AYpeZAr+W6JuvR0maRdfWMicuRbvKiGveBVBT/I708zRgcuEzrMfWtP6+x4ZNHYNZMhS9z90cZU
OqLw70KbYkcBtl2z4NWJCdRXQcU+awwrAT0VL28b8mN1181G5qeySD2WET9MzS603b6Cysixf2VY
BJ+/aUrrtHoED6iyaHrfrV+teK8FCzdLmiyf9b32FskMdeqj+oOEeolGwCNSV4aMHtdfK2M2BUmW
BQA/0F43Sx610e1j0uYkFhbe8RkaCCgmw7uMnSETSWpMqRchLlWkVIzZTzptQKe1zxPSx9B2ijsU
UPDv7cX9UXUUHPVF82zoEkHBWosgVBXU5Ky3nE2UywR5n+iS85PgbbTzuy9glrfzo4NLbMTXU4Z1
mZSJt9HSlZEyjnpp5VSfNCPcNsK9B8BhpkqsT27bVc97zOIwxBL43j0xk8uwxnvyBRqLCeJIi/vp
nRF892MvruliF4x83sD0whlJjTAf8e+urJWtp8nbfULhDN41JRtHjs939MdNdFrGFl+NPiFVfLXb
QPLTfQDCrz01+m10Rd+AC7rfcmxWiKH2KLbfzLE61CusqGS12cBE1ccU6+DtbxooEPtjtWnjFHC1
VRjhepLv2owSwt/CHrFwz8Q8ghLT2RHfcYVh6OTpHmoJBn//M4kCyga17IzNObHNgCsF/M8fDqVy
GgLs8shjpb1c2WYX/V51g2bODseS152o8XDc4HZYNpWzGW9z24uacU5LMpVmmf1eu2cFOQCzmm64
PXV9tuGlpSAM4NKl+3Ss9KA2Wr+UABsLrZj/SfUmx0Ph+MwM+g8f+axSx+WIVuUJeoLNDw87zDHG
B9uZD1123anVAyKEORFC2Ck7jJffnyGBcoZUpTxOvVavbNZZHuM4wnzWvwX8L5CipUagm1BliP1J
KUjHGG659hKz+AI3838QIRF5fyPUcEEQraYmsC5Thz/fPOnXY2TG22V7Oq+q4jaLL1KF9Pt1RuNQ
RW6MbHbMmnROt4pfPFAXlYmHm/CI4ZORJ5W2SGx6JQ+mil+oG4q6GwHswmoUZs5Pr0lKmh4t+R9k
FXtA582AT1CKTc0HCXVurumFYEG5tJ4luWn97UyKMx0/PbjdoOawRnEClXq9sSlw8OFYLEgGocea
V+DLt1t2HcgnBUMSnfbakYh5mOY0XcHBD1cDFwHQ9twCXgvqmmOOhGd+8E7RcqzxjkXhHxYR0+1n
y1fP29nTYePhuHF5L3/XVveTtOmrLYY9E7nscGbrRLZKq8zgt+Mb9FcTunaV4qNQM2+5yTsBOy5t
+GyAwMT0dsRECcjnt7wNsQJv6jieI390fK4O+8qKhJkwOKuJzx3QHOR2AN3Cb3TcX1BA0E7OlwSP
Vc9VqFgMZe+iL/uaKmpZyGnmK3iFs/gNmbkb8sDDmqEFYLvmutbqpyq7jbpDhiTqwlUyMlUOlXUN
njEDYWBznZvwL1ESWYN7do8y1eZckP8hPwMyLmUJbcZWqkrrAAKja9hQt+4Uvaz9pp1e7HHwWVkG
Eroq2O/CBoCqcQKJaxsOi84KEY2y8EzJw5R6i3R0a2JHn1LsSi0eeU3bkkYV4Jf4yQRQwJ5anqXS
Ns9XvmB40p5aQi5nESNfv7FlLpdV6YfnMCSn96yZJnPHcAaRo0NcNHDIW2T9eNsq9nDCOLco6oGJ
tN7CXySZtixJOUGMfjNdk/nLQuJEtjGS123/YQPmRwbfNhPtmB+E7nuBwNsvgppbpPB7cRfPInG9
xMtt5XzuxkCslcqp8zhwtWFe/lKjPfEVBM7z5knpgiKmAvY55ZXV8t96bDwgIG5pJaaElCvWzi6i
JKmxblOI0Jbq5wuMQvc5kJVZO0QUPgnsFKh0jOBy3WEMr/kp4wfSgvaZNtKciETkr0OgSI+LCcCU
EiWYbFm84b1PsGdi2gMrH9sn+DqBWyP+iCj2yVZueppHu5JCDdxnHmSep9c3h9caiyqfa/xI3uPh
g0xyg0LixPG0peOtXFw5Eihv3K9Z92Q7vAdRB4/UDF9du6nmhHQvkDUEbZcL1Y93mNZ+oRPQBQ7f
Mo3Z18IdtQHV2aJYJM/Y2m/sqD2heNKr0vcjrDElXV7gwhEGKAf8trDNLBo9uVnTCIC+F3M9Gxk1
XUmkcv6koy0kOf4SorgAHRRw4aoNQLJsvVabE3nMhnS3WVAoXC154J5DLSH2R+tznvePljXIbCjz
ifXSlID7GzsmARTauRXJpcR6Ogyh+oag/rNdVhTrLWCmt2KGUiPNHhO5V5DZRUbjbWo3b499WeZF
9OJfeTHcyOjAbLpX1Wjoojb127VbhPh78tLlz13NHkmmIdTF6LwbPzPI5CDxHorkLaAMJkdkgh3L
hnqQEiJoqVTwcHVj5kkUQ+wjkwHMSkHTtgvWwFQ8nDCr/5L9tt7CbuHCn9GMTdMfTMq+XooP/Paw
7tqu6415Tt0MJUklUFrwAEf8MvykVoaHsrkS24KoZQajj1PLQslk+Dp9mTT8Ng6ZVBC1r5C7ypKb
vYb1yJHPsqjRe6KpPvAunY/p2nncb3c1ADeVc/67Lh0eLh+HNiS5vKMWtvd9+J290zFeJaOMwGxL
cafjh7pIM24C8AVjwjH7h1MfPdspd78U+lGN23xbQ+a1wyen8dHvsjCRmYm9ESxSLMXOvVDqOcCT
qXjkLh3JkFCg3mjkF11mR1c4T3jGnds1fY5cXcqKCi2lCkKOO85c7HEhXOJX24i5Qtc3qEQUNtcc
nVVT5Rpk7t2SCiufOy+OjNs/pFdIwpDQm5LHsnR1Sc15zMQPp/IWJx+Z3ozqKZFg3FFryzWooXID
ralyqZ7lsMuNVhYogeR8p+npBwb59RXY4oOTh4u2SIOeD1ei9HfeoHi6gqrHgW2GRZkA97Qr1xhS
s+9idQ3TYIC/L+a38ZVaOq9kESq3zk8G5NBaM5wvmE60abaN/uu2+wHckjYlnPNKiimwOjSz9xYn
Wj3eLq+PUvL78/ex6hwIWE+V3hHWp6wnRgBeQO1npww94oC5JdPcmDeLa7HvQC2nN/KnRnrGT/9K
FirVREQxigjpLBgn9cW4ou9Mr5ShVt0d4bELzclLqrT5/qFUYiBrwdekpFSUApYRyr4V5MHiD5yY
XfRvIa9bqUZqGFSN2CtF36m8W3Zlk3ROj9qUmdtM2XVoUSXtKmqbDE2Px4aTx5aZyidnrtdXQ04T
Upb2+zixukPlayI/Zkm5ZeHwBigRMD37CnJ27x08bypC9zMQtBe8cqJZWDhcLbZhWceYn/Myzady
gMxF8vb5dPKDivlrHppFKzeTD6mQGzzqkmhcYNDLb7sUP12mGz63NZScktaPCz4Jt1o7Pi/SZZDo
VgBgXkPBkoSQ++djS7+XNm2Q9N0aUBLu0YjK4qGobHhjUwXNr/LBaB6x2PIcZmB2v7291CQ4K5rH
jLHmGY1rOJTLrEJT2XAs0c6WmYqKhcAd6DX3IIxiOc9iPljoUscf7xXkMgicL/sAc5UWtpLbjiBw
mqhYr9hfAmEFK6O1De0yTATJJinwEagvzSRMlrVTPZ18qqQClPOwhOmOmOHxKjBzX7d523IG6ZqK
G6KNyYkz+MNjxzFzBdCRiKGuXKii/MfIQ6o7vWfc7jWgChFGVoV5tXg/Czx+tX2BQuppEX0GyL+C
d+r2JeJtNA7FC3R8GSkb6lHy1ODF/IzqbOtcMFQxzJjWqnsnFDL33ng2oU6Xuc+OyCQT0ZAW5MqT
RlcXcy26HvRtD01XuxjM5RJwNIK9s3bLl1Bb1+Wc+MdpLiqsoMfEwo+VUJ3TgVYdcas09CbSKJaQ
1j+RiqX5Z/Q/sUzdxYu6GYQXzq9/yZxy59TVvUB2mbM0NiuViy2RwA96AsMQFV3fy6fvwE+/v6XO
I3HLIe7/eH7T27RMoW/L6JCDlDtSCDdYNwQiwbP8EWSnXbz/i3m+65/S6zvD/5m6cc9hywzLol18
/r8UudzNZWIWtG7vhN0EGYetcyJ/SwFiQeXu/t5eiPBX4rmzsARtm0ysmEugJOspLDl7hIKjsNdY
TqXtcnKwwiaknCnyiVys26AjwelWJmWcj+dExI/5bLmZ6inIiuIJGgKDdm+XomFHTjg7R6Aap4B0
i/enZ9ueNetPg+Fn/Ou+z6wn0uj9ygZZ+MAV/Rk7AXr0BPo9ee243VRSzDirVfhtcJ0EmQ60Obd/
yuLlI2vrLfSo07RnlN/BHVWRRH6tlK1bhFEdYlVHO7ks2iJKkIXQQGraewf0jpW1Y/kN5bXeo4Qj
T5EqUpC7/WOyatO62o0q1fFvMKNlnAl070UM7mbgOGcMtO8n2Dojqjp2pWIkhnr89Is/WT7HyI+Q
780caY7QaHAPCqK/cSvY8iKFWhlIqrlcvIcXzBdM3pY4SY+8wHV3dwMjh8Q95wWFI9N2pPEY5lgj
prHejNYzaRsmblkd2UUEgMvobAnPO5qid+/bSZlhQKx3gzpjorljkgIVRqVTPZSEG30IVRTn9un3
5upznmaSx+alAol95ljNB/paDvz04NbG6UJiqYsJII6gFZfbikfsPvLXD9m5aN80PL6cDLQigIuB
YMC/PvvNzInr7BxTEwOP9hVEaoclOGE3MzOgi8oTk8aG6+jT1J/nNNFpNvVrU1ofY/Nx/HaSl5Zy
RqREtzQC6IgV0jFSGiUPlOy4Q9d1+lZ7ngBPuHTDPTJHhrKXEWHwX3fKy7q1GVIiJenrwI7bu6ML
tE5ugIe/SMev2Q/L20J8hDl6dHPJTREbPD5mtjaAC54IYAdLXU4oFJLnVjxA/YfaHz5YLaLj4JDn
0BjYHqPLEuhO3DgK09IbtEZvgVkHLsvfcxwevYB59dYvImFKi97TSIZLZPjPVDDhMSMhJIjFOgva
IMPmrv2zYhnEf6aQoS2Gpf275OdBxRVFemCmqOFnOtw43GPrrYWo7chdkA4K9HgWK7t51uA1eHQs
CJcZQzXyhXRs2GWBBOkPSG2SIvZhJvIR5i79WgXzOpkBw37Wrugu0cpKemC5Vs5OJA0uV+xEkB6k
MGUcsQ90uAI8DUbU5mbb3bAayn222qgdGxP086tUUWrsmo/dzeEstrNaC2soZ2JxYEc8FUrdrUYL
LBBHPr/ZRFo4RYDDnLFkLvpcA4mCzNzbVUAO+GdNCt1Eunchnx+VYOhs/BZM/J2cJFCQOxMzPVdL
QT9FYIUL46A/YVQ04FFKKp0HWKl3Yy9VfY4mD4j2LQLIVsG+CZGSj9KtJbsZnz/IMkW5+soY80nI
3bOBQJ2qg3ys/rWVCRtjN19R35d5AozetWQUxn8IcfSTxHoHGtBJrwSTt1iLoanWNxn1eky3Fi1j
hJUOHePZWV6FKahy6FAIDjzZGFx4z8ndlU1gl/patY0+Vep61bJSN3ZlvtX0l98wAIw+0xjDmVjv
tae/HFizu82tcldyJ8xKdyxQc29u45sdGPFW7249bx0QSABwsp8xJ2LogWyAJWACfVMNOvtjFRzM
hRrKC6yBQXCyLu7vUNEXahRfoF72qXg7d56y9GgPYSPK+i5MYqBhQYmrAxA/Ww2Tgs9L8O8Cfwj+
WXxt7ertQ1J2r1odtH/cao8ILdKlVrhQFirU8MLeEy8zrCYOgeAUAnV6su9unC/AplfpbfUVlC28
oq554WfoPSVRdtyjRHAxndUcdJK1KyUzHVka50SkuyKVPwoEV3F2c2++4u3pu/eHFSFitxK4YEuW
K2m+OQ+O570YAX8GzkGorm6iuu5nnpoWcGYrtYcipqZ8j81zPHF+x/vFLawyvjMyR633NEvq6wPE
zoqnpbMy/+ephZbgq+/NWn1vRgA+iUqwd3srQxrowyNOBU4EaDDFRBdQcxYBrwJTRsTIGD7Ieyq/
QzR1Bi17BEiCuWQCysKvdp+qt3ukmIgjVzwZI0jgREWDrNARALdXtxeg6zpJ4a6uC0nBv0HHzsKd
3DAl3xN75BkM96qHzl/COcJnuP+N8N/fK8NInTguffkrcX/hgcu1Zfiwhlf2srON9EChzvtaw1JF
yWPZAeY5CjUQgNUtUWAXCw8PjxWYJwRTrgcgT0nl0shsRRfWnnk8YiRbd1B6zVdKAo26ciDrwLVX
aqRC7fYvEFYPLzBgxE3/1oKu5Imep1Zax9n2+3RHHLdq24LsOXoaKkdEi9fBPsozWx2ceDZDsDlv
noOyd8iL+xNX3ifW53puZ3gd4lmSU8C73Ezs58dBZ4k7Ii6nRKehCfsLcalQhXSKYLO5++9Hb1by
H9T+HYBKsvVv8VTQ19xhOvbATOpPDljiOFCQCOEzoAwQgJyMKcsfHhH6pnmul8ePFu4oK0DELhXo
EHdjmFEv/uxsKD+UQKCzVMC6ik1UoGNLlL44xDtpHzKlkmDCFhOa48fPRqS7HV/RpApbhJLBBNa2
HhSjdd113SPGIkmMAoDUMnG0CAwbXW7MAHhk4zsIyMuUBECYzI71KZapgqloioZxwuCUM0Pkc310
jZH4UHtoZ8zO4bq24okpfl665+ZXq8ugBSfvVZdUCJggFdspFa6VWliN3CK++BohZfsAxW9hoC2j
TE56GKnYquSIonx21SxR29YkDrlzjbRw2CH+i5+A/r0zljq0awqZnqj+i0hWZ4vP+99isrhY0RzQ
NRJcgKwM+zC51Wu1EBPq6G+xkysLxLAUw0U98KkwX2W6XndOzYSC6EWENZcrJexp8UJp70KRjajr
4RZbBkdQ+kT6vWOEV+4ylF1C4xSVyEVwSNZCjvtQ40CA8B7BZkykF+seqWn+4Id/qj6EGdwidx3q
B+sBQsVq5nPZW+NThmYHDdwSa327rFU29XQF0xJwKAfp6H9baRQ/LrldKUSzFh9M1wV3pZrd/SwI
H2+ZV3RdxJ+IcybHB+hSH20pXx9Ih7B/o0x8pSEmNN9wKwFJapStW0PdvB0NJ0I59H+3yY/J5zRv
0kUTipGX45qBnCQHLCQGvz+HzGf9HTCdJuabcCQAy4X3YRYVxF4aWyeQEzWIleZmedaN3KBsQmgW
iBikfrl20JXrsOQIQktX4LhBdQCAA3LlpdDvqt7fT92Tkr2ZoiLGojCKrUyVLO1uhY6Sb6kI3qQw
Di4RNri9X2xZgk/nDxp4VU1YEtK8R3L9d6Wgx0rmzMdNEs58w8uqa6LGu05nkKX6rR84QFBFD9mn
WX0nUgvKtmPUN90pma+7xC9rCBhWXCUsFVf8x/WwERwDy78JzKtQD1WAGTMEBKTly+p4xvkBxg8Q
Jx9yt0LMUhpgrvJW2ZnO1VVD4EiLnaFaSD0wfbxAFZa/J6C1KjCo4rq3VEpc/MLsrKU8HfxVlQwN
Eem6iqfuaIjzthVihS+xt9RJszpnCop4Qa3MH6DcdD15N4VO1X38GZ8Spy2EyX+tkHvSrLS0lWpc
P10D89fbUG7Ja/6CSLJ0wwpq21SZ9LoJuQsb8V9ZRlaHLH2zUIyczkhQWivnU5A1y9sp4gAZhZ7W
8fNYL0zabhJXIHNTz9YQyfS6Eq0mSCpG8uWMF7tSaEpcjXTi65hITf72tw6kN07G9NcanSTjGGIS
8i+IGVKpL9jPQZStyEvYCY/jvxJKBMGARC2emtVC2mr3n8tauw9IJ+1skGq1pywcgNJRK+e6hNzQ
lXYQX+W1h42W+d9oIPtzXM/+i3LNr1TZqtm7GiIUyc9hV/9EpWVqUag3l5OzTC7gkr2j2pi4Fy++
Wcwkih08moTL1D6177Rg0oWiCg4HqGjFlLuaoIFQzeE/eETOgpyJKeMshvRe6DhqwEZzMSowQttG
WUfAukBRIBtmmlOLexYXpA9p+VAmidV3i7Fa9ymb9MrWo4TVO0RSbJPcxahFq083rZm+aFpZlGEk
HaXVeXC8bMRFry6AYLj3f8AEUfZMl79RldMG3aqlW+9IautzL5uvIFCEk3Vvx0azP/qCGem6Sz9F
achvvjpjHsVN6ZIAcgXGKB56lNX9WItclwx8EBmoMJHYofr/1/xCDE32DexKCa/pp69GZ+mOMC4i
n3bF7LFObuXWmLreSsCtjV9+IpCWmuHl3Qq1ZUkw/RuEhNH/phERrhUdbk8P+DqovTx/FBf58hH6
gW5vo6XRQCki2KmWv6U5utQV7r4kyRQqWXrvwqj5D0xjrNLawnLppXekirrJ/O+W+oUggQIDDOUc
Q5RtX6lFmUSC64kBY5nERlUn024SMW1ya7/t5PD1V7dJ8Wx+3aSphddPSKrC+NnLNR+xFNavly0Z
A6gsBk8lc0lJb8ij/kJ53YjRpVUFIJC8zF4TY7LR7xhlmL+qzmCkpnv3XQg5sf0xcFWA/9DjWXuL
BzNQ3ujjiByduD4mojXFZWQPo+t9YoahMq5OBMlLuTXUwtTzFWrbiynAsDY3WW9AODpEtuqwSigZ
aE6KaxknLQjE3tWBkGC4MIxculbxUekuxqmZEyfsCLACCSO7An10kGniZjfOx36/1spuuFeEsl57
hrm4Y/DaCQvaSXMh5d96DAE6YngKOvJZOpHpQlO631zgnJ8pekO5XepfTCPFbI6YhyY4gGD0+v+j
QmqNn/1yVVXklujYWGcNlhT7sk5vUqIsgPfxSIQwutoZCBmNZDs60ScojrrP0hCfiNJjYNv2EITg
4+ri0PnAeUr9EOwpuHSfb4rSgQKQgBDDZJx1zULITr5TcreoryVY3Xqr/1SwaGb8mXLQv3qdeF8p
orfQObasCE2RTHGw9je8P901KCmzw+qaUQTbZ+ERNa0S2Y1xk4NUrDeqHWIzhxmkrOP3uT+8RCF/
rPqIOZnPSI+xTy/WWacuEJBD0ZGEuJEzFS0p3F/J0k1TXfXdLe0UQ04fejmYsjaSwbF7qYOnWkzD
+WBNa7klFlBH1V8wqCtddzQ1WlTiKDufjCCTulksIzZ9xpkdHMDjgx2pIr0pw9qZNElknSVKU97a
Vl+vOsLc2144+P7h6OUnptOjvx1gHvx9UBz3lQ1Dn5ATOhii2/UcmOie/lMFdXyGnTN9wG4w1zND
F/SVTQdgbwjp4hgas4oBI2w90XEY0R5XcqHHCLI2LGVieiaSZ0b1sk2Ui3xH2MhwEu7UtJdc69F3
WdaiHiw7xttsebsltlrXJLHgnmEox7TUD7Ie5KGs5aF9ec81TBAYQP2GEHEeE4+NG1g3fs4g3As/
F63ZeO2AQtXjYprk0orBSu7UhvSlAESl48c7l514NC6c6dlho08IVyZAKv9pC681NlSmANRRt5Fi
gRDfR6e833cb4QM/CBqErmdpPwAfWAe9Em4KnTEa4sa6F2BAUrzZmJ37yjZtLq7Q2UufIGzCAHNf
ML+GuBng39sk0Dv53ErY9yoiX5X5Nu7uTyrx2tHy64HMMs9TPtmxi5fieNlTK2jnrpPcn858WES7
O3x8yjarB2ZBEDGbFt+NLLpIzkD5eC2UXgxIlORfPONDd8HcID1tlZWk3NfqeJKORf01w/mMxIZa
jOtMXj/SbIRuvslnJtOPg5UPChOl/i7aDRttb4PTJI523Pa3a0/lKLalrGRiYGncsfYMy2ztkEWO
YKa/Q36POAL2xJK6/KTzmU4yMlSn6uRIUj0YM1RtaBbvo5DoC4WgTXS1EtR1Ya+WlS/hYr6E5mRw
/X+zYrfWLyv2e9kaQk8H66agQsaoEyFpxGZ281bxVqCnlihM26TaX3NvVD3upFMS2KFgaekD8VDs
sx/2zxZ8VzRc2ug32uLg3s5zPMN6d3FjJ/eUtZ+osEaWb7bdtxu32s3IwCFvBg7rP6AC8SoVtF2L
rhCtHEWUBAl5IitMKhT6WXxsROzfEJVSxdA75d/+H1FtvCgu+h06hiIMvSJHspju1QIcrO4I1h3i
5Mrx6AbldQcyZkedTczTOMwH6Rm5ZWgEZ+lZ7WtEAmBivY+lfBb+Lk3ar76cQpCcrNT2+t6kFjNZ
M/bZAzYFjxTTsc+9YQiqfu9+3Av97wRjRHrXdEZYMCcj9Geiis854R4jzZApbgTVMG52j1yK88r0
zFpX60W0ykMs8imICt3+3PfyhCYhEE1DcraYyTOCm462Hz5BLPvmPAH5ymNI5friey+LpD/m2icY
/xt2RaVi8G3Q/r13DrGG9Q3pY9cGA4Tbiuhj3q0516OhMlNyG5+TjMUZ4EQIdvgn3tveDbR75WFl
0RzQeCT9mp1BKKdcA9CKshankZTqUlKaQs04J+QEOKadjnONxs3EAfLcOoKqN0IjuqleTrXNNMmK
94ckNr4EiYHeHTY5HCZqSfhJ0bOPVftvxeuO1EChrgIPY2y5XF+9v1myNA8UAdQrjFr5vELyrgFM
Qr11CrExZN+w9b+ZOIFFCGymF7BIK9khWRXfvel2XnRJgIPo0tFJH01oX1rvi4XYhyC/N8CqvUK0
nX0R75RQoCumG1ifHOul3d+QLmwcc9E+h4Lcb/RD4s0Dq18O0rwAP76wNIOARkGiMltPO6J7lDGQ
3yUWXm4OFdga3iSIP5SVVpbtLkvYB43pu2ZCLmMFhDqpvSHrCws91qALwB82otmbg4shCGg33VaB
7MjPLeA3GIjkZXq+oMN+WDMv5M4ocndvSIS4GTGascEsAZIFLgbzf5ZKD5JstXbD4ZlxR3p7mHjq
7xmJJZaHYH9x2Os4BEZfDXCWj91kvhWvAAyyjPLhYPq1F2BXJ5FdueIU7d9nw2JPUM2KOIYh6/9P
eza8XHDdBqS9kMhfYD4tf14P+DbhvE23Pr7HqPONEpkId1WgLSel/BPNQv6ZgSbo7khg6ZPkckzn
RE7JGdd2hyyvekuJvG/DLy41a8v8OGrdMn5y7dS/8ppSoF//wWqV81DeLhTwvGXJd/qPh7YKkX5h
eYxFhyG6F6QW1R9Haaa/NYBhe6qOPlCI17iXcFQ6PRwbU8Rq8jQkPQdEnQsw8YmDDO00O6SNL4OE
lvCxkw29sRq4yNuHiq3nhO3myv+0PtNBhZzCx3/U2FlL9DXi248ltZvs5S0tQkW8qHFRJcTvlRwK
yqh/xMQnZUEfRIlk4xFeELdAeLZ6/ekhOAf5w1f/20v9FoRTtwu4lfVpKQkh0DeMTKIBA8WYsPSt
zN6L51loMY/Vej09sKo4aLMWHBofCwJUG+AAMTU4OF7SyBeLkL61ImLmsY9NFlBMuDBrtRZInfga
X/ey3SW5lxCUkyOiPP5XsHswpI9ZMHDf96JZsaAKNY+fmE6CLjS5prX8Zjbec8lY5LnJk7WRUELY
TUw5+OO3KOJFZDd+4jBlWyHZGjhu3LRdjvmZ6wdftk6AoGPu9Ob5VtfcBebcvSI6/cecMBOA59wb
o7mQUSuCqvCw3/NsRFiBTw0hyYz8zTcitSKfjSv5b4OErn8KvAGoXSgRB4tDTHtf7l/5wcqox7Fh
VuxzAxSR/u/ODlNyU3oYPyZEH3NJ1qD4NGwCbu/P+75g7ebjHC/6V9v0rSFLlnNTsF9O8Kemsqz3
tTAgFmiRXQ7B2mSxHHGumjfFeogwjHnHvGXdP5xLEfXN1hdZzfmypyxPh/RaKllXFcGWSP4aHTDm
9XYWnFSQmfPTdUfe5uH3PtGdAKdsCfprVQ6MoyijOhSOBfEPBuMZN9L5hi1B2VQZbWXynGokmKXx
YB7Z5STctQywoilN7FyreowY3VUHcLn67rPY7GjR3zday6uGQ6ZZBWdNH/5d3wgBtvCIyd5UmMwQ
K8aLlp11Q5aY4mBCpZcvH9uyOSY4qBN6ZszuZZYHSvlYf2NcwdmSev5GmGuyjPeRUjNa/mYsqTRc
echdTy+3/ArWqBsdC5wOPLJjuaeIg53jXRFotySvTZcQSvWbMqCXgd6hrw76CVFW0H2U6tW2hyPA
hTwHuFHHIVr/tT9QSM4FvWPmRlfinzpl8K7dnjmHZiJEj//PHCGpeqymphVy02uhK+brz6hqtMz0
CmMPZlF5O+gvm//ZvJlCh0XgZfnUXSDBorNGww0XiOHyqS6+EuVkZ+GK8DlxW8oEPI1KzKaGXPkY
iy8C01IwKv3uDT1qDfz/7HPLqtynaWWhUOftuWgvljxNKDfeXR4taBXBrq7/rd5jHQqdiee17uDd
AY3b/4ZUz3BiHo6paKjT/FhJ79BefN593TfUcxGTlcpyXa4N3khqsebYtKK0DwEMfkLKUftYfKAs
Ijw2cIIy64IT6TFrgca4HJvXe11TPD50VoqXhaeIL3nTJDhr59N3LIpQ7sInV7sCoJbXjFNwbOr5
tS9bcwAycXPUfKDuPC2bjU9ae7st9jpkjpCaTWcBEO9vLBpLQ2t/KPCPysJ4q9sSQUi9tN7rH1GE
7WUHic3TrHLX906gZjEofo1O6hlHP4ueW+YNgmlIRX+igyC0SPQN3jUNIItzDJ0I3TfIlpry2IGj
lupp2CgyxkMGWoghAvUOGYTaVQv5yTGRkRwSZEM5I5QB8ipAoeNvqJiyiIoojWlLyUHT8S1/8vTM
HdoBcgez7zSWQB2RWqBZdlCVVW2Apq0gWBFpKx9Pc0tDxyL+w2SWLIXalhLAEhS+6I5xoTRdz5HG
POqZJ8z3VRK7Rgkuzf5tOSL5GBsh+AWtelA7mi9iTAPgGnFTtSDEjoHzV38FttfC3Sg10t2qxWpC
KQMViR8cA4Kyrv6iUILzIRUQh+vQ0vYxWMkOHTGNx8xFPZ1sdoyhtRnhqb9bqBisjpXB81lwEHWp
CVsTQrG5EZOcXK07zGlC1Uh1MIBeRhajYMkmf+dQsFsNbq3ZjjWTdv9vJqa3mfUokS+9D4edRHPg
fssA1sRs6MzWyzyiBREftJe9SRfzvLIhqXL2nkW2xFhZoMwu5wQVDM0sAhpIHANN3AwMYaHZSQec
XvkrGnb0ywUSoA55K+IYkXtjBgWPdmOh9Rp4MmgZW0Xl2s5gbHV5hk9iNQRewD49BKAL55ktfBlD
l0GMYg5BCOO/FnNQhdMBioH1eG0hCJa1k9rJKIzzVv4mx2d5obB+JYzkBWzCar+ZZJZNumptFxPd
QmT+BUQZZRKJB/0D2dKnquEFiW+rWFouLi6W3GCSsdlN2YjSbSXU+d6RXJMS99IkD1Yn9Shd43Gj
19lFucQtgFaMuJjWE0hHs3OSTFvXnuGTs8y+XobiKvbA9hzDW0GTcr8jgyPSIh/topjvpAwDpAKU
xGy/KahhlZIobVFSHUXoMNbJnmh5YXJryJBAQ/kftbIp9x9c/uK5VxzBp0X8OK8PVOQyByBkfQx3
7WSda8lZb5M56h4xprpBEBmc0h/+8+Rv+6jdIgc0WRywbdxiDc+9WgJDYYvHRRprLlX6xiddZBYO
m6573EExBtk80lYgmxTkLBBIj5bE5f4YZa+Ubs6pXTKAO+OJ9Qcf7y9J1n2+OxWiIN5PF4ODH+uT
P35aJPXEL4gxD3vlVIEgW0pDD1a+2nNGMHgQwuM2GY5p2pUTKNVDWdOCPjTGoW7HfKl2xhHdrpQ+
6LuAbo4NhsFCPSiQh9W+Hz7j66yR+o5K3OCRraE3AsQ05brVi2oxTHmnQMZ6DgWufH1IZyuqYrG6
KcfaBgcsHc13OKTJ/OgWU+nNOI+4Ly0hCM6emruURYveN3fyDs6GzUSZNa9AMF0WEpfNzGxjFq7o
N10QStMnkbzcRdu+ti3x+1SlVRG0Ab+UENwNYko/B+UiMpSqAj2xzH9xFkvoAb0sHuzKBjVgpTrq
OAZicnti0gK0Vh2FsuRxORIXJNwYtkKNPFQd8Ap11N8HecDoBa4C6VPhmh9EIrxNo8RDpuOFRbBR
H7wtyKC/ad1fC4oiSFrHMJ+/rKauJKdg3Jke8ZkInQQj4hFxZ2N0j721/W5FRregEg5aEOOzkAGv
WAMemLxXkX73rMSStydPTBXhzFq+DucEIMKKeqilp3G7VuFwGt0XoBcKGoX1vhdiWNsVKACXBnaw
UyyaYGqW9c+w4siTXDh+Qad7QWsmc97NDt8FGmEk7ewge5s4nQ7IoHQjyxzU093S2UbtzjYYFGB2
Uz3ZqpqqAIt0ldi3mG59Zpnetp/uuFNRkJcFqZcqeHxezKhLwms+qUpoF/c7q85Lcw2dhOLPr6Hx
3nhtDc06IcVpX2PjmPnZFQPBPcBLrPdMR1a7I8o6ziHp3muUPjiS0rVuMD0MbjgBuWMBkCS943C7
FLzb2/+70mlRmlfSOUpzj2travThemjc+gVFezzkdTnLTL2uo8COyQGyKWBilOJDs0EoIniLxhb8
FJVbvgQXm7fZksSRPb+4ZDYu9hR3P+FBFxR918SzA4Lgs1DiKB/XOM1XuLcHZXtGhao64vFBs2Y5
in9w7KBjteaSQT5EwcKjVWX1Y0qaxsit/2Yn3tQDqLW3fhGRG1TUmBGCUFpvdhUaTwu6GazuAqdX
mdtPsGRgbS5CyfcALHUSx7lClXHAfFAfOv8300Fty58RS7TqXvDWlQykIjlxShs9XWeXNOqnXTWZ
OUtwxM7rTipSDNi1zNL/p59jrres6T6IV68hxzOt16BI9FYEZZJWQHvcU+5vgXyw/Y4ygFAPdDfA
QrtvffFgXrWkETYDMWx6hC2zwO7qAQD8eybVq7lW1OuJFA14nrZl+pCI/C9TZffEkT2QZUvEDT4L
3FEl8Y/z4Y4wy2zkaCtP5KQCB782chZIL3Sp+mAt1H9C21gbW8P0mZFilu4Tw/am3DYRvZlhOzDg
am5HUZL3KSZfCipDbmjGxaUkXeI08fhOFYlO6s7jIiWcMo3F2IUhCRb0OmOBYac3rEsKuGvPcEzH
VbIYy0DYTCzmpvhcwcaTttz0clWK09IRcJdWisRKwSByU7EGRoSWFwbNjkfOSiSm6oAcLxooay6S
9I+3blHGemGwLHNSXJV095RTHZB9cFm4QenK5RjP1v+0eR+oSExabN9W50BQGduxleOv5P9OTST4
TWIH97syhPW5o8EvTl97bbcpDpHPo+Hy+NLskmxj4yC/XPayUS5OWrYApuhuj6poKa0F9cN6FYVS
mqaN/MlPDeJVVGq/PSOLZuTJdcWmxeScyeDUwSehmDZAgVM4aOyorAYZIh1LDbgjQgHnMRcigtv9
Ikjd19lCfwatBaCWooRc8M2SItxAJeTIEnLgbnponj2hhLy/2KY0xzgPGVbU+PuZwgUTG5jYphSn
HRYR2n4m+FgI/TgOBizrLH6FmOhUXyrO+hew4JQPHeS4NQkOXH3PaueXH8dTUMizcEaY0pjPWwMy
XLAhyCZQZoWoHcVdYupPWWSWbB7aGkTRoCUoc6YlgWRs5xkyXQWRAwjFn7BBCeAGWTp36p27qW49
9SNde9dEL2KwXUEd9nxICOU3wCofLxU7J9dCGzZ6xqxadfHtDLDuGpEFUiiyGRSfFvx4wh+qZQ6k
mRGs3aCQXDFpcw8fc21asYm3IRNJmjb/LbNeOVCAPITNnAahTvirXp5C1xqlEvpnPsUwP/xlpXoI
ttCZWTzZ+3AnBIKnmK7djaUaoiYISQk6v+f/cM7TpuPzuaeSkNp/+r5G0uTEfPPrptxfSzWeUZpt
5NrpgZvoP3O2sc72RkO0mE/qJfwvBm6x5ehHhGizQNRn6zEsmpKJWqFCjC5MN9zN9WBttl0d0EUA
cD8bYG48Q0fxK82fOHv/HUTRn3M691p2voMg0z0ZrwnQSI9vS3MoOX/DrtYUks3GOj7dNXPhSygQ
Wtbmw7JEo7p8G6KtiteNAQ2d6rL+XwO1z+/Nrd+NTUP3W36icIV/fNG/PjXQF/QeCFfPvd4/YHKA
/fWrhS2sU2M1N0Ks+DdcsJnghKbTAFDLXkzPQ66IWuRzHdtCOqgZVl4HkSTzWseymXqyoU7HNFc8
gRjQgaISkDWTpgHJEwlGv6VBfpcpUUX9yyUooF86sZdVqtgQbO5OuRrphoOtsPkTW40BXTnvnGcc
CjNA1pCNGiHoUxBhqgnb6y26P2I/cayGcuKzepWDGTRyVcVokL2Ci161mYiqQ75rH+mEKpqhetIT
5OWRY1HFqmzA32KDawlpalJW/8814fgX2UvYplJLhEnBYdoPQhwkg9L2YJNH7OZvEYgBt8vxN/jE
ZMy5zxtMJfBB8c0zOsdK5mmj5oiYrF2UgmagqNMYKwwXfE4jdFIPnZOAHltRPRgRpOUeauKvmMyK
yDezsV6r6ANwhMAAMiZUkUqra6fwxsioepBDga4tRyQx9t81OTEPCQmrCSrVndmGah3Kd1UYKmOp
83VbiO9l9Ezwr1jRU7dm28G2NXeYnxxT1v6n9d/xpsnm/eBK4cH9w0U/LawxXnTUF3xBk4HgZmad
+6ikezNXdUPJqw+Y8fQMWj8tgj+ZQG5aVByQROLTHSm1v4O5CXHSHi6pJeAi31VuZleDEvYSBTNO
XIfeQfPC9J+NZR82XxzkWOI4E9GJ9Tc3PvsHlz/SgqmvhluIEgnK8kPPWr83oi6VQ1Bq+LzK2n1Y
YwmDyao8xUib47z24hgMwU+0gUQfLq3Toy5gPs3QvkskK1MSHiJtsKD3AuXjScNLUDlD7cxgebE+
OJaLL7Tw0e5wDoPlT3TlLmua3UjisIjfxMk/KLuqaaq6DchRMaHVwwNMplF4272+uNqldxTWs6yO
fKxoFcBEnXl3uySGPj3wi+r6sWXroSsixFZwK0FwogB/ip71TZXLTWATBQNDpwspCwyOWYbMDvNf
stv+rtfa/Yl7yqWisdZfkI/2XrBFEL9r4h1efCsTyHNbx79d8VY7pRYzkcnYS9i/744+AtKXq+XC
bdDPtl3IYXc10YyXU7JDZhIFLWLahyXgBdFkvLedDQQGC4gubmnmbEDkZBqgsLTbdF3UozVM17N7
wDkxUBDGc6l9q2Z8UX/dlJoIHpFmPkHMPLLeOyYyisAsPrVo0BTLTjOL0GEpLXaxyWP5QfRYss0A
X9tVBBBxvqSnkUAKtzPm90L3Yec0GpQpySrDPHA+WSoMsq3IfsPHZuWlzLNsZWBvtQmZG2mciSv5
j67xRGf0kDjl0Yeb/DpWywIFCgf/lWVRnNHaY4Wp3EpJV2EpyhjkIK0h1rZ2+SiKSw8XvivCuMhV
YJ923flCaExws/QyvMcvFxbATuHIEASn0evPU/zD3VjejT43ie2avQkwvh2jNgd2vc0GonW64Rfg
cumUed5LTgVTaKxxJFh4HTFaSOSK3yb8iArvrDgJvbLD5AtmI0/HW4+IftSvBoJtCPJn1QB8rKYo
UWGsB2rrgK9Mu3IOn1A45F63WexUXId1uq8gV73XUUeCIyBSep/7MVag2bo4ZIaab3PadioIeosg
SKG6ml3tAXpj5V+FFk0AnjYuIH74Y0kpFyUCuMTZ+4UkG8tV+uBcsXUY2zb/ZJSmT9hXnHiljrZo
YTsC6I6nZ6A4s+mIaQ/hfiryYogfpn4keC2/GULQYNQuGsLF+na4FVzSEVJgj/DDFMGmHKfZ41kT
hU0h486y7QFhIAfSYHbwkUHzah4X4Q8MIgNwhP49QMNke+mGwEJ5noTgbBJctTsbsG5lrx0kft6s
hUFzj7YFDqHb0dOBpLvwu4t1YIVqQe/7WRJtJKjLlSu8+COYV9IwTbpPVRYyQq0VgC79tpgWdHVN
AaPKROXagn8F0ofZS06zzTRshHdkRdPQp90sOgXplPQkt9/7QsckBsM1p8aXp/fa2/4cvxaNK+Fp
FzSwaZJTEfvetdSIh3ywJ5copRofZu9JvNIl29jUqyMFNc28rSPOmM9W5PojVt/CjaxS0R6Ttl0l
Y+xTxSZm6y105k4f8IrxJYMjZ3aWeY57aZubGl2ReT5M8sJX7y/uAzKXCH+1D1YGCJTafKG3cRgx
TRT+kX6nSl+O1VT9UvYyurLPUsk4vCrV2MS5CYrg0pxdvn8h9oFLrsVmBR5rKYS4LXEPBcUn5x0C
ZqbjXWTrrSMzcwbqyHv/HAybYLMYuJ9lu+uDjTxQllJHtSvtGqxoiO3KY0/sJANeJ7vEymTkJAfp
J3dv+ewERdFEiiyJSCd2IvnmRT9eKpnWHrf4+989TVebxIbDHw3jlkm+dythtv6zdRm1PxSM9Aom
RZG44IBrJ7JiJUDZ4UdZiFzdf3uJbUrExxxPTwjqkbNA5HE9hHWJU/fnwd7nA6buBH/XILtRFBAX
yNeMJ24PIoL/FOptLdcIrZgbWtR67Vru7zsmMncKJEqhm8RL71wriSC1t1GJObwEa5vT6Y1Gr7YD
IbwQmMrPPBF06M6nCqMm9cPzZ9eyLreqW/AJSDdY4HCxMILI52MrcEnWpk9/IVOtf1f9Vmi5QarZ
CaaIwXJIeCzo+eFA6UA9qBm1IRtmW2P9RHGEECalJRzoXSW01VUM8TupzZBMTQpp/mfDs/MuP6Ni
deRXDdt+ft9ljDb5RCpUhaJnXrEIUpTubjP9vlOOptNzzMqECKLbm8zmQYD4AjgeYqusl/PEZy3i
/QueMq7VBqj7Ic58RouA+fg4XT8pigmXvGOTmwkMo18y29oG63aGlxJ9C7esD93/gX+OrG1APuUc
aI/CHI5zfpBZft8BqIPm/Hv47qdh05kD+PQAoU1WkyNK7Cnwxp3qgXSgDEWdQ1/7lr2t0AfXIT/n
0E3AP72WAKyuet7DhUCdbnA4R4j961yTmU1AfBXvgnpXfrKPPQjvenHFkMsjdsU89vsxt4IxbQLx
upx+xqYcGP5ecG79JyET5vpyOS6L/0edxIDh5pGFS/4G6TznysHmgwwI9Z5KA2zDxeRWi7DKThtY
waVxulUE57+lHXTAfErZJbaoSAqAQvWEQGE7lAkiMCA+s02wCj5wBqON2PFNMDbUZRcy/uEMvrZ6
8jRq+isGqXYSRfYWIvyxTcCbwps86b5+a0k+iuu9+okh/9uWVQiB0Ds1zNiffvpXQmHZjoIOMxFE
CXXDnaDMQECu0SVus/N9SnSjuD4CCqCq8Sp2mJwpQ3SffCAwbI39tNFeGf1mTME8YO4KrfMeeebz
dLQegX7vyM/JW2sdDWwccpJWHzqKkH34DP7aL2tvZtqhydLLdozq3+XgZ53aLQZlTnswDTLVVzsJ
T2OBX8nQJmiWaXYb7evPbc0l5aXMPRgzxeT8rNBxzk2nJTKN8rXI6lNzYjq4+5LqesZv2aUVzG2n
7OvpmMbkArs2KcPftaldgn4DEi3omLCKOvkCTZCGbXquWPywsEGRHL4A24+2CFtLbmHVG1cqB9tA
LThkVmd6c5RL+Asy/F1Dpsj2j+IgUwv4rM1pY7Kte4WK2S0pIbN+Bp7YGRniumLHli521htO4Q6g
jW7z+u6Z3T6d/foZcPSTlct1BbKYmkiMVRdMZVh4276gF+y5BCdTA4JbCJ1vrIXUrFVYPjo1rvuf
R/p50MocGi3S7Elo0FAbQ3Bf7NxBt18rvA/w4J4SF2gKjo1EHCvLrD8iDQ/BXBtNVFGW6qkR9pzs
+vuYmCPxXqfJ7IWQQauEc052czk90rxvqCZEDNanwLimE+fRQtvIHl4FRnlOGgMuOgSeGGkd9/Lm
rG9NJMWa0kqTqKlSB9ZfCeSfTg4cl5w9/+v+06jRVTd+h4rBvUDOl8jV8X20yYWbRGzdsCUxfN2c
tLHD9pz68omv0P6+UbZmFqJye9JIk/u9rCCoW2Cd9ITiZW9FRp/G9ybqcfkywAaMOHUBUehXSo7z
nWm/3IyTPzAT1Nkp3ps1g8jMJvpPELy0mBY9WVbkDnGjS41nxENtjSiJ7q08Ztn1dAKFb1dp8PFg
lCecX6QUXSjlnmkoVv0AOPVlzD2NZDwoan2bggbPXJiEueK6XHqV7KIa1+tmNUjVQkLZGhpu4fMG
Djn/RIoj0ty/Etv2nRf5VwrEkf0E8xxwRR9DXn5xpn+nkRwfG18RudZwiR8w+BdvlMzs2b6k3b5w
UBpPicDVmsSDs+78wmg9GPPgN1Yp4Ko7Xe1/+vlZGfUURs+t6ph/qVPjcpaN4ZjaiNBb9DlI8/cz
lul0uszar0wsw3FTkJPszGluFdfnOSLVehwHgRvyUryA8E6RoWqd8AK5+Be0s3EGvglF1yuf0r17
VHbXOX6oUpvS4OLfVzK+d6Rannf80Wd8KaPLUjOEDVv1iR1XLv06y/FVq1zC7vQ8Pr9llOLUqB7C
/T91pIs3i74Z5Lr75TgR0450LXnSSTF1fLvzApAxMqRDHB+c4S8tTYR5uc18VUBGH3CEhpOe48W1
2iI1WEqxyjEEAaOTuv7pVEYzqj64jfSmwcmtfu6NP0BJcbRrUzLYvReovF0lWLLqfwFmV+QSVD6p
1s4d9xroosQRbgGOX24bo6GC8BC2PKrzs+W1t/LnUSQwekP+T7ASytNBnoH9Ep4rQ1P60AWGaQlw
qFU3P96POzY7KyTeejzf0F/NfHRYyELdoLiOdP/IFboIQKQ2Ab8B+hznQpHT2Ek6rk42+m9U7McK
5H0MkGtc48R5ZIQOA1uPkPbjwTRb87ozdUvRLvLxUel8b8en0srebMCzjxYheeqIqF48BaF1gXNi
IuHkc8IB8K3LMwtNJmjYLLXuQ04NKeUzK1cKtN332D+ywxTQdNi/uyKeg2m3fDYm8c9EaEpdbPhM
xKwZxZ6GuCdFpoaOsOTSzSXQVYZsfRJe0SMMtXnsrdn1MqV9mIq4DJ0yhz0C4vU4YtAyWBnfcvxk
ajQchQDNjDtXq4yV9Oumf2Jn+JL5ptWw5XFQhlfsN+Cr51bt5vo+sYe4/STjVd7OHbfvPsqIZ2nY
Yf8f5EUbaKcRsvB1fcol5k416RTvdI1VElU15BLWwRnl5WHf2JEOT0TOgLZDC52GmYgKu6QQdwlC
3MzRbMwRPfVUxhId0Y34ER8J3SD7xAgTl74eLjeigFeCi+vQHRLgiFyC4lBK+K46Jd/SGjzakJMe
1ekJWa922YqUyb9mf05szRS9IlHv+6hySlv7wXv8cE0G/ZYv1A08n+zZcDpWvpRSw8AMLbOJHTIY
S9MMoxKIUW3/hqhCueCKBgGBYXpeLrd0xeV6dCemwhoWkiMJdLFYDUCcH+GaPqrioi4fflTYyIyp
mFKV1q4e0rtd9HtQ2mtDKFnDXbdJKC8LsRw2dhXv1lJ8L3dcZL+Z0d077+rPtGjbgAeL+8WdHUmW
pKQYiRgoiSil42CUHLcCKweQ6fKe1iLLnmve7382xtAT/wGpGnwcjC1JJGaJfyCNeP3R08AK6Xc6
Ja7FkT5xVg0gSjEKbposULYdAFduHizB3C/UY5fSxTNbYzxVZUa1tBHM4p/JVA6hfItqBLiCUvPP
+gGfjWmLXS/+OKZMOFsW7WDTvgcW4q0HGsNA0tBI2RtMjoGfy9ryTicZlB8uH4E2H3LT2te+NZNo
Ia54l4v3VDUC6N61UGRJSxxSckYiaU86ft9pWIUJZhmX8crH5uHD6zrC7R2cl22NKwzomI7n49Bl
Tsl8HnfZLEMGlkxAzQQblAAqqMhC6lKO2gG9TQHNhq9GZ1uQcKqyz7wqzn+40af2luffEyzs5pdg
0sUNQuafyhykIJD4KqG44v88AZsAFgSa0NitbHPHk+vf5XsYLZIvCHk5F2QHKKX+x7XBP9Jfxyew
s76ZrEhdjk0XMmWIWTy+OmiWqRdiHGX13q33i+KclxS8s5f8QHTbPdzfiVedt59MEItoJZhebh+a
v21gaN2yLWkdbe1U1PreUx8KXYgLPPqkiXpvM4NQ5ASU7OZMzC6Gs0fd0Y/mUchrkBSMP7m5ZhvE
lEnQb7vs7n3Kmr/Yg10d4zolucBNaOH57GQfzJOh9LxbVLjjghX5YX6eksv7P+NfpRg43I6fb0Q2
1DbGasb5TjjbFSc4UVM1dPatDDxrOW5lnECmma3/98u5v6911KVNq4lTIA08c1FB0OOAq6yJxZy/
S/jpkJESa5KhyEluvanXkc8XdtIMroxD2GTudUhhs8c6IIhcqMzMbEYJglEl80vpfsMztQCVZYeh
83kCGhu1RN06e50RETyOIXF45Q5YiD+DgLwt3MHgRhUwjze2RBufhgmL3pItYGD3BwEANmdrPIUe
GenyPtXRoBKOCyptQzxpF5qu1AX0JSvIv+8x2Zvq63JRSDoaZzUJNA9wNju9swNX/gKXog7011ra
LBcatfc9Pu8s10a8ns24MFQn+G0qQHAyErzROPrvJt0ZS9Xmrc5ADpc5Xp1XgenZUsXxwtrdMOJ/
0gCkql7ScgqrLsWQvs5tlBwqiD2q4qHHjkEBKnLBdH9Jr9zgORgAkVmKvY3oW4/IMOe1/gut2PS/
zust94rxHFfLnsK8ojHchQWxivPDa7Fn3exGp07lOmhrPxhVUwOOsn7/eQ7a/vSFdGHBu6c8rkmP
diGTz3CMQlh9QOQi5DdPoYHhc7OPsyaPPDZ0V6BDQdjOyKU6OgaMPEQ0Px8jR32rjKZf5TbWwv8F
pUuaQio+1+DHAUO2uKGaq5MNWT+Ec7EP351KFG1ovHrdLij9rp1323X8eVv5XhCeeIWKjM1VYBk8
F1urCENlfHCok9t0P5mCpUSkVlYt++C9cKmA6zmroR9U7XCqzEXHyhqsP9KXh6bZ8fzYOX2TpHtf
pcdjhmtClb2HB7s0bxtMBCyFWKK16vrJZSyIvXo1JyS868QY25t2jR/mYRCwCm/ZaDy1HnXqygZJ
SYAJRf/JcoF34yqGzKWTtkn4VtmGTEla+6Ub53H80O4lPsPOlK5RYzS/b+MWxnYmVrzMMfGUdeN6
XNp0Gp4fC09fOzZSneEwyh8NKaWeIuEvXhO2z5F6Z14Co4AjJtQVPmYMBvxFkOYejUH//n7JpU9H
8fbowrs8hUQkzzrcTjQrhMs1aZSaGDIxumIvGy0xtiufEBdDMpBmV89kIfWB94X2dav2nz6c8IY6
3aY/BbXT64AI+7p2oBG95vYoAYSYb80+jokjMMvDnILrXKwHsZla+S6VZH6WDCM3prUu5uvhNYXe
7aZ0wqfk55BzP3Iza+yS+fobLmmlKlGdAJF8IQ5POKpSawfG27GJSBoipKI5stcLeNF4Ct7TczTT
IyUdRZVtB1fw4+rfFPJTVmPWb3KCxw0it3oRtTgVcCiqm/xrc9vQaEKEqSx+/DmqeUxpVzPY9eUj
+Y8Id4oBEN8au/ma21q0nPsAJlTwRU4n+YzaTCbtsxa2o1756AqaWbnn3qGBnP8SsRJ+4fl39AmT
fA8+LLGfKMJe5HD9rZttCUzjyRo4uQPzYS8e74uHGY1tYyzM9xiqWpi4XccoJQ6Gt5680tOQ5jvX
cgIX3QCZ3zVW/izyEak3hojmGFnBjf6XfSkT/iq1y3UrOOAp2yKb7x2Wu8gDyvyA7OqP6ixV4MQK
C1kjQ8WxSLcvuKcidsQJ46GVDgLMTnIKLZ5/vJ6ev0L1zCBdGm0GThHP+S6RjyGgIP3gAhvJjysR
F9IRkhO4jE1exd265dA4HcIRA6wR/Db3UOAd15hX7vu4qprxCLY84WXWAo9TE9hKOn1kvC6XCFRh
/w8Y7H9Jv5jsyZo2RR2izC6UdEN3Qx1FnwVE4OXedL08sHPA4k0DAHoyB7DN0gdVKlT8qxhs2VZn
fPPrPaWzT+6qQd9AzTExV3ndyxMIEcvYt/qrlOZ+p37EJK+nTYeAcjUXB/eYnnNy/bg3WYo6hmts
Xt0a7FMdpn7/lhvzfiv9APkPSk6N/huGZWRUGOjXZB/UYmONo/y8MlvDeLQSsKU1yj/hJBPnffpc
uRHiEDGqP1txnk/zkL2bkOjd+anfGTxL+lyEjKlSHlVYjjANEZI9cwcS6nSN/cz68g0Wm7yQnMRG
IomsfuUIIn8wQIp6txl8+6FvBDdTYsKbRyfttbOq+nZ2toceYtGRkNGDqQZCu7AB2sPwv3yqqsJQ
WNrx6uVsMll31ATn356cO/cVrI2Q7gMyXWdQTSTVvedXqCqs+RaY2Er509RtbR/wJWzeO4ARRQ+v
PouBhhB0OdShwXQMovWrIGOB97DexCQWig0EdTL+4Fm71WoGUZehnCmfP7H+PW8eD+UjRb284Lvu
dnT1E1dr+yGO4Ms6Ahw+VguweF631lBSrqWDkZ+jdMD9GE8gSbrFWhwzN/kclF50MQNbkg0DAqMq
KN92BtjTZDXn02J/JZ2cnsSfIfLwuNgD7l3F4vPfjgt/ul0cpoZAn7hpY8cpde98UZJsP+mwm/xy
Dw2o+J+PQz7qB7GorZ1x4NiRPIBc7/Ls6Kq7D5KawsKGDP+7bbie2LaDgAmV6LlPYGG5aSuIWMml
KtDEcVar/f8g/nQxg+IgdbnJ8V0FdKixw5G+NLlCHsZrMPK8+uJSI5JY6oDDRFEfipCsbqq20qXy
aD9zVFh3BZ+itK26bQHKB4jKDaUKlqBbbrTBObqCqPfTn/ZwoQarNfpY/WNEk+AzRL+xH8+nmZCR
ZMi0k53XazhVNXrVWyaQhMaK66IohrM08laIBEGdZ302FEjL9dBp/lj1IcjxViG1maZX+1fxQwbS
z/IR2LX/8tP7jgdcMmiH0xzMff/xjEgfA8GZf56i5Xwoz02qJssJRPZEjOFUHK5ruCmHrsMA//rQ
HCxUaKGSTjkJUm1a2VPWEE+5SrSieq65wcRR6c+q3DZPrMjScIeaJUXjCpc38AKs0Pj7u50CFeJZ
RC8CEDy9hueEYkKn37I720VQd4qL59b0OPFZPXJCpQAzit/NpXyojMsQMMHWah/pzx3cvOY0x1FW
aJKuhzU2/a4PyiP1HDNxW8gNO7nLomPouARAkrgYLc65L48url3964l2b0WmiUXouRuOET8ca5Ou
WkgMXeTSQaAENdj3OLSO3arhOpZh5x3/MiissysPQJ3uzTpB136TFphXs1cob8Bx8oNXngVwRIuJ
Or7TIfLvkw+P4HmyigrGhYxiWjUg1ZBhQPFqjIwm4eUVIEzcj/O0LbeM/yMyUIgfPbqkxqnrT67V
DWMK2KCZUL2JwH9hnW2cxtiHPm+iNi1nErhBMyfJNtq0PxGVd7XZYk47L2WlChYiixg9XXpFOA2J
VogmHEMJQh0dq1fAqu7sW+4W7+bjNyqApSw0Wc2qqjUvCEQhupHHZw3yFJVI6LSStBZSS1QKoP18
B958HDe9b00N0qbRM2zWsxLoy4D9LV5XuB+vyIdi06XL2p8JmUY7WeSNSYoFJoND1MsTqomfofdb
7idH0JPMsbQqu6maN91HhbYspqo3yS60QoHjRtSVdnrE4JchLzRP2LeugKVzNDtoUk2xI4jzIabD
afWhvp0L0KVKs2vXp4TxLeOZ6iitfURiezZ99jzNYqXRK3MNO5MwX/Ii+vz7d+3F4Ud6SNMQ+FEV
LdtN46s4ZrU2I1ovyoZxqwIhhnBtt0jorlclbek0KbxS+T75NwQ4gbeK9oh/VxX2pGfbKKwnFz+1
hPnJEi5uoOr4FLCNRcf87CnCWCcR8n1rlzjgbmJ3Qk9DsFM6ClkKAAsWB/OKTSrEQa6691mGn1NS
yc8ugDNYeMyTEPs/dX18dliOCpHkSlZBNQUChecstqj60YYTw1FWHMv3TArLw11N/TNcMMWS882W
HRPCNAsAsLrxgpC5+7B1PbsrIbJ9B+6P8C6Ogl9PG1TY/bvYTEM/P5z2+eS5FcAqIYlcawWNgHPM
HjhtqWAtIXp8VdXQFeKC1GI+BgRUe1+UzE+dgKnbNQwNxG3g831xRa57aT7bK/Xtcx95asIRoSdJ
kfjdjiBfOIhP1fwnYEnCnDlZXI2ZieG/VLq2a0DVHFoZJx91NnXXgucN6OOnGqAUxsCbssxsl5UP
gKxgtgZqiuRlyEM9cpseupQldtLcC1IFxqDsW/LwrVQHd1SDjvE3/IouJ1UzIr4N2IbAd59hVEdl
NsTX7Yjq5+XqZNUy6BmrijzAHmKTpp69prdhx3owuvgP5PDa7w/c93huIHe1tD32Tz/AzY92MQuO
L7W4Wbjisxg5kp8UhZA5+HU13S1pkOp9VlAQnI/gKUmtfTcvGY2ZonAsxAbIazyIvIg4bqINJPYA
qJg5D8RAnX5de1vFz4lFecGhfr3HGFjjaNp5snwTl/wFxT2sy2A33A4AOhZJBN3OPXTph9kT36Sr
j6PLewUw/glWQAHJf44jqV8g3ytsE7/nPpchHZqvYyGmO/SO69cqSvuInn1HLT60BliMKVBCIaSD
ZPQ6qF/LuzWyD41/pAVp4gx7YgapjdQT21QnqUTXDdcUZ43ax8HTAkYvpDwBSgpYziRcdOcDqyjb
GB9G29XyMCqi+R3GlvaH+6selUz15XgM81YYbPRxjYFV9OMx586N7yabW4f3tdonJz/vEYC1BmpH
WFp+4shXhSPNToTce+AzG5+NaMg0itkJNzCFOosRcTv1S20Gx6d76AAUvmwMXr/U8qaMnkRlucmQ
6HsSDo9ZqQneY6V7RduZ+Koj9CbT088FSknEhtXHSp+Hc+oiL5bANVP4I88dDkDozmXru8MzFFnk
bZr08rAo5BRWi5VjBJzTcTShqWN8j4JC7XP8X0xpm1AVmQaY9O7qJqrQzvMOMzF1ncUVtndH4mc4
rt+ERQ7xnegYqewMWV2uRrNUEkkMavCxdy7or1VsheQNK4a0ix6iThBwy25ibEp5mqu23qER9Mm0
s60ItZHZBICA43xsBqu8fGUqjB3pcaOO7XU/rOAjXVErI4KNDTR1ZMwTSKM+qHW+6KgYVk8Hs61W
e2rv5EYpV0+DR2KXGVWgL5M3dFBSoVvj2RUKtacfBNiZJZ3nm2kPNSVpzK6fCoxGZuOoik/fVMT1
UkA1vhOv6hZOQlf4Ejb/lRovUapJak7gN6cgA/AR3n/EhBOrenZsx7TRQC9hNmjQU5d5KzFAjMm9
oR+vC9IdP63VoyD3JUxRez+vqYm9UGJAFLxpgpk5sw1rOWuigcoie/mn/QbIP3JF0rbsHZkgS6eM
IYqYL1KdRZBe4skKtH5L5UmGSOu6lejhnT8lPdTmGzTj76VmTmXNMzPPLTC6JJKRx4E4SmZmsspU
/r7KAWua7FJXE5wGaoUtAy6DMB3s5GM1uo5n9f1VLeJEt7/jgjbqS8Apdqu6TXuLQGLLACX3aTy3
Xo70Qwb0PS08aVIDQ+qFwnAKWVfATm125vcyRsS/8vFLPAhnH7dqRwCSM2JuvLvTcSuhWQUo0BX2
gSGSwOtNxTSpFXYgrGx7RXKR7DgnL/GcaK4oaBqPJhuOQRQSJw6wxQdColsM9PSX6gbALzzKtHuk
jelenolBcWJFZRbeZh8XqgSPx75RsQQUW2UlbpDgybrOYHCk8G8VtazNw4AhgeRMidbKfcaEUJrN
rfJjTqbdl9xh81aFGr/FaQk2Ff3edTYNkeT+JARv1/XvO9Viu318snQsaPXeeDWxz2F5GRRNR80D
CDfHYqg/FeSvV9TtLjOBucDR52+F6uL6v5fJElbbKaPqtjxJp6QJilbw/e2HWaLh5Gl1m3f7xgni
AKuRLXz5Dai3pqMN2l0MqOpQkY9k7qpVDXgXlZbIcdS1T7v9QgwAiJw7NaVXjKZAJJErmZL9tqJs
kF5lzojkw8xa7LolksPVof8YbtWeyI0AtV6hbLgT86LdxxV5ayKtGsIp8CJluwZ/ZEAo4iLpe9MA
8tk+VIS2vsFn4NIDAC3jKu6tb1Xs3XhnYE4+YXWIQpdidslYsBv6lzDo4mbikZdOxrbeP3dtRQk/
Ft2AdhSovmdym31xs7IGxxsynlu4AtqlHdlD38E/By7sehvPIoBL1nEoBKMiBC8V8ZBdBGPO+u7i
9TEnm8nsX8FcKK5lXuNsOdHV4O0Rr+pkUPV32MwDGMY3LiR/EihnIza908ziUzV6P/sb3GykO+sg
HxD4sv8DmTp7WhfaeeZ1rjwtwQnNE0f5XXs89ASFplfi21MIM6maN4hYsFRo79JnSF5+XzRAJUGr
5byQLLtaipKzA1xTQ64eSMI9WV5S3Bp2BUVJ0+H5FaD3gyr4O2GKdH8N5RgEzzZ8qzIlW+7l+rVA
wMHkfGbIQOJrJxZRaEZuruL2PW5h6pB2gYiqr5bwOfyV7kcSmPSXijErCP5doJW/685JsTHg/YBD
2SsYEZCfBtpF1eYuRq1pcmSbbEigAdc2qMoLu+DJO7UmmAfca+q7aHf9VYtoB8Ls4cMSy79c/BZB
bvg4qhvKQ3voaJV9rnJuKA47beYD1S758KbCThV2foCfXyWZvy6NLAwV3qV/f4ypnFfNJ1lZ+3Mj
ujlRWSTInxO5CSN6ER8OxjijGJPqG4wONpo2ePECc2rncdrVQdIE1RpI84vyeqFRvgpc48goiju4
r+840NhaL6XAL0jchyLS6weir7s7MKEQsDqwQ+QdAxmsUme9ebQ06/zQuqvPT9i8fIArqAbx4DdU
6HMO180TPKv2m3psE+8rS/oYdZ1Uqlc3Shkr4J2soZQOQtJU3//DGFw3icnRrXOyNUXi9hxGlWt1
1iIdlj8Nk8KxcGX0A5f9oVsDLRdqLueJ7TK73BK6d27K2a95OIcAz/mHFbwkCv+k8bTmEKQvAruu
oQn5ZMLoE1slu1N6KQFg0c5edZViHrcR3guqaSE53rxnsZzkmCTAMtq0Sf1kxEEqxBoMMng+M77j
eBCLDLNBmTmlD90yvf0OVseNnvhQ/1c0Tg4RSrqFBqm/RgcG1ejEr5uOKDOnL2BaeSNwD2Meq02p
9EO2prq1YWLaURf0Q9GT+w0xinzc/xF0t0v+4L/NWJ3W/0zLyHun7MNIw8KMwdK4ocKjp2vIlsvr
i98nAAGDPiaAVyTS4FUor82iCCVCJcMVx3gK3mn2KSxGUk9+NDj2OrWsb5Bw8ksbC5jCUkYSGaOr
bXYxAX/GCz3YjMhR/hCIxC6tHtgh8AdMHFnIWkZZk9AQJ0xo7bqYEuqv74w1m4uwrQ30HJCZ+OwE
fdDQ+wF/heTc49sg/9ZZ9SI2MX0IzKmYGoLHm0wPtCJ++15FHqHifRW1VL+cBr+OdtgZg4nGEjg5
JbAmc4fXwL0jheSCzEzVA95OPl7tgJlWStCJwMC6H9J4dmmtBEHW4dh/LA94IEzhosZOZa5lqNyY
yX5DIG6zBJUbyF3wfOcTYPlHv0GlYI/cefFqZw1kTPvH9s8dWq8mlivGVrNKhYstEZcRp++IUg6w
sf4mxqLKU6paIvMzWCjJPmbITflucHzLj7ZWzq08d6clKagdXRQ7AAbaHFehyFa8XlHUC4smFFY3
1BQPjGVhhohXgbEi/I+tsKKFbYLRuzrR3yqiM7cQ1RymrKIzotPgYmg6vPT1bwt6z69aT/9gu8qF
ikxQb7uHObQTMCQyVKMqzLWkEjBkIpYI4Ad6VU7kEnBLv61169KnnpvPHaOkxlIBArf5NRMHZWVN
rEcErtYBjCDSeQ6ZlKviOBQ5B7Td5ig2J/8GcTopZFy2kbfP1+lh08KdaL3fVfNO9x6v+QLbVhp9
AHIBDeLkG4iWYmgX8qQY3MlNwG0Ce6tCTUdtPuTOKMQPyUd2J0IsKQC20c2O7jgO4zvrmognkyqD
pqn+JMhS/1pSLIwAuQ6IVYWg7i63FmGB5NxlUvxz3i1Iu/6DdF/C2mcR4mAkyDdUr3mcbZLjbvX/
5vxgd5DUqMcZ0oZ/Yms/+3z+98gm4cnjSLrIBfzixdGLir2BEa07ssq+6pvKYMxchdFyZk75ReZS
Kq1FVz0j5SotJGKjzvFjpdNhP2qmcgDXYkbnm/aMSHKSv1v+u5qYmCpt7SAxPUUxtYRlAdSJPhIV
Ilmgzhi6xF4sGxUV+xOsjeXSgwvZCN//k++FSVtHJS9et1jBPSghcGzb0M+WxXUzcxefPi+jqJW/
p2htmrVXCZYEjnQGWDXvTPorjTCggURKDcTx4miMdCzfUWiXq4sDyAPnEGBhUE0JPq6+KJLN1Qwq
m9ZQqEfMH5tbfybwBcXgr89uVImCl3mihSjBoaLoTYV+SOSXn42ERulqJ48yJ8hiUXZ1qCOeaswC
d5QON5KRYqMZbg3XnH9HJwOext0H+qr7oIAZLfYpjbGqmocqmcyNaep+0df5/JSoWss8cPWxYaw1
OCD4XcEs/hupRQYFSBs0yrbC5N4NOKSrA1uPDV0hS4ROcFwsc/zb5M86jh/FGjerRIhwk29AtyMl
K8uWgtRQ0CafGXWNouPVtaiZ7qipjt0Q8MiIuBo9jXgps50Ql2E+7dZ3qsy5LD2eIWAorQK7M0Z6
ypnN74r7aFmBx1Ot+8gMGYysqADklaYYF1aAAxYF8PZLQfmBVw2LLCbs8u1ahsXEvY8yzyaoWNxB
aNafGtPNrAcCu6Smd4u/k5Hk/k7WUuQnFEy7H4lXUvj1OzMeMW9b8JLWV43F/TZLmzdEzbQRZ9+B
uebS4fpPEQ3XzJwDMYGGKpDwqPVuMLLl+WlFW5MBRAUWqQmSF1lTFoxL/RiGt6WKNlC/wg7UydAo
8ip4oBRCs5QTFrpogOi6j+uGS5lKZaPpAYojBpAMWr9boPGqtMxEw3ICvnvHGBBBfOtqxWdoMR8/
qrlgCmZTVQd1FKv2jAl2s8AaC7MpOnaMnMcQ8xv2tLo5J1psS6VyK1Mj0EVqQFrRyrnp5gUBETC1
s1SldRsmOzDW7xfRu+T35XiKMhyeCCWszye4UkH9FTjeRK9lla5yc9LmbdelQ5lPl/fdNhBnnCZM
3iin2+tbXX4Z+RyXmNv7RgUXFdqyEtQUFl5UcFRQS+udvI4Hk4U5vYw5rNSQTYYD/d/zFTNsRu/e
KFcXAwLKl8nqSgvDHWdsAM2m3z2tP1fzzy9b8iJJ3bx1nW1jOpPD1QFOFA9t9SseAuVWUaPeYbSH
7XWXhLqwmECDkyn+q3ZBpPEG2HuVAyqIFjZ2B2MDj8vDfXct2CbToYDV062+Nq27lfsrLJH+MVat
JG0c98J+vXGzYNprwydn5h5lZP7Ph3cif73tFBQAekW+IykwEvOn2i3fYtpeFWDZQRrQIfeXgVnm
ZiS9TGwnwAaaIu4gAa5Bj3F4XKpjoSe8UdWy9mb8l5iLlEfXKI35Uzn/l2deiWoxLgedLiEaflzk
/Ufd3bFd1LgZBlNJT9zfFrhCe9zBj0oLnTG82rDsPugD3udadHIQhxaMPyMq3u1GscjaXLj3VjvC
aw7ejwOp8n+WBaGX56iDdTZaWGDR35CXHUpeBv6sdbsOoc1GhefGfnAFAUuNRAG0+BEg44yoCvdd
Is5Y9OfaqfLBWewzgMI9pj1NQDJFd67+X/LjBYmoT7bwiIplTHoLdUMnprxG2hiCJBHFRjOaygxL
/605ODWR0dj1QGGkHLWeVtmqsNoky8yWTg+lKI6nTm4iHnxAFsjxpTkK24+OrvcQq3lPN22iy+RK
YcAtdt1g5z+hmB9X22MrDMGkuafSWfWWbCknZUp26SvP3XyC2VxsJOuZyFs/bGsSDRyoBwFruzgN
3WTuS4vSY9yA8uTsYZcM1RNnqG4xBRUetbg0kmC/HsNYM5i5Rc5m4+4o4Ur1blwSwL3aAuGuwx6l
M2DUTVXOye79gjPIjQmOVRyWuTK0ozCIY4d4jhGEkS3Ma4w1ymBFzoBJvlT0Wuwd/jk1+fhSCLPI
y3mwzxqyE9ZA7yQV/CxCXFKtLND/MhJLzFp/3A7xGJzOZaZHWkCSV5KrnaAhL5nFTWwCDASRY2gS
41BJa+z+20DNcmS6Kzu/f345qbkkPERtcqwlpUBbrxJ13lm6opq42TmO1dSFtyILgHFRmT5ROc75
80vYzvHyuwDS0dsN8/LeIBmZC6SNVCF+s56EHONxA+O+Fl/sk93E1ekP7Vm+qIfVRc9uMcTBR/sK
Zep/cWa9SWwYPHFMv7xC3bWNyziidcDgQVDDgX+hxrpRV0ED+xui+vCNJYWvSmalCquG8gE9DtsO
kTYxMw0ediM+RqcPUJY3IH8xQclcjmzJAeEfMd41k6nbZc6jy1QpNPihg5V5Jq0dqJDhI13Jv33H
jVsszBocTGRgTwervf+HcDdFUjCEoWNwUOAtrUfevCg/Gh5BZqDHCBiWlHoDeFgXxB7WSBpbZjTW
l6lVYjdiPwetL4eg5MMQ3goXM3t+JysqvzDmaKtxS9lQRSzSNPzQzIA3fAo9LuDPhXi0MrLyx7+L
JCBXqMCGkr/nn7HrOTfuhQty7mTZWCGQW5l8fJ06UwbOmw4kfUui4UgfOQZDVWmUWIlM2gEAe+AV
MBgAAH4lCcO717ewchmbF6/m2NcXIsgGs3BQXC6OEy1yKX2hnNgvunV3TP+YbD6/jk1J4C+Cv7r/
RHW/74BUDY4nNzbcEzlKG9v6X2xbEoXN3gaV+iCvF6uH+AvML4mbro9fgeD3UTfhoBM9hXhD7mkS
DZRGLlaXE/+l0rLH0FeXNQTaYhaZlE/6Adp6hjvfOuxFq0R6d2KTLTfmu3opHymFOqY/DcPdAOda
PFCxwZqvl2apVWyIWgwRDalHQigE5oNFefPkcbEBe13ALSqxNrdhSP8Q6cZbv3YPEfwMLtnz4dmg
DtMw4y11uaDesdB0cq5nzNWrmQN2aYqIj6WS8NO1y4SHlAx4U+gg+umwTEZNNbBFAVUTa+xSUAbG
Ba6hgV8xBodZguHqavnc1uVpyNviFncpBQz9/ml2gJ0Yw9KYOB1KULQlvDdI8APoH+boKGPcEVsR
RU71vOkpGVDQppt28Izh6fVpAdrn7msKQg9NUqpajM1qRzvSay7QJIeNTlmvMEaY9FREbCa8/XTq
Ix+AI3azyJH9Tcjhzc9oXQr4ZBF/HOzrmEwzf7K6ISoUAdFR+3FcMDLF8QMc0jViBnfo8uEXGbuC
NqHi6VMLFrkCutZliYGwCGTte3LQLotSZPnXaig0e1qHmDSXdd72b6NU8BFiWnafDT4/JWUhR5h1
hDYUpWFowpOPfhYTMSgN4d5uhJrCRFuAmyC3hQLCy9QgOcdXO4yBcOQkMpwgBpuXJm6WUkoT24Hg
Yp+0YdU7a2WplF7cFzEsexooQrydQ19ej/F4EZ9Lhsn5mcKaYlCXwgnWfZsmq9+0M+u1H0PDZTTh
XvWZ88mIFQIWaEYh71PUtqoDuh5uwflmGF0vOQZTW93535p7HZfQdS6O6lI6C88odIXZstDg3nPY
9zQtKo4papSCcAKgQP57YShWB53oIWlWyzGpOBfyIbfKhtDfEP/wVRNGO1MefT3Tus10BvSDiRJF
EAaeD98WReyumkqJur4e/kjhV7up37HhDZ7hkllpZPYIS9+RIhaj/PRVKi1fZHRdlAeueO3ANg7i
UEEQ19PLeW0hLuHRKrulnNj0bCMBwkVwCUZN3g2RJ+sxyTQIgUaQnlV40enJ19WZzSXqb75PgrR9
eUCbBrX/KHQ1xD0grGP6ofRCYRf+yXMLrxSHmn4XDumVyKvjO+UROcD4TCbI/+nS+ef3b/CS4UGv
Img5bl14SyJiwCbt7QhIgbKm9g8XnBDMAEHOCMx0TR4JnyWOjSKuVC/ylKAs06BEi0qdz3rhbpvD
l4r1ajC/MQtcFSgK9SnxV7RK+T5i9yk87Tqy2bGymNWvxT5rwm3Nrwazi0+kIu1SKsI9naXoAD28
Y4QM2dnDvvLSfd08PK8v913Kbrq1B9NE8A3wQr/RfG9qHY+YITq408RGaq4vMZtdTty+pirRvXBd
OTEiaHf8ufgRqBLqde4jz2rBT1rFKx76msXAi58H1yTc/jebBksfBVk5TneDXyXRYWt1Uv7DCN20
Bu2R0Ff5Ogvmg4tipPhe8yW8W0WxaWVecFOWlm4i7aWieCc2kFzkk9dCrhbSL8DTJJ9ZeErgtSyJ
HHlcBdXlH5wahjsE7fMGvAywu8YhYPgTIehqSC9VtTqHWRAMjl8Jh0r5IcOLKs4swuQubtLJKT1M
ZNIt8ebpDXX4zm1QhyS8+xVr6etUXUAL57PvU7RmsL6GbEyjYEtL2DZBPDBO5fOdTTzc5/ndXYmP
gMgrTJA+5J27zhqXYwHxvo7aZRlO+tHDuOkvAGnnoCno70dHvtxZF03yNbHtO+VPCAE0RWF3pkcm
Vqgn42N/pmvRMFfXiCK2C8OXk1Molp+4nYPZ/UxHz25t8SAkbNR+jMFjc4JRGfD7w8P9vvAWKkXq
eir5GHvv49qBHZil9DNwFOL0o2pT/SC2qiIcdNuInMr3AyJa30b2/hjWTozQcm/rQ5QK+4ZZpVYC
T5xeUq7IZnAm1oaK+wA6EJuVokICdZe1dpOdYs7ofxI8yPwnuq8mqfLTTotF6CAjgWz1H3ZDmkUl
PCNQWt4zcesQbqn5JT/+5AvJ8CNasHvDQ3IWmZY3tmQPHnogn+DEsAmkodEaAXzJc5Z5+92u6+kL
nmjjJWE4VOepSewtbxegwzAVKpeytLJrTOB2sZRqVly8P6d9hlSfZ5BAMzbi34ssPWc1FCktw/6q
Uco2L2MtIBmn6Yqxet0gWGeD5EE5OtyYFvqhXR7dPAVhe3Pg0HEjHnindG6/kE46DWrB/fL2kMwD
mFysc2LX3/jFtNSp9p75/cl4Jn3PCNFWFYI+3Gw9ynJTPn31adlBEvZi+opqhsm526SoUpjILhg7
bkCBP+0itwVF4h5JghM5fN0JV3CK6ccWJvdIpauxtVIcjXwF0tf9IU82I6mMFQkxVCKAr5HTBFrj
mpBkHOHJZ2hCh+EcIgfgWfjTfHvEKZtXmRJ6Fr0frK2HCggBHQLLxkc+0ZzFeLxEW5KK4QzT7C+Z
8W7GsDp18JYLp+MH/0KBFMzHEZDLseWEQOqFmVawShR68ZehTykLleoVwIBiL34Ouy119+PTXGqt
opTWhHCjq/tl1aVJ3nKoV1YDOEOSvMX4UOECEH/3IGvJW+oo77D2gGp2van9PNU4fNd/TcpGrCqY
wQb4xEIQ0p9BQlU21is82fmQF3+fZN0PLQfelQrFkytfz8YD6c2kBV2uPItbMLMsIRP8eQbpLVhA
E6WeNIb3ZM5C9eMZgBbe+zbY31NKr//zejsPhdobxX9TRjMhJsBiJEF4qIT79sl4rHFZcqFLgErl
GclA5O0qqIxUFchY+bkkhkagJIo/bPhLTPWZoV/CmrMhVlMdQY+Hc7ci9Eogw5FTNmnVSrjNIyhX
BlpnteGVkXA4CCTmtlXA6yKnTRAv6VP9d3XRNuOS994TI1PRowa+dn6yRrRdADsRD9h7cRbsvWkD
chD1/ur58wD9hl/DMRHaSGL1D2QuxMnAEaJp4bSSJPw9yFfFHtQMGdUTjeHDKR3zbLD6aHb2k79d
h8P0Z0rYkluvWwFbEERsV0h01chzVTWdO4IiylpEeULEvm6CTxOAFuxj5hrOwEM9P3Hp9zoR53gu
FMnzAsZU7BF+qRaLmqHkLaUVnGKPE5I0bJJhmWzMHBNhUOz3l25A6FEN8pcL1/v/yGVDzRYuLKAT
MH4M3ejTTaa5O2INf+xmUJZG/U1Dy+E0tccQwi5Ntqiij9Ry0KDMA8gqWgtKVJb0VjDoLUYtvqe+
i6848LaQGBjrz5nj3eFJSu2NWOaI6XvREYZp1amujPi6ONcMM/MRFfQ5YEdKUzTtJ+X4ejpPPBW7
Xri21vnXnQ7CKZaCpUH+GtUglEbEshLyQxgKDEvR8IyfrOmtVCiZt2NFHfmMHGyjwN65AU4WeXNX
T06dgccz9Frj6jPLhFiFdtAgX2bwKrUu1loPIJPi3Aik2H0GBUTNwieri3CkT+GTbSJtw8803Eu4
sZgwJuFJUoJJnG9M+Td1m8lWg2MBebNC8g8x5isVACRSJkWSTrdG2SJjO1mgJdoepkRe6t0QWhhL
0DkmTGqXKR7iUHMUO5TWWNQNmajHv4wsMExWhnZ+397ftEJn4md4mgZKYmKK735hpGTpE2eMlX7P
2n/U2/H1zR6zwqSFOGityIsB05O/GucsoCyL3szaHh8qFxeCzhs61DIQtRCIK73hIIERGUfAy9I/
IzLRNqNn3Bv3mhWK0aAG9uvdWVDmdk7HK2gWHCrG351kUVelU5E2tslnF0EN33UYHH/ifj+A336z
A0bIp2p72zcUiqM2hOCJvwYv3PTSfBGeL3VJwtzwGYPEO17iVu+PYbWGLoIloZjzjD6CcqdKShyO
ZdgWHbPjgpFoZTfOLLLEogtbaVHvd/H77BnJhyjROT55t2L5Rg6x1vplf8tYkl/Tn5FPYjsqms5Z
RUYCyD6WEussQPdCrvyRLPh0B411AWxTO6+B89z8ymS68DW6UTgSttOWzOc5+L2YOs/mNt0B8QcU
R5v8xkuMzAfFFhb+ReKxUZX5gijpMPeewHnpz1NK9ZUpU5i8i/Gm+momkWxYKO872oTno2GZdm8u
8aJMUF9rHgpZkb2JaWq/1oME9MTEwyM/MxZXnuXiUkGLlbGICWlyxWpQdfoTSq086UrZLcjNg8X8
xXhRD4DaU5T5CvIpDt4SO2Isf4UHVCod0clTdBYaxUi1pfUnA8wLusAlAdzrPaHFdP2zFKOz3mTV
IPx5xY2EX95PfU4NrSSLW11yN7tViAs68ck3/6B90wTf/98rbzFrY3M3d44ysqtkc90I+fY3LIuC
3mi1P3nVFCAomSqaQtoPeU7M/RV2a7bwpZZdmtinUIEHz9EtF4iJ5LMYdu6SVOmQ9KQC/05T7AqK
1eiq7GKaceDL52KUyz/FlGyuWmEsbT0em6DBhh0vkU8tjaXyejtI4gH3/rxa6V9pJzsPnGr1XsEc
crBVUf8FSwTISmkNwBo1ieZJX3ilXC/IUS8KkzMuftSe9+4pA64+6jv4YcuFxsmdMuKfBqR7wW2s
eCTyoSmj+K9X7LEAMxiG1ro7RejwYuEP/JxQRcDGaypuMmdQZX/+qfWHy3tYRvgzVbEyhF9YIMmJ
MbtmnwIhAtMlMcyj04jFCD7ixv8NNmHbeE624+BMcyKmX3uM60epXCJvt6gRv/1ennNaT9wTwjgT
OaCIKPEYG4xW+EqSn3ZHL7ZxJv8i9tqn8P3i74P6F9F+7WqgCg4bvvLr2FAFQ2+zPVSB3cCYwgbv
XPKM/qQrDRLeUbS6KzWG05dLoFy3JEWWmk1MNJVS8eAQJwnZb7r169u3Irqbc8K+34Ci/91Qq9Z5
K33qtJpbgLbLYO18Rilhr9XuXfLniZwHZGNXMUL5FbIG5mnsb1qrwxFY8/SqZr1BOwZDGSiazxTz
EMQqYDuWIn3AypD+OFXIERZE3bxlP5zkrAfhbx5pwthHvdCICU8Ku+5mRNSARyotahyduDFqwwio
grvDpbPSIfzF8zO63JMTvVHGykRgQYxdB5aI2+nROz8ZAM+s3p9tSYRFuvEiwRk6zeJhLViDj760
B7CbU2qrJ5Z6aUEA5aUftBDGt/NPRr0YeMW+II4jMqZjfgb5B0yCVb21yYZ1miLnG6U6j+8hfZTs
f3bVMrjksPan109jkMxsSrXA1V2Kc6tJVoRl+O5rCnZWQe2AsA2m5xwp5rDlO74cPulrVmqu+HtR
jd5m2DQgnTE7xzOkFm92E0CCAViZ70FmegX7GXQKZrlELCgSntIiSd5VbTJDpnrkZzeWdBp1XdXd
Dy89jINK9V3IiqW+1kfG8VmhBYOez8VRfFXZsWpUfWdZXoBWoaip5ucAXHpZHmp4sb0ZgJcYZtNs
pNG9A5pKY6Jupk/xNZt7BFlPjRnKT7EImCTmJ5WPfMkE15/WW2t3ixkUqbodYchsp2NaPgcYR6cG
Jp7DP9gzA8scEe6hOWxKENQgUldrgDgGKr7/xSS0TvipSNULQljw1qp7BiZLrD99gQHyRiu1Pxhy
d+v0bXJ6oyp2XQLh0TX+GOEjVNmMVISLtIcyLFDcqri/utK304GqrZ97kmM4z1AYdDIJ0H3XfSH/
ix3T1Su53RKZBoGr6QDPuBxbrszRe4qydpG3ezP5a6CpmK287PFmgsK8+s0yAk6I/UUKgJdpBpC8
lYo2/JerNf6k/qMJ4CBlBnJ0dgsv75d5woOOhJ0vonMyrnDToQZF0shyR7WK96QRCJ2Qz79wD81R
2H4xYhzSd7E9rLIMWfCqgeSrsCdoxWcm6Uiw7VyOFOcboaeIwEG9nMWaFTDKdbz6lO1eC+oDcXtd
NvsUyX74dBmQgdle3AHhvUh7XFSfkXLZH3SojPAb3sIlMpu2aWgxD+shrNyG5Kgb9L3q7/CLV4WM
dZh/IYei+txJgW4MuGQnlTv39vBNJTQLH4YOAvnignCWaj4jWo2/y0/niZ2BvimzLM2nml1YBIq8
qkGaKubbmXzGvJLpRRAAwtD+6tih4giNzkCPOPc7aJW2jILrvfIMkmLkIoCYCnej/xNBFmY1MJAL
j3lENj2dTcyBO3a/ZTwNiK4M+lqGU+H14JSnOPqorcCVzmScGIzOmUiMHQq4Y9/otKJuRTIiQwgN
8+KGJPjTCRuYPMLEBeny9k8HdF3YpKtveNUUtxBFynfVNYtPHl1/LzUZnxQ76gnMVL7ODSgzebvA
tcpcztq0ClVxdtQUamtOPeezDcXZp9e8zQTNFZFzsDwZ92Ro5aA2nD8qCjIu9tcl49Hro2zn354n
kZn/MRrtyFqCR4lHxmoTnRr1rr2FDKR0hnn2CYePhNnQdSG4LJ8h/ewC0rvzoCvDyQYq/fLOuDIq
zOe5bb/PSf0ueUAXyp1dS42zgYyaNCBokHGM3CrVLY9sILUGD5QWh5EUfQRz4s6F+0d9+PWS4vfS
uqIY2Q8Vuye5loa/5NLW/Ki2fXpNul3vOQCeE1TrAs80/klV6RAk1sZ/kttLA6FXVN/MB2mVehJ4
CV1Z9FxIcSMBJ73iY/GkLaW2AjVmlRWVWKknUmTaw21zziHD/5PDrrhCLssTN8wcXkRzWg3wKe0r
dG6ApqKJPBJSOe2nG4R/Nt2h2C5OtYyovEs/zOeUADbqQyTMtWS3PJTseR5kGlizL5p8st/vFonX
IaK/1Y+oOIbnAznk+XD3uUQrz+Ml/BH5IWRITbjRhs4GSJDiGBV2JXqDFxlpG4xRVE4RaoTAh9dc
3o+33znxTNqqdqJpkHxfShgRDjTAKeeJ+livWFg6ahiMucv4lTkEJ4ywXPMwFlyITPnxQQ8X514y
s+eqst6EmHgNVetDuFtYr0Y7wFLI7JfdenNYNgxjGvDw2nfRDAk1DnpTETUJW5PDxZ38lalcTAm+
lVm8aXN+EfxhY8Hqzynig1BY5TBVRlpGUjw7pVJ9IMMe+adAgGst1EfbjXWyf0u8QucdiQzv9LN9
pdJQcQIiFKKHQNn6nADsE0thdBELg/AHhrbnBiAmz4EIBeW36D8LAwstiehOp/T5b0rL6Rw1b7BX
prAdFdBAfHk13w0X/uyd0FcKNoDubDLisyG4RJH6N9ZNobH4jCwOEEWhbi48wy8fIG9mwkYJp9AX
sOi6ia6Ooam3m6zckRKMrjaGZ0UZspR4HS+8vzJxcLXIkRKS3Ig34mZlf3RxH/IMdcktw/QIBhRG
LcSs9iyAfbaPp8KjJ+tLb/D+4lk5Z+pj1e3EFnakcIyciw52xh09Iwtkc/ZmdtMIKykprNFCGMsV
oLRuSPQZke0/qhxjd3g48wj0iUwhA49VyHodoGyFUx//OWsn0pmPeXeGlBSC1Krd7ZAXBH0hyAA8
S1nZ2e6CqeJtpkCNRAUCTEzwKcRLF8tnztNJt7KKus0QfT2T4nIGocTkoHv3I6vN6i5tezN11WuC
JzGHUCvQR2hIKH8EZuwRU+mCnY111uF79No5PLTTmsFj2JUDMbesNaFbcaMOTdcTB4GMvg7jRfCM
h+YQsmBO1zmbAC2UGG+3bVbqMrJ+qVdFG+68xqI82sOUljHnkHXdY88EYbAJMlAXvlrd+Xb+29Ay
xKq6xNjTAusIWOoRBc5qpFqWaEpYbYnzfIluseciOcTAdKtL+7vGbWYJj5GTcRPsN5CyiEnsvDJ3
MXpEk6DUTIVM2JY4Yy85E6ameszdPtgZ8IgoHhbtwPEF8eRVWu/B1hcTWjo+RU718OJEVS4Jr8pm
gstmbXaK/b+4OP/o8lJH97DYWKInDv21KtG2AFsSxragc4Sn7gX+31pQjTDWm+N8Ob4zmu4bTrJF
By3LkoMO6fQ7jtkxn00vxET5ENaGiYYbA/j0H6J18G5Y43j6qI4aiIPRALB5CQKnqRlti+4zEh23
Osey9g5aXN+KIFvJ6TvWAbfPLRiDm2moc/url7P3TP3ZMlMnfaU3XbEsMCP0RHHWrPvsqli9eRfz
i0tNgrggj6zqcc8xx/DGQd8m0h4+YLEugK0uW/VooddVzMxuCOJqtLuJs/gp11QBLdMKMJ/hv/Cn
0Ie6i9McSnTqRwyG5NLg3AaIs4Id4IUCfcC4ivixTTEZjpHvRZOB/9lT2kk4D4bDVpvOHi92DSru
9/yBzLSqxaNRryl5WKZCt3v1zgTLfOpNhSEwez+fE6fcmsM49wBSo35Gw/KaWL2x3PAF4kslSLSl
P6kLjOsAtY8dAN6RiY3EVTNgBbsahOFXvfbCS69Zs+84M26Wqi4xr3TOe0yYyuo1pNuQGvTknVN9
Ao2BjOcovUvPfHdQfeKK8UBQtXxTzZANS0SWTG9lHamGeCs9MPmVmtdVNhGQiTM3TYDhTb7BkYIE
7qpKyvQxItt2ATUbKC84uHBsN0+TuBcs530HWzRn4fqwCgEp18no7A7qwfOUx3MkBIdkSVr+6xU/
TUPh4yElppDCFqRkMq/mDTHvmucl5e+YgiOYpm/FEwii3aeeeTkgpc7eKj2rrpiKTDmQvoOWR7i5
jKw4hPV93zustL2L+m/rmq1lB0f87awYaAXnDTs0F3mwbBFkHhZVPFGcGnVaigpEex5WkdWm+nm6
n1U9XCzKVuXIaNtcfZNuUU9ievn7QfScDh1sddD0mqMTR0gJec9bWTHRMNRbqgHQy/03BvL9kwki
eFItvfsNyxoYqXpItWErVLFwdmmiGlelDL64fH7u7SxtNjp50ezrgWcHv0uT39smF4JIda5Pg0Et
qphsqtHuIJIWPgDw4J/ufxuqh++w0MyZFW/Q1EwUCJnt2SPsSP7JdI3yijafsp8IRSMlgxYu8JUt
cFyNUu8775VpC4pcPkgC7owBfL+2lNEoTUUz0vZ2iAh9bmPjAPQ2UKnHPOevcxs4WwH3yZvGlT/c
9Oe+gQ1QXMS6XiDy5hQs6SyBTM4e2cMR8M8EE0vMj6hRdAexo851ViLBQ10WPbv4MW3zkup0yBut
ZgJSoD/XDI85qGQdPf9Jc8QGREY2OwLJ9c2MivTTSueSBx3vQECcB8RRQIz5V+zBZPX5Ofe6IEhM
i+GTQnKkpu170Rl5Ol5UbHq59rv2QQTCiJyEDrO8wBbVuhPFVq5uXhAm6FmIgzL8KegDjhGT4ahW
suzEQH9ybQ0OVyEP2+FMNwP5RDaZ7HNVlL6lgPuXE//1W77um06BKvW/KzQJe4DjO+HzehhEhs6z
T+v6+mSihk3OZo3FGNAYAJFVOX+iznUhOXr+yvD4Ouel7TBINRqDgGduwqD1o3eKZgPoizLSCxmB
Hd0QNe4kTGs9oiqQzDnwRK6yEBE/OZb5cbiNDhy6JHUpZRQEnsBn0706/XjfQOfft8HMyiDYL3cE
878Vs36nglFOUEMEEE0ytGQPZI/Fulfclt39VjrKQ/i6Em22CY4mHejOtDBOqz72tLc6JczX9g+G
/6ACXTJPQiWC+9kA845ZYqoNx1so6ZH4ZgzRqqoqqS/mUoAmG1jG56fhmflv0h0JXSRRuyC67Jfu
Lpn0aIbI6Jv9CzoCTb5btqJ2bhFJJd089lYZN9fXO9/DNvgw+GqkmrKsK3gghriaNWKY4DmOboBE
403p5CL38KfE1X/Xh7TdCdQU6cVazw8+2elw+jfmYs136xPcVcEL7BvLl3/txZ0PKEj5scUPmFrU
nBJ4WzK17HAK3atkokT8dvRVE1nv5nOVUGkyyTCZu1nXjhfeYFFs1xchbBWsKXk0WYnI+vtJZgOs
apJnx2xdfZQ6PDKNpET21jzQlGjLGClPYSwg4HY2oOXSibi/XC/4l3GinpErGn9LKR+TVidQCdNF
LOlu8+x9ULWwC0Y8otoheHYfEodpCgwZL+ZiCi2e1k0+iW4gJZ+DLOFl9mkaTHZ9lH4tPadbVps+
FdI7RbF+nsOwjNH/mcwqyw/ViG0wkePqBZhe43u5f4eQzkkwA/DqOByJjcH+u6eGS+DkthdKXyE3
YXkFMomQHRz8LwKAYx3AbXNOTZ+r9WHvEUarMHy/v+Dmypl/Zogg6tdi9QoYNL2cW8hFokaUr6sa
osvR0eXI43Om9/b7ioOjb0oNc65JHebLIHhE54sRNB10KAtWgLSbpdDGYcOWbozKJECLIbnpC9CG
NCC/mz776+gT+MVAXLcaJEipsgHej8WTB331/SRs1qTp3TEZSVsGatELzcAOanHVQV/3oMVj7qUi
J4Bws8VaoWLQ0GJroI1EnV7iNVqVsfyeHzbSp/4V7W6Z63OJ4jiIRloZXK8s2/kTSgKlQvVAinED
mW/RypaKO9lpHEzhq0ck4KIWLa1NJG67jA233tet9e3BgIW/IBOCy7ZaM3WAkMkW9Bu+RPPx4Zhr
Vr1H9S3pOYIlCZvXRRdlhRYIWc8+ahIM5/hmjvBWzAertm/Ok2+csO0a1/pLI9q3noV1mdOQ24sw
O8x6FgRz7Gwm09+OtI61LJAGMX3QzGoZ2lpyvS3yZolk7H180/kcWrkOJ50j6hTr+g0QU0Q7txCS
DDd7h/rBnBbfeEZhyYRkwJc4MRRAxbd4k2EFUbwcwI4HCe2nJVaFGBoaaq25vdC8dlOpzOnGDDJb
fONcgzQr8JoFBan2Prsy0dTHYiPjxBcuC5mwT1Mdz/Wbi8IX7AHGE+p4PEOTTxHkpEuYKkZiMbuU
SGzn+ctBBd8vIE6EX+Q0y2MQEixtOg/lMMDmWvrIastZiePojSoRmkxiMMlhmTFS3FBkLr4sKfjH
TFg2sYInZdJ/piEKVgVX92S7Z1Pb5ozAfA0ypoCVmoqxbJcSr8uJVNifiebxHtEd3n39e0+9QKrB
R/SIK2MpJ23TAktCHtPTHgXtD+UZ7jm2aEBomd5ux/64GAx4EG3wKR/dwtUIy1xA+LzybvBjXiKC
czSX+UEU9iddOk2/1qBNWfEArW86zyu/LRjEK56KZzXXA6v+NT/bagAQrzTrGFziGJULDKfzz0iQ
FHeKDMQZDzS4NNnu5cht37Np4XNZxH3AbLzyELA+0qRn24y0LWkSRt4D0H/5BVA3WMBlVw0MDm/V
Dm0503JiN8g+og8d1j7lWigVf5FsOeN6Kro6AgtD+/DweHouK0ruLIE8ynU9ud9S3wbROzSIZ7uk
RcE2BN0iZ0dND9Tnf75VxizXmIVjSV0MN7Y5yqLb/sTvHu+5PU58BfpEmoX7r5xz25O4FaWHtw/z
z6H7AcqohOdWwUkvfILwPIRNQw9nu4IJtrS2XxRC9TYfoNSBsdt5ITuTxsZbTfTYrPOCE4Un2H7z
wifUjeZGjBfwsUXfkkQ3tEdCc6EIAIk3uM2jFCfSHLpV1T1EJEWgkIBXasoHShqQn14+MchC5WkP
LaqJnfu8lEl6AYJhBURmxN6XRhskfWueQyxnZQv1pUzuh927I0aWXwjXR4X7FmIIPY+3oTsEFYKH
6EeeBMXrFRCJR22meR1OLHwOvFkw9Vf2eIveXIhTx9RFGbxpENpdCNM8xC0x7mITlYZ2Rj0jhxy4
AKeaMonjpEdJ05ky3RiUwzYo8xGa3nJA/wppuueJkAOdUQxDIJy8j5k1QcFN58DcDM6oR2uWrPCG
PXkoQp51Dk1E8EE4lXyk7qhQeRPNr8DQ3962sPKbMwYmhA7aNlRZZYrQsrq3gMa/IxyazScSuRjB
ND+bz+Esv9dk6GVaCdntk5ecOXTnI24ptdDAC6/svtmUPgh6JscGlHe250Jjj8KohyXv6Ttz36LF
CbktU/x2fOfCDyg6FXymIuuwIrCu4jgqAzjWH0+wJgLUGDi7yqLQU8zadPpc3htruC3LyXX8MfF/
Q3mknmiXZ06WF20eJd0btggSAlITLtYCivo41/lbbPV4L7+ftmI1mWxZPuX1WPgGZQrH/v3el6cY
Y21LNjYaYUGsnCHb/FhAUaVG2/exLUmeKF5sFeIasQPO7TexYu4qWwocxamYFSwsUInSpwx48pN7
Z+Rtke67Cr9xUA/6f+kTDEUKrSIvjLwNMeznTgFwRxL0Q9r5P6juSHUis3Lys2RxF/di0Zkg4Nwa
9gRC7zkHLuwc/zXAzwWn/tnTLzbNzB1IDQPWox/5NR+1IfI5jJ/k4elfFY4svtheqoRD5WhtZZhV
SZ+D8/zbh90+diGAFu2GybE3jbL3LImu+oL9yZfMvGE6nPD9QJSxdY+q4mBPXhdH9FpUgcTDa0nJ
HJ2lOHxXm5HzKdqJNSjYkW3XB6ElF73AWMN0Km2qss789VmzWi37kaccr+EKfUX2Yni+axivT5vP
/2rYPL2pDySfL+m9O0Xg7JWLkZz2XtkcNLXgVQuQ/pFKTK2I0qgulCTAGrGidReWKJ+SuJanvnBt
FrzwrMY5kk6Kgz9bn6WaHaPoaZEu5OZob7VURWzQLn7vMST1whlJxDmT+heuEOjubYPpBjUNRS/w
hz5iOnuxUa8fhWe/rLiMWfqQZOFAMZm/9/oGeOiNGh+PrCXcl7l+/W2t2YTP0u0RlCyPH55SH0BH
Yo6ecyCynzTMOOA1LCwDuDmMkQTOxnSZM4fQxNvf4YVnB1MEE10zHKwefFX0RmExaEYKe8Wf25P4
nKzkojMgbsQenoW9bwZ03OdvkM1NKTxhKtcz5Bo8EHafEFMocr0aGmvaGQRvgEcF4qhdg8EZUesB
XLMIQW6QkLwe+MF7NKOF6b2hiNp1xlVq/UOzk15hdz4BRreqZD8PO4IFnWpGqnTu+mYtdkCVxkxY
d1fZIxCvvtjHxuWNL1S3K3fLaeWSSJRnE25AyfHQ2h4dGeoOU42sBh3Lmim3NEi7Ly7yB5D58fNe
DLw82BXX/bQ8ZHh9KUFGMmQyDDm1/pIw/njw4QYunQrPA3uJGSTRUopwbQ6dIY85JpX/qgtNER6x
joCIk83sg+/brWHmRBSyX8mE7a7A9CPi7WGIWbqHZ22b1gBp0aMC6/LeuszYm15J1xEZkr+rJJ1L
YXe5af30x1iTIZTMK+ZgUJxgxWSa8azDbpSMhUQKiS85AZzaAAo0DJrb/BK70e+4byHDrJeQmV7v
943rXaG0flQ6R1h+hJ8G0pZgcqTQvG2GcBb3VAFJDH+fFL0mE7B7W1b6gMyRK/vp4xh+6q5wQlJi
wK5nUd8ViJHdkeJGMbB/hQFY+1SCXOrTkMyE6O2CPi5ws2xN7ndLAg72sCSCReysklvA6G7BjjB4
u/EgB4W6KyfvP4ncS/Y1seTVeedAIIx17fjdQah9EiVqg1CheE9vPrDf1i0QK8cSze3LLaw8cDnh
2LMi9/sCYAO6qrDzVUIh6/Fvbo2j+musNWVMXJ9dSr2OKQPar1D3lEAK2AVcbCdG46Eu8+8CTDRP
St2fh2n/v0GBGmhuEA42tgAd6I3xpxS5QqG0f7KbLNrxa9CvUVPPoQcb29aMHVY1ltBRF7mzi3ud
o9LUtT7nMPpgZ36fafqLgkgTZfgmZ17exA62P2E6CF5PVEIHXyH238v4tfv1YsUbsO9RL97fcRS3
iq0h9Y4mOf6nr+MNHhU3DXTcpdJpdcWilDbolQEDzR6Bis609mia6yS/hZ3GMynl0NKojMRn19B9
HEJ5qabwMrOw7g+F4O2gyxCpoFbLdRM/e8rXxLk+XXDZnjHMZmjT8E3rYG6G9e/c+z3YQwbIpmXr
cTBRaKWp8pa9FTbdTpPywv171Htbs9n2fw4lqfhdi5uV4OxxrD7EnzVVPcrRXAmyWPHQ3JmvV6Md
oL6qe7Ev8/bg/EjZaY53SBlDR6IjhJb1yifaNJvgZrQvbQfXLYhnxfS0F5GE+yE5zSURSoJ+7aM9
VtLCyylxEYOfQE5bOrzVMpfQx16IRJrpwDJdjjw7P6zRJXtCCwBwd1Z4T/9a4W4m5QjSKfyvwBJ6
/KP8wD0P+X6lw7moTWBoZR09kUC+OTXtkPet1lWhxmeyBXaRJN7nDxawiVa8N1y8cGnAIMdE7//k
FNa3fhbPYHumSDurNtkLieerfKnND2evMCuB+VeP7FbVyNtchRXr00ipZpNPedKMZUpvxJyvBLnu
b9nemtb4ZYlQXlrDQXoxdzjSY4HPAXdgsP+/CPhPiLGTTEgCDzPhC1BvL6/LT03KLFs1luVLrwnl
3j+XoqcTr8UJ/0xQBupLTk0Kztpy6ltsxNdkm9LAYX0fnhIDwH1NhUism5wl4lYBnJKj4iOJhgpk
W2LHw4X/y/ctohbu94q9cWn1DUAYIykZ+Lqz/wFZBfv7OP/0EuI+fImlx0jBB9dLEybucdbSZcat
VJeNJSsr/fO9IE0XgX2ANAC0MhsEcj1IUVMgAQP2TkpPzO+3/ENDJ7nMCUFnAYUvM1ajcIXvcDlq
gCCxImbclEws/IRn+n6DKJKN1Cn7WKyQB3/GQia+515wsPFluERoVZ6hpDVatoMy+613i6GmJd5G
5KVyWS3sg9NiElaD1OC1tmFRHGycZDzjyAB7Yex3DF3yjBWILz1wTrLGfimtQathd05tiCzyIlIH
jWL8tXtcM2pJw4TqueT39LIoqSdKITfySjpIRZmDYunOJlxPvF4hU7pjQMfJTMgHgkjPP458eYL+
vb5XexP3BSlsmuBJyOqV5MlCaIq9FjMZ1Fx6xw9E86wMCx/o/NsOkvMcfBz0RxXxMofHNhvAMh5e
ceHuF2k8Fl3rsFJcUT5f9ZCutz+Oc0D4q2FVoUL9DcqJY7SKP4P8LPoLCPnhwaBnhAklYidMwMRC
vkTJsrqGMewNxYtlG7YYcg+V7Dm8camhGAeP58sFKadQGyXDF4uU62KVdIypYAUvitBXmQC4Zh8d
TuhCOIymCtdJenqd11/6H5WblJcLuVr+h2FMAHLeB4erpStCo2cK+jI3rhH301Xyk88J5aY59JXB
XNbSnPRg/jBHww7g8VKIdi+vcaYIeV8JV2oEFfXz3V3oFRqL9JFCNriaaNVohqBNydIt0T3LwVRi
rwV1S2fijF6cGhIc9YR3xGURaa5fJyYeZdNLTEiQM18vtZRCUzZnHlNr6K3vWcYrTtLRauQ6Bg/R
rpZvtjFLBIDZAms1u9GPtyS0sqxn7v8DcGAmsWyYNK3Zs8NRotYymss7OCZdRZURmJr0C8tYFXwT
gIhJOuvhGeByuHqfdMO5k8B3x++F1EEAJLYMyYruI0ynlQHN2Nu0UXktmfG4vuUP15Hal7skOKAw
wKjWWUyTydV1zATvu/2i1KeA64jiEFWOR73ZwfLgH2LsF2slRIQaB4OnYa/OTBpMsAkCUY2v/iph
2HDRGbYzxYKqQnNXXI01qkesPOkM8T0Iyqz3blBvMP4ZlUDhQw9R/DUApJGb2Fx1W5aWEQGKHzz7
IIACSE0bP7ujkY08j2SapeZFksiKEBEme3rB3TzN0h3BK4QgyLsomG/7v+yqf8MEuAyqqfx00DVW
ClZDuQqh8zc89nlkjPHMwP1rSvMeFKKbAZMwSUQTkA60bEhp26ZS+d5gkE84zMewB9PHusMElFJM
psjtRws2AuGaRDoYetQPhfDzqLVzvF+5mHu8gs0+xUjBZJruRXv0ypFHFRHyFcOvpdahPxzCv9yP
+5l360kmECdug7HljPK+2fSGKojNfiwQK0MsVCPy2CBzRcpJ9aMCPcisFTF7EnpX+c7z55r8krte
pVTEXOaEtiVan2RUk1e2ZPthh866urfjSw+fMcQ/4kiJWTnSUtJisoQTZPA2Jva5a/MtLxp+pWA8
21VBNRd4506ShYMJ9BrNkVRZZQoh6KH+jQAaWfqINQTuiymUwVPvj8NcLXYIV0RMFO6BxbghXwmX
zUCDd+8fiWt3R3zcdmXCqOSEGBxPLVTiAnD1dZPYVNe6vA32C2H8fdT4goUuQQ/vFNv4QHW5JaPb
gGb5TiLAyJa8++2J7QQZTf/b3KMR8uxsGWn3qh8TL48e3L2Oni+jMt4TNnhAf8DuGfN30PaoFiFX
kjFIRmYBtdzj1X82CCLYH4OnqIXsFzlaMv58+MbWbSg6NW0s4eX+qNOsk+E0NvKHlzmY8estOok3
xfDBHWQJyAr4ovSNxL0LPRQKaHmlERn/JjVszF7XxbAKaHVoK1qMOIUSU7LyV4EcbKTZzaY2zlsg
NMe4FEL4wIkHdxLuO3RY73g7Xsm6KMOhlLDNy9AI73T8pbdtnBirAJTmr5yFhBBtK4pVemSM6Ndk
WlIal5hFGWlaajlgiJWuD4qvwCRNV119dpAagT7tjGD2WytvMVKYvwBQigWodKINxblNM07AS4rR
vLIFprNL3Ec3WEbjPZbSt+kVguCYYi3DegNrCcY3xn3wUPNfvus/tt5SPU2J8EPRGxqYx93HY4jT
aD2IMaOCru0sBQQXT9OR63mIk1bDor/pp3L3yF8ivyYVqEGc0H2K6rtpmALHfURqssCsJRxWQVLo
bqDsmmjGW6Ra+Xq4x2EMbdRNcdAHA8x2wqUKLkpCQBJgL8Eo9i1Y5Jm3dvytLgI2g5gNRifzke1h
3om6+T7vyCIUO7jARCqc3vu5XijUtRqhp5FBJPtWfzBYobxKGxV9lrqLqymysr8jdu12pV1DZ2Tf
/5sgNH5TlV7ZLTURYZ/iOUJjZq5bYrUrvwfCNxHGJ6UZu/Tkd9jjCrnjFZwHOcxXQaMF3g4/bJk7
uWN2mhN7gSDq0OtnTeMbea13vEbwv5FwJv9yLkJL2OPOI9FB1e4/2ioO6xOu8VpXvmKq6aTBRvOT
z9STzasYO/LAB6A9q2fXaqVMsSYGQ84cEAc+u6s2Umw3kxrLr1Cs56Z9xfNW9Ja9HMRmAWrDko82
OTkHmhVU0MjlVbbAcAYXAn2QPusfrhW2dWUAa+9Gs8jNH31KmE7peQqruT7RThtKkX3thESDLY5K
G63/Ye/2nDbJ59slfKvU6pntZlmXvGm6PTfUGNHcUST9DAA3IUR+Vig7AfFpNXIJD7wJL5jg45Cn
093t0oRHw/LfDDfL3jnunarAdfdnMzpnwstrbq3jzjEcRWaclHZBDVHmHWU57aWVjUf6OWBKUIhX
rXkyvG2PfxudtyvTJGuLIdijsV7wUOQprx0P8fwOWFNaHteaOmXCIxlR4NIg1QVRG0ZnjEFeGJuc
slJ2WipujWrfUz5g+cDrbmdJz10q+3sl0o2wFR4V+y8iXdfYijW5KKarG+SMLZWhCQg5yRcc3933
iVz8+ugKJjS1fJDoYUuGRA2rl+5f8cDmDWlmuwLYw9qvHhbawM/17h/XUfakRaCG2Zb+bg7fkLFG
oiSQZ/LfrCPgWVlPEfyhBFMohhSOk909NxM0+oRjtVC9XQExa9afbUaaM6xYTF5EvIKxujiU6bO6
s87e1Kah0vf6kiw14OSQ0F6lcR22sUR9QD0r/3J3ty/tYfId/xO7TapaTIm1wLsdg0MWFYL8o/Qn
LApR6OqYGbYA+oP43Otp5iuRcc0khkRo9zavTbwrflpxTZZu5av+tIC9dWCg+LhSgt3N6fAC2S0d
tOUgKTBL0Ao6qobSPKnR6LjTLFALVr3A+tivE9rqpoiXMbvFNYMyHg0qn4FqfOosqK0Ydslrcm/T
oHkgQqUeOJssfb3tyixIdEIWERwfSpz4lcz+IlkgPew1+FlosXY/jo/WmrFluF/dgxY3KMJnspEC
kuf4X/7gmPzlYWYW9tXAA+PPOL0uWBckCQc03uU4ddEQxMndVHCcZjEyEd/LTMH061z6YoPNOm4B
vwgQUEj9vsu1m3xSYkAMA/lYxApDcKdb1NTkV9RR2JS2AuOJCNHd3800Gtdg3TetiLRP4GR8Kq4d
9PM8pkPF58T4fncgSzgFHuqQaJ0qHTxhWVdZLQ+TO0PVYCG9H1Q+PL0JeFMFPEWsOrdgQi10iUw0
OvU7BrKe/Y74+hdSpMcMF92IVrLWET6ODfFGYiKh0WD0u9/Ns9l2/0hB4MJibtqirJuyk+olP8CD
Ae0JlZ4+LPiBckxXQVN4A+J5/JBYbVuK+vvEteMkI5/drzpe9OfdurooNWMucgrwiVJdw7w0XjMG
kOWsGaBJppzWfvWc3RAda+dO4jIkFHR4p9HSGkdMW8vu7yymb+23exiAqPqteTnkgre+9gknGFpp
XCzcrFpvG4RKCQHNL2xuDohyxHXlMMPKgGoimSnqEeVJlXPmWd1sjK5iZUQWkv6QbmwX5hoHTeum
VWTf67dqcCbZFXkZ+Xk3X10iMDKdLoub0Nx3MxA2jEzBxuMCeMkPvDVRqS6kRe+wh8+7DBOCFpz0
wEG7T0jCgu9XPmsM5FxE6TIHv5JSfcA/UQu18Gnbh2bvwZ+t6riLeoKez3O488xZIzOt7ZVQO2v3
3RlSjwTioexRYxJAuHuTLpeYlv3Mg4mu+K1Xwgyusrl18RDXLZB7H8271BfB8AzkaQ4QHHcR9/40
SdinQUd8FayGxd300OzZJyIz0sNo0//m8Elarb/4PtUhN2gt9ztxDj/EP1EYA3wha38XAfNPSPuD
Xj9RE1QW3J2t5efZ6JX543FST9npRAJ+saeS8eql1njzGzw+6Ah8bhWkBxXCUthHZnEC2GtP6SSb
P4MRHMkfTUwZahO8n4tZ2bgjKYv7DR0kRQz/9fVAfHohKAkBCLd8b7ElWdmaKs/3cAZ3dfplEmwd
lnbL8hAhrjyGJ9PCyK1cDXZdYJ2mJjLC9lNvMtmgoCAih7bU40P1uDrk3nI0D/U4sXfxMzNxo0D+
5hKbXwPwKyaBfAlv/JGy8l9wWpQe3jusUxxTKt4P5poRYsNhmJy6ss8c8k7hulogZH40sSdbOoHH
vwdQjDAdwZwriTeqtdW6/1AYeT9ztMd/j4Phj8ozAfu4zbzl8iWOLdX7eiUytH2mf6zTNEcRay7j
KeagtPoMxE6+Wa4uPP+4BoN8RjLiatl1HLZN9wYM9vud+fG1rYRQQpuQO+DfJ+NLVgfsMdzQHF3i
GxyMeaGwXWQoFP/4enojdpPEd/d389CKq1W0LfN6NH8kgqFq0CckbDLUII5cMzFnK6KD1o8yQBI3
MPx0zTtd/ISdTXODAI9v4ltBD09FPhhblv2uL8gNk2H4NSsJKPaW746GHNBi3bwqkfP6Ce4f5EYN
g/q9DyI/SXqjXmv4C+vCEXhTLwqpVqPOg1hAXnMiXsOAdX6s/zdcWUTwI5ThVV8X39DkblkqyYvx
OH/Lcxp2i3IxjdGSZlWvweAwWNO4KbjKpiwa+RWGVn5axkvXKrVs7DGtbf2H+sk7ylPFJH1doau4
dkKIG6NH23ywePBclAGNjRktqm2vFQMCRIyVxeTUOGbC3Let0LHRirfEIEUnO8i04Myf/JAYjhvM
oTb3THMWDuLU7sbhLTEGSqA9ArXjIMOiX5ik3Mk6OsPOdI9uGLfeuo0tXHU5Hjp4IME7YwRDJxD9
TB9Pl+j0DeGKQr6Hw1V++eUzp/6a6Nu0FSvLxMlQQktKMEA9p6SMEqHsALLGCBq6Dk7RvM89hmcv
zYVfFOq4GqYvH6/LPzKplh1ArllTo46MLuPDsfryt3pur2368uBeeCdl06yqCVY7M7xedAo3rOqD
+MzHmJ6F4jPwoqauVYPXKxlisdAXomQWbgNtOalDq/HzSTSACP/nZ9Qnad/u3s8+NdesvqjbE1js
WE11ETvG8cUpHg5AmHSpGPJ1iAZEE2RCrn/nEes9v4BEVAqyLO4Mb0BNz8YZNwzgnCgVjdeh6DGH
FRJuqx6BzMAGmkOOgoD82XSXgUAnFsTLdcssSsHjC3WqcH7xf8i3UOLwlScu+xWpjlF43T3XURaW
6rcUHApJyzCCon2wT1Nujpq3jEONLECkKwr4QvDk0AwKl/8Pc30kze6obp2bCCGdeCy/IB6E4VS/
0M++2xgNZLKDPqdZbwF3jOrb+cxVcvgJ7Zpaek5eCcBAA87M3kt6nEjVWCXIz6c65cWkHoGUfQOY
y97yl4iDbI+fWJ79JAicdeM9GHblnuDOfSGucQSp+10SIFgEka2HAliEcLM4ulqkTQf+gqxHkLpM
ex7Vs0t0poiPTdslMm0d8TLurcneMXghfSFE+c+jE0bjwY94Qd1KQB4sPXC2SWTpEEy/EhyKLupr
Lf0gaqCNV276GHr9uhhj4b/oMdqDpbDO41Bq+u5F0cAqQvUOAMPsK1dd+jGvj06K8MhmOk60CAdO
jV0bEs5dLLVZFr3hQkxr6bTbUZhUSRJaAeYDx0aGC2XMDiCqp1KwXjpxTw31hcChZn/2UFTgh9ab
g7NU5tRD/migRaQA9UTQaN9b2jUhr8uIitlb/9HwWyb+QQ/ZKjW+8k0dyXmO/6S+oNcRxHgT8XBW
KLcC9rU84ruNlTM5eluMW/GMicmS3gdfReHIUHk0mO7PA778h7fkgWvoQM3oqkwEpumYg5lHODEj
6yb/i60auas4g8M2duaJFp3Kmf3XPV9ICgdJKjkro9XhBJIZDYqRuK4hHjTBVMVNvlZl5JNfKx2d
+pTpji5DIBAi5iZyUjn4pVALHINOtVyIKs8HDI/cKxp1X6nFdF8COydSDgOAv7+R4Uzff3NZ5YiN
VFhetG2xGO6CgGzciP/PVLncgYF5MR8q552gisOlkl/mK06duI2H0xwY/gOCiYxiGpYPk2MyTNVA
vqgS1Xjx3NoKK+g4/SXc6rOeruBnsC4BV/RYJLP2mUJBs6WmoV7npdcKq1xZX67b7MqD/0J2KJ5T
H+e+dUXDrZTpSx/GKyZceOH9L2rUMA/CI8OtoRyCx0yUO8q7xKazjXx71lf0CZBpEk9lfjStvsv1
795GSedbq2Yabkr7y4Ot0EanJuDSGXg7idZIURWXF+mc97OoS10rc+QyrLUEKNdbDqWH7JRBjKZF
eEZlwenh7fKwY/CVzvwM/LjWFFBJLxr9hLFH0OlbNnEnGabRMrKx9UF01QJ91vekX5/rPe8wUd33
LGK4EPcITvrUwBvqeR1uYKwkrvygkFpicoyVkbtJbSXntUOYXjJKT9SBZOk+X4NxQnMYup5voREJ
aFJ9otZ1fLpGNUcvJ5nZP/skCcEzLpO/z8lY3ls2BE6xfHOVRRdUbaEjMYdpCesBtY88EdUyV4oM
DrCyCOqNTGZRlzHZIFDutKdjqENjiOpT2bPjSDkShdJNrL/I0KJW9p4Hmx6OJwjrpC05SGuPQpaL
Wt2j/GdYM4gdHkQ9sanuvMMX0p3MRWAdJUw/VeJ4R9z2XDh0RGjfbEr3wSc/1sXvWlpkCArCa5jP
FrOYeGkV8x6sRVLN1bLdIYDk0QA+REeVy99sR2SW8V+ATnXzTKqxLq9Ai2Ctfly6x/SqzyZZoyIT
rTc6w7o52Fs4kLxWncx4UXWYj3AB7kABN0qj4m/IUliWZ6rG/R4zopAgWmwYAtj77UJH+DTRfbPx
P/mb5wWFeGrKqhOjNcvZFs4NDueOsbgMrq4D5fgnZ9fVeIoHhTmWawg6mJiuribs/HJ6/dAoOJeu
PAX35aG0TEZVPM7S23ug5C0oQV4O0gnqJsq398IYGvcHOkqOOrKgtcc+Shu0CeHS0mlVaaa3q7UM
E44IAhrjhXPcFn7Z6Oo21KLliiGB+SA/gbfSeChzN3gNv27dmZLMFQbUKbkVCJLnn2TRhXU9ZVz9
VzPgjrR6L7ITX2u6IJbLwyakFiZIDN12d65ydmZO0WaY55ZVSbeICdP2eKRnhHkK7F4ML5J0r05r
dkmCwifwBMxSG7m8EzQuayw7Nz4JyTu5V9f37j3JgvUQ6PWTlO+x4qUaWRg7uqKSPNMAhX6lXory
3rO2RXLK3rzSV0wMsjEbeLmU2uSXiUSIfR/QCa1a7ZUSYRtC3g0BMAiuTFfE1DBPAgTLsnu+cZjC
7+MxqRHb000vfITRvW0uzOZmNcs9dKzffegrNa3gCxr3EMGUyLai5r24Qsg0f+6IVejp2rJT74xv
x2mcYc/3RPXXZWMJsrt0KV4pXGrhpzKEIw3nn1gWv3ksGKkjWNh/UtgO+RtQeAhYt4FW4w/AZ371
ubaEa5Oj9wK5ZH/JpUAjBK488wgzTUnF16b3HxcPaAbxYWvmhTwAKP4vH4tCLvNdYG34wu6DaYJ6
YdmDOCyXGdmW5M5DZC5XoI/MlcVnR/hhgbP35VLgBDh2gjrU8FcmE7Uhs65NB6SRX5kMDK0Q2Dhc
oy2THVwolKLV2nbcwjZjKsIRJ9OyM1Z2caM1UkaVFGX2a7hu/DR/kLS6xTNAFf3uRHgmI7jnj4Fw
S5cTlM/vJv7AIJzJndG076U58YkJod18DsuUrs7Sl7I9HsUY7t2AT84okbveq1rty5tbDgUjC5Wx
hSqSBo6Cs0mqVwGtGdkubNl8FZskVhUTlgYNRhm5sCivmqECuwId9Q5E7RlAyqvkMzxkREsuVOvb
cOUQKQ7x/o7IiEwTIU/chIv79VzvTdxWpT1w3gjQMS97F3aBtpKPD1O6BagsvdcoT3Pb4KePeP3h
e0AMOzhNU8DN6E8EYGS+LF4OX5zgoe3A9k0/y0BnnavHQqmwLDmL5CW7g1Q+Kj6gv+Mk1uBFWhRO
OP4M6vCN5Y6oMhO1uAY6/+d//qVBTgoOrh070MbczTsJfMbVo2lUQJ0ynCgibAOVSvbRr0wwaF2v
LEw+tWArbLKQOzERpYdH07cxyWBf5FQDHaQ9ae9inPO2wsQMFdb8i0HkYJVzyuOSz/IFxtvm/1nO
V8QmdmvgXFZn7fnZQg4S7D+Y9y1DjK1WgXrDCBRh0w+XVgW4ZVjBphILZRFHgXreKnO2AKvicX7l
KcNdjerTenEjvMDzp1AhCryfEKZFItghhFdm0jptg5f94K6nAfQjpX/9UdNbeJBUA1Ney5FfPFhn
Hq0bB5d2cAodrrU91Zv+88o6duFpOmw1VYrfgDigups7aw40WNGv7lsAB8MXTBX4TrBg7YfQaDkB
HCDsCNJGRqfW8u6Nrhzalv9lsNGSCj8EOjXHXx93aSrlEF2OvOx1zTstAtJZ9ENQk4N04mnWpeRv
7UpNIodIxImGcF//2mr+w15ht6JXLfPfc0oyPlG7d3DEij5flCGxuK283PhvQqEbMEHBR38WMI1m
wjK6eWIfMXsp9oz76qhnUPq2Ms2prRVsUSDtc3rkK0Y3rDGSWmw4ld55K2x7UjLS/lAQOKFgWKOv
8dDjI2ghl5nw64vXxQJ1i+qYxFY9dCByORiG3aHWyruWyQKhb7Uo1HtrQMogqXm5ZPS6lMWA4y+p
4eb29UVxgDILMs1IxLRb4TUrA77Ls77F2EO/callrmKbQ86j3ZRine9LlLbrHV0jNGWnQnbsAYnw
Uo6LS8nkTWoNILN0R1K93Y/XPFDKdoEmlKgCngbQzKA5r6zH/Au8FiMa6s/bNllYizLACviebdVE
UmBw1AOBTf+8tE2Q4NV9CMEo4FPJHm0T2jNXtEmwJtGfzTuFSzPWdOdVhJVcxiRQUht4Jo2kpXJq
kFMrKraILqQPyXEpsbT6VjYu/TJXbWHw8rooSlT8SYJrtREVLekVZ4UI+gQFX/VwIRfZOpbgGhVU
w1pTzVC9o0VTaVRmLW4SEMQELex08Q2YQxVj2zKK/4B/TkOTnJrgHBkMJQvaqR1OLCsNTTDLQk+L
IxsaCCTXSy3F49v4gBBeF98sSZijAGPH/bl1mmhOwcG9hU/94QsguPJDFy68w6HGuUuTJ0hCTYrt
PYdjFW79KJnfIgrEUgzBGSyPt4/slT5lH///d9qlFsVfVXyurcXe+MEm6SyjXMlMHwb71ziQK3YC
bckGVrQVVRuGsX4MxnKe2Ovoh7y/DI7gFZkgHq4ZwTiGUr6k07OvfyrKPvFL09Jh+WV8NSIelwSr
YBGDHqKEmo6Vaey1PbGXzu7E4FJWmX9U6xVyvEQdstcOhuyojL+szjrrKfWPQ0fLCkXd+W3Ilrb4
UKrCNv1sqNd9E3lOYgvaP/hnngxWw1OcYUhRwP5M7PXwxi9vrHZONns+0QtS8NTBFgYcYXy4cDJo
09kFxzlOO6z4kzov6ZT/fnxFp15EKAqvozlyZne6ID7BgG65r/raztYlpjCwwfcW+sDIrOUJRZ+u
jOZ9xXtKt3nOLYCBpRlgfm80DlSHrL1f33GpQGvtUX8+5U5p5vqZclbWJ2wc5/WxJHsnv7IlU38W
nFwQbiT+qv4CRVRCy+fYcN+NGaOAc5GBRP1auqwTMIjS+nvZ7ED0cea1vDJBn5q+gkT1Gx7SBMIa
/0GyvfmkE6lCi4FkpIeTmjflhiQstT3cssuRcgq2yjKVnjNUVQO35UPlr/T4yqEC2t55Y1LnglCo
wDzLQd39+l6KVMmM71qCPxPHkdwakZNp4WHvgDjYYTLiq69XeWHJn3jaekvcVIvPie2DKuGMm2H9
cB25HM5EhFp/MjYLHbfHFvk2gVmlLX3XwQzrlCRb2WmddDUDh4XalV2WuLdbViiYLl5WkiBd741P
eJJuO6lECeKuR4HJlvl7+LlhXXl315+oNUHatnOj7/lJHUewKZ2EmYU0leDiYfUTt/OcxNg+haRG
8O/B92/LlvDlYnlpQFWmBFo6bxXRqTCDBZqS0Qj43S6s8KSX3ATRCPE7774/i1pCPwyjOEBuG8q0
JRrc20qb15dWqVttLFXGh3/9ybBCJNeJZXKLaPYBy0ERbudinzrqrZ77K46huqr5ceeM1Ho3O6w0
FRsTOi3j3Rl0xXzRp/kvWM9MC/BwLptEHOVjRgPIUE3L2695tdKv0e2and/SLFWGSdh4wwMtC51v
nJvA2jvncC9DrCRnKm21ut21OXuBzrEGU96kafzAObCIPlLMenR0l3y4vsr1sgF9/+h2RSaBCnnN
FMgSffkYOn7TRlTiet4KpbPXG93Gp/LlwNnOKrZNhEuVPtlncxzSlEhDXGd9COGCwvLBAqtHI16t
+H0KvzFymKipHNrgmxdGrf+oZceeD3QeP7EMVZpZYVjN6pEp2iXZjoeosJlIZhKjdJy8upD5ROD7
7jOBKbodCILLAQ3e8km1wqmPlCLGCrjCfnBH9EmjeH2T3Vepo+meL5AX6VKkehTgC4ajbNJ/4YGT
fSovG5Pb0ws4H2qHlMs+VuYyai4+ScODo1+9LHctKcgScn3I5sszLEjV+mvlOg0dltv9IKRUnndL
aDGM45ILjU/Gi6r7ArIj5wPT+qm9q9jbOl7LhGsKu2gGBF85b+sHiUh7QZpH2YAXUuMztYExqDu7
e3ejJUeD8XY/FsbMZviZFklzf79XrECJ4sNFIhFXQg3DUP1gjxOJQ7auC5232dZXgHMhyMBUeVAo
/pAzTTHYwUHU32L2CfT3u5PxZSW0G9/getUC+/HjLh41GHJqjW4F6hN+4cLHr/hxjzQ1fBhyYQn4
UKIAorUbo3Jvyk+gF4v6qmI9J+o0FGaJD4c9P3QdIgBqIoqb7XhxHunr/35yIkQZ3f91xAxuUhWA
5mwsKE3hxJYt/EZ3UJ2xCafVF1V3iVGBrOgctdtBOjA5ZAwMwNZT/A+rdu0biI+08qacDrV5fPrS
Hs3MuHmqtQ4TUSW7roq7TAvcAeUIHWc38GlFh7SazxbtesDK+G+47Sn8hyVEwATqFHqA3I4Wm8BA
IiKVB+J/Q2+Ot0n4q42GLELijS1UD4+XHoqAiZHu8iJ9jzKOpK798XOY2DwQcfwe2ML0A+7T92S/
8ybIOhAGeW/fn2NE8ZgS5K9Dl4Jbt4MnRZtH4d8mHchVjMj+rXMi1FuvibGZhPnUKcQg9uA28UD5
SJNazzASKbWAZHiGszMqOlOQJ5epdsJ+JqkP8vVtKjFZHp8v4ghtCw8j1QOA7HC9bZUBRgoaR1KX
zjgd1KsYH69Hk0h3wDAJNRbb1ztRza3Db6qNyhzQHFJz1LdnKeK2mWNK3YWHry+fYqguRSyrGo/u
24TLAZrGKRF1fN8+xtdq3T2ZWNnyz/sCsXUmf45b8Ovgo04XuQYLoge0amjZRQAArz8/Wa5tfVDy
JQE9PnJzNitfMnZ4LeKBpjW7rTKGLfy6DpuXWYByLCViMMc6Etn4W8n1VuU/IWlg/eaUTg8zrovM
uyoytQWJMZEAX+OSX1thVkXWiudWzQz3b+eqB6W01HffwBCQHzFCQMm22YMYQG2GWT9T7/is59cM
myi8XQlXGbqxdgi8oBDltXRyQ3uv48SbBJXH6dx7v881wEySPX5t/Ep3UxoD6WqK+Ji5nzhjaDJY
vD1IrEabRrS8pYJANBAC1+4yeVqXE7MvdvvLpKJmo3OZM92890qBcUE2boOIWY9/53sLueBHmGsq
5bYHAEqXGmSznaiygHceC0MnLdY0cbzOj7MGXC+noOzBMTJejG7mZeAg68Ksqf87IeCmHHktusSp
VM6eoYcTR7CDeke3/L11SUk2DM50xC+yA5GztIHOHDDAQcUFf/qUKs+dKons8KOabR0Rbg+vtaYG
pUrFzIX55NoCO3H21oKtJECIVbOUDmVSTcIv1q49iLiSCkasu2mMbrbQJpvxgNVi/i+L4T3mV6V4
vf+p5WVFGZ3FZa/ptYm5tURxBQ/ZxmkgpnuYXaIW46ICwoi3NnfJXzcs0zaJ2YaGHVcI0sSOSDKi
hf/J430mL85EslVl99SWbB1OSugZjjEiCtGS8dkzgIwPqrGq0m+EdlkWuYRm6YeYkHMMmUFE5dLh
B0N6BoiYraKgWbJ0tBvRyn559H3JCEkdAsYdNiN/2xoNUBKYRhrjARxEir2cJYJGfwaOhUom+fKp
OPxgRmUjvdA31RFtJlVmEzhAKSGgBIv2n2hB6M1B3mnfid4noFQpzHhSG951dOq5wMLsAI0QfFJC
w2caZ6Xd0ihP59LIAselw9QcfVH1z4O1W9vGK4GDeIvsSzODtoPe637jLvXFPWd19I2BA+HHzQzb
wF5vN+J39VdfbxtFesGH2M7FMMZZdfqzJ/PFQwJXa6wOgYM+ogazB4LKmfZRRWx/QOPSHdsTRaxe
gw6KIs4SC10WHFf6Rrmdlyy2O84/TvKMcL78+fnYiIuMLiU1Ax9jw3NSDBv4oqYbQTBJ7qy8O5wA
WWjMPVxlg3z5n60uy8PRmkscTISTHRiyX1ShONUkrcTJLeCZKnvp/f9vit2YJgGPoJUnqgN4bIAn
xjdVJGaGymBBVU500wHby5zwREyooUdlxzd5ntPYkkGdKMCT8WnqGL8xuyieTTPZ49Oe19AiZMI/
WUq1jt/L6FD3Sgrk1EZGt/fZlRLbxv0DwoatsZmcKIEOb0BV2wuMtsvlRO4tVKk9smnumTQYVvTh
/3xNqIkYc9RZnt1YXQ6lRNtvQEPLZ9ZuahYUTghRXk3WUvqdbkXy5Qe1g8tIRa1wzUVGDgNfz+G1
K9SmYD+zLjwH8nYVngH2vTvSeSUTTZAHBB/Xsv6AeOVZSEbTK7/8dAZg0Gi9y6VWdDBuahTMLV6I
V3dGbQ8BysAayfzuzQVWSeUlkMrfLg4yk1uBxUI+o7Gn58Io4A0UvVkh6o0Fg5hy+UxHFRndEXh6
Osnpa86eK0DbzZ/DrC5zv6vzhQhT/CtXLtmPcjWbi9YRI+uTnDX3pfL7v9fYZJ/tKpwIMfR5PogC
1lIYWVFK/6gvbhzVIy+6+JKFtli5wZnLvgu7RG9AQEHfbDP1vSHDjOtlknCcf10IXcdTY4ujFDYK
eQp/BJy8wzSqZREqT+Sqdf7uTeAV3saRFi2Qwfy0DTOwoPdexnwfhWvHBB8nzkurbkGLukyZF2E1
vFTwl1KPbc6QCoTkdLRVEdPkzDQAqGuumz3EnhUwmxggwugwoHFLTzPdMCWnAS9DkpkiDMNXyMQz
FgYWnpIvnAujzA5NT1v3M6B8Z/AJRqEd+i9JSAyu5o8sMK0mA42zMxjNyQnQvRAsWg7P5Jyhikp3
ADVycl3k08mOsDXWX40mlluzF0SxAQH02O0rf3gr17ojlcqRlKpr+0xKcD62KuyrVqEvjQro08nV
PQ6DDwjyymXMecBpKx0DH4KXO8ob4JnSNymBSXD4OI+dRsCG4DlcaspC59j50kHidwioieHUiCz3
Dp25MBI6c/IJMdf4DQQTekR88OXej50ff78md2wHRp6yaMSRT+5ILPVblbBoyu2vNvbxuNAtnR6t
5SojIJVSL6OrftwENk5YmzYS3sVTOXGgJ9xxcz1Zx87ebs9xe0Q5G39B2iiJr7Do3+f2utWooOYk
GYeYcWNYvytRV4RP2u+McsYVZXz8sgPbbKxftBXAw1+JvM9ByG3e2olyouHBhtTIJqKPm1r4PX7O
G+H4tNqrS/36BJOYrgYWbcdGBrcil+y9g3DKpm8MifSYfenEL7V0x2zOCckriwLaTS+XovI9/vPy
XTl+rCGVcYnowvo9tpN2XZ0lubyHZo8LQ8xlztUawbYXLhnFeBgbxDrqUQ3t5iAncGvJ9mhp25Rh
ZprdC7JGMirWDlbw3lJJnqJqxzRFaNQOmnh1X7VTWcYBnIWv+CfTzA4D1da/tzoGT9sjeyRcVai/
vopXfHPny+e2eTM8zpc97WkOdo9KlN9vpG1bdoYcdVPGCf28weE+/K6cCmOT7V+RSWA2h+APXILh
rY+UZqT69X+K/ByQJCAUWHuSGp4jvb0fO48Cy91rKTa3V+nKCb4azirZPcPzUb5dCKekEaQTlecy
LO1m0BC/fQ33wIQ5RHyqar22Y+qESYxGfvRzX5Mhi8durPGZSPF/V6NrCR4SZrhHSW3XLpwJo1Xt
Zb/H2UIBqfovMb48qcuScLVifnkU3XR9z8qvLqIGKXIubD8DauupPCvzvnDkSURWHxkU3Jds5zEy
Q0ZwBmSkubdIqacd64Uk+7dDussWT9mjjsa2RMwxSep1Pz0gb/vintyPGYHY8CdUzE/s8aN3Hifl
O2Cne15/HCSofC7z3pIYxqKN3cOw5LMFoqCKgvC0m+95PUkmqY8HmBHUxDzW8ovTxOhm87YVDfwc
67K9a9OmT+0yhl6yignlOgfWDFrpdFST7dnQK+vllYSdlJ33v4B7e8iAb+pTioI/Qkpfcj0kI2kr
I20Jaqa50EHloAfwDGlwiZyCgjCVwwhes0O5GxcOPw2EadkfZhKP8A5Hz6p34fOrsQMv0UtgbWE3
t6Sj+U1OqIFKBQ3x2bkavSOXcOHOYZ3fUk4lIQ3xv7+zBZImuIE3pOnbo2ETsKoCfzsnmQ0VETv4
t9FOJ7tjxgq7fgWoG+Vak5CUpFldDaGDAyOzfeCYDA5eX/gA/EaFtQcY7oxkVLqVeX6BM8vpLEZg
XFLHMHgAgZPD+vQRpxRV9+OxJf2zPweAx1MhlF3MXvxprD5hHb21tDfEH5JmCQsmZGso7VIwMPwW
r4ckkZgx70kVhosElqsVH/T5jxgygZjKk57FlakwycAbTczD1XxTMvw26zSEcmVMsM9q10ft9buZ
Hlmauf1oACUifhlMhOibdwTArfjbjBS5DL+BQlIsQziORVG88srKbPjEdNMoHycjikZAa3FJ9PaG
QaLHBj04g86LcZnTjeGXqdcDsR3gepXrogskTK8aFZZ5YJbmIKSM4lALbZ7MtrZD8W33avCRlEug
W7G5CfHtutQd4SzxJdybe4OLtwPhf+nXoCKLvehInkwg4LyFjJpwtumR3SzkxdNoOa+5Fw8LpZ9r
Q7DNztoOJ9zwUy3E6Whmlt+KVt7Q80uP7FxvOkf7N6yQanSTZ4tNSZPThqAqldoNnc9nKy8Rz3Du
gSeGJmi+emvGUIaeBXhKm5XqmQtoSOrUrx54rX56rUHlWgu0ETMrO4PRl/mdwqWbnKZkDweUrLWj
rmN0//nt3LvXudG1uqlGoYrpwO0licdxNR7UG9Fh2ZpJpUHLXTdQt6FvssHFv+Y172wYvSB2ljxz
eHVUvLjbaJpKObZbH3W+BTxLBdiqR27vnAYhTPD/rlpCWbCZE6RolQtlGu7gWGs848N5Ldv3ERPl
w34Nl0iSoM47ajCdjQQO76O0v4zQJokUYNyuaKdc572sVZ9mFVRcLa7GtZlA41+KXd0AWjEg9W/G
H2SO5FirSx4hUIQse/700TdbVVZHXyzIZuRcRznCUxm4TRjwlSAZni9Dso5ToZlfYnjdUInaxU+i
BxikrkuMaCnitph3nrc0P/gkInm//c72qrrwrxabAHHVBBS0zP3punSAHmpIYPk/1CQANhY1u2Sr
1Pmd70PnFAL+KVLaRF0XW0OaV0Ou3x7SAeN7OHgz+qHEVraG2DlfWZQmiKFRYA828GtT7gxpk1JO
m0mmxHSgXdKO14uAlLPUvjUBR1hLCFyNpfzEUbKNj726IQg3Ii4S8Mf85DNZe8Xc6W0VS0gNS4xQ
KVeKdSgdVzyVAQ1qwTXTdcznPhMRwJJM+uoNaGPsu+VAZ6prWeyDYl2VxGxu7oetiT3GvLN4gY8Q
YIrSYTbdHRz9+myLqbRuf3bsjEN5IcFcGxULx4jOK/EtRENDE/TDRdJ0heCyOxLN+g59v+MjelAQ
mbscOk7Mn9jgVhjVTL0MNbmPxK7xdADARwKIm1zx5cecvckuyDw1NBzFkT0DsKSaulf4nmyCvL32
PUL2z89hlFIGybi74ItlAcb1ruGKOFmowYp6+WSSBYjyC1sRbNMs3qrAgBwJtky3zclkcuuP2jhz
fn6AlFTi2pgeUIyaLsEskYV04bJ87NEeO3HaylgqMo6ZgD4VmFmgtHcUlRLao5YtK6dxpWPhMCst
lf88asDPzUXcGbx+xFVnStw5aVBwd6zJXD0N4v5GFTz74P52SaWL1y1WRpnG6kGOqCOw02qeB2nr
Z+kjj4WbMfcfAO4YWu7iVUGf3zofCD/9Fyd6zkYyjrponF2Rbj56bWgZ0Um7S0K4HP94xvmLl+P/
6ur/7wFBLKrYiOC2jK3Lx32kvs3DGVyoSNTmB7LIf6N3cqtv//DTOlkZfKSfa2+afjwI9duBXpod
o/YSf/8hgpngzGpNIrXQxhRgr+LwoC3q2hzqjlx1LXiwEHEHhRb6kT67FmKzbp48ZStd65Ootv42
S29H8ySHjpMBn7WFnkxAAbv9yZXfOYUEJ+csA0cqSQsj3yj+Q3zXokn3taAUYpoMSVs2gHakFVNC
rgluzmgwLsu+76NXxhmewfSMVHGHSJ6pV2tBP6XH1TRev6Eh6TbfGubZupa2/H3J6/nIDTn8SsA+
6rPXQfEuOSVIpzBVL/wCvPNTudAv7bnO88Nsv0Dbg8hB9SU3GdVpdu+Hn3qqsqeW5XsWJWb6h1CY
crag+aJJzj4beJvn5Z+iU6IUwaBsy9Ai1vkRG+MEQt29+cKbnANpx8Ly/mYQLLyNLBqFj1FXyXYg
4STBu46LYcymO64Cm0yaDbSEXQb5zB5fv4S8aWAMp02DsvQRnXyphF9aSGdOuUrPUmBK7MT4lBYB
Wa3cZ0GoiXzdO3R61JUDH1EJKWZtrpIGpXGb2eeYnaJGIgfJ07wWmIRbhH32b2dJQilYfqt/nDO7
dYaS3Q7xxyPx7TKcSPYM80asH61t8kFu6L933HgZ88yq6ZYjJWgWbEjJShC6UxJ8Y4vSfrZDTkD+
X5TB8Ru6DBi+EXO1Bohmu5wvRI4Z8BOHoMB72UTAOOxvm9PmTyiUgseDOlB+K4s7Si0yU8j+LVMo
BzMisBc41Q7G8a6q11TlWYEtKynow0/IzTz8PuQ4QGtWL6/jxym/WvzDhFeHjgdxXVuYlSjK5bnK
y0Xla/lACwJw0Pl5IO5V7wDf0HkIQzOVY4hpGXESGxiSslE/isvqM3jBVRKbjvs8QT2QpGfrRSd2
gxKjZGZ7qZqB/+RRc4oa7WkagfgArEO/NATDEDkTNdViSjgn21rYygGQz9YhrzkYiHR1MjJDBymQ
YDNcoXIwaieVLAD2o+22PbrCGyf4uZtCEdkesv88dajv60KlY7FYaYB7CyDe8mYUkpz/51Hkg2ni
k0KpNb0RxCLhIJDCK0m56bNNabm7rDGhVtM0jl+gedov/09NdsR39ukDiXKmk+Wn/vJwyhgjbF+6
Z+yX4VRS7hlNTdcqUAPPRIf18YvoJUyMnTjhvQElLmCJltEqzHdN+JEbmec3QvND6HxlBc1h00jD
nr0VV1rH8pQgQNEevuOMS2lOcB2FLA+uuz+iMb3/UUyRHOwbirtLgQ/d6ly8mftBE+lYn3URvhJh
LIZKoGRDkumu60c9YeIUEK8zbtjSfjCGQRDvtNFUTrKTia7rrsPOXRVf69z+HL3pFsa6Uy4Or9X7
yR1jABIVXq/Jz7pCaSu56s8DNEPxiRSiuWIjZMYHIKwLLfrJ6pcMwY5+igckmK/9ff5xHC0C6UnE
mZLMGWad1YDBYn4W89DAcvzqGwOFcknjhugMEQMdEYFv6TSKW2eP5uXujjSmJ/c0c2ocV+SkSsSC
ZQg3pZEq0vhQSFrLfRDwI/kXTPhNTYcV4P+SWKB4f+6nlaMy6Q4OMogn3gClBPCXSMTozxPATlvi
S2J9K2GitcnQTmaZ+E/uiA8IoyvBoi2Uags7O10MY4v//oksBT5I81ItUKt1D97gEYFMZf3ijGsi
TXhrjXhl0lCTNQSZFgo9SV3XTohJp0e8NzS6aqNdesS2txa58UDYHeJ34N7cXIU4nK/x/nQshD7L
qi/YB6O5CjgrxiECTChTzrRPVj/TdxRvM3jzA8yqihIxQyurhb/dvDwDdope4VPstSfMv2Ogdfnw
VQzYooWxR03DZdqR5NNGFIlH424qPJtw+EfItS7BWQFsSHf72vbUpiA48LcC2ROWb8QF4pSerZ1h
fli7L2YQC2yVQwrg+j0Jc5NR2xhjIRFy6E/aYbmWVzIIv7x6MBpzDzHcOM7usZPIPKKkImFfCK3q
wZHRRXx5YI/vYNck7WKIi7GJBkuezka5hhiZM/tBIv3VrZNXEiq+1i+Rioog3K2fByEnUrXDHOYC
314c0IFOCksj2M0xp2/N7GyMBQ39MuWS5mXrEaZCoKqQ6dVqnAjygYClj/Ht7u/RDElkYMZHifuy
26Igq0i0CxJkfPPJ5HJGECLk84mRQh7J19tjD0D2P9ltSos9Xp9uVgw/QVCqDDQwgfRhfmpUDjBR
rHGnuCzrni4fPaefnk8vsZ4IQwkbMC41jclS5CcFfcnUOKA0PLhFTCIRF4vDNNof8D5i6jJ3I4K9
V6gd2Y+DkYhFOwFeAURZxwWA5zVo88rofLs1N9yIOGR8hxy0OVlLSbnRcGZpro9m5B2wuqhpbyHZ
Ad34F48u2kY/z2ykcOhpr7GNgiPncIiFRqG8Rb5sSsZtGi+q2ujVkntydQUZOHxfb7NswllDzEiO
VpvVGnLe5PeRjAwSCn4EeqPHQ7L4b/xDTSUIjggsAFYLwInxMDe3/sFSFP/YAsPCdMf3dfnMpHcB
FDcFiLGf7URPOllIdNC8AAc6PDTRSBXITFPYrICFN5R/aSNVwJxtm/WQazU5C6fn74vRCKtudi4w
eBG29IMj26VBgLzkIFJ8c4TZUnppqR3AtBpziv6uMTdR2C6QqRXrbeoJoMoxHQh195EzBfbbmIzf
PCXLPpgpg96EYPTtLtvfPK551BtRJ925ZDC55KFH7Ow83tUA88DuwGdVcecsPIHcpsY0Aym9J5HX
gIq0kSnOxWnxrZAviMFkXaSmbzNpqGtn5yO6Vul0hK5t6IahIcGIrwL5xbi2eBIOxQ8eCiSp02oa
a68GUrrQIO4Luu8Otv8qp6QSzOtB/eqcYqSPafYIG85JIQl4C4X5fh6NgT/nExR/E9Qo5Sc3LMWt
t6QZdmg9gy0USdnhsoRWg+t8l/3oNNcI1vt0DTboGy0DrM0y4Vzlh2qabxU+nqiwaNuDEWVdggrZ
m56chFZdSyEGrqgjFac6ilT5MXNJinoLKDrcQdlCKlttgaEjn/cmUAS9nz2YIcsqfnEW8Jbo/kUl
3qAHh0F6YdsVY5xaFNNbih8Pyk1Vw1EmnR2cF8EHOqVt9XpiXM2a4BevITa8atuR3z0uFS3NbQij
ZaNpsE9rsjdZGE8DfENsexks6nQ4q1pw4hVcdlK2/DJLBAWzLeSQ9rixOWD44I5S7GITUgSuwEUr
oOE4hlJFxHjB4fseoKMCG6WJMNrH0CRfkP6hNj9HqJS+I8xkEBFJp/GoNywS/GF2NPW85MG4TcPT
9v0uylcQyDuNcQqblioiM/bHFUgO6abGoWVqUv2oaNaeRw9bdlipTvyZqGNeOxOaQRLsMQMpAX28
4qTDcnUxgt12BrplhjQD4u1cdWOaRXqigrGzgkWvlKYnnJo34O3TPAU/7b7vB7DykXBPBxYMIflx
7xoODHWrEoBgIet39/9gcEH3iNUSWun9dbWSWs0KvAh5V1XbRxLwIn5NUyHwQRjRfzO2objVUY39
qX6cB1shf5kdteiEIAKCXgOFa2eYCzYwqbTUY2OPzZCYXM/9L8efOLXb7EremIXXFNd5powBSCkm
QEo1GW5tnUP/uotK7FrOX/1U77n27T1onH3iSyCpGQK2uVqPPEFSXUn7QBmZ+lcb9XyXEJMI/Idm
C5aptQ/xBpGFGFlqtT/VtchGWMgzecGkdCVnDqvQ68e1desgPFq9SsekURHjN6ZHrRYxW+DSngDj
h02pYnxCegtBLeYnaP8Y7NZTYnlJvflI4zBru2nmB21LhoUO0HjEVTm61rx8ffNDfJtvuc3e2Ct+
SKcDtYREHyfUkr3ywV28uUKJRLZCdooaFNI3isTVPjB+0QOBAJ0vc5+wPrVftEll4cLEOanlvuGE
k2N2a3GN/pzQGiBAipSyutrzV/Np8PE4tYY/ONvnka/YvfLj7+y8TG1vvW0PxbaZF6NyWR/2fzX0
kvFGmQhej8EVYSwp3MDxYXzg3QESQu5/LLsXQJk6UWfQy2ACf68tqesSypuFijitZyCdt/Miy8KT
bYUBZ0Mm3OufdYb6NaZfliVbeypZD9fkuRpqutfwwlI+2f5KpWjY2pOoXyRf3ykbSLAZfjpUVrlK
aVBEUka6wyA+GkibPJF/ZQOj7klA9OJM/03u7XJsjwkPHOUvBdpqqr+/HUM1/wxi7OF6qT5DfD/4
ELDRQ/Emr4tzk5UGlLNVTxeGzSZQdokTSDsGSILGADv7LaJeX4YfSdiSmF6Aanu8tiKP0EKVvcip
lz/5pCvXLIzLX6oTogkC5d0s+qfEvmoiB2qaXzfsGS54ENTQc3L7+/rxc9FFHjfHTt7tBlXsMdBe
Bn1lklfxPN6yc93SPy9ywKYlX4KWReYTKPKIjHysyibjOkcLH4IzskuycCbkkM0AmUiWUf5+asoj
xJpBw2zmTEoVV/SsW8WMDpyFzXlFKSU6LKBqVPury2avUmCmrC4s+HCd6Y/Odv1qlIcBRdwuR0ES
7znYvldAme7cv+BH9fVlO2dpwttZVrDOy4gcVoHfbsGqL+lsd+c9/1v0gffTAFIeQ1gYsfOrCibt
g7/koesAyp3D9MY1SrecpoiF0v233TvyjzFZu3JtdPbeSbnzGOSANIK31veUKGynLC0ijBGsdTaB
VzPT18brbolFvJX7fUulb6HGTaYyislivTrLoww4ayKi6woaIISr6s+YRK5PgAz3W+bvngewgJtV
4xNxXj7qaxZ+DpV+ctV4YgaZXwXwkYP/V8xZyPL8YPCsqupCO5KKAK/75ysQIttfjVkAiwWuTSlb
hjD0TDCKk2p1uNac3sNWoQH8euuwOG395SR16QHQ8Dy3dx7L8Z35l67jJmXxd1TAIln5hulZA5sT
ia7g8KZIUbitlquTT+7ySbf4y0ge6BoNmc2WStPUgMgIb+AlQnOzmHp7SA37HjF0JPIkNo7YvImQ
259aMw7rb8VyLwz3ltIA01OMtW+8N9lyfdVMgqR6CLkC/aNCMbnNvp/C1HrCdhEAbpYuQefb6rs1
QPXvGsRSfPYg7cI/Hs2dQSFyhIhvFe2eP9C/cz84SKnXJBbIBOwTDuPG1dUqnkYkE5Hc4aVU8Yaa
tBX+T3jkga6a/bxy0AeLIOcOOvy/vHF9ODIPgrl6YpIIA7gNff6JxmfWy4AUs2uTuLJ/EIerXWQM
yI7XSZMQ794reqzQSyIGIc4XPMguQcqUWjY0JECJotmiP3neAjT09RTEEF+uiQVW2crcCRx1OzLK
8OyvFnUdVRiU8D9dK3YatJ1OIktzaO96ze0Z1AfMtFzl6lFvUj1P3YiU/R0DZHTTH/CxouZTxtzu
ShJYHTokeAL3zq+NpJcGhjKVxa25H4nhrFNGynGMtzmRNwoU+9/wMJBV7wwN2N9E1mSNF9e5cLRe
HrgDtAUYGMCjGiDMTYw/+CpZalKeqfLhMhsbxkvvaMtw9RtmPm2nr4r8uDvqk5k3Ajw+f4SK6swH
k148d2klU9jkBBGoF7az9KZ4tWZn2T0eTOW9UL8CEZ7Ll/XAlLJszSENElowVyunjJlFJepnuKZ8
+s++GyN1Urcy8L8LGVbioDO/frBdMdt5CZjNUrT8JL0MP3W5pDBwYqjwFzeJ7/exO5YAEwxE657u
2LWaYtM5ukide8QGjK/G3obLMOay16HWH564yuUN12w5KDiwbSrx9GaM55awBUXNjHeKKZqcab3s
QkEun/UcEhCvpIcLwGIVuBYLLG7Yl4MtWXqDsjjVQwJGPCJpFxGI+LFwecfUPWNc+4J/RcKRt+Rl
x35Dmq+3+GsK3fLSFBFwb0DZfg7ai3xphkJnYkS41OgdbdQ8KuIeUXZwVPGQFt1cZe++XZmIig+b
4LlGxe8TYLfOOOT9GSHTeWWCjyKNYRa13nIuofNbVAdVh6C5+igcQFRzrljsM+hwIGDMn2GuolGH
BvhS1SqEjjneflddf8u6pl5eDW0hK/1p7KbCuv5eanaa+sWVpe5AaiVRWnvBEwvABZTQBSdS0MPd
uRFAAH7EIG+5WiH2JOZEGY5S1TUoVmtHHYEg5fA+gjJWGEN8cnBzApjK6i32EAYazyuOgEDkz9A8
lbO1Mg7egmBJw9fJ10U5XK39WtIhNRmKkXE6tHxTnOz8VkPynY5XyDy04U81Lmkn6rkf3ybR4b23
7IkLIxhDh19UbN0FihNK2gO61PVQfDeqqdSJQdBAwuW/q/QPv3t4v6Adg0AwC/CZHi6OciUBHLZZ
93CiZJ4FA6tZdlN/fdIJhZfFRcse/TICQ+SpzVUKu4kX8Hih2k0Hh9CQhxeZBB94hCCTvYE+8uig
GMhAA+z0RI9ChXDITVQAJTnPvm9IjOyh00i0KBUhN0zkFkhwnz1oUOX4RLPI0GFfVZDO1s/5Ea1B
1CVE0cKt9lA5Q6XuQ0/8lKALecNjQIlyUPDo4LGwMcbuKX7JyuULRKC4QYgRReLbPUfTz9Dm7YDQ
B3/FQgv4Ftfh1ZrPkTRqHulLoCYsY/waI7S8+i8s4poIMCFDJZbfFU8pm5E3K2n6k4J8eGrPf1ye
+Ima3yw1MPwDTCEB1MScU3zlitxxjaU2K8JcJeIAzYmrdgMg4ZNC6kQVptG4D+0avr3NW5BJa5jR
M39MgrVfanosP0uzmxSMiK3oNV9xSfK8MD+ViSYxRp04v6K1HQFOgfcO5LXfZyvF8G40oH+89BD3
6scTSr14ZhRz0X6n6guU2HG+iNB5MV/O54loHJktKLv9Ch2WyIxHXxJh/8jETAAY6jTVBfAmfc3v
1MzF+fey/syrbu7gOKlfbDgJ77HJ53d4eX2KFd9QePvz0aARQUhtEBYxYh9r1xfporY7d+3/W1cO
PEclmxEvp+9pP8RO0GT9vqHQKGAO0Yp8O0iqNxWAqzFkD0ubTiGL/gFVd7zfzXxfzHwX2ujYDWKN
jIzqi7ASjswsIJsmPOwNNl3R3A0/ATod8lG8dxX5gWZPeE1byJlek+xw2lSIDLU1pAE/TG1QVOi6
lsnWI+xbEfzSl2RIXByltl/M0RwSixRiP88gdbT2qzoovWV3CaQBYyaTbs5RRcynuUlpNCOqtQ09
HKXRk6eWakKxuUmtNfrfbkAbTEa/aINA5sn3VoSm2lMPkkYHmcM/yjS0PF9e2odh90ux1RqndmuX
Px4RXY5X6MJfN/luKWBluJHaymh/5SJbgmSacj6uqcyIWvmT6QzdAQKlbRT4BbMGGlRLWdVmET5K
eIHTCeZF5tVR1fkvd5PGNdVQEX6rlccolVmBSP2TX5sAZxZzzge8kEFxM73b8AFRc53mFwDexAOr
iGjtQ6omnJedRg7WMbyL1LLVpRPLdLO7YxFRb2Q+8uo/PluXg9mwJnXIyTYA////xFzqucDHcbne
WGZKPF7Ocr18urBJjfKG4OPn7BnOWOix7rRJ/9Lj5vC0lYRyo1LSw0HpgTOaBBFV8LN1aYcXQds1
q0HQe3c84KdPncxcq3GzIkRLFt6duSevxtbdDFIfg19yceBg4ps8r3GuuiW7F3ObsKDNBwb95Y94
hJnMBzkZ4vFLcUVNIgKXBnRDfHejQpxTbw19mZfSpLvkWFpNL5mRfUKwYYT2bRnbtiZLtTnBZ1uQ
n9nE2DTaeekkqr8moJQehhcda1IiPrRiXzX9x6nMWTAlsR2bbhdVizJY3C8lS9WFUhrns6Y60UkK
W7k9CphWokRO71gDvzxrXTluNfFDKA0RbpxaIpcZWdXly3bWhjCiXU2OAbwXa+PI8OBTIfdvqQhV
3Kcv0sVTuGc6FyezcYZnz+M1FS0yZ5MEaKWhS4Trurt9SaFEsXO2xwDZad5IrL7qZG5f8qH86c9d
9cL4CrooO/o/PJEDc4TkBEJ6gBOc8Otj9vSptlOXsJSGAA1SMjwe5biH+7DeVDKcArxO5KiDxla9
swc8KvmEiXjYQ4qNA0G0fwQJDiDUqtYvZi4NPupWXObKW+UNVXORXt0v+OkOZvEambqkIomj81L2
r30EriKeqsnhVgyanT+OtZfoD3Jx5ioSESjFjgo8ELk7+tht5Ev/czCuZBnF+6ln1Rv9lPI+IPMO
uRP2z0b+I01xYoldPz98ciNYFnVc+D5hDerW7FkS3ZUA6IxfEtgt8ZoW4EhWNgIUlurkQZq5jtLc
KvJTAnfeXD3nZ2EJ6Bv64MEkfs+yShCYmlipWj3hwEXMEiQymHl4ADgDYcEZfnQ7dvlvOPS56Cb4
3ovlo8YLHKwUCv597l8hFzS6RBZkDWf67LkB14uLw2q1Ewo5H8I/4DlxSpdFUK/+aeepUskGfP5P
vcl/xjCGRC79bo6ENf/RZFYL7j8P//dxg7qr5t11yMLWNMHAsxeEr0H3c+KtzAXEICaCFbnuvTT2
V8syixmDibvSucQrbURQnoaMcmg1UjaBOE/ZgR1KeXdO1uVGPqI33CJO2imY2aV3OZYn5EXsduPQ
nv3shhGfMuRTbnOBB3BlCvlbI40bDbLkB71nEKA8nHyC9qNhk+CiE0kDxkNRfOvcztWcWxnYRLfd
YD7EH4Cr2G6z/Mp6l16R5xRAuvoUx6FDl7mOLCdNRm3ijuyGua/k27etz3rONtkhqRXHj7YzwJaX
1BNE3L3mOUT0beX90ZvGH6kAvkG8wKXwQRUtx3V8xhESsT7dljMadzicsDlzHt01DMPINFYMYyx4
3nQ8F5ydMSb5DaRVhufrVWN9GcNXRdm4MGVypjDD0vMrCn1roRLBlvFYjWElYuvqPnz80WCjQMku
4mySwLFOcsnrZNgBRtoBXJH7PMfyGOyKMrkjL1+MWBTD9nJje9DjgthTwKfBQAsTQVcCTRA9wxk7
qSeNh/Pid58iUe8/YZkqQVZG7fANFXMgw9LBW3vDtcQAVpwA0gUWMvSDsca4Ca/PFmF0xpY0LSAb
7bIfkLfRHoMaOLPtSItSEKaSQQTDIoGTR0sWZNQ18TzcpfjLQFGCEXeMkGbXgV4EoASNvZlQOhc1
K4GhbwbDLHxHdDA0srtmmDQz+hYeXAu8W+tyjvSCvkJ3eYYzsYdykafa8nyEM7SorQ7TFYo3Hh5c
XzErydWyuY4kvtUL/oDsDVBaVJiSrmxOBSSsBn6yPIyP5inmrizk/08MZQEN0Kv9nsydtZkJwbcD
3ntgUP57tLjn32m89RcaneJYMDmod7XrRNt0CmeC5FGFTbdwNCnpVkUaQRsD0dOxubIxLv5p7TyJ
P8LgD8E+TWRcu3fQ1+3M/Ki85EfaIhXSEYTTtelYTqKFoOfKW/szWzK2s3FhRpWcM/AdcQYWG73z
wWu0NfBEzJSG6VS0G/BF5a2paXsy9QTxvWT7NhpfmVBs9RDk2d52L+Y2vZzQLpUmFZkenUXgaOu0
vGSBQjI84LgmsoR9PUgHC6OTiEK3mMatPux1OLdhyNKxdj6yYTzfBEqQASU39YLzHr+ETbTV/GH/
85YBCgJ/Y9hCKOTbZLCQAwKjOo0/fEvz5kko/1J0q/LcVQ38BbgcQ4lGTHE0z/SqyLwa8v/kxayY
NnqTCfMNexWYxKi+xLvOuIw/m9DvhIQZvFmrm8g3q+oiXdxyfWzka/Af2uyLLdWCDXlkacTVXzmZ
AvuBvprygUnISV4SzSuUnt1RKa5AMjxXUcL9fN8yzaMttEQuwTAO5Eyhvs8330c1x3xtNilIqNbk
F/Pm8EJFfC3gkZbx6rMQ6cRaf3/8gFN3alwZMPJcneRJGp0uc1EmGmhOYHF0a52WpRhtHVbIF2uz
FBEUQmAuR3dzdVZsV8ZBkEeDCCsFpXttzkOhky7hyUFNPRSauCRR3obAI/iT/TJTqvVIuq9eV2mQ
zkNwAfzobCQX2ZIg8DmXi0v/I7BlQsJUIsTDZAFDtcpuXYacsTDuadlJfBIKPjPR/UdGevint7S5
cO1gPzInzWKfMP8dCuATactvn7144Foa47VwpoSFnekzKOnKWmPtiGIo8ZA/TYNEY7PHW0tAhoTt
oGw7f12uvC8Wc8PHvXaCfPl4pu7dljLAYAUzWYDzawV3JFO9OPmDSCSceaHLifte66ShsLW/45+3
ZKq1ofl6s1mXpLY0Brtl7MZePf7tYlJn9Qp13dOZRtH3a6I1aezKUXqnSg/BMQAh6p2T2Kme493G
5JlHabhEFF4nVYhA8p2Txc0JwU/kjKp99sh3UQq14yMfSxgVwxBr3CFpaNbilumWsXxUfM6Ep7kq
kbGkogODoxeFEpC8ST+ksdDmy82cA8uEpQ1HPmDog5ZKjrbfor0IvGThnAxNptuiuc3PeW5eR9by
o4tfZIDRk4qCShybcSUQtQ/tTZ0QZYWPB5/HAWdtUnrU+WMOFgSaUCnGOrVpjWiLs9z9XUip9KkH
wwq1LwVvxgFZn+yY3qnC2Z/AgtnX1huJujtJSCat13SqtOgG8ntZl1CDDh+9BPDWioyxGwa5C01+
tatmoSWgZeth6aKS3PFRA0AkWRziZxDixRa7CA+kQE9UOGhwhqrv+7utWuwb35AQx7tyNHIqr2o3
/QJOwqmZMoRQmxeB8dYSv8G2IYoBxU/RibdUNOqghDDONY10muGa5x6avQuEWVdCQY+cFb4X0SId
My7JX6wm69ikD0nOHBji3ET1i+hGPhV9Vk9OGWYRh5tcuLMv4VCSXpHVJxf2BtuoA6Ek4BCkjEeG
OQc6cBElb7s4daaTCxTNRPVItWKu5XKCvPxOfpAMo3exjPZ03aJSAqwRxnmfmZekyCcHbrPkEQlG
WcnUJQdBh3mypQxVa4yfgZhyO67h96LTHZKQTfY8SPz2uCzNYBnfjDbhbKvxK56n4MkGvIOFpRay
QqGFwdHejjSNepKRccHR7kUAXD1n/nTazr/g1QdVNP5NKg8zl3QDPTbBZfKNHPg8WhZznRAgYUbD
0N3NakehB8lXKEsTmbM6V09XR3iDMWZR+dqnuXLyqflVKOfh6gCiPPmIKxKPfa6B41pJXU2jYtE+
TJpcdbj32nXu2spxSSWuN58STmB8b9NZUzLWlsMYIK++pNu2OdtMAp9jSSMz9gSTzxyNkHYC4Fq1
qnLbcS2NIsyBmH/xnu1GWNqaUtWywOwpGkadeIr2GN+p2gSz/qRtDeqz2nLmmR5/NDsHTIsQNrzI
MEUQJ9CwstGu894RHn2XFbUcZCOm1IEqH5nDDcdqZZN8GHgbAM24uamOxwpKiusw4jns8ra1oZoZ
ySZL9l2cSRFDBS2BKqgHmesoetd0oBIfE6NNwZpTfglotiF35oX3vV9nqoX82ghnzngHddxKtzX6
0QepB5kDSse+keNbohIg2i8RHCospdbLUlh7gWu1jOSMDxdEq5DH0BlUrddaOB2eu0EGaqTuJnyp
/3211SKHUNrWloW7Uukt7+6q3WbW10G79JlHQXEqvgxoviFoWO43QTDkshKQT5gcxCYBD7dMR/Rr
/tjrcAZ2n0qgBLbb9zZCYyYKewx3dXyvGXArFh3I+d5NjDSQRzC3odKeg5eO0LfwVzxhBqz24Duc
YYedpyqto38Q/g5x+Oa+IIWgGcIsU46flUvUtmX1iqz/tysgtukFN+obO4+CtlA14JZLrENmSKDI
WWXywVrEdx3dmJVpgtLUUg9EyLOB9+KNrY6EdG/r9mpxV3TaEwBgFu0O2cTiMUOQ1LTJBXEnpTbC
GoyKyhXWC+ywrISQHaRXUvj59WD+31v5ogO/dkPcYdSlMRfNA+it/U6J+6TVtVuMRRYA1ewkunxm
V/NOpLKk0kfxUe696wLrSOciS7m9/hJBRWTsHkcErEYI8p6JUdD9zuglkVLu34RKoxJs8sevV2Mw
NH1z+zMJTTU3SdXFiCk6492DXeK+Cmj09msqr4/3p+ip1nAkqFTVYouYZ3NO7tGRKtpHlwKzHpNS
GF0Iygf2mzBuRVsp7CztdQkQvqt+LNFgeaHhS5WluyhPv2L9/7UItIpR4SFEJuDIwXKSKjLHdoBp
Yao/ZSbwTSU6jAeJUw/gv3W3NFWxCmPd6YhIgotrBoDVyOw6+NGdzPLYG8bvQlKp1b3yw6ws0iv0
I8S7IAcvrPxRwG5uXNHhDOM2n5iIOUi4xjR2+ftrt8fGC/x1+DbZnrnS949/cccfAc2D+/rEovgv
68jBopf7hiaHDOyt1VzP3FRfC7wOc2KGQ9n4IP5b3d9r4dNSuyJD2uKIobPHoDqEHx6oF9lRW/Sz
lUApFVSHRdK5ae5Ddz/3AXvEezyp0bLKBKiv1GARNbxW3Czjtk511fkR0jyhqQSU5cdB8xFFiIhC
xoJsfrEoUhmvjIBFj0vNQi51GJipx6mvkdmF6bHBdzGTJmXIdEA9gJUwapRJuVT25zv92i0eQzvA
UI+68C4qB+fp4S+SXjWmKzkcFm9hFvPXAq7LZdIAaOLR2PTxpgvZFSbM+VqFd5PGN8q2YXhdfPhg
mk2pLnYsJN54BpyXiY7+4vnaz5+dss00kqACa9n6om0qGZv/GnhY+MhJe/nvB3zcUprXmeR2dRuj
V90Y2rk5E9z5c74wRowa2tAkps7YGfzMPsCSf7IUnJOXrMZI2O8U/E8455neEAjjQaR+AdutRvPR
7FcJAK0PsIGgYlIXWXroBjE6WAtx4cDH9MkQJaeMH15qcC1dtjEgUDQHITKWg5UAy1ChtOWvEoEY
tO7fsS5CvSDkh6Kzgu59LpDtGba71qLvIc5vmW/pRjrHNM+zjKWmHmBxgqrP/rQQP9LgSf9dQEEB
sceeWvUAo6M2VVikSlHYXh1VZWvx1zAAIYoZidydwegYk/Vf0ao4tLH+AxuIYtAlQMPw+tyOxNLm
kIHxpSVobmmng+FbJBKDz6mLk7BSsKHLXtD78eGg+M3Liji7MvpoO8068AqJQhW6L/NwoJrXl1Cb
EEVr0qx+8fboAa1MxMRhZGv8ynHqJbvVI7I+Ay2VwHHcb6PYZHCr7510Y/TLIiJbLjXvTT7f4jrq
adnx5bF6/uJjNFH3MAqYBNzwzufwzHemZGn5nLZbb6cUC+F3wz385QbNmyUybYuvN1CVU79FGLCr
pZsBOepBWX/fODksyWALV3R0FBfFk8m9VhjKZLuSooF1mdByVzCdSNz8DaVzANKqQLsPcH2kg7wm
berJ/4euBV7txxner9bYpG9V8B5ODY2wx0zqMF3hsTF0Lhjxer0z1+V+HnDMEgw9XGvxJiNa+6vU
PPk8m5pnAVC2ZwoBpgYYtkwMLM63apKA8720Oi+oXf4Ege0z0uwvnynEwh/EPw31n1mnHN6Ij/9u
tBj7fIRoYah+nStETy3mp2uRfzgcshKnBwlLV5b4OLaWISX7D2jiLTWmaWL4ehPVsNK5yQ7TR+ki
Dmr4nqxSxuJNkV7CrjJmc0K5UmyjPsFbahePLS9SRQoU24XV4kX+1yfHj/w4oh7nAHAoL7mZawvw
zxA/U71GR6BPmEMAaZUNYAYP/faPR3aklwiOdGsKGGgcM3XGuWrs/EvXHqmqf1xNcwhbrf557H6I
rJlPpFtfUUo7Gi+p15o7C9r1YfbVZf/0RyraOIyF3XyVd4gKqZyESQpEGAKZxP2apNOn2YIzuWLk
RcS8S/V1b2vvZWsmA+W3wkuihn22wgd+6HbP9PEWHvaG/+eivDVNR3pW0W7d30c/jNp1w8dTSJEy
r6B+IrsDdJU2ykKiZG8o5X9giOBGuJD+QNs/FxebrQ4W+G3WTqDAmufAfGZvcA9nZg0h3VCOfLUt
/LXkBEG+MGPCZAClM7cqmyP/8hpbXxPDKEbqEtvWpiqOSVhKiQZdp5vQq2vU+wDgKa5CREDMlXGL
zgD5SeCxHloE4icTjHJIs3/6Zl3zSjCx0JGSQRr1y0jXz0EmC4z1UmLCW7QLALMGiyC1zVb8A1pJ
R751vhqBfYOGwxzcal8Do1cutoVYphOotS9UjQ3RZRDFUusv3g/pDtfZuCAw92hgSS6GxlGh4ml7
j4abLbkGOiKN1ghliL21+HXA2FCOftqfrCqTfIdXfVocBDzSImF80UmHEZRCEXu8Al0HKBWAtz+b
Rwdd/vKOQmnl6bBm3dtygsmbDDpVWsS2ijUYx4etHLqKZWOwO9qkJAZIMpMcyIWFEZa9BtC5ooyK
ia46CgmSu4NUvI0IpnMaJb455SpNhVwZOEjxYsSW5isUplxm98mo7osBCj/7XrnaopYVSLFqJt83
YldQyQI3L5o5+yopPOfw6r5VL7ytKlrYfBb32wscP8Rqn+hPt3VGF/f9BjgGGZYxXfgkQ6HN8Fyl
YwnEr9ANyiyJzeOJRDFv2TF4LyWsNYjGsHWq5svKlaHWs0derz08fA5OhMh1yzehFBXvDyo9wWoJ
w1a/d24E0CVo/GXzcrD/wHOf13SJejUV1vz3YoCyzi7TO/6Oc2Pr5gCSaf9Smz5Rkpjsd17o8V6g
BNtBsHWMW6Uv85pmShnyQyp0jQteZeuIfZ/yiOZHjK/RY1TMfwHIfdq0jAM0iuhVapvf3E9cXjid
TwYJAIZBKRR/0QvxtXrE4kET7+0Pm5LiNLJNhtW6wg0qq7t6YOgap0QAP4ZLqiJzBwNeqALaYfdp
eAymE3I5gOTGPC7lpFaOcPTXd1NWFvDuv2z6B9pYx8pLJ2EJAiR0PARuqJvfVmBJM+NzAbNaW2Yh
67e2jGBVgBxL9dKavTTjkAUpQYYg3wZCQOZAp2Jj4Xi/dgl693YlbZy+wwcwkXzoZR/twMKErtNb
JsUjRKlR0Bm11+fE7ctGosoix9g0O6Zy924X3jzwZbeLzOSZv5YH68jNfigxe5vI4KWhUZpLdANl
S64jUcJu19N6YOrEs3+rosv/5smmdSoHX5blG42gHR/dSlmcGpqtte74WRvk3rEGJXb3LO2mUTd8
r3AfRhRSqX0lu2hXnd2sxNKVcv5czzh6UgPgAxp/khuGiwoxDnhqIymrSmf7SGkGK0KR3+ZeY+4N
AQaI1/he35jcEJ4cJUqJE/ggMFsVHZtHg+kg0o3vmiPCCRfcRFVU4OhyQDtr7JUTSYln8RKR9raS
GBpmGKyG3bS+g2agVPF9tNGnJpCTCFEttp/wyFdz+Un6fZU2Q+ryqlZJb6Ba8/6JYSZZAKPhtqZ1
NWtHnTxLqmBaHt23DN8pio1MYE1S0X6Tg3K2F6km7TCNLH8Tp8ILfRuRmSBpqbRU4NnPBqgRHsoN
CCzK/U0C3gc/4xMiB0A+Y/LnGyQoXEWSZwA6Ste3siHmJGo/ndOI54pe44rM7CS9X+yNYB31O6PB
zocJWyjGLbnPAlWBdphglBE3qh5htsbb9BcYhLyf/HR0pobQayBmdeH+h7n4vEpNJnlvAVYhnWFe
AeYsxamdUrwWT93AV768rBgLDWm0B5KeKXDJqaMci5xxRSnt3dwfcrwWGO5z5uH+OOKdfLFnzeYu
AAaNQeJ282Fg+iKAR5vjOv3ttz8OJgTRLkWSPh0sml7zuuflaThkfGP9tJDiXxKZRA+RgzZTy/C5
OkdwW4RAITD37cmQDUX5TIPI7VUkSNcQ0yETSVWvw7BCsxqDqNftzUNKWAkbkpqlsMNqe3XCz7Yj
2v6TQUEoQX515hYQYQiEBxJmpI1xXXWZKaKtcfgQZwBQ0nbbx3v2TQYnef9l7pSEsc921NaWHl9C
MSfykob9C48GnJe1JXAvPvJP4WVy2lMnZsEqBjCC9GO9kvnwCwZEGKXaaAboE/tLJW7+bW+niody
zYiEdxlavne7lda5qc92/WWI6pmLEQlGZqK7Rg8dACL8yRJyAlKPDtn+yXq3epdS1sHJV0iT7qL1
yWFocblYMqFHtzS455h3aDOdVFvJeHTiwko1FAN26njxFGhJdcVzGvJk19xE3EcWJQNnTIzrWHWV
bfSltEiVvAPG0bn7PTGlZOWPJh9oKb8Qe4tmpiq0UgwdphxSFp7PJUwZ41aOQIvgp+p1kt1/P+P1
Ol6ghnTszCGgw4S/9J2LxOODfHX0CUP+Omg+vU1wkJsGBrhhR9dRoXxu+S9BmBTow7UK89pcDrMC
kegOhfMBDiu/X8sI2C5lgXFZjtzlHPmCsNfJ68CSQ6nOc06rAjXcmLI1oNFgXfu2Fu2+bHRsbxG+
PmGYoLjD4Fo84fB8MrwwuTtI9dTHxt/6cyTsVJlBsoDC54vI2NCgFyAyB8vDagH0MxIvr8aNELxH
9VycDKhGxgj8VS3xyU+qsdzDSrXwTFRxk3eSURA3O+dnFdVkZDCVSFgaoS2tPk3f9PHf6P4tjuHp
+V4bZCTu5yjeRynd2BBePSTBj5WGHZDeb6QwBAh9pibYnM6dT4oKM2oAvLXhT2O5ki/C0fZM35Tb
SfivcaF9Uq9xZJ7mglYd+jf3yrccjYSQykt7ch/rahgr45i9Nik0Ja1Argw/w9hkSEyaBqS6okJZ
6JQ+gMwLzYAE5U5bUyUIMOIQDDeequ+tgUkrTsBD9DIVT9Oi9CK+vQlPNCT1d6FdugrU1i/4bU9U
QnX6u0Z+FjrP3+qM3X9Xbek074g2/vjR+lT/vNgEErfnF2d43J89B1TmjknjmL5SJ5RwwoibAt2U
dQWi5Q/YBheBC6w7mkgY3hvStSj2AvkrTCLAurGSriCKILMH/dS997HZrhP8YcJHeFudUXYV26WJ
RndMjyUbo7i/2QOpI+p/yNlQdaczK2PwnXQ2kQHlhq2eS6L1tLWJclFKg8b1+FZDJ/FLIr86FA0K
9L/RipxETaZZx7o/p8wBbUW921MOo+cX/HRF3cmYinxbEVJn/3Gj5omE/umM5mhMvRqJb6xD+dUd
5ntisJGPxjwZzGqnf0tlBJmHbksRo2Pn8dt+hp22aPz374fQzqd0gBw5//prpIfJrT0aCqIZ0oPS
JQJNqNniBAa30ATB3hVQ8jmgozHrRnSBD/YCRZ7QUJET75qbwG3FSsldzGzc93GeMgBBdTwnMofz
vH7tRdCm7w/LNxR5C6ZDOHwK1ViEQE7dK/3gqJb8P+AQpaajTZ6y8nAt4xlkW8Lirubz0e+vdJaq
qGO7Ld7naJvzv6KzHZSrY4kZT7tp2M20Wtq4OQNgq7hXOYHwxXsh0l2KZXMBA2Y059ndNlO8EEMg
7xVVFcV5mJfrpboVbOvy6nt9o0E0r+Kmt0ok24my7g+8uRIMiSaJ3gpczfX9RdZNqlLk24Y5eGap
/RfwH+Jggnf6WGcp2xWO0Ytx8aHAuFWTOpw7GL0Vk+fZiU9STo5Qvfi6F5pKELG6zL4f0YTuRt+W
7zfRDBa3ZnGmGcLyzJo8rcXKGBoyX6U4cSpW+YSXXPf+aOdBEYbtecZ1honAv1L+yn/rMMhZTPgP
YSMJVC22tNE0T31kjrCso3nUZkvXn/0Jv8EsSBUDr0Q66QfcMX2IcjREaNwo070wbhv73C6kwDyn
Dn/kw04XnnTUrYZp23SRN50mxoGAwr1PW96R1S+uFm9HyK7mzfWmWacfkvTsaduTOi0bQarF66Lj
pi41PpNAhZ3Jl35jeGnWMkfUzJbLJty8HQdFv5EgY8A5FLEuksl7H+fiTQc4HQSyzjwd+Qh+EL+j
pr/CLm3QoHdBCIyPWUQVoPRQ8GODrMxMZ1lP3sd7pj96AE02s8txxepBZoz1JId63wxpuljYjQLs
PR2ael0/eUHfguTLEbKUwzwWJTChdMnDYWv8iE25FD4NYyfzDC20yQxhXB9n4IM4qvOfwhPrPbQx
82tYATB3t6H+NtqXqbKazBnEUkN//JVqtFRfQiDO8cD10XyNZRwpIpEdf68LD2XACFhNjdKbrTuc
MYU3QXraDd8odMH9xtM0pz+7e3eL28VlXGJ2oVNJL/ydo0c25RacIXcyipZeLfzqn5Wzzuaa/wmL
kcC0lKUnYiHJ64cCqV1UNSdbidbMy574XRQkT5AWR3QAXtAxFxL6PKd7O5pSVHAYL7iNcGKmWC4b
r+arYOAklwuIy4xjdNHJbPKbQxC55SP+zyHSH88b8uP0sIZK9K4bJbDmiJTXzUgoo08vgC3iG0Ko
NadrgkbIkezraYOK5AbqI8lT/uPfpe1K48zlM9X36LpO3mJ6PS1zBe7F163RAQPa1tn4AGjLBL9Y
T2ZYOISSdEIZDlcHsVytlWdoj8L5SFja2fjUbz41tHibUWmzl8Xr8958biHB1NHO59uWGIGVZRUJ
wz96+7kkUcnzWCOUFmaOzp1DLMGW9ALrjCkeWGj204qZxI7wHMYU8Z19zK7n+3rzotBAULiewBXY
e+TJtQT92H9DMuhAy1peMCRqODBxKXRCrCEflI/vlOrwv4Nx7A6/W0zNn/MmzedZzq2S9x8JGMtw
kxn9rNzhGrbfwllixULum9E3Af2JpMsW1LuJYwlVd5UEcCqFRkwdgNSP6iblMkslAj5mSRyyzx+/
oNFANxDPVPAjznWzGSb9mjOuxokg7dZZBedsKjMRdomqOFuAf6u5np+JRdA6jIdGHleyGbMYpeMl
pTiwzSQImE3r+oDmE9QprGphhyLhvdGIII1u3q+lX17oS588Uhz+IGenxJh9JfoDQptOgXBGVWBS
IgyeJsXMX7CbG9vvFPooxehkGEJJ0OHoHu6p5OUcADXBIWvVxczOYj3oGorpokDY5K1SjgMB4gZh
/kR5cSRN+fzh8nnVx16kOfgAvVjHtxSO6kYCWmUOKhZK8Qbi/lt73vsyAj8Qt3XkR4dQXum+RWxf
EppCe1Km+t6SJvzH3VPd3tU9OQ3kWBIbbom36t+iy3vkPuM8pprNaLmzEK4PPquysT96Zx6cY3+D
WP3QBajVLKGNHYc3JxSHmYOPGEJS7bMxcP/HzbcvppVzc/fy9zqD900BH6sMWrSfaZapKMfw4IAE
YFE7DT5i7a0s74LPTA1hKj9c2tepWSUAo1pMnfqDA7dMSp6lpRLIHdxUNBH4TR0ULDVVNWZZJo1w
uhdMadjL4rg4GDq4oNnpb63tPQuzZ8FIKlDkbz3qDe3S5AUWEEQfNmjqxpeeC4MQYJxH9PME7Wmy
PE1jwvZ/zsH2yIpyYFyz/pIqzshZt0ubrrF7Ny5A4wZMWmu+LokfO8qSIF/wDvd4vjYzGBL3WH1u
sS80o6KjPc4ZR9gcu7yBOh/f13uJNWuWvd0JmHO/ApPIu4Ay5Ueab66CCYySsJmxOFCVcXjqbF9y
zqbLKIwvog8sWfn4j0dH3blXK5cVK7ekwmjVy6e4HRFy9lU2dNb83dUrnOdzCav1ysUeYHHD0Za8
3DKFvQiv7AQ7G1syyOvpfbQK4Qkss4jbkRMprIkazrhA7eTuswpSoB81YDToj70WIVvVMsoZQMZc
1Gdo3NjMjp1qHVFMDY8GzM9nMPvuU/nHSMmeahRf4oC+j5VV1JkpHKYjZrbABfsrrOvy027Yz6ho
9xllMlrvtHUbVhS3EcSgoGY9AQF7VdRSwH4NKDvhpChfI5NaYEmCrqs4r8bV1ZW/0/9091td0V7i
YpkPjKRRFey+vZbDzsClaHMszNu0LdnORuNcqWOelHdel5EuEtSrzjTKNOfZhDCD2hte9jQ0peDr
pHe2BamLLdvFAJoWdSmzviKN4md4ycpyp0sZ5YFDNYSJ0q0KYu/X2tiLvvxqnqjZ9cKTC29M+NQC
XLbcUCFBgzCkeSxkriH8zN8eQ5OCThh15xi8y8i065vu2IsiLMLdZ1gRMmY80KAoHuBHiK/QHvth
8rZHqv5k1+0rO3KJiXe7OT8AQS50dB3l8FPj9RK1ToEoKI/VtXd+w9LY9kV8dYkEzgCSsyE48aCS
YKb7a+/FEkLW2ggFUhvvFc3GRc9GWAOW3Vm+LaeAcjFbi//W54JlevQxKB8sUmgs2mIV5scwFVzQ
Qi37SeNr0BHPyb5Eg8aF5K+pC5tIaqmNAP9/l9/Ta9NTCM6IrMyzVawhehnRSA7I0u+Q2eVfb5nr
7p5fjaZozbGR8+xyOQZovk/vuorObxXugO9l2cbygNCX+0B7hJ/SX4nXGzy8Kl8OqsCrKqlEieJ5
580VGjx17sDF296EhD3EBXzPmIv3eVbENsEZOwl8tyfPmwiw0HhTxBVqw3DsIS8vaK20nj/K06ID
6VQb9r2U5Jsv8isNrBDNcwewqojyBIqXp+uC1a3wR1Qzr5PZSOZifL/8BNxoP/9tHdNVSh+vwtMr
Vzcogbrq78hi/xEFKLxaR67kWAIy7iqD3/ohbANM5u29dH6VnISbfgjnPaPr6tqWOePFz4W+Yo28
bujKSZ5hyMqI5Hfwu0vDt5RJaXIBQsEfPCqtoBrT83QbBbB//gIEz9IUeUu8x8HZIdGTOayxsnvP
Y4fXMH93urD2M6yzK6r7mQE17eZOxhWv+2hq2geAH2B8SQHcTW8DiP3upemNXyW8mnlylkicRF+B
sLfpuxnp5fINQZlwlExNnjWB6lKw0IejfAncQgy1xrC5uF/Jt/Pz+SoD2AQcUtZ5DcqaLD8yIvPb
yz2Bk77KKyHyGsHtsXjyM0NwNi9bbtsNDJwt11cj2z++/lA/iinR63vzufD092LoCfLvhAfLJWy2
Dhyi0vGgZCmG3uNppKc+/dHsDbdwa4d4xL0vq7vYiLgdNvA5zwMoSrZcgTbpkhHh1BF6nzQHOYRO
V3HDIrsG74rBpsFaFOU2sNb9ISeKeAkt/67Z+c00R19lHETvY2aQb2+w1ik5DTKa70Z3pVpVNNAi
2RNstUWlIQe5vMfVOSH03kkF85c59jCFc7Yp9dActLiIA1dv1nunAT2dVFCZWTl3/GCcLNnUJJ00
OXs54Qv3vVs+Cwx8P9b0AU/VMhRZb/v/lWUlbbf7Bkq+y5Jm979trb/jUiJFjsSM5ARPyAJ9dtA+
46moNEaNuDfcgte12hGfoaGxxGM058nfXx/onHvyz6A82tPiyn5bwM7SIAM+5rK+hwJX4VHesu+F
7Ov7ZHqDGG7fUg4fzbd18KdwxLyITGjuJv3Dd7hlH64xBwhvq7h2x5X9xhdICOEOKn5mzOG3ZkFe
BvAJv/L57532OWJ3+EgoHiGMaHutxfHb4wdxzAYkO4mPo17oAoksYdyyaeQKbpjjFklY36eQA5V9
PyCzI3FhF5ir++bqqdHTfIZ6xhlZBFxuVgYXbGS7fS7eDQ/xIF1XdrJs3ze01Ly/hR8dDQjg5RDd
nYr78Is2U7nObHKkIydazOTxiHPb2TGQwU6OjeZxmdkDh8jj6fgz9QA5yqnWQRBlcvICIM0vYF0+
Szj2W2oPKf3x9AAO43qEXKXyoYv6vuGBlM6tP991sYKRWI9xSDpavODj9es49/cRyuhlrdVkvAGr
1Z0UGC5oStdrd54mvdeLP/fCyO0jEd0NMa3NYY5NigEaMVeHBQRtRPjhnaM79bjJ3z1vrYbYGdA0
HhgbCtEJnJsIetFLumny4PKBNoktRPvHmKjIBIHgMR5ScGN3Ms8ZpdoiyoifMPbnrHt1YjohGytk
+rCcUNi1rmKWMIulUxUh9neMSTHIw8+roTYCqpoFvZp39Ri/pFJgvj+t27M5AFw7oMPxnpR77QAD
7r4b0mfa9MjylZOCC8DBHBL6i/CroxNVqljmwPC/qHxO9Zfvrt7dvCzrD4JG86Nes5OdJ9lYN7w9
UjuheI6urzzfjWqD6WmAPD92ffFfXq/H82EYujQrIXJruXOkOKJxucxXn3l2JTjH6AFhCBEtSh7e
CfjQjnwlnlweJNRNQwMq99An1C5VP+p875RPLXMZnU7lQPAdW+WsGdbwLp2RTmyEuRzbl5Xh1QFF
mFyM/3gRP+riBdw1fwM+YJw3GdqEYA/I1d7esqfYn7Yki/1EGkZ8L1+UC/sulIfC4aIYWSqpVoGI
zYiY+bP3XoYp4n7fQ5raLJk+JtVFtyqqpTSbbBs1G2nX5gS1TkFadmrccIGyM8MdCKZcDj27jRIT
Wdn8O6BvOaVIfGX8lukBcBI+n4gJdtuiNmky0+yXePmqqSsafC3pfrsBEozMfwB0s90sOhLiLILn
XZFseQXMsOPqZJcagYwKlWIR2Ld3Sf748sR9CxyBUEoCkOcQSPMPALnOHtjgBBNbLdK+sTLXM7Ho
MKhcjAcnAbJQsq02zgaJTRX5MqS0Mb1d5TjJzpkCMUIS4KZKLPusuYMJESHD/cB0a958v11RdD/M
Y8DmUpgUzad+IK+OtPxakgREj23hIXkc8C9mv4hIBgeFk5qMQUE5zc4XQhMQLdwDpozP58UWAzcj
epH8CwXST3jL0sg8iAmCqVgOjCWoThCinu2swrM0JhioNnNZVYxYbU2Kd7hnkHBqJVuNA5VIWCUh
nimPC9uo+qD9zquMdrTPdrIgwz6+gtJbW8VwKdU0ufDbLAIj9N8u/W/TpSaV2UGlo9Q8dNGgesKD
kuzz7cqEItWtzs+B1MsqxtJKJJBCVJszG4SwAal6YrGjtrM8AZxuAQ0WG0/Qba6MTsypCDVLQUXV
22ESu+mNnhRLdfh0Xqdfe6rCywVSz0DG1N7HeCj/HiUMoSXHwSXQMYKts0diT8zjZJ+QtKVWTfiI
uyz0q9AsHICMyZp9G5vlS5kB0Vm21bcTsdLcFwWgQJUn48EMrWtnlQsEofOoeoPnionbQly8cGy2
MCrg44n78b83/PHtwQaaMwoJ4g1V3pXQ4R36uEDXe6p37fkEEB9vNJM5Q3skiINC4A0NyNOmd229
GeYvEM/RqQIGm39aLoY3+r0pP9C1Nj9tbYrAhHvPZ0mKiemDz5rCkP+OSXzYphjGlQM/3KmFxc0n
Zp+awwxshZP+5bTJ4g8np2r+uVKpLKpobhJyu8Noudf6vgRZYHxw+631onn+7lRXmaWUcmvCNMlK
83zIWEI3Vlhh8h9ARdxIG6pgg6xdlv/CGWidcfryMKi7kZoQJ1byhGUXPPeR15Xpj8qIDJ6KoS5x
zreO1M9WMw1A9P2WGSCDwfdd2zv/2PfY9sbnSuCnlknLDBGEaglpmBXwQ/W+2cSrAkdxqkF+7vnz
q/QAL0w8/rnGSfl2+BUVbK2CfaHH0AQpfIMZHGD++jbkdCsYaDMvbJ+MkviqFeu1sAlFzmPVQj9Z
fErMSEkX9WnthuuxEoYJ0Y2YUpoB6e/DFUvnru3zpRPJ+ISpxWV39TNkepP0d/mBcrDI8tJ+7hYs
7bZOi0/thBZBgqCyhXneXziBTRydUZ/PRyBtfQeU56WihZ+x/LCOK9nsskIsC8kKYVxNTkaYHXF0
nB8XPf0SSMUAejwCILhQQ2Ok0JwRUR9p31eHBA2q2wxBbJblpGbFjRZAace7OnMfxV+wciDxPfyX
Pyfqm6dqKHFx1gqCcb+6liW+I8mnMVURsZ1lB/U4oJO3Ds3adOJPwjyfqVQr6DdiBahofJ2Ccf+I
c2vP2AbZV9qk6eZizjQp0N0UKEm1ZQ99iIqb1L2F107iANibliAXfqEJdkot0W4eCMYz9OSS8A8a
bC01ctbtdyZOac8+AGTTU0RJSuS4YY2ESZ3tQBnAps91bjVav2okTX4X6F3bcwUlKElpCse3L1YQ
mdYEluRCHGWH1efPcZT4hUptxhZScGe6ikmFfkpfjqDlDQ0PgTUlsYgEsbGq6+SAsheaL5wKLJkw
N6CvYjallKFWjn17tZOcD9XyoP4z3y5wK0V/qkfzsDO/d7xvNWRr1ar70oqW9qktHaqosUEGc2Wp
s7ipZzCK3ScMffC1BisbT1HJJNb/bzTAYolzstytjQm5BPkNuwhshy2PrKwYXendJnIbUQMbpB3r
Q/fZXhSqYSnso3HPSzWH/NCrAEuUZCa+wSqPZGRIGhv4D4NjccReatrZBARE1lpCgEFXD2mgrO55
sBnXegdhCIcAqCphwgk/NYUm+80cRsb5HDOlv16W8oQIPCrRtVb6rQQF65mpU0umtbia+UeqM37k
0SgJ6P4OIiKitTreFYeeuBShkxYhT39+oSccYi4fCs0fnHM0IJTJSYJW4vmSErOwQnduKag6QBER
7ZEC7J4tUb1i/DgunsWrHb1HATJSwpWoH13ucWFgBlqpitEP7d17OwLsHsGbQlG4qO7lrDferzNW
KbGbIZ7Fh+072d/2G///FA7Eg5ic7xSW1UHD3Po6z6h+OLGZkyVCA87dQhTOm/HGdLkD2io+CSWK
5JJVqYwAu8WUUg3oP//UEnbjbXkCZ81daW/sQzhxm76lDiH8M8E2SwyDKiFVwHmzkL/ojE9ygFNi
nIUW1/97LLMud3Kv6DKcv2mNzhW49FqldnXdP4hOb0pwUUCInmdupTgS6bf12QFtom0ggt5fRvRP
gHhsarliGd/kQI11ZRJlF4BJxuhIdQRmCXQ9vLqEbJpbVq7h8XBOTd4BfX7BqxvoSO/0ZWrSPVFI
IvxXISyDcaCE8YsurQI+D+HQF00yuL6sm8jQBGbZ70reUQZIF3vQhFYKOqXDj96pEMwafzYZSI2+
NFEUcFlU/eW+E08SYnnbayCWaX8divbGCBDyQzywe7AYwVzHGeKKBNTcOJqmnSgh38tXobKQtRD+
0WNB910vNdpShcoQl52xHTgDXA3GjgrKlSdLWPGX7U98hcZnrn33g9NkfKbZGFtTW7zMld+fh6gU
SyJlw/dd8bRvsMYrBaT6/Y84rceOamOzVhkjM+NhEZLq1eryZ0g6L2T6jXgWmssHVWcvYMpCJ1uZ
Yz89CaUrA5s+5Vs0uaf9eIOnwJ9AsSxt7thyANJNaOK0YfWsESRYwjqU57Riz3sZfmXd6OMIWmqZ
O3/cyWKPgN9A1JcluQ7StHOgK/dcBO4TPypLAVJYOedErFBEZlvaqhQGojag1hP2LfkL8zwNsOmc
85oH2LIDFeJBtwm54luhMp9fAXmXnSa8F4kCJQ2tjS2U5fSy93iyIpX99dY4NiSppj+nK74lGEa/
qXDZlmEEROOG7gayKpRBZI0Jm98amzwwR9cPLuKz2FGfsdJL93meystvNPpGFfUhSahZrVFed2I+
E0HM9hyoQh0OlTiZJkpI7owznlCnzvHO20tAQJOK1WMtwhMP0AHV+J/JVsJ4hdYqAzUZSHWeKDf1
ErYKHCPK2hkvKOjtbUPsjnNzM47hf1RK33yDt/UHATOVQY4DeRuCx9IwWglDOVGf0BNa09gvNBV/
EAOxvMtKIH9I19Vr9OY3kd0EqQ+85Zr7/DQOx2e+vrpAYK9AXenmPV1euQK2Hfcq3hv2/zyue5g/
7EMbF13GDwnVuKsZ9gUBngwNoh8s+W+tjvFtzSIQuN68rTlI44EsUHSLV9u6qreP5kGOtZFcq091
2pP7dR9Ly+b8U68g2JYC/C/U4WZAdO4DnXTsTJgQapteLcEy9dJ8+QlTHLmE0RByrcNRuDg9iZC4
zYGfaJQQic3N2SzCvTShkQtxTB9WH7CJa0R9BJvuveIDzZPSdVY9kqD+Cb1RVzCNTLLRbquD8QWp
35K7KV5rZpqcNzDkq3jdKgashfzXsc0860HixJEFQDfocQbGlL/0joiplDYTKxlYKIMN9BZJiwo5
5n3vDfzejpM1rvTGnrNBSJXEp/UgIiJO6ZV71pKRbV8n11VbVu4lgroadx+Y6Iu8UmegwjVluk0U
Yv4F9aAXqfL48qGyNYLVQ2zXnmlCQ6Ayd6N+fBpyYT0TLQ6WEL1LdsSTAm4peyGEVeuuNC/yQ5qO
iGyoz9zDXxsIsXOTzCKwEOp4oLzPD93VYc62nbNwGDzVuxXpOUoQQUH6tFA9c2L5pAcPCvmn1lz9
/zwaQQ8klt73gFRYK2QT6PAc8ERLqliXJ5zf42qyvyoUsz2b81Co9Xu1pzcRplaB58wdezC8BJJ9
pMmtQp/1ytXau595u8GNrJ8v7K2qwX74ny7r0Jazg6AHMKbH45zcb6GeDKUth2RtFlfJKjgqbZ2H
HAjq49ZJGN49DUNtj9UqbHLbHofjX9KMewKqv/WtYdhjUPb6RsFKs+qOeV+jiYNaG5We1bvLgSin
QFFxIhbhoFPQu2iKYIXwXcPSZGChpd5aFr6AriZWbcczCI9G+wPeoov61uapgtPD7yUvEvQuC/8P
Cd6/zMstktDCfrCkHmFsC1Bec+VLx9WSW3Y6I/um18GGmDJ091ga6+tMXiidPcO1qpnr408Y0NiX
eTvb5RbhfmvT/UKu/1A4dNbim4yUchoInX7iZ9USVY8Nw4HzESOUGNJ4arethLRVaHEs48LkkQY9
9uqDDD+kQnbgOt5ABrPhMHHHl4pkTP6Q7RfbrCuG5d3624mMMmSR6iJpdVZHkbPVWSHJKIUxp1DD
ZbUaaoj5idpD5SWePKMF0nRKhH7CocS/0iYky6271g9Jg94XeFVnGNO9heryZp5mCc7ZmosRvTVb
qnP+mQyNgrcU/SfdlfLcRUZ7I5XlGGtmBNFNv01PPXuPA10YaecZGM8X3UyoGFNrwb1VG+aEDbfB
myeJeY2Ze37t2fQJYKn4cClZ3RbxyyG5XBcjwuh8C+Lf9NPNIaf0gutty4qItGakhpgM5TeXS7Zf
KGoiwi/+fV7cF5/f8208pP5HCf4suzrAJAc3/zKsI8tzyuVWQOz2KhzbibuYJSdIsj9ItovmHqen
mcMNhWJQ4dRId+52eLN26I82/eqgF3/O2uFzkND6QDmD2kGF9AN4rXFwkO/lPP1yA3A1y11Dqqmg
mC0gohk1wL8+U28im7oSZzO+V0gg81wLZ2XwTkw6CVNwsypCgK02Dy0seDfgx9ddQZN2aEdbPHP/
4gXBO9KmphhQEf0S8a9bENHE7Mqd1Za4wFxiK68W+Fcb8oihE3dNWMLYoBsM4DZ4wHgkzUcl89iu
xqunrLGCvJyqq44fF/Ue5tUOd7IpTuk6fT9Q3Gn+iQ/R8atYrY+qdPdmIBe1q6ceWuYA0otfeoph
inS3LWG1PBCrIrux+jOyISTJmjP+LWNVufhzKLRlrPHuz6T+oxYKNd5e5IOI/U93MRtf1plHw/I4
0X6Iionjag00vebmevElJNzdHObfPyiVcLouXhfur2R6gCE3DtS+sqHAJoLrMru9+YSP9/DJcDO6
qosOqIAG+7mWN4ZOWe4EeQ9+5q6wtbhCAzelVxDBywwC53FLv8Htoxq/qREJpHZsJyRebkCPyDrL
V5FYm3Aebg2JEnZkBZwHVRbdQgsovxRcOGJXqX23Y4eeErYpOYOq6sUnRSs3h4Qko49sZNTHyGmv
BEiW/qjwnKGGAaHq/KRVC6p7g1DvwFlXpG2g/N173LP0G2pYtT6Nqiag96ort3BMD+UMmJ+K3H9J
JVkoUX2+NdEgOOVqP+HG5+1MbmYdSomBd1tCV/b1TNZdtMCQTWIELcmfi66Y/peoqhpqju9kGCqd
lfs+YzVpF+jlpgggHH9bEQzHREisx3Hi2JTAugv7B/yaciVdLmbBuabQE3nsIiuvu91/hwY1/bKD
jEI9+uxJ55t8SowW2wxPM1cq1r1vp3DqjkMWLkxWV1wFlP9oXULPomNyOBe3pyrAuiKay4nu708Y
cY8jkEcDn14DpmOT1LixC8k+zoDOp3VeU19YEwa5cnu1UYXMLg5M/JO7UDR4GtUS2Jv2MpoRRT3t
BqiQufpPJjYe0ewv/xvxdUMZJjwviu1DljWiF8fzAB+fAdAb0z3zuk+pfr0/Z8Wc1hm2CzzlGDkn
b2zuP+fUnTXZ2vZapQHvkIYA5EAVj9jdQsKhJRH8jJgZrXgoiFgIFmCcepDeioW3ooMr+xi/WLXH
PtDmYO5zWcWPLv4XTPKCYT8Bly+4VqCgySb29fY+FY5L7uu1T6nlMPnl6wWzTauKOvDNfUCu/42Q
3P4hIgDbLMP3J/1Lj9XdYTomKL+cELJlWs7qqztvbZFNwh+1MfWe7eeRbkpkm/5y6VYO6lSwRNaA
Dbk/PByEZbaHOMRYxeErOqi2z8kaFGjDbClnihGqBmYjcrK3pOl23QRdOk8H4vLtGVMbNKQtnqQ2
ynBt0MUCZMGxpxAf32rxyj/8WWZkbhsoK2oYUI78yftDM0+A9hNyvOahT5ehwBKHiefmexkvkxF3
y8aGTwnbJFoIWbU3Wj+GelvIhX0bw7/XXcY5cMPFqh2El+/GkqlKJWlQ0lwCzNAkv/hLm8OEeDqp
dhKZpIRIXcgFrbz7Hn87hl2lLWQQThMH252NmUmxleM4JPLNovNpIpEs+xKLsNCLWjNxSbInwfzA
zXZrG9ZJafh3VWf3yli66EGIVuoVBuHe6AXdAHK0NQi7s0uAYP2Wb6/J583L3W4m0s7hBAJTWEsA
2b2A1ky0zr0MfY6S4M1WgzjwxTHInCgRHCw3htUirKS3QAenPIOWqSt4Fg1Qx1XQy9grynyPf0uA
9H8ZdP/js+vLKsDN2b+IfyDBXymRowQeQM1ldy0Nsl/hWDbh92QShakO8vt/uJDD6/pBYOo99qJC
Tmr36x8e3GXOJrYFklZezgV8nYvOkNHpR5wb7aZgzqO8VdSNgI5gcQ/YlmaJ9d/Jg9Yy2dmMKzir
wLFlGvjbE+kwUY6n2rngaqxfMvgH95js/qXHRpgrNkBecu/f8WVDOLI9xV3p/626M0w3YWEOd8SH
n5cq2PvOZ4QHAeBq/e0V9FpkCD/iVV/2zZauM246byjPMiZ0rgh1ciPrOccXmazEPnFny4Rbm6h+
oXvz7AA/3/vFChZacLOCzYXJI4JZ5ZZncRIA9ATysCWLeM1Cb92cAz54Fe4X0tfIG1IRmrMtYqRi
qnhu2aXgMJyWVihYpLHsBCrg+Pz7o6Tws/0d3ht2GEPASqhaQ8aQdogC4bIEsAkZnx73g+4NMLdC
4CZ6Mj8lNtEHLaARtamz32N0l4lHkcdnheVodIJOzvH6nQJJ1hwn372yWTR/OzeFvXouocNtp/e1
ZvNe5uR9GBCPO5BpDvSZb7NBwkBuyD2JHBSOq9qFj32wNk1t7X1oQa9OjAuYGsJSUM9UBDXt5bvp
NtYflNN+4Ec5hmOPw8C1/GCWRAE0nwye1UDSBMdTLyRDAd4Ij7cV35hsHa/T5E0w8YRO5oUsIUeT
KhZyN2XZf2fP12H0h1lJCaAv0nTNhf+82TGzi1/40hRVrworpJ9TA40JTLQX11pwABxdOH/oAvk4
o3J/wp8RJz4wEPKw7shuYhr6TjJO7FNcBPKSEXYRAdnXjGu+xlxAvGlTGf7mj6uFnFwkTsxoqSnK
hF3Kj+8d2tn49w27YpWp2llVWMAyKqHNsj/UF1I14X3eVz8Lakprvw2wfIQO6VeLhYfZyoqezHW6
U2T9PL6Pnyl97lm9x6rJYHSGfRFq1sK8ffIhFZUIjQw4AUK7vYzNn0Qb3nrrzznHv6iNPgptELP8
QryewIIWsq32y5qgyqikPe+BzZs551nQc5nO8G9njP6ByGbYfavPziLnRnovq35/NdBVyVrDYGIn
3+1kWJWZHSxFiWyIghekjygRk66j8EeIbuHevoswtS87x1h0/FzNfIkhEz3iRyYnJpZnqJiOVq8c
vs6nfww5KkpPSzPg//SPW15wsgrb1oPXEtEHK517i/umBtWbgKByMbMVHPPRaoZfUC66Bx52NAPo
KaQy9v55Q3VUK0n/98zFu4d1mTDOV8VagMs9eiJJbSheBK1z3+FYZwv+CzEN+b6nGTnnXrkpIsSk
5Z+mf7CrwBU1RYX6co+kIdBfyXe+pDOPydqeCoCJUo5Ny56a0LPAw877SyJ4L5ZVDaFVwrbqMFzi
4qsWzLNyxxtcs7raaq7pBJ6QycivuhrZ/ltp1WKDd3mfF0exRK+l2It9//OE5Ooqs+YiRrnt+nm7
TG6U7lIBQLFAXT0JqrJpVDydfd1e65tZFGMLm/wpZbHxtdzL/lND3N08LF99NsvsxyVXabx2sn6f
qDvJpkzYACP6BH+5d0a4RBfPLEZzCJPLmsWx0QYzdVFYIdpphG8QRyLTQAf/w4r1YbdDz2ER/41P
iw0SxhUwoB+/ZjrBFVvx7CrG84kxEYDrD8/oO8/CvvwOBn8ZHpLqeXbTOsBa8Fi3yISk6k+AxSD4
A/pIhGbIerCc+1+u10vhZEzIwk/Mng1MJwh7dqm6za6BkkPlCNDbAPNV9hmLfAWAna5RcrdXd4Uw
Q+TlqDV5V50XXK81qX5AVXkU10SIoVbygszzPM+ljJtZlrMz5BHx7Dulf/CJFZ+4EnjEzH7fYSAe
k+cH3tIRLS+eJR99oFc1gz9r6N1tHj1SkIJYuQAkbgrvC7+9NjiV/5TIfLpuFU/kActRMCC8hMNw
SywKtR96fIj7aHqCWrFjAhWOTIzw1Ky2rw3sS00HnDxMAVUymLljNjmCewpJc79/meWH7cO1sUGU
mDIcojjUhZgq7JusPOHiERfrPSmsJKDokZluvE66BfnHBCqo8TfcmAkUp2X6gtq2n2LHiP99ofv3
sTkY/OL7aKY47nDVkkWribcnUWdEKcmY+M6ATjvlMWfK5r/6RA97k81PJpZ0AEc61vrZXMoWsQcm
Ewh2IIs+WLriv8pFq+paOrPOOiY0dMubaVp5fs0EOFzoGkrbm5JsFYp81hJTOnFeunkkJ6aVuwGK
7OVSV5S/kbUTE485qvA5x4M+0QoGIDpF+tGUkMmMm4aQ+n6kgBQzx1ckkynUNl0SRuZBve75vnI8
qAXiR7h+p2Q8ptm794EDK8x2sCp78iMl58Ss3keY07QI3D2TNPejkNVDLHhm0IP5rZ9mFKuzJw7k
Mnx/V54wXlrcxEm45W+1snCGqjFbsqkef2LZu9qi+pkIy7o8w3CJKCzqGgoIXkgaSETBcax7RU28
3bE0R3ddHqr94XUGa22/HO2+fUDKOVUDBnucAqN2Y6dHfQ4R5sTIZO4Y4dO9AwX/ShgQ/0GWbva0
aZRyyHUTMjvTsYJLvV+MLGjmORZi1GdoIR7lsFufnN1U+WZlC3wjuKmGeQnC8i18D0s/Qg/PMN6O
0URr1kxvHoEPD77TizzCEgrwTCMfjzGuzDUsAa6EvmeZlWCfkg6S6fxNpuSEVCUBnopVPM64YfKT
uNtg1vwaign9kvpWPPzoJQOhfjTgjYUulidlUpsAxFJX3cY9eFbdZvn1caWQtnmpAKkK6BhcoOip
zq1ETxDis/c9hcxQXzaTX169MRq6Pc9Ed6w7DYEQvd0y3vhrCbfa/HRDea9cj51W6jwGKzoCRFPZ
24bJ/GsGqY+EeeExKeg/94Enfmkzi8tHxD53UaYLktBc0486G+VTiQSizqZcXVCmoUbhTrVI6hxz
pwEK4DmSexjihQyd4JKajclWrfbpE5pg2Fqj4KWMOBqDcWosVQlT9bVL3HY1N16nOoWVuEVajwWo
orFQoB+vnZs0f8jlj3iHxNlUwqjHeb0F1HOCsL0nqm5kf5qmnEBFa42JWcvbyHpgIMtJyuavYXk1
iULuDOduENKaUu9Dh/bfjwkBtrD2ovhWT7vbaAc7TerhI4z0Ob54kvqbG5AV5GpYsAg6UnWgYL2t
veZaLZ4A542jKybrcZ5wBd2ZyN9wHrHxxOdZ+X4Gy/8coiYPudR6MqwZqLgoYxhV55lJv6JKTeX4
gmQJUbHeJTPfm/CeTPp08euKKriTchmy9wqC4vcjPV0/fxbijLLcT/LFu524ErpswQ+1EVi3AT99
bQzpct6O1Jt+nY9d4/ajI83/Kx2eOUT/qdPzq317LlgIVyAPAVtBiGa+kP7Y2JPekDKvnyXvMXc2
JDhJlsHKV2ZZNfKY1NE10tJeTs0NPuq7T9G/f6QJnK50f72AsYJtSRRYHx3yBl29XLTa7alvpkHC
7ujYPiE8yOpzKnyYsB6AY4CuJdq1U7U74S4CtbVw/6IGhSKCOxjaq0NmId49IZSd5f1+ulswdyk9
vLurnzW7ErXeBgflCyz03fODi+Nuqtg0f+pBvkd5cJ62Xu2t8udyknrPtIdzWhtu5xHe0kzKDWBJ
qGqFWMEvUclRQRX1Hh0wj1YR9ZqAJlhsv/K+dE3spQlyQ7X+wFSOyBtEfq6vRDEQYIzJq3XUUPly
YKwr2WMApv5bqRxBf/DDQYdbbHC77HOCblyvDAkzIZnVPlRPNr6Dz6UkI321rjrWuogc1/wSscgP
4xhMCxkXeQ0D3dAhJbNoP1O1mumfcumUK3r8DzXoPUJHoobWhhmaXVLDjVwDabWcrcfsRY7diDA/
Wf4PUwBH+V8wsTLbs5eEsnV7ghPVjcEmDbIxiDrJMeMKSeokc2QAOF8DNHkTbMfB/XYAri++Glkg
W7e35x3sh2tSKvjyUNCnvn2UH3/j3q/ZRKxkdeLdaSJFN1hF8SKp2duhYS4m7+FDltUAlqvpct07
3p9A/zVXHlyK9+lUQsup8gG0aDVLXzfWItWCnYNnDzRzjvdY0t+1JKu1z859V4NUmG1imivjfWUG
pQdyGKu0D727kOxMacocRsYPOGTn7PmFPq37MP1WTteBWQyq3HXWARq3tiZscQwG2/3319X6AP/y
zkZvrxnPm8cRPwyYtlHUCxFRR+wX8sGakCZy2Ek3XXH42vEmUVWzbObnboPZmZZzdQaA4HvKtzau
eP/s3wcxuXDWvoUeMca4wuWAsWw3lEMgPqDwYxuaZoKOwMsi7//IMSoeWs+U+lMVFV6Mk2IIl5V9
4pPrjcvO/5hv4ooPURptTwgbMpM9Bou6AhRR9wE8hW9EL2NhDz9yj+D8aYRu7wCMbJXd7dzZ9a6y
ZiMoSspemLV2qBmfoj/c1iluN9KNIrJ2fKC3kl2WB6xjttvTXl9A01hHVnrxF5BSTSgklGEATfLT
opHo6M+8Vd/uUCZbzuGcyWz5fXsbs5ZHlYHfbiRsw7CSLF+trnRMzYiUSW2MY2rqtMxZo8KuR3nm
fVqmVpMBZw/shIZ57/hAn8TSf/CMByLX+x35C9NLWO5EJQ+sufI9QvEkj+NOYfTNHcJ5vkYsWc2t
V2g5Gh5HAqUab04MRT5DrnqIKMJLsb8HcvlSx+T740sxuo2s7Ote8e79Lsciylkcj8+OLrsoM8qg
7UdXyTBLBcDqK5tKvmVQTL/q3GvkNb7tkovgim/+7FRP6Kof1lCqpRNUCA/Cb5Dy/25GLj+CaQri
tQKxrvTLJTsxOMAeMfcWBNcoYIbeJFHBqRzly6X+d4MIom+pSNbZlLFDeDw3OnKocMGbOA83TY6J
wBxu++n8o9iubDjME1x/RRO8P1mNRF4GSvcYIQ78UV83+0wL8YQnHmtHySrjBMl5fTOY+33CH4oN
fufq5ct9AQKCnkvJr6L51lEysLZwhBEIoQ3HUShiNsNpDWSFqc6zGMTiBxraWGj02afcSY7YSH/3
pJDp32jeSzlCokiyRe3PrN4o9xGbnwE4WXv1PvQ2p9niYACJUjG5415oQ6GmQx++1lze19qNGtC5
bxov8JACcQ1c9Wz2DSzJ6oD/InLWGVQdkU9o9DhZcv4nMPb1RdA5s6ZU1o+8KHxrBaLB7eIWCBi9
AgZTgCN9ByaA3z+0vcJYE2JmgsqTsHQo9bMEUu7JD+KPuw2ewUq+Rw/dUdQlEHKpLmRf8D64It3u
H4Lo/8dB5DRP2DKbbBYKHXz2lLHDmigFgORnECkjUehs4Fo/81rjW82ycgmf2YAZHTFnwLqcCz6e
IApzAcMPsIq17a4D15svGZjvRXsVInRZ7/5JiYMo6+E1H3iZElvqYg6ziGwamN/5k5R1bbt2/8TF
4kP6bT7FT2aJD6j5bhzdqz+2np6HPWG0qtwGJMwvhaZzNBsYWz0VnVJhZ3on8MQisLMedrD1QsDq
h1UXhYFKIzKGrHu8S0IVK/EmoIVz24WlG9IDbOvJpnytwB8ld8VsJw29He3/903Kl/oypxDlWI0A
DBl9/M2TuThwb7SSQDLTdOTzq4HAgooOGRIPGaic7uFpD+JpyaYOamnl7fd4ROvTg6wUexeOzYJc
qKlL7jcREo4Df6RdPQhwlxsd/R2XkZfZCwzKkouwcLKCkQqoha0xrtUmhHtEAvoPnMXc1NC+Q3WT
XiTiQBSVAELiAYY/cAlrxH1OG7arymwm20//lS50A86Txn/+176kH77l4887VFFFBEvL9I1Pnz4D
bR+3k8FGRj2QF20YuyNaumNdLocCj4LQkIxmhgVcFN0iC+C+fLVEuR6JJQrZ8ATK8MqjWjbMLpac
YXrhrJ2NguT6lh3Wqbtn6j0xA/fK9difzTwgL5H+xfUbJpasDuBJR1Dkdp0E59ky6UN9FyAd8CjV
6f+BChcKRu7xXtIyVMItzbwpnHSoY16iSfrjbc7R3TEjlr00AxqDtcFIsUYF5DqsAsmQhZzwzowu
zMvcWhkRMN5JNVN5rFyJp0Qj9QESaZSPIDSk5hymd6tJBUFdID5X07q7AyLJ3HIQ48DCFj2nUH+H
/jRaIblP8kNj5DnEh25FpVt3X1s5N/lgHPMha8noWLjOOoeCf9LTbfGIj0ZL9m1rr6pyudaJ5HvC
injR1Dnnt/qewB3oZJcjfbr/YwEXgooZLH+/CSvI9JrnCzLN7kZGpsWpmwewnGkYDlltkVpZIaQH
tmiBTlq9eXIIg9ycoKrxt52SmVmdpXBwJKrSQtgsPyCc7ju0Ha6cxEEcUs8h/RYEmyzl/38xnw+U
2R0qDTgJC+etXLFpuvy+1ymCKKsQyzx7ujVhByBmLTxOLa8Dorg0zEoxDbp5o8kWmQrwTfpPHBXi
4ScXb+GMN0dcmY5KCyDclPSKQuJs/PUZAVDZEhggJ4xnmwDHb8Y7Is63GNJ5mBprLbwkh8ZDmEZc
8jJgLL5lckeSbBIcSTbDnYsmTR0kHstXxub7Wo1gJ85wuqbC8CFLSLFqfO2cI+0xVWaft6154ZUX
Gs3M2OkWTgXaenSFORQqr4zxpNlm0KI7wIkFqaae67obZCh0VxCh6pKD9f8z3/TnNeH0IJ7lHl+8
oeBMp1MLY1GYxyCF3ykT9O815b+hW+f7C6dF8IZlxVfQ8lb5oZNrBXrrouhXofP+HfEbqJEITLPi
YsEOIqRGizn5XX0nqWlvYB2y9+vjC1U8NuF1duUttnWzr3KAW8BQ8U/oDcfzWPPOAekA6+hnDS29
i1VKLqMvAaSMdlOQxprSbIqdH3b7A6A76w8iXXMcUo6gGFpYRVU0y6pgaqFg40ZSNAKLHuS9uOaH
/TxUOFbfvXl8uP81xC+Hz5F6UMyMd1SvsiyfqXYtpFytybasAcD5MQ/+daj/HDyod2wUfvOz67aU
rbM5HvFnT59fwM2FPxdVWADc6TFy6qG49F4AJ2bciTzFoLENsH7U7z9cXefCUCakpp6xyeBUacZ7
hqTfCpvGs2BC55dcRdmbMEGu4ndD7yuEt4BLvj7kylvTKLYLvxG2dFEwMZassD5KO/06wrRgFPay
8zMoo96BPh4Q9zek7I1bFmgFEVVnuAiZeH/uCOVOjDJDwhlz2pcFF6NEFwrj7FF5LqbE6d8Ee2nt
kh0ymspkcwo3IqqNrRDWGSUBlq04mFJqmQXuxuQYdmp3DDszW6wFEuQEC20t2YlVELf/pEhTWtrL
E0JaMSFcJsqavxZTCZ6k/GlChcQZweGIqX10Uch2aYrmq6+8eWELwBE4LLUa1xJWtL8XOkeJH73o
XtAqCT+0Wrb7G2XzaAt89UE01iyeDgJ9EfwK5CbJ0eWiRpd7CXXU88dRudbjPKZopL7jnNz4uCkS
Ws4o/06dpfG/1XBU4bYnFp2w843s+utIam7HsvEHZyM0Ot8goiIIWpvbd1mNWR7cRveyBQaFw8Db
GoZHOQWhBjjOXyWIabfYUMFNvGy/s231fCPhg9nxxP7pDDqV8MSstaUJng3/T795alvdFHaEWwow
LYifw0cwXoXPQ6ZcRVOjxtWBOyWxFi5YvLnYC1nI89j4CzZct/GMid1TUNg2t9k5+OjT/KhzWSM0
tXgpu/B0FRrhrcwqATQ4hjryg0we9Q8zB4dSIOyF5Q4bbQmMk59n7w6ZL+o95/++kjDk+nXKgJCe
h53WlEXkvyy+e7iVXU/UY3GaQ4PwqHP4BS/AJkrPR1nJRc6t8YipdkP5EoJm1anZGdhJeJsUsO5+
STa7m9mwSbW5CGIUn/XzwIWZZVKnhTrQIFWj6eVV7Ox6V54a3PdtueyqXB1OYVse5o3UITjeIbTg
1Cqg9KcU+9c4nanpkAI9XxuKJa4xw6N44toTxM2uiVbtvMtgvu7AUiE2+cvTFzufOyPSaDQjB4dy
oSazJrQoxTrrRzS6YekaoRpJ1kGdoq0QjKWzfM+iKuCK0tQseSZMWW6Gj1unfOOEYMQvv5F1zZE5
9VpGNI81EysMuyBrn4eWKX+aezR6epTb4OpdUHg4ROMrE/6B5TGoJf5spZ/gsbWhITQvPlFN7B5P
/wMFbFny8JOSMRL7ka714F9tn7cpYrEAG+k2atAT+XVWiXOKcHyeVC5uYUmOdNFnUDNDt1NPyIb/
tTCzhHoRJZPzqW6SpMZj/YE6c79vG4pO2e9NBMkldjBIAW7WLmevevV4oRajhjTnzbNI9cymNver
P1SR1AcOJC45P5hllfD8V/wys7yfV/mlK2ud5OqmlAd5Rz7MPuIRTqSYxj2YctxuGjz3adABEM6b
msZXABkXumVoZkAiEaxcVp6YebvLG0774oksnvfvZI2R95xNlWL9UUod4gNcyQ6BB2G7T65spVA7
KQKHuAk3VCmieRHIRwqAO7vWVjVd8PQKtnFN4ahArPjp3VU/p9vW2of/s1623jjd+am4+1hHZu1e
B8p97XuL3Xf5/xkb8RY/lD+zWxbxnH85rOsb9QyyEN05RaVd6sCSPQTFZOLvI+LxB+4wwnzDUXgG
7xyjYM7POHAZIhLqa+7FJPxqu6t6e6oodN7nDGAyLMCXibWnjacuRMekS6nGgKds24uBmvEGTLL8
ELKFCJnOaPfRXxVjSCk0fjKwTZUhSIYs7Xo/r7S0UuG19a8ZRAnJx+cEjtKbFhuIVRuTMvreknN3
fuZC9RuKLH0LsKDaFRQyGQXVOyOwK1zG1LBNo6Z7GMDDI4fqb87+HpzN2aY2mZPZxRs53iYIwsjl
8VcZqt3opJRI7OF9GXq4cJJ5DzdswAq1m5Gi3H0dBlWOKGmlrz36g8DMybmkjp1oRNSKIkSdfFVL
LG1PT+tOzg5pnUh3mO2RP74vhdeg+6OL5e0+jCLG6xZmHm0LhvtZ/Lh5Z66iVxWgCXQ/r0HBCeam
4dCAcBQudGlE2w0/K4S77uRc26WXeJBwx7szzRr+7Ly2Xx6ce7Gj0ngvTkV76MS/shXFMDXiY9WX
j3ys/H7yWvyP5O1E/v0zPdmcWcP0dZJdEdvoh25nuSw+6jbi1HTAbqqVz6KvJcdOSiHx+9F0f7p4
OPwRHrpwMlBM+UHqG4nJ0NikT1RtEicrblYWUDGv0J8VjhXXIZNhWyk2pT1FmS7oscXkziAeeetf
h84NJKMf+kyZBlVfOKBgoSnntbg83dEa7TyWMjoRed0D+MOZMntKurR0pqEwbgY7xQ0yy0N3Nq/r
949Xdvc3ccshTZ+a2FWqpTI+8S+qf6s90qZUmzf8Qb4C/rgfNBeg+pqJrBtzycJX/x8sks8Vd+ci
BWF1TcCo2M9cjD+hgpmVA5dtCd+tcdB2DvqMS58ua5tMTJhhO2zV55srLHQBx9fwovjF8rTnQ14S
cG2BJj3jn3ucFD6pLaY7L9/7jAY20tYcV8s3M/fBBERRywz2BiPu1+EDSSX4QGHTIq9EopS1y6YB
Et3b2v5Ft9QZU2meAfj6NjcPDzpEDNVokNay/RQCKE2vWlNYQc++ptX2kPFFUcsvq3cYvMYJ9w12
yllXi4SqesUlbppG6dGACcUiv4z5Bmm4qd2KxGT45pPGDIK8mJo3wLduPDEqjCaDoa4uwY170fAE
YUzlONdW9FpiMbbA1AzVbF7D8laGc7l56MunJIQLa1GbcoCKpHcxyWHdYygb1Rsh+IEsezCmf4hZ
k48hUMBIv0Mfm1jVky6GmGzewNfzGOFy5ztDGn1stIC/Tt7orvkpe0PZQXcD7ZuQcZ4e9KTbPuUh
G++edUVS5UULlPKX758+M33mp08DBJeBWxiDdWzusaEK84aQOgzQM6EwEC5LfyPjPGlrWy2SHsNF
lVqExiZh37sRPKOFo8eqF65G3/W2mTq8EIxv4IzDNY/TPhxBAy+DTmz3RQhCJZ0t9pdrYoGz1yul
F/QxrvtSQTMV08cd+tmDytZZUFq++npPnSjvx3eBl04iEgEFHKS1y/+SVdav+3ddamrbaPYimCl3
dtBcJHTjvncVTCnQqIC5BuH4V1AwBlACfdr2iLTc35PCeRKv1WXgWMjXDRKu6j5PNc6+t7CIdt1g
21mIeOpevBTM5q7XsCOk1imGJbcUHqXe4Lg2sSQmlJQ4C/uwwLeyvZyXqREIJIWhKeI64m355Bca
CjIJTzIg6Uzc79If9NnHri4PBXuJD0yXSpb9dii5YLY00ItmbC198bLKy3+dlanMawibYzmxvX/w
Cp5r07d0b/mpMB0XBrrcxsebwkErr48JTbKnnnEjF9TmOFBrFNIYTZb4S6M+lm36HUzb8RMSxCOD
X8Subi2G7CUPn70klGI96lZx5YynRZ8ZQUpndi9GYYIudikBZwcwzCTI/c5f0XyY/oqUOstRKbmx
Ri+9z8GoNQguYJE9JaRGiyVkBu8TmUT0Z7yW8omvEsyX7GM2ZsiG1sTJgdnPc6oB41p7uIEY+Q3B
REoa7VcaJ76/NcNHT0qhYIPHgkMoscGqG9XrCJbCN9CFDfE5PrVJqWzJmmanGvCEtFs9DCJKVnVm
15zySwXbMVCia4lA3ZK19NxJsSKKKysinsX6vyAms9jQR45H2FxhaEzyl9Vg3C5q8d2CCZAq2ajE
503u67mcBprJ8dEkK97F4k5xRFe4xo8Esn1lKmHXqHw9gTxJ6I/2H1sb8NhIlpUqGM1yENOk3u4Q
MTTn5bpICugv1pCvVQLp3SDO63qY5KnU/4er4Bjyn7cA7J8a6TlMkZ+x037DtkBAz0GhI5XJduG9
RlCyoxDLcD1D4suf/NYQjmOjQIz+g/0cxWKiVfltFqRNqkmUXPvoBsl80h74WVwwJDVlM+58+Ytz
0McNd/U5ogqTUqa6pmSTpcrCFJmSmypsiecrAZ/1IazSJV9ooVqqaRvESILE2w20ZNS5uJCbbZTF
vcjkn1TO8Y8VnOUAWy7TwxP3ZYeouA3YKPU6LAZTCIT+nVY+ctN0rM2qIdPl4fyibIj5mwF6L2yE
3nRV2LQK4kgr+lS5VVp9GrjSTV4R1JF486rigBI87xt6ShPRDKsr9GWiJfFTV/6UmxUq2mTHTXbF
5B4Bnv1vGh7tV5+JN+n/xpYB64l0Owx3Y8cuEoeMLZ1Yd4IG+SDHSSCgEruu9zqSLMjnhHj0fgfP
bj34qJpPAX8YKa7UHdxQwcsUnHUbWdiLyeDpB5PrS2qXAFBH3qcSkX4D9lf/zUM8gCtsjbNRv3UC
0GaEJDuaqlIYse8a0+Z+//OiNEa+ZfI/X7k727a1Al9vNK/pPvOnwpntPs7UnVDKVGRQzV9YPdff
bcHQwKWgJlt72/DF89f7cIRkSZIz3hiCC29skTdqOsrHTUXuLWz9RoSe/6Z5t1DHmal0GySxyebz
hdsMI1GpYIcnH6Z9crgcJIts8ayHXAzy3jlW2u/NTNtSzxIUINR3ropZyaNE0vAeP1aVj0tmwHVW
yWiPmygYPJj5qqI4nh7RD/ujGqlPQvNf4o/M5/lJbjGUvtTccFR5PDkl6qMURBAuBQLNXlFkf53p
t6Gh/W1sBL+oAzbcs2J5cBJtPqs9INaur2iQ9yqTvdDeK8ghOn5j1efn0zIW9dvhf1/UoVnvDO/c
CO/PcHxTR8IODTO2XfhMAUL+TbT7pseXVtGds7ZC1Fyj6+k9uBO6E0dGn8GzmVebFkJO5Tg1Q33b
l3WKxSCSX3W1r+SJ97Zy1ISA1zuftdMohl00HAbVKHIrhZFFRz+Sxxh5Igw/8aOQOFxLhdWCbu/Y
D3tjB5IlTuhy3zC4Ud1hPhzV0Ww/m3Fyp87VpmD+4OSOBVJeBs894xuWHF/iuDu3jcvoYC2GUYz8
7F3Y33olWWcmnn0qgqOOfbaG57cj1U20mN08oV0wRQ0++YmgzOzQ74DkwXIOL30SnL9Yu7VfAJ4f
S6MSRiVYPpADC2MOjmpPleHfofowcXCxoH2FU4pow+psAkFMSGwdwMmugkgHw6B1A8FbBB5Rfd1U
r8xdCBEPvTLEhItUm88GxDAppH64afmW/1gnfmGKxeSvznnkyC7mDe+iU1X+r1TPH2D2h+n/dx0B
+CaWCKHtZ6Ziz/8TQXmlz/zywUX+QWoijtaA1Z/exCeLgwhCuaoybybXJzha9zUEXxfmUw4UembL
cF1E66ZXNRXRPUM8BQV/YauRhKbri7ovwnFB5pyjlUFAqINUPdReogNNqjBEJY05F/nZ72N9DHYQ
gSUdlMMQHZwyQYumYyJ/R2JUdQwm+ycDpbqSTcki7c7H9iLN3bjVutmpn9rJSSWt+Vcm9UDvDeKM
/R1uHl98CPaOoa01oBsqMA8LXjH6/KFxxJzNhyNi0Q4cewkdpTEEQ26vmPaBbz2xFP8TlC0MPRHJ
7MAqf8Xv6t7VQxHVhen360no+P1mK9S7P/pLZOiJQpTAqmWft0Ig9oPrUyH4z/DwCAl0ZfeXrDwE
hQdTlGDjhNKi8YjjGgg1a71h9iyrZLCYUVJ2OsoCrGPjP20mj9TOPQqOa+99s1VIN9vaqqKD3Q0K
B3IlV1lc1nheDLwJgAWap2Vuu5WYhoqzt+RBzSM4tUAil9LI1kbfVlGtlgSNJ6t1cDVDpbn1022e
aVoSqOYgTmsGs+9kHIASXcRlO2M7GUKmdvpuR2iIYcFTrRg8DHaDEW49h1bfNLyjhAwnRBTbEc03
YhKhkWvh4ks/VSM6ZIiThUVUqSt/J5kKKr+doSNx41RSmK7ne4os68i5QRJwefYTbgQn/eMqEMyf
ZXLonILk31pN7vGpyUExfLew5cbz3cH3LbljFZH5Kg8+nVs/RhwVRwZmFqSGE1Z8vDhh3PI8RVaR
ljwR4bq1/AEW/F8AXTlUN5wVbV23R7TVWAx6vzzPKgItnqMSbhQ7sJRtfnTt21k8C9CCxSRxsq7s
bs5dfllWKxjVIjz2dWisw0yFwI6npsrHQ9rdLOeixFKKgnalbiq0eY9VISf37KBlTCecnJobdf2I
VcF79Kqbb8rpZCNxuXPqig945f+WDpMzRsMRHEdxb1VovFeQin+a/B2iLSGvF7RSUbDALyTE662V
omwq84ug1tREr5FNF4b6ZH6x36a5oZQtDqyO/wyZMlGxVCH5Pmhic3BqyFLqSDHzjWgEgnjYaPiV
o2fcUNXEhWYU6mMNC3Rjq8YpwTSCNzlpiK7k5jhfdtjuXcFJwBHbWITBrphEZv64UfDwEvk1n3mS
vDLrTcQX/eY9c8cR6zOSq6LSU4OJpSGOydELkEiR1Jd0ovD4pkxPcgwA70f7xE0tcPE4z1QV0Yrm
D1pCQ8xjkGEwcBews1EaZ+HcA0Tq91Jh1xcaQDlGHFD0FlefmLz5k2J6cGJNH+CNWFd7gPTLh1De
o0iOCkINPdP5AMPQwMJZaIuLhzSH46vLzIo6lQvPBBCgeoJerV1ZnMWn80F+GAY+pEPVl9sc55D2
CX1YgzgBZOu/rBuZmQQNBfifcw1INmpamhNd7KAriwrjEEWyhP4W6/rGzrUxB0ZRkQNArVmfB4YF
p58qTgXSgkFsypNFH2IeIY0fxd2Sf+vgjytBAv7VKmfzkwnqDvxQPBZ75lCKQHcREUspS0CMw+Ce
uishBqbp2ca7ZvGwsKRChnZ1lKMK6DF12MWfkuYcUC79O6H6zkIcWoKWkUlBDJEE2BqtkW0FdRcM
BjgTlr4jWwv2ZkXABGgWpZaTZmWEg9GJwRv0lh6q2YthFIdmk200dyLZ2wd7DYrU0YrZm5JLM0hX
6f40XOfwTy5T8kwT/zLwqcKKfS4K7G660zYkQ7f8QeNLi/F/FqG2r2YUH/lCuylAfX99EZVDKTZE
XGhIckN7WwGvReSzayyKZnXSl1C/IltpHVNo2GxpYfRXL2KMXqUVbaroF9SLpHOIxDlJLC+jiF00
+vbGqCism/tlrRm4GgpU23Vd7Kg8LTTGdfs593dk64urHTf0k1agiFOeqxqEfbnz6zAbGZFlCNIY
ijYkBUIXvwloNNLBUDq+XyBxWRA2eMsNgWbxI7eJtn6ct7f1MD9ZOtmIppK4wukVj/fPbUOPX4Cm
n0XcQsdhefJ5mzGsWVqIJqwdUU7ZkgRjZd8si65kLCuAq/o1EjlzZLNFI9NzGPmcW2hZRdT5YoCo
S0g3n/m8L/RtR99aWuJHu/SmhbIykXWL5srDU/sg9kVZOK90sEYqgyYwaPJ14gmqV4/QoZ1A4vho
8+DRR/SWvdD7L7mVKbSIHV+gvFbdBgQZ8PmFnfMESW/OwaAMp1W29YfI8DjOnD/YRsDS2ZaKJKP0
Yif9xJaBBcNoMj7UBZ4B0looVZVhIcIeY4i+WfqySncFo/SmdBN9PC4GKJAX8J3uSNUn87u9/+VV
HUfnNKup1JWNzpbIP2e38tQjUGJBALBtjT+9Frfh0OPj8gnktZYTHB5wG3APfxNaWqFV4EwHoDmd
V+9WKi7l4MQb75p0NV8eG52hO2rc66PC+CgRkpr0xddQDH/5nWCBH6OF1XHJk1LB1WQLlhNKVuvF
LE4GBxjBQh7xnZz+dXGvEofcAC5oMjmDGsnElU0K5+t2HwD4HTsKUCMtJaHmUbKq/3+Dlpz6glO2
NlNEOhm96IAzPlzQNnruwAg/IbmcuFBQUOeti17t4u2vSjLZfjC0jzWYOlBvQ/B16JqzuRLxBX5j
g3xPxjRub7/pDcbXXReyL3V8PXT4p1p9FGoiMGZ0pulv7gf8yC2kCOkz+0zvkR5IGRT6UjZmkkXK
JJzrC4IyiYSZ9UhbxQUmh+epPCqjlAs5+SkqYTROk2jZFxfpGYCjGwwun36l049lyzBgDBdk4gRk
lcBHIn/j7J4uVhqRDJKF0/IQ0eeuf3/YK3yHMvdP6LYJ77/rofQwjPbGsSNaD7t5oMuhVvczUXCu
R9BGWUmAwEGXMS2xy3uXWRYHhTFrAFbQ2iL7Zo4bR93HLQgz8h4WQaI3rWw2oUVBjDahSltskbCQ
ZkYlV//ZDGWtu8W77Ppbr7c57ZjiZUNAKM5K71GIjLPCmrRPt5ZGFWKi6SJXf3iYcnBs7Ndc7ORZ
E4n9owguHk+zATFgJwRhqsNPU8FNALFY/PZ7WlWSiagnkhjqVm8ThAcsTeo2ERS/sRn/rbBdDusH
Eec58m9Q/VldPgHl6WhHSMddL9Z7wOd9Rem3+Tnnm6oo54tYfZBOelLFzVjg88+qFuGp4InORHvE
rehOXkZVgJq9FQWgXoP1j3jdjPn7NqmCb660aGTpyi1koPn7GSElOG2xvWKt5Q2m79rv3IOkvLB7
onk0rK5PAUlGzMDEK/JMKdAUUgxs7z4URwESnn/lKmE4I1PlGfD65ugttsOUoafMnXO6vZyOPA8c
XNudmxfdgLaqfI9sLyat7cfPLPm02Qy/pIQO5r1mI6DYLl1VbMXT0eALhn4OR0gOdDzpWcbGHtPR
35dykvV5cPCrBBIEiBWEIktP7lrJevQGGYC6z4nnWQDvJ0Qvxi4ppxykEPotfehgpfAYNf6Zzs7x
/cJdIlc4iG2Om/1ChPq/PSNdp2RMMXc/q0Kbx6pkvVzK3xdrn7hUPf4UnMLPLjScRVAeB9GwZiYI
DaT5mH4S3xkhQKIG2E47Dj+VSbYSIkBp3pA4So9lt1mxUdBSQJsLF41pDLI+cT0Bg90sIPP4IoEb
ui2dFKUSEZ2ELvbA1eQkdMQiA17ZR2XkbdEkEYmBdTJLGvOQRqGzd3I0ZY9VVjRqKKQqFOSSAnEE
uGXgj6GynHvn01U3vL+JEL7x0Y70pUPAY+vnhWGGqz9Km2K3FILhMz7+yPixTWiXgkbe9tvfA28T
rV1JzuOZs5nUB6R7TbE4kcyPv7gp+R9EEfzBJ6EV2Bu1CHp0Ytyavqc+zGMTD/OLfOlG1TLPcjIU
X/sM7+6nIc663MTLIgDtebaQkYjWv3Gc3A7eak47ekk+X+FvRNO0e1IUpCDe96LeirpjY0FoKG+G
c3qt9+KNv/tRPbeKNWJwhxrL6IKYyUNCTjDazRm4Yh4feqqGSwzJF1Wqn4FDeU24LNZZ/TGm8bMc
/YTnp/8FaH9uOdho0MyEXcWnLz58OgGtBsgNxRUQksosLMe0wKXYeYPoXhibPmShftwXigZVvuzK
6SiJpoT9oMxL/RSl5tXp+x7RJIQTMCGHTj4HDU96RS3pP4bqFvzH97WpS3zn+pnkcWEByv40guHS
P5ZO6Jh/j0bw5E5AMipk4ClauduMoQt64xWrr5KXQ8GYm9mor/ij/mQyQ6U1nhMvFuvd0+NpyC1D
ogggWn0fh9HBD2QnEujBbmUk1f9RQu+3NmmdRAiqSw9RMVi5dylwwhRnq1+wI+LlxS2mXLnJv354
JUDeLqYOW//MMOvRM1CLTL2mtE2TxxJyVWt2kf9OAnyT3BQjWK/k5N9Kekojz+lVQmgF5q2oBh9P
yhndpyWNjnmrdMMyqVA78lrttg/oWtsKmQUg5YxvSnUyXoDHVbJaB2nxjLZ7Z5fctGEHRfKMF+r4
mfezoIivNsJ9b003ZR828iLEqutuqz8nbpi+XOxtTrpDvX1ZfRHd5r8ljaKROJH54CDKuTVoUf7O
FLQn0NKQuVQJ2IdgpCyn1XZjOAfaTuA6W3zdfeG+Rnte6gFobLA8QPUvkPCJLTENKw5Q6JS8kxUb
+Dr43UKk/Xoa2mLc4cka3WoN+zWyhGyIzJO+EixSu1sprlZHmr0zBxjjJPwz+8FzoCP0HfJV53Le
O5SADDf6GqTlySO5i4/ElN9MrUS0srgH31/uZKm2sAjYtLyLKGtBqNOUqzraQZcSfcLxb+Yhce4r
I6Q9xJzB9fYKilpt59y3QoA9yuvMliWXpS9RbOxNAHK6Ccd8a2Ew/jvjAl1Fwr2ehqQugQ2lFnNX
U1m3Qb0gmChZJoCK3eZNZUuxwIP2/w5ZwRRnzW08kKBbIt/knBR9lhoF18mXcUHqH2XcYtOcowqr
NDPZLETv017TIOsc+dr4SwOVAJbWHHPOuxhNoH5IFGrqnxn0NohemzN6cO1hIv6GYQj+xGOasJYR
KFPuFrlnPa2CG3Y4/Hbo2Q3CwEffAwwoiDhRFort4cW8UktqoYsufCWN6MQng57seVLnID+JzMOm
XkW980jBrS0llo8oCVqTVzPdTEHhu+dot45kNum7ty7SDsn0PjsZWFnQy21bGiqV3MdsnWaLkDBS
zKOHU1yb42Lad5odYHcKC4CrTfx85mmAooVwBzPau0myjEDqqrkeK4fJQzAListCJJ1tZvR3Sj4w
D20Rr+GMaAAM324X5/o4EwGV5TdPZCrjj7TYWY5fys1jFv/ChAsREJ/86tdJEv0oNMf3dg+i5VRK
ZwxqAarhJGBLEl7ytvq2w1xarHHSkBQ4MUycC2f9KyWjx7gERus3LyRm0iXxINcDMf2raoaR0KKd
dH/YlT4KAkDubs9G4EOUcw1t/Cq4jrosALbEVTduNRnbXIMqTvHcufeKVrWFcy/DGWbYICH0TRQO
CS4k9mr4OF8W7eYV872OiHbF5/ZVoNlGD384RtDNRrDnBcNYmwXs7wP2Ftej5oKAy+6NdGaub9r6
aiZA/XzpYZSa9gnH6rTEfytRWwPi5MVm5xq7FfiEMhuYZsaLG9EtBRsNEcoWwRFC8CRrhIwAwUVY
e5hZ84YA+d/N6ws72DN8/B0qXbnW3vzv/oNqxxUoEIGqW8SviLiEG9mCtExQAZQluL97ZpbQffx2
ZgV/53xlsQgB6mGrUg0UljX2OOpFnGfl+HeHDhLP94RDWR/oYG08zmDNF1UBrjlNcA4kX0kO1C7K
cg9i1dqrrVrFYb2r8YefjDdPzH8vcJlW0NJOQANSN9902r2H8hTSrQXpuEMBruZJYvHUnka1NSyE
bnaVTxQi5Juiy2VzO0qcGOmcNn+PJa5rfKRXNc5Ua2p9Rz3wdFxnqkMkuaB3du/0W3+38Sgb2b42
mfUBWhRmGQx8cMG1HtY0da3dbLPoS27WRBLotIKPJlEV5t084dvyKUttO+tLulACE9U6Bowin6C/
ktMVUT7bOQ5q00QWK6CTJDoq7ZQ1EbgzZVVKxsf2E5yaUlqxndJCi6io7xpsr2ocDk4qxjaRAF1F
NBwq6aaH7RUK1x2OQm+Ah1Pfj1KZ8Ts38Yu+hh/GPtYzTlW/LlBuA/DNDTBq8PkX7pLEm+J24gTB
4OQNUI/YXbwVntmL8z1nZhfTUN08g5uwK5trGQfP9K9PSrrGLJXUe/vCj7c8KeRfkU1m40icXi8F
RM/CPQuy7oGET4PcHdZI08KScJ9HdNjPVHA9uvBM2fOoj6eb6AdKFNF04RdeWXYXXRbeAgFkVTa3
NCnDWomTp53X2ZJSlkUb9PpasH4eQAh5hqt4f3l0hs1B31YyiWg0tZrtw/pnZd0bOalSSPmHs6MT
xu91Y55ytj4jVQ0StrI5icvSGiVZuJIpnDTJQbxxrONLcCLk4aPSOgA347A7ZuAbnlgF5msYszLL
i2Ehlbpo/iu4OamtBzA+pgr33OqjgvpjsMOfNURhZWBO0Zat4fa9Bzw9AbHGG0Bi5/ynZF4esqGc
rYWHqpQec7NyV0NhqxXsXuPSxfmpwweXG0V3bI/Kk7tWpEH8HHIchU5NojFmizo1Teyd//5/kDyX
am3vG5LkZ42yjj1cV2IxXpqWjSMejr1yuV4NzSzy/CVq5H3qZVMEjD18t6BKAV9MMFWd0xOyKuaV
j8YurJjTl/13nyRiS8JmPR5UazwG1PFlzMlS1CmO/ifEeHlrxtVkFTjq6carpIl48DBUz4X40MTa
yj8ep9N+FgbN6ZxBIbvUPZ0/1rKCiIExXOlVx6pxDGzo3dx0Uyv0GrHgi7qqFp/bFjntp0wzi+2O
McsbQtMvc5kR9a6HqTNR4w68tIEkLTqwKZC/HNyurk6SuAxpQ6Az8f3EioL6V7ecxiIIC4YbcSOU
GjfGLmVeOJ8vnCDx09HJryIeuyajKVKUjMMdOUVdn2BdS9btKCSLttSBIIr+J3oaOfXZ54mMvAQc
XXe1BmORmbmMgQVa6eM1IU7sedmafGjJtb/kVushTa9e17DrWUntOdiwZlwOzT/NaFH8SSoddJpl
TP9koTSoP2gg3S9N2W8McpyCq4Q1OSicSp6PC0qxk7iNUUchCCRepBW8+mfsvJJLGjJw0ll4CXyd
5ARDYy/pAmJMj/dO2tc/Cr+F12Q9VYdTEzYDihcIPT0D8zcwTyropsem2SgQDPzuf/SgKgFa0n2q
Xv4jiW23LhD4czdPeqfSDZYE59ts/4MzFD/dka3CJQD+ti2s/Yxe1NcSB0SCzL1oGBaP7NFVaedL
zNvoWV19a7+y/T3JZFaC17ELr6y6m2fVbWKK6kc/zgWJ9tUBYNfg3j4tbKZ/jnLrC4muilMMODIt
BuCs2/Ts2dSv1ETgdTGaGUjSTdQlIwDkgwbxUnwzB8mJXqVuAE7HkD+CC08eOWu42lPX25AsejMQ
k2H0IFBv1OdUM/350t00GDVc/RqtAUzlj7RcCqysd2VHwAtWvTQhPICk+SiCnxG5v9Bi4vd0nb9p
HIUN3vz92qsicvmqHSAKd3Cg+SPgL5pdxLwPaGAL7MjVIgy6tAV12MDBi7yrq5G4+AAM8BU9nyBj
Yf1E0IQoVOGi4V8fGTqM9VZBf3VUS4q3gBTsyRtKJFlBJPNVYrQKvqBDIMeN49Un6NiHkBEzm+R0
8JkUlgM6umNaT2u4q0pEBVf07J4zg9lgADkh1K+Y8KT0SZ1hL++C0xZmhS61XKnZsuAtLlvKsYpN
BpLa83MNBY4GUGYR2slyhsZqoDDFNTbRcmwEqsn3boc7wba1HYmGRc1Iwc/wNUXsr6NyEPULRLd/
89W8l0fCm6daMz0TeLAcWuo8dxAzQ8FQ/q9FSfX2OD82FkN6eG7CvXRfKhrCg37qbYGBMsnz8dmT
dQosu1kTsSVbjX0uVKlobvWJvu09fofap5eyF71HUTc2h7jkpR3f55FXSaew+SSbexdgQX5Qkkqm
a+tHEeolV3PKZ5GOOGINWf7oyKII5kF3KLtc3niDl2MaxWiuvByqe0yB0XBsyzDoaIzTgKrMMid2
XYCcvVum8CMD42o7M6TqFfQ9FjRZgDUAOYp9kvjgtf3yFqG8SB7FJU7hXMmWpwyN47QIbSJ6siWY
4D1S2WXe5P/fGwHQriSkf2zB4AHewOmuiVT/0ht+BEBmXVVgrNrdu9ZMxti/z+h2gO1sgHMKL0rU
W5xc9IzHwp7PbXE1OprpcHv7HY7t7WCQn+7q025rCYz3vXTA50mkhqFvLVDuypYBFbqLdCgD7XtY
kv/yXe1D+18267Ply4WZCYNiHyLZxRm+8sbSVYdDcrwl8VrWChzDSg7lRScUIAm3duD24adRbgmg
tsC94sB1OFZ1CQd9AhcxRhG9Cro1cJ/nt8lzbfCmqenrABtonj3h/FjEotUkFFjp2K/0zsg9srI0
ipl16zWEH5P0EYs4jbiCkPejTj92jyaAXv8sSkWny5N70pGUzJxQYhWJAK3WVi+Ff/8U7RMT/iNY
XEWLkfBrJxK0IYsUb9sVke1+KzKJKX8b5o17D5jkbuF/vtL8/u8IgcMbKc+vdParaQckElJYENn9
52BsTkbqpobAhA8jlEBBCuoeleDv7HHtuJezIgA1NNDmu1Ip/f4NSCAWbYxT9wWX/GRkj4o7Mcrs
rjKzL7e1GgdTxquO58y4X1aD4n+H0d2+gwXXKKguposWnpReXSWdDbGwX9Bb54NM0TWA3XzHRJbK
u92/m9be8DkLfJzhtgKy7fZ3qbWVz+dD2MO1ltCOcRX8WK9gYzVUOwqYCgaE/Iltjy974//OjFov
b3c9W8OdoZG/9oDp4W3N20DVoWkXZS6We8Yr5rQBs64opkP9utHSPG8GXyfQnKhxvpBRCy4vrY/N
0JngODbH8mPM0zyRNZPG8zayS5Eckezpal1U8VusXfqyCKb49NwBr1d7nQcp1IBBAVsDAi94FzSw
FYaoBxUJA3LellsKowlQxH5SBhXsP375hbdUMnY8filL5t4e11dwTiAMSdUMMh7z45pyfUEn7O6D
XsrgC6BriiL8pYBqMDt8f6COs44noEEeYU2t90QPXHpV09Ou6zL56onZ+rkPrGKzDNjURV8gW+zS
bcdABOQ1Pj4To2ZKrLf1bpkS0qxH0FKrGH9t8PW9/khrP/yzq6n1QpSpayfeeD73DhvTU4QHEy+K
yC7rkd32s4pZzJNKpZ6tMyLCfoMi47fMQCU2PBUB1IqLyMUdxi28WonecwmLsFCgTjsutabcwzr2
s3YqGIYJGT7+J4R5u4QnBApYhQbopOKxWh+Q8QW7nCDgzB0D8xRvCA0+Lst+SM9DKgWttAYyWQYp
T7OdLV8zKSolLRKIIg5issc+dULX51xUnXUJdEZ7t2y84X6SqXeis9DNrtBd3hyR+mX9UIpxEtGp
qBe/Tps3zKadYDtkn2XzbJ8p7sFFU0Ot84ZD9zd6XmbGHv1u/L3UT9SbC5P+5naBzQ66EC421cil
atQ+S05SSsBBiVGj+naLBa+NrJqdBRf16bhDFFIuHPVWUGv4o99244ACwqdHeMBte2WKxo8Uvx7p
G928prFJUvhSRUhsGMnmtNvvCBtcwFOJNkl+O9FNJ6DlMJsHgMcwqcM+bHbArjZKguyPZ4X+f/Zk
4ZfIwECrKlaUdrtkHFu52wykaD2j/6e236yHTXdzoIebIhBQtISt85qpqi6bdHxjvsqp20ikyF2X
DeIa4GGHh3paNFB17ZMbIcsr6ILi33AI1vGxUt8TxbNcaAat9LX+xDyi6ab2DxjjEoSfx7eTcjU+
PHSxX083DWhXR5NqXlQa+Nr1EsecHsBYMueErTFk1j7NgJt6PhnSrWMkGfpCVLqKI6D/mHW79j/E
FlCqb6t+o85mvOrilPNiHzha0tGlIseGoCfVeh5lToF6+EZkICMqe5hjtEY2f5aZniXKZlVG6FBs
gbF1J4I7/I6sXG6yCUukHVkKmc2K/msrBlR1Rpy2cvpGBdA7CdcIC81A2TJR+ScPGdhV48Yo4us/
NDJ+yvRMb4+fFfPtkGhTwZ9AKNXMtN0XanWDP3wy72eAbYS/CkvsNyH4Xws+0MpNEWHeRSpWkPS8
Ekyx/mmAI6PKvg/05Wbbkvux2ciY5QjmUNKM6O44JBc+YPZ7GViiPhalVrnqv13dYs064yNnQ1rQ
xrrylTUFs6P4MMlpRQbBSiJXKVjE9ElUlH6uEIRy+hlDxvmAKjpdPCcWR4f4CENxVP42+c0ggS2d
ynuLxlKgvRBCE/jA+9Z14O9RAaV9ReQVf26s+JtBE0lPvVwqHeeCY8EVz6zxPCDE05dvHpa5a4Eo
FFgBw+xBsghb9IF47yyU5+7D13ypTu20tvSjrMVKQJOttN/7dZk9zst9DaL0p/RaHWzwdfzVFDV6
PvRzLZxdSdgws3sdXNbouNNYMMMiQoNVVWWdKexLJvFCOnUWIY0eZbs4IsuqlACRqL+0fdEeXaKZ
4P9wUTGzxklHu0EVusqaQfxGKN6cGRlc4Kn63VH7N3oKAS62yZ9L52EpRgWMhcubRveywazjnDp5
leYsMQk9cfZB3SXbzVGi9QVBYLoLFgP3E8MWl2WU5Bpo4J/OCBYfgriYfXMqkAE/H8gYOLybT8gr
vsny6Wl27ZcIICLEwv2VXqJIxS4H94CpMgHqHKUVN9+MR3c/xNTeUtN3Rn6qutH7kwiKI7Uee+fD
aAtzJ0PGq9FHgMGrOdp08Don4+OoWe4SeUcBM1LkgxExoce5OirTaPUnEWRJPKR2j0r+ByY0LMx4
y+CxZClluCn8PbBuZ6zI9FjSFWmkIJCUMCg9Htqk7yV9PjzjNYnsKn6iocGeBEkIIPaXeWB2vbaz
QvzOXidUUfXnSob5boa9/EseoggVlB7oTWupJrvXqzPD1EJTCgzI2+LQUPbjEgzyp3tq8mgCHsKn
ta7fxo7LtXs1LIrRRtwpBfAf85/TtIl8z2LTeRdu6bxzoWvItkAVjlDIzjjyXUMbTU17WO8I9Nkd
u1ynjphqr+wJX6+ALJfip+vOIcs1P4qnnW5esr+Ozb979tbMxFUoEWriwMDK3Yi12Uikzs4q6Yp1
86nXlsoDqYXC9mQ62IlEd9WobkZZ8LMXxVLFK1D8ZxjZ7epuyOh45P+qMGkRivIYDAQqbTbolIge
avDMsm3POehOzVGLCl8I5/FyLRctruoJ+St1HcEBIf5eu1Ul4JuQKjQILdOoD0KZlJj8aYMWApVH
yY2WYEovG0buh7M2bd1RJMwgwMPtbkqy2r7EFDTguWqYewciGb2oFfwCYXx4xtbzG0Q93vAjRQFC
LkFLwEMxnpZ5KwOfyjw66mmt7C5gzDaEGboP9N0t2b8589yEFb/OvcCmQ/TREnVO7ZF0Bk1ZLlG5
eGKobnK6VP1icFGsFqKCCjbtORkCN+H2l5TJlJhPei1+sN4GSPEvvHFzln9xWJZ5n4XWL0p+Ghtx
nSI0bK4UVXkdnIQSg3RQo2NiOMi6Ds34n+WwETAoBIsVPf2PKVfV7pK0YLIb+TlfNK7oElDTBpjD
yVChatC/OkmrVPJJ3ufuCMmrPJs3IHhS9lGTPrKqLna7HD+fPM27Bnao8MH1sUkFppYePlZbHmku
NEaZGflHIsJFS9POpV1pPldhvuuPZUUXnBZkH6IZ3N/5WgwCFfNN/avdLqGG0Ii9bLd79ZPbEgo4
D3IurKwGwDl9KjQGbUZOzfhDyQeCPxOpkI/QqzIAld+fpZDEygPZm9/xVmJyF7nIfnkqlcbH2gz3
lDee6yTEWhV+vk93ijRcnzc7RvXqJHr4qgLRD+WpoGFp6RZMRE6pgVbtAnWoVuOtEnpcXTtRtp2U
v94MoIolDrVgaV8g9ThpMoekQ0ICKsasv74ha/vGQkQknGd1vo85hYqztOXiVqMIlEj+yIlk2Rra
o9qdeMvRU01Dj0+D57OSxAuqrhHURTmEs/UNIo4kf24MQOnKTtaCG/4tyjucndLWfuoryQUk0SCJ
KTUgkzyfb5bZsOFfp4SJjgEPxUSiDLvCkM6Y3i2+F1q2jCVDnjlo9ZuWJLzJtmB9v7SagitiF8Vw
1aBG6cHPupx/6495MTUChuv73tb+ZQJ88MGJnLxN9pIRUohgIV2/0TXOJXzh7EXkDy9J7I8SiJup
H4JFOA/mRHCiSJAO5vLRjcJKCWXmXj7Edg4zwxlb98wEfetqsVP0D1TIC0PXw6vG0TFzMCuVg2lp
VsJlHI3jqUzVRRCjKlpnQWWgqn0zZ2E0BcyQQQkwiIG612P3lSaVDnAgSVVqI/CSNxTg/BNdm17Y
SEXEALn9r6vqycWQuXDR+ItjLZiJxxRFj0fnsfOnYTqVFeYXEffJRUI+N++RAGjv90Nl1c1rlOmh
bgJ50Kn/LL3GZtLaiU/xSxNwfbVrRiWODku0KQ82c1JI/nWQVsmANHEe7mAbfMiqvWCTdSzap2PZ
ymBdHMP9A7mzGrOwLx2KAvaNdRQumNeOHogxBe8xBPv3T4BwmtyxA0WxvX1CkCw0ECofJ5qtGoOb
KtrrnlZ+y/kSEw45u7D9+SpSFS6mNAoob+BKrUTEERywWwMpafwkLL95qV0ahTyKqmK8Sh0M4lnK
aIy13b6F+Sn1g2BEjUrkyONJ6bAopQn5xQa82rpBjtYVliilhlKecCqlD44Ak5krZ9drPfg8M1U6
o9O08Vn3aiCGvkBAMKguf4K//HpHv5qM7c8T0e9basJATxZAkOxEHn+BvRWsZKwspVmhUjFLQtMR
EMDBIF39uNhKn5wQOgb3maVcMr7FJAYsBQS0Cg6/ukpvEEc0IRXJxVejLsOkBDjSusx4mRLfETdm
X+QC5+UIwZReSK6vy7VYwBSoS7k/ITINOL90W3hoefERauUpLeM1GA+cesw1om7Ly3lrdc3Aw2CY
5a7XNAJDHUhjeqf2nJAzau73MWHbzyudVOJfX51hrW5GEcSYNkA7+TCBSgEa9rIS4ACXq6Pv/sBM
IcFY2B52qcKIpPT74wiLoA/0PYGAKRdLcX6zBdZCaOeVeBsq+ZXMBCDg51MXwU7kl7Wkt+IyqlE8
2bWl7vn2QyNmx23IhYg1ZhE19PKHQoYHbngOYU8EuHI/GSDqbEQukLppbn8UZxuIie7zufs+xjgQ
nSUbZ8o0OHSiWtwAATJOcvUol1nXv6Faw+5C+YFDLCGOs40ycvsY/bwTT+VVEHNePEJX/HATPe/+
qT4KRpTMAKHcn6Z0pvc9jrcVn36vr9+RovXUmf8fdkuvbf1/7T9OSnC4TTW509fPot9gD5KNkINw
Bur6fn4lgLJvrG6wzkFecsx4R6hnoAzbO9m+i1JT7VAh7/q30EMaDrpbrYzR+neNSHr2NMF7rgqS
Ir9ACmfePYM+jOgEdbaoZm2FDeq+w2jLBP7ZZ1mfzDgxRTsjoBEz97o/UQD58vbZf2z+r6tYzVQY
gcPvL6f3AUUYrEQQYAE8Zdr9WzgnH4lTIdTVJd2hf0xj/5BgRCdyFBIVpsSQgoSxZUMm+rlIIldc
Nk/SHgn4zor5l379pGyVcA1qdeIe8HNCoxcHV6xZUluGBZpIQ+SUL+Fweo6vY4LOJDZHFJZaqdx4
Y1rdkBqDULVq7EdAnL8fUIElTa7d/vNKL4byxn5ZQeJ1HZWHEHHS9SeGun01jTllWhSf2o8Q8S/g
8YhuLmPpk+EUk0KJhRdmT+2R67T1SY3RH9WBJrnLzzhzekCMEufLqYG7fHJWcmnh5MBIlpnIS07m
nQjiMEkDRkKdwWLUShCB7fS0ZH3m2Gujec2GYM/8EmxKRhzFkxktUCrMBKxfnMZXOPOrrBTTdiCQ
EP/y9fft50P39+EyDgcZLdq2Xnh8RrvZCWeFbsSSTIcMBbBk+XMje4nBjLEV5eqdfaVHQ+CQZcYA
L/MyBOHEecfVZET4TGCSNRihOCme6THnXbIieEy8OBKfJAQ2mAI5zwEmb7m79g2mRs9aY7P9Wj6W
jAf8ghhDJ2rWvbqJy6BHUS9cFbUBzSQ/KB27Zo1eOeokrnETmDBPKHmJ6bf8EArLYFo42YngU38D
4vhGdSKoyQyj3tE1kdMK8Qc80ujVi9smjLR+so1Ky1o/Oklm2nOECfG4yuYj3czxH2GpRUt1VFFt
OoYt8Hkw9NlNPOjMbCb1yGZy/DBuWgzB/+HXxoFbHy5my94CLSG3u/dihzufHCPeHhYcR6GVLVms
rvAnF7XjGy1x7ubP8NUkcUvAt4z/2MffV1jK1wJBg7bBLxhiqHWBGx9KuYL+Dm7Py5fGSmDuVMqU
rbhQt4Ffwojgqo/GVoCe3n79SUez2Z0mErC9pDY0M2JpPBmHheYCdEmLbkcmisBbyo57TdIZaCMC
VyDPkXStz/nlQkcDsoIfHMNZluUXuWFUX1c72WrgSmBIpttC2v4X5IDn8doWNPN69Cg0LPO5iHe8
zLNByLboeSZ6l29nvCUyNxVJjyjuPWoPGNDcR11zbDU0BnRNpGIAmwIVWk4CAQ2IvdkOLmv3Zluw
qNolHRAV5q08E3Kt8ZEr1GZpL83xcbgHAURjSCfCJKgniXjHCgYTOJhcX/4t1couP22T5+OEpNry
wwsmT5xnBHiJ2pqfx1xtx2WAbJ6TecSbOAGlOMjYNf3qLSCFhzh8dFERzw1+nwpomu+Tv53MM5PK
gD0n5fvSHgcFWn2F4jAr19ZUyGZDjcw+56A7KAqeWkkiHJC6VlDXOlaw411eIZnmD0nDuUQWkBfR
LSxOgGDNeuJB/PaxlfYClyQizRmRXdz+Hyntj5tbZ569FJpym07AjuM0e36T5d5qL2MdND2WWU9f
ATe3pi/yaTT9wcE6D3FS5jJq3O82lLmk7U3ObGGvQe85MfuMW15VyqWKFYhM3RCzDXEmHAdfBLlU
4wz61w4rQeCB73cV7UhTczMeZfBEs6nhAhQEmbzYSSbKYnKKKOrWj0U/aVRdqbEU2iqWyfIQnZz9
lAebuh8hmIRsy4DfR33HZY5WwzaPWEf+qRAOcPmNa3DnDx+qi+iuneIr1wXNTBRKmBQCl0glDYEW
3+22sMCXBjwq0EqLyb9HBGVJCUrI4PglFhda35oHyYHlRzL32CUHo3uf8XDqQWkb9VXY/y8V18EF
oEgUcY5pMIjcCmIz+JJnVF808/8cB3DmUbV45nFZkWYxFAAheCex4u3nJpgRdLOst55bL0hdKjZy
sVvxmkZM809I9xdLcAtFTQC6pP4PHVc4dsoylmTP5OYqPfV0QdP4GGXu0m2/r5tlrJLYeT6R7OPq
C5qcHKG6d/VgHkj8MQvbx87wFXSkTPa8vYOZkfT+BApv5ptNqeV5E/jhlh+4ttr20uJwwlybbAY5
XOaaTv+O7R+FL5mQ+3iJrIsSoSA4VybycUbpSZ1LCzloP3P56+1wsCGx/XC+rAIZwx1uuASoH/0m
A9rOUVUYDOaMYv5I0tFGOLxRzShq+TnNRaR41Lp67Gwl66mGH3YRAg3fy2dopEGQQB+7wD4bf/BI
+xHpy6rHnCJpVSeN/0dI7syqdpWvtcXTOS1JlBQ1VYvT6HZKBYpR8tcr8VmXgVjrfJeGV+dFIZ69
X6n5+pCIp9wnb+m9IS21QTn0hQQf5fAg7SFFvIGzPv7D1brUkCD2DH5KcH1M8hIv85DidhXifGj+
CBAgvEitmsMNuEMm9dzOXCR4ntdmTDqRdmdi+erVxH/co4mapst85ZvhjPtPRRlDymMXwptN5jlC
9hzbPIZMnWrapiY601oUg7/MqhAg6HlD9gx1LWvtqU84gaQt2MF9nmW0vH3MAo8W+DfsiWnbV+X2
ZUd/RDa7aGGoz8QPmMOGpV4c2XNhxxM6t/rmUVcvhFFDgpYfHsJ2M08WnfZd+xUgCQCiomXFh7kb
NLHVKzYe45hFY7uplTmO+XfEMKqNBA2WqLCJmoXcA4OFGu79hIH7uD/BIXxkiOvt9qTwbYdH9rEA
gwG7YHmzCK9YaEnB2wwaHuAD27DaZwZAPiqKVlW/S8tiyFplmqQ4hNPv/5YZ0kqO50ybK3zm8rFb
EQBAdaj5PzgMX+mpLR11oSIWfA01OMIDnlnKB2cy+FbZhamUZRuSLHEOJMpy73j5hXFQ/rZ8ZSfS
Vud36+5i07DtUIbjgy0LNHNWi1jENGS7sbHzaBIlSTZ7Ay0HYNeiHaeuo2QWqJRPHmhN5uGVTjx9
JSb0kHUWpKDBK2ESBuRV2GLmXD/U9/IB6IKWMfYspgcJhn3KIblvuIhjDCyBTr0D8wR0oRebnBHe
M9Z/xtoqP5Ji8prNsZ7L1N+DnwsibyVuwzbvEapSKBfSjCGDMkR3vnRcWj2aXb96HrZ5fg0d98WM
MuX0jXQhWpJKMpKhqkJ2lPsdSYAPOx2tYRKm/uOClNW5LKPyqV80vYbd+B/OBns3aCnyhLhD5Mp3
1K/d5AWDbwacJC5bN2xPq487e90035Ir456TifYqdcpmbmECSjdsIxCUjTEinMuVS9ZLgZeT/sc8
WAFqyQEyKbQBXMHoRufJqt2TlY1zmtohvuCDyWEPUX0H1qqtRIEGwsgTh/G3cKXeWOvAOHyYD0ZC
NUeNAwf9mo5triE03XW4kuAxDOy5e12B4nyAeDjPg6KTcUdGlAFAM6wu5NIHWfFn10pRUk2FkDSB
b/MAEm2MTZwpuff8CffEWBUvWz7SLWVbaIb0rPOaVOD8YFxVW3qrrdboRgpCFeXzpRe0EsVmOBqD
IyCc94nnEYUPb8pEj0V4EmGANM2smSz4WUp3hF0k/Aywft18uHBoaAJvDtbBGFwD0OOCpwsm2xEG
zy8EGsCnpeKzeKLq1JL0tq4Yle+zrdvm14dGsolAYkPhgn7moFMImkrx2NXj7RXty+6f0ojgcJeF
/aXCnEdIsNm1V/It/Ry3NGjmsqrvQ2AsaixzQKx5VJZ97+uiZb3NU3sp+vHtoqZDZkkWHP2DCrFf
Hx6lweNjHuJaNrz2fP6E3jvm2iubuHewIpaTKj8BYM3jAUiKKf7eXcy6C3jXJQa9nmhtbyRUx16t
B65QUziai/TTesgSy81o9JvpmlL34tsxrWmfjNFdDikN9XE07zlAwYDewNOLmCy3TsQ+lo394cZE
GJeFwlX3YZipf2LdXwNKU+ZwVpm++kf7Zq5J8TwJMcUAGfbg0cDTEWkclCqjB2/CFpU08kQXavi7
It/0IuFWI3wU1TVmkgFGAIUq/YEthtI8YQcM1SnK+Y/3gxnZcZnOBJfkDx69gBmKDo1mQ3rl/46T
eYISTxk9CXuhWFAz7wZBYerqTf4toJ+emkfFGDidV7vTW5q1PN2ZVxat9JEqE9yBiN4k9nxV1XgC
i5gjI4nviwMbkG/HxTM2i9mnpmFNamJ9e3sbnlrUYw4d4fZ40AlFuVscDdCSA3WKsiErbkyz8qDJ
SqQvBcSzqQRz/ocBTB6phW4mH1PONMTYAmqN2tm+w77Oi/5t7THIXBOzyo9xwVn54vPAXugL7JPV
3Z/7DwFATiNej7q1L42EWyPnL8CfsbHtYoLf1DyksHlO4SqglyCnWqpOd/3qOcYYro+h4NxrxTcT
g8fn8Xax96BPn4ISWzvAfex8FQPh1Jpk2iKqvOt+X+rpLp+63308/4HYWau4EccyYSjVnDaZEUeb
i3yTjmfj/+OlXANreyKhzbSKWgKmmwuqKSXcMgne/C7H6U57WiN5W1ej/UObG53980l5McP6xACu
v9lK5M2cAOc8rTodkpeCbh2hnqSsg8kkrACr0P6BVwWuei13cz7feKaICOnbxf0xoCConOLGtwx0
01NsnXPqqx3oMzfxU3E0sECo+wrFXdpGk/DtsjleTHLnJJ3hMrE978Cjb8d3fAdB6tTKe6Qae2oI
MTSxPBytXfmNLVmxVQPLKK+nsNoL0+mPEJLo4udDYAIZm75Lw2zVrqHZkk31o+7R5qnYGLtRBlBW
GMobXAdV/beXWyoBQapRiOeuQe3/thJV6CTyHL9Fs+uISosyNXGXmQhZ6LcQuE80/Cg0LY4fLrnd
IPK9oZ8cDkvjYXXb4eonDgZmHr5UTpGBW5UgAk45R72Jn7EjYvYxaSMyXL7VP4A/7BCcujgS6Z/z
7HZUxYeF0clX0/QTT+GA9DV2bXli3gYrkmQxGc4wUbR0gD+U0Vl6UmlBO63spsEDd3ze2xNwh2Pg
sgtxOFW8JVFzXiE3BBeCxANql41vtnMROrFIDl1SVF8+lxviL+DMdWbK+QT+TUViCOAUdPGl6zEm
xiOz0yEj/WEGbRhsrwsAMrZeGTvbbCQsX4xGiN9sHIUCZe9iUigg1gSTOV9JJOKg7qveBXfiM43n
otQ+dbBOVSI3ky4TsqI1PK0uN+pOrG+E3RQq6AkEJh+6PuwCo7hVs7hYDbSysfRwixV1Udvqh8GN
AMWAkA7ikI2zKPHsrrhoU39gzXKJTPJHtRJJ8V1qq9/hqC37tcaSIV/Z1TPHQtIlzxdFDLGwf0wl
f3tv9RodVsKzwh+yEC0zkW8TPRpIJjg3J40EszQfx8VZVeZvYZk3w6skxFR6vxLn/jAjspDe7bR4
7azdLv8nCtg00X9YgQ1+c25IVs2kf9OG9HeKSbK4+RRESb5Pdrx7zUNt8rlbjBgfNdIktc1DR2vx
wys20EzH0jwkijjoo8sTy83kYhjAgPOY/Q1r/dd5jmlrZwoCTCTlchWanu/rUJKjJzezfMHPER3H
VQ0jvc4uecyK7oABNoUWgHyUwZU/PQpFFgRkD9K/OA8bC8QdUyoBHwCxdh2ihG5I4B6CxoGk/tqx
T3gNAGsnl1T9nSMGbopWMItINNWy+SUas/GQJ5hxh4518o3/d7+q/zKAQG+6k2oN7UUKDxQOAXsk
MeNEpY1sFVYT09Jpc0CShRPdxj0NlbbxyQR5AYtUJ7/d94KEKyAF/pmepL5Z1yNou9XeL9/yjE2u
Ky7ZZEovHwHDEwDTu5hksNhYD3501INJbeJ9G9tp/JhrZLdcXl330KH0EYn8uDH/HTbaqS+ND/3O
eku6UIBiCCyI+7EZBnbdnAUdhNKgMKe9TYlG5aGzyTEbo/148GuFi5UsbTxEnSlq+sntFaYACUEU
T3CHoxrmjP889J6YiCXsPWOkZx5ki8toZNGbclYn7ErlALyPaYk21EO5pbNPn5l8feTR24+l5DDz
wURsWGk+1WDwMM7ZrI5S8QMMx+1xayCreS2wuB0pOaJuqaZUBrN57O74W2prYEOtuCnAcebWV1iJ
rf52cZa2Om53xsmPXZoHL/fNo0VLQ7aOEU0pOEfUMOz/u7s6bD3HcfWsNuDCHD5/fSFuQbLEJ8Yu
JVOB6K5YkvZDrjDOdkuRLjKE0QspALpBis0PFeYz2RQRUPMfWJmbfncjqPeRRLxO/0+HwnV/v6Qt
MwJjLdgNCEZu+T3+eaLSgBqjrBy07Hrkt3j3NUDoRaj47M3y2v9+G5n9CKhb3ojUCkItl+Okg5wW
nvW0Tnw5mze8+xlGmLNTcGlr14ExED1R0hciGHwdO+m2x93eZ2PlsJaXfuExL0nL5jjuQnXxC5rY
eVh8Gp5mlgLgEtzTP5ut8Tystj+t2ZE8OkFIPAj3y44KF9DcBd7oOiySEFoDvfVD5JXW4UKxLTyW
pcYmyCElLU5MfMP/9Mqcb8yl2ivOGhAtpbj542sRe9goXX6W5agw2jyEOyBVx8gYHXO6aap5Zfny
Mqi3leVyxaK/TlP8lcftPwFLWFImo1IDnM5paGVGPFGDoGg6QlWCMwGxCe6WK6vvnzYSbsVQpj9+
2YegMqCm/qLgToBtJ4vie7zyQkC1dEXADsY3iza4qGq4GiYycAMmd19vgzj0mWg+mYr5H0VeU2B6
OHDBYjC1bP70MhRaNosioYri2kQTkg/+KRhruwfTEtMD5kCkr/AeTEOqq2jR7XLI4QSTnW6ooQli
SjyQwy0YeBQHvIRSDiosP1f/doGGeQ4OHDU6yJ6Vbt7/RzMOOVkDVW9EVvtfkT0HgMvA2MIfp7wF
2KSLJgMDyrGm6SzunqHIyfMuJdnz3jIWhe3nV+SKYSKwdlLmt6EYzS9d1xPxsPqgSAf2wtWyeqka
iTPPMOQtILNW14814VGiL+ip91RQ6XL94yNGKZg8J+89CwhAEoq+FA/EG49UBE66e+nqpt6DlVG/
4Gr61e0ggcbQ5Ax7Mksuf8GSxFypaL+rB9rxYSA7JbAtN2PFu02X/8+wAdXXkoYtcbJf5yo5P8Tx
VaTnV1eIy10NremISlCb7C+RgwK4jU1qQV5deEUFQ4I7utUpaN/yapXi3qxTHj/hzzw/8SaIO9Sx
C/Op0KoSqtxCZ62tFV/FP0wR0FNTYOsliFUKY+EmqkotegEpF6f301V/qeWgsofr1rj4N7cJ/YXr
bg7ee+P2oYshHzB/PYzpXvteuZDLDyII1rsgKW/jPAF5krqdgL6V1I5wL0MZnNo1a+/HBISlbsl1
Kt7MOLOtPehQ6NCDp4iM2g8gdol800JwORmtqpCA2SSPSNgZpt/t5FpFWDszomp3fZMYZmmogIgw
SwE/aAcYoYNJB4xkCIcatC8FlHxsh5QxqrnlLILhZTs2GTXSACAzLdGs8Qx2RQAGkXPeajjmHkeO
130aCJqacfrhM9Air/9V7eQXOQ2fKpfMIh2ItAtePETHdyhOeas4ysZk559qKwHJjdMD7a7TRhj+
cQgixcLNLrXkG7BIZXH/u8Nx71OpD4j/K0rN0kzpWR8puAqa4CpN6DCmjPKpzYABCVY6BVp4kiRj
AMKUZA2pnPQ6OY95upqJfk/7AnAXlfy6F69kGxzsAiUdF8t2JKD1cbXT+NYjwBufpwqd53zhBJVP
zGlxeaq24+VvRyZ3EJWdpP7lQRM9sZa/XiIC7LwQJ+oLk/7UAbMbprXgaWKssuli5isrKrBPOCMm
RZ/s2z4fajBiHP3nVPTFGLzrBxTPkzsliL+k4ufySa/PtrpV0mBF37leWbJL8RZ3Bk4oIebMC58a
jbdEmcdVzZHwLyMOHvIC3DVZ3atQBecGtnJ9+FbGpxNCxVP8BroGD7b7AszApNoM7S8GoZspslMh
Ay1XACP+BK50b3cwCQb8E/vs8zmu0fk88KqtxsPzyPCzwAFPq4xRTwaQrhFcBp8AaAPnwBFUDdB9
4YOcz+XRHueiIVWUYkhXwaxf9hzyH6HgiHV+PCW2jDpebzq7J8XVM4rSKFjpOyEph5ikVR0hA5LX
umu3bYjNYaccRpt6ObjSeILccVeR19uDg9r7XuUbhHgo+QU5A+15wzxXhQw3i34TEoGdZgP2Pgd7
fFDCbEzDsQteBxmHhqWEGWTYq4c58VD1uTTfZyOxXr/Ld/ug5Vtrnn/GTyjQCKA1Un79HzEnfbFo
vj7IvQOskqjQEU3lIJa/0h0NFmztZUyorDQSfFToyeA1v/nI69p6ALH10BpVKOWRLZy53u32LuIm
D9WBain/j5BUBqrvf5u6SO0NK6ziw94IyeBTYuSlV7d5e3CNtC9fsD3MAr7JGNxYEJKAVVO8asIR
v2VObUxBwJ2fpQxWMg9Pgn0wGkUjz161MRLTvPvKakkzY55JoETS/j0IbgMta63pr6Vnmo+LCRLO
/MniDormwID7K173tBeN0vr5NY7SSq/ruiM5QNmELkMx6A1qCbecW3pzglFcLPt1z3K67JtWeArV
SVsD/kypNjK9GWkRUKs4EOsAM/5N75aGfVADBZVgpx7AJ0KrlJUkGaQDsLsaj+p3dUCIB7aQ3Ct3
UWXkhJPEV+E/Sf0LI+rNMTQwPNS/VYGVz/kc6WkcU1haIjBC5y7CbRQmEK5Jpto38Wu6+k1wm0i+
qeTT6giIDA4OJK/PA4uSU5RfQ5GqIyd6uWJoVz7WQ4m5Mc9YxGDcEGqp3yQQ96VScR+VFwCSAq6G
OCFRRj4412ktB87o9cf/bEd2eZBOblelYTlRh9pc+kfWFs8rQuDDJyvBf7eALIp5EVcq0mQgauYB
8+DA6ref3onc7akNKlC3Ph76JO7on/q774CnAeOdKvWeqffAWdsglwxWzosNnrnofLs9AjFqEO7z
uSuDuigTdLjtD7XV2EJFlM0T2kRv+dMv/xu0nC1GuPrivHzVI/rbDtIM1aNpNRtUKNOKPIds47C4
jH1DqM4sQbe/2gvexzYn/U4KakzAIy6kSmwwTuVOV2yd7J9cHaAI4C1BkMWV/3NQQEuAf0uHSG0Z
QdWiOEmgG0ArseUjO2DcE/d2KRnP2Bgm1dBW2X2pHdeW7HW/DDbYRLs24nXxO4iYXY82jBj1un4d
3QUIFzXrAVsgaWAsdMEqzoXlNahEE23NHeROpyPCyn7vdRWWLgJqpI0Wkt3onQizbEo9UvsGisda
ue1gPA6Jb1fhyUoIdJEl/iTdRATxBTRCiHVfzPQDGFGbDo4ni+z5i6rCLWtDrKXPotLtdphm4cNt
C9L3EdKG2xZ0Tut0BcdWA+n+rZR5BtOkFGIV/2xTuxo01drXj6jBs/baLWpmrHbsEOzEzXlXWX84
EfnzLLljwEzi3CKqHHaxVXnxuGV+aZsUtQ3GN5NwolJx89K/lwC6zM84WymPxj5o2GsuuLDX7gJY
Qxb6VOJ4Ea8S8Qs3y0JpGQ48uOdMfbJ/oa0EyxVrmVy++Q8BKKlgLTFceYKgttFJGhZBrkekyTbE
8TodonfwArK8feah7oRlFCU22xFXRt8IK4vCIhI3t5Mux9giuMdaeGfoHc9eF5amyjqJRWH94RBT
KwcwJAM+CXCfO5qfxPXjos/SYDYxk5o0kMmkqcmNZ3fod5wD7gVHB2eHiI1Vo97EwkRMvc9HahYR
j5yPyZLDl6f/uLt9bb+WG6KG6lVXlnlfu27O4XdfDqYnLQ92DDYRQUKBTsoFVSGtAgSHegGaLFlC
K9OEVlSg1DSSsjyJfZW+d5Fz7aq7+SZ7BIFBL+qWEFRQknKBGvJO/60J5/TgENPYgQAz0wBQz115
3OXYApXKayZh5x3Pi0/AQUc482/u2AqPyo2WZs3jQ8KbUh/J9Cx2Y8KCovDye4zT8RygEMRsOF1H
MvUsLTGu581yx6iBtwl3RTmpa9gwEG0MVGozaqRv/q+5UXtC6NXd9eFw6cFlWqi742SrYzjo4YLc
d+BRj+5SaNHr5Bj5wmFI7RicwbUQRgqSNJJQwNVbyofaaTZqFDNPsNENc0pvUNAhpc1QEifzZT6Q
4OeKfbMO8h4wQ7/2aKQJo9v40DmyYUy+jQEVDJGOgBe1qjNFBy7TMwp3Rme3S1KcR8thPzqjt3bW
hYFafo1SCDI/qeWxAlafvYdjP3FprBf7gwpLTi9RGztvs4zgv5dG7y33XpassBhJ9ZIGWU7gFoAn
vYLzIRp8teA+bKLLxPmEP7vAVf1Asbouup8ZJC3WlDRQXCjj9ruCbLC3I/cJjLXwjg56BvdK17Yo
x6xaeCVziHxOQrpgMmqGaLxJKzNtk5gkyLTF1TlNxevN0mO0qWVa7w8Nd4gBo6SCFZpixt8gndUQ
Qg8fcL0VWMXOhsJtIJV5B6PsCGeQGfMtrsdAh/dv/mpdtfWtNoLWQhBpbTT6tUZyUgy1A5ckgpbF
eeVhn72xowALONjc8/0OFhXtHUhbV7+r3I7j26VqgMpjtSbujTEmM5/EFvInYLVUoyl2/O6JFTNf
3MfdV9j0qAIYyyoBIPk+6DtErMDOLRYKDPcxDO4Fg00sJx4rCfNjVyISHPDk6X8RKnqH2quvEVov
WtS2mmt7Eknoqb1c0XKYUH8vIEAIZxa/NKKVlUzn8zQdIr0fKQmVwqhLbCIOHJoQzJJFzaNHzfjJ
tcbVyqAyrxV8MD+xVGS+SRa7UHPNmBPSTK9OrowT1T+V4kWxeYyu3qR6N5OjjuCLE2luXIREbKew
0aq69w/qeEAqFZBtqHVaviWdzdxa6PaHDku1eleERXtMolqfzantoy74SqjsrAFus4b1sGq3RXs/
O2PoegGc8IxmyJTvfhFhmhVpi6uAXHf9YYvor5RAPj1IhXFqWu2yKgHQa1ZiE7HfmpcCdvQ+ZNSJ
YJxeEqAFR6Gc6SKg3fQKRa2KHKT56t/j/Cg3VjqIpLscW87XHCUe6kMVS522XGPkE5lvMMBpVlr0
VvDkeGLpAecOqy3ym8ngjjR3idLvJlsYclGarLnhHxAB1C5C/gKmY28YI5xouzvJLQouH/oSHhkh
wgowupscChWhmdinw8IWe9gimUa5KFV9t+j2qNyB3J1U6LThb/q9xfD7oCLwYgJkjU31An3tO5gc
SevDiyMrIrMqX8kvIE91RRSWndrkQ1zZa9qSqI04H4kpHROhARlRhnh2h9219jayBnYFqL5sesBu
lsf8KTTm7jnSt/4hHA0J3F8XeqRcLAtjRwzn9+Drv7EDgfz1GW62g25wxeGO+mkGWvkGc9HwF5Gn
pFf+NHNJK94biYq10KLE3ZU1bwzT9rqD6Ps7ECh5OZokacc6EOvnrJio86bDDKtJvWiLJFZCFiZr
r14JdizvGIZJY4728Fwt48aA5k1M5ig5vpfr4NAUurXexlqpBQccIYXUX2X106+7dfNlKYXFa8i8
ohPDgtdVeIbZYLTQIhpYhwjltcLOPnaeaswf0a/X//P77BcWc31VnFw+KP5NGrmH5QzNKd4xaaTL
9xPX+iGP582KaM/+TDhvV0eZyEjpiNTQ89Tb8QL7UVSSiY6OJnYiw/EChwaFVN00AGQGyIjjrawM
eqKE8yl934nBRmyRfBSLbFkLIhCCnQIuZp4/ApMoHAY4QTWuejYc/t2UtkUoOn2mCpJJepf/Qdzr
6XAT3LzzgGWBP7LjOA4YpIBHl/Hyl4ZaaSvOwEm9aAcGJT/XO9/nuIQuKt9Yc07Yiq6nglsskYcu
FfOWMSpaN3rGaW3bode9FsvYNTk8Zjin1XtVTHYLXBUtU/6mPg+grGmbsj04jxxaoBfx1iQvxrUk
b+NF3vGzTgDf1e79MRSiifJzjM4TGkRxbwPS0f89sunv+VpNaahB+Yeg76vppK641BfOEkYvJhFl
rRnKRYdoyCHAihw7wGydJUGEiR0cd2ACKN92bhO/f5jIPAxBD4YytHiMQd+ymih3q7q9Ov2JoEWG
Y4Il/9ECeK2QKJs0kyCO9Ex3ksLJiTc5gHnp8wIkXW5xfaKDh6Ms43Fv1cSPwjh9NNaxC5COro2L
KbiJ9jt+cKQeSKJrF0ggwxFckToArDx0BBv/zyuJ5AXKtWw4d9NLFQ9nl7Q9YwsXDU29arqL0WgL
+ef3HRQGuG/pgYYu3NOrb1V+ssUXHc2axBIxCNonUCAyVL3MJi2DnRF7xNK//QSlvyZbfCJ2RO+3
Vt1U32ZYBDdlT8FimwuSHLc4/2WLZW3GLW9MeiDt3xGNjmDZvQlvJ2bhOn7ePu7Cq+zzR2NBtMvD
0FucvHxN2kL5eKqWLONqb44wEkPRgY6bDAnpQXqxNjlO4iCkTO+NjoaEdu09GVfnEhtB24mnKgT9
vKbfIBS7Z4GdweGfZ18YpVF4BYF4ifBlAzWT29EUBA9eWxGP1DAtwYzowDqRNdKnVb0p5pnBS2su
ViffGUvKOwx8dCiszm2uyRAtt4zdWxOgIr7ifc6y8sQwNAViuugiBkFQ1npkDJbMxlfUwaBBPf/s
L4Fjs58sLvxKwByy1CJIfJ6qpwnZ9JKzoni0ZdLJ3FgpHkzx54+gXZUaQoT6UunycmVWBq31FzM7
pKePER2KbJUiC1gk/7zoJVFhGkobcqheJ+RVp41QqTuUbWF+cNSj2xDqazMn8mjwLWeY6awsNQBH
U9gaROtno+K8ToGtxox+tfcJcDBHNCieGuxqxozvSC6JFSzLf4qb71p7pWttL6zurXPlYhs1D+bt
zSyKE/ow/lrTjut8OTaQ40q472rfMUeCEFDpty1T2gDyf4Y2o6Mc8tryOuIxm0Krd2g26+nEizXJ
G3Rw2sAsrxyr/cxcC2wAh4C4v5HZNzsBM4fA5o7l0vllDZRDW0YPn1vfOaP98EJVQnVnHijsA5A2
7ZlkReslUVtaA3d2bGuQkQJOiOrlRJP+uASrHN0bzEKM8bg+8ZsacEXZrVK8XSOoIDYBxZuhxTwX
INP4zf9MQ+KK9424fSvBgHRNBiRQExguBuIQuSajvySDydK/CMi/RZ84+ik+UgQnzrxLliPMI901
xDmRc3VfT3r/s0oSZuYgomn01VfNvuhYgGbWGBZsq96UiYK0fyyqtslVtewTUce80VF/Q0vssMzm
KC00lpufsfL6vO8+pv1j5HyDKcInvgEBhXgfGevjqEc/8n54yUVv9DOWXDnQDkF42b+ckdfMeBYY
jKpbiGwJVbUT29EQH5gDPHR0pGXVfKRRgqxV66bayBqyVq1bIhhLqAsksrxktcXovGfhVFiP3IT1
TViGRMxmZuFew6s9IeMEmPfUao3Hx2yhN1HRH2/WHCea0PXFv1JqscuKnLrP2AgR7MSp2E3c2qJc
nBJOZq0YdPo65GAOIaWOOd96co7woPu01QlKlop+2yUwJd6S8nEo/DgugR28q9qofoo33V7dWU6l
/V145X+H6UYK+i6Srv/xfhEp+1lXLzeBeibwn3DAsGbCMReZEorHhZswBUn0Dij22U716eh2jbFw
3YIhqBx1y3Nho/vrzYnNjujOD7SsCdZsxxPxhUgy/Po4AmNJ9bbu1Lt6FCBCSCfvoNvdM2ioSWF7
9rraHReLgm6af+UZogSfUqN9LXvH2BFa8bNa0Tjvw93KrfSgNDVxmtvgmMKdKqthvrpdHilF2Wf2
9qU8dbtxZ53QADXGOnOpbE6EJ0SSgGe2ye6XAzqpezlgaxUK8HmGaul7oAHxl9eOLg2VzG0AtgKf
v3oBTflKaaylYZVr8ZkK8rdDzm/nhBh7ZPVCqJorZzRyaJyMPcWnzk+UcU4Mh6IJGR38GustgNQV
iSDPlbZl3MfDt5trIWJoBNGC2Ea/2nHiaUX/hJmOpgOrnHX+e0EbTIr+mNniVB/6A2VvyO/elDOv
B88gTsJ283eeaWc4gTftA99aZxXnkY5H2Gcch48sUDongxUEbSAzba0JTQ7V+NyHxwIw7gvAbkrc
swtdo6tcy+3GIm0m3/iUxyNmPx44+EWDAbE/qgLqDhJVn/pwqfEA7LpT0UmysYsdbm6WIYRCNTuC
vs0y/n8WYhpf47BHfacsl+bbJ6vFWG3LxW94uZxBW1iSEb0aj3bU2hAY1pehGRNjUhzby8HQhyE5
hf8iIlwwpwDfI1LE30nL4t+sQc6aH7an3svcWNm/Kt+mLdt9b8MBE+zSS2uh89txUGStl3CD78/e
8lm/ZUP5yXgjW83J7vxaSxP9yTx0Lhmy0KCYxFwIeQCNVhUYMpJc3pNXGzX59kaUBLgAaCBF00SQ
f7y3qTHy4RSXaDtKEwsm8VHo1oSEeLcQ3bxNl5nPbd3fgW8np8lzAlJKdTadwwZv50BDEG/u0gLE
YncbbKmGWq4JwK7sPm2vT2UX/QG3Y8NDNLhGRWG/+YJy20xkGFtXLLBNjM76I+Q9Dm9jS3vks9Tx
0MECvaRKrJvftp7SZCRs1GeTEP7t/4elEX4yWONuJZgLEKwG5dR2b+ZgWKtaiwUVUG/zv2PbqEEG
DiWsAt7CLMLzX9qPO0iIWm7jDo+nyaSguXejiPArJSM2KkchTm069SUQIld5B9PHKxfg7mF0SFNm
tarcaxakBNeIOtrPLgDPpuC13zM3zSeVTF1aDYrC7M1uCC8Ggpww+C/5qfSoI9AEG4PknYO3GUZZ
P/G1azzYPfKWE0SduKatNLyjWOFEvn2GehKbu/Qw2FpGk5xUxc3nR88QXyGY/ocveICbeZiTukdW
anaT2OzasO1Qs6o0sVnZ2TIFR31It7mZtEButaxr5FgSqJm7iIpCVcslac7fUuXVDRuvVY5uYiVU
1Q3FUx2j8ECSwqAtrMQLTC3eP5rVKY+iQOHipSzG/4VtB8wvEJUNANhsUYKoGEVKMnqOHn4XrVQM
UR5Vigd0DlneZoOS805AapleC2NWDf7y/rDTLj/UMqqTVAc7yWz7TEFuB4ghVDZRa/3EEAC0/p70
da4YHU6BUNguDrLhRCTbrA1btULOHPbEfiMVzmmd8/oomO93lM105EcQN+g+psvYIVtwZ7n9vgjF
3jlxO4fjktWP4sPCQLjEB7mgGt9eyX9S2UA824qzGyNVn3Jfv0NVpTIbcr1FPWIxoxceifdZTX46
bIPTfXiNvPer1hGnq74YblEdzO/dVQZmBPVbTsk4tC608gzz7QikKQp1jg682vKUQsU1/VFiL/py
K8fL4t2bIZz8oVSSF5FO1M9laTj+Bu60VSBVJ5Ny6RCIe5hOG1zXstYdxf26lkDGdTcbnEV1vaWF
+qVWXlC2DfW0723ICtkLtk7f9bj3R/ur/HmyDGoOaQmWOTznxCqznfNZh7Z3iCLteOfs503yvjXi
XE45jSsR9mp4EKdsndDuY7TvaWB3FFflN0f85+cdgPsl4OulXKIesPJILEjSmw7YjsHW7m0Lx5QA
0DvaQZEEjz+eAzomVU4y7dziOjVoJM24U5WqaVgsJz25w2SHoifGASvLUmgpylqz8sHOGyj8sHih
RjjQ21LqvOdvPUoOFWUv5pZzlew8vpkghX4ETiJsH+3iBekXqWaMUnYXGCVXcB77fhwvb6GHjs8J
9SJTFeeJSJ9P1436z6pUfpuMIcJ6LlkERxBAIGYxOTXifXfG0akOeRHLIeTYXHgdBF+Q2aRKFmm8
p9ucA+2HwqIbSgNjrWCzi9aNj4rFeSaTOy5pUdp9PVgMwrmlBh0q8M6lFGy7mFAUmyWcW4ExLWSk
hI7jyDZ05AX7YB3F46fVPrT/FNbzx8t2i9FvzDpXQMTrVw26i6uhKCorm4toflXwbCs8cJ3hpoaP
CRe0ZuGsr5lXCo9N+jF1p1tS7niHZ+JcuTzPOzfIyybzrz0J2AwGUXXB3FRg7WeRzVyXDB4F4XJ5
iCsxhIgBYcwoCS24OM7Cqb8ztW2n8hwRl6X1sC9BpgpnD+dMM6K3hdmZmnXYfQT2AkWY/TB8lDYl
+soAO4GVxBeFr3eDjxh0mJ8619xEkENh3qDETnlm3y9vCWOeLvXMrbHJa7YyMDl9sG/USdLak+mj
0th6YMzfYRr3WNEHuy95981GrcQu0AjEzDnvOkYj1zfbVcI/CBu/WZ8UHZbfkx+BOxmFd85kFkwX
eUWIXuSsCa504KJrtmZttS6euJkCoy2teoCibdhIByI9q4bCTkTSKXWvNHSrOhUOb+idi8yaHgaW
7uR4MdDx3f+dQ2jSoZz45p0Vf9d0wYZ68+Ifi04YTJsqVAme405GvRceWGfaWWp02DblNCxpEvma
jFbOHR9TBwfRbv8eBHb36rDhrRt1Iz3SJbYPRjGRM/PU9uPWJE+5YBSKRqKZk58xjP97iU57riiM
fF9bWdEsZfwnmIK06WHoVhOmtVSPmH7kXORGaWg7hCK4qSvFgNcZuG7w/HuCkFkoUjI8w27JvXII
oESEjKJ3zUg+HxTHmxs93HBgmSx/R2yhaJelIYgGjVBnFmO2kEFvTMnUH8HBfMxCKaQpcccezCP/
IsgpN5xp4pk6JMFILi+0OOJmhJrSAs8UXEW3isxkB8weAQSYeh3SDdnL9B+x2lydicIwsTCiC8AI
wch214UDTej3EEUZfAesMHwYxYKg79gW5cB9+NcZmJsfmVEK27ty1h6C5ME/jnK6D/U/ypWFSdDa
GYxvumCUPFcwJFl1A8nonx2SnaI+7MBlEPSwXLnbCzhfnV0LtKy9BJbMPm9Y33sYI4teLBDhb9do
7QFid7Y+HeEXArk7g1wo6DWjtncYrzbr9iB2XaYMQTurgfMYxPPsu2J+dFEMl9wtSkap90s9qppy
WylMSOPBTk8fSsNmsE0p+3a3ZJpBYT+r+OfrGmtavuYoQ2gJ5xbUOX0pk8rmizJSZ4p5/zmyfo9x
DVK42OOEnYsui1e0lImTw4P2K0Qp4/DBq3rGwqr2U9eA2f62DPcE7TQR/m/VY77pujwaR/JIXkvu
qlDfeJuVwB3GoiyUql3e74fBzCed0UL+ToJcGSPXFunf6yrLZI40VYUo350F685/ye27S2myhj8m
tQRkQ7H7dOvqPQGsjPrBem54IdAllCbmDahjqR9An81VUkvlIVnIYbySb8X5yuvv8rpuVWEyt7Tu
SRDy/ddfP4Ad+PuxIQ6FeLu5aBzCDtV4Q+jOAVLa9PzNRWgyxPWHo6dnvYtXdZ/qKarAe3edB+t9
dK8z4JH1o2oD/Di25A5UHl1Fn7F7ZkU27VOcOK/Z2juv5d4HmbvR+k+gbw2L1ayetuqrqW7KbMK/
iYlQGOTiPYkDZgNcI/vjxdMOpZlX/HzXMn7UOWDPZIGLdBrIdN9ieECPStsUOmb0+ZRrNg7kNOVR
JK4hpXCF8N9BUQ8+HUHGSgN4DxJ1O2ywzl3pOxzInrxXETBfxP0cfDsC1CQs+meFsLMo9CaklZDl
KEO188hcQu5iFkplIoPhgqrXKs0oAsPG2hq2rZZJhPVLopHkclyGL73HtUYtFjl6u4tjh5VLJaUR
TRQ+XLJmdLeMvXq+8SPOttp651+aCvinvnXxPy1b4SHCb+bUYedHO6aE+HeHe0Hzez6BbMfBt/pe
4vKXkOghhocMSZkr4bsmF2WiIgrtfCQeIfpZIezaUM6AgTwCDxPf7IJBfshyxM03Hf8ZrWJXayyv
SfnqEnr3wlvegFtexaoMHf8ek/q4i32+Cm/JNLEXtOQ2P8zaBLzenqBBHC/qy0bpKrj/FaskXX9T
qZrFnBHMLHXdU8xyKiQDydQXZIyoQbwgwUstlw6LKdBIkAWobwxMAekX3QRCnrerxJOpRuyelPQR
mSSfOqXnHdfSDWDjYl+7koVGXpoyoFpltJvVZJIJZastZmi+QDL9vGb9oiA2GvO45M/tKhNqSQhZ
m6YwYP4UT92vqiDsU+dc4g/j8MeJWqPUZKCupUVGF1OJ3g7GeMVfOKaGJIHWnc1PXWjtnKuLTw/l
HOo9SucozetyjiNkEEamr7bZtIN3exHGe9Dire3A6eyTXaf3RAxMzusX1O5ZZpxpdFqjhUQk3tEf
Ls1iKT3KFO2EYilpKkrIdsbwkrs9UXKC3CkbDY46m/tK4vIjwUE7c7cU4UxeDHc51ntfA1T6dHos
3U7ELSVogal+casJT6I7sVPSQ1oDRNHStJ9tjs59Ctu6zGT233hA3HKsIZ6G2S62KN/2Dsx3AeWp
qu+WBySceQ2G0c6mq+mKDK/c4+UErT+uXU4kBUUKo4YqzlMUvWJUPhiUrtmjRXJrkKY2su5tvNGA
AjYq8rvj9BsosKaQ299o+4MMtl8aWYHyoBc4/dbvz4Jm+QJqhLbvekQISzv9SwG6n6ImT9w+OLmG
l2UWTrz8DMMHIMJV2jL7WCoPZ6HtU5m0fcS3DpKxIuH4LEVU0AAdJk8WggHq2DSb6Q2omKrKANrr
iiblNpSg/Ec7za5E6MVwAKqLo0mg7dRK/dYZPc83Lhp8bnc7q4a/7lpyPPdqGo9auL+uWCuqCaar
CmDiEwnwMDr5MvV9zVNC17wDT8LHgK/1TQyswf31FEjasFS5p59J4XGomytwJCuoZ3dfUZGh9lEu
53Ke6wLXgQmvkSzrVkZT5XqZIX8Rf76fqtMBcDg8XJ244jRT6fVleCQ9xOA3TWts1aA66W5/01BL
0MOFAUPV4ZtMBRTSRNbF6bMxa8CA+cZZEls/w9KkAQXmI/q/wumi2mkR0jVAql32ruakJH+CA5pi
TL1OMJ77tJ4Bk4hdGDkG7hTu1jhI3Im2VJBc2Vh+z0n+5ui2g3wuWJxmiTADeKMEHkOdA9Gwcijz
cRN0fekg3evIVnsfSp/iMh/951xXMbi3AbpwwA8R+Gjgp8AkMQRsXG7b4sMYMM0O8yOowQffRuHz
T67U8Zyp8+Ob/ES23hKPkyY14LtycBLOtxZtjH0w3no2jfNWvWewVDw74y3qQaIBpeEz+CdVexYK
w1OCn435RumqkQ/SovEQeP6bzE/JZhb1lzRZjzAlrq85k1IC139WcCo9NCrRk0mvF7OfiPhi2Kmm
c3yW1Hp732VQ5I96w9gdFLylIwp/dMh/UYrGBWUVVVjkjtJUKAinT1WzVTgQP/rXR0q9geeAKhL3
hs04+w8+kg1t25ytGfTBQQVuclNolSOwS3fDfkitBu6Jb8qRVMFfLQvEG9CZQfPP5gWSI01tBK6C
neHmysZUrjE31GjtBqvnQyHGAkaZz5k1zlnaxukQmazpu6mzoJz+z3/PmdVn/D8gIF0gaSJfcgtn
gynpfKWQwVrcIzOfLzIsxMBdjy+M9ob5c7ny6Y4Uf1DopRbEeb1PrmgSMRcwhqnJ9xKjzw/kPshT
JEaDDqaPITzCFWCMDsjcvHxBXEuz/LShXjYNe5eDs9qnHmebKG8YxJLX1u1fXBwz3lRPyPHTi69h
rbBp3Z6QPsgYUj9RARl5SlRVUUEdLIjhsl+HCBRI2UQVmdli3pc68lDyWz6fFZSfwbOf6RX1clPT
JAVmiryv/MSdY3aIkWpVAstQFo9SSbYb4R9ziJms+/cV/NKSZn4vyOmnKd7CR1xLAozOnHfpBt8j
3saG/FBqrchViIqC95/Kg98j8aqjHKrWnMjfeppxyMyAovzyGgsRMX8U6vh85svcbzLXGkmSN+57
aPGrdQYzkucwBAY7aJZiVqZBFNhJTN2XAu6fsU+cvPYA42eDw0aFzYVI3Fta4gjWNQWK5xamrxv2
mcZ97W+4hwEoSyBu36MaX4yP104nV9jRZfzN61HerWOlWdvbaVJK/2xfkFWp+8A0z0XhlgRg2NVa
47IGOccdf5ESh912dBGXWGEFjeQWX0Bpgd8BHgnTA+uVXYU7njC+QtSKnoOsq6TlUM07+sMNin9i
6EbLoVnBUK1v+df8v+PPEhaUteXHUr4H80Q4/Q71QxRHwS4OkP7Wj1i8rnTpRKIzXrYZHCUACQ6/
D/V8DNF80rK6BIiUsXALVHtvHZJzvfrv3BUlpBTAoGKCBQkbv3iUYjCenKMcwG24Vi12xm6fM7EV
ocXQQqNUeOhaH6JU5qC2K1bnJL7rbj+rN3tJ1vQE5eh3xhaE5D4orApmsnu0bg6Qo59RNiLdo4NA
0S/JWH/M00sYhyjv4OpW9tY+dHVVDFgKbAf5yfFlj/5KLhDINoq1Rnz51LMtvvbOk4qtX4mVNzGb
kPQab7YucASuhpcW9NKRjsnX7LJi6dplCOytdrWkbjyL5Pa1fsoDmgtaArDa7Biy3HtvsuvcQImm
htnSPq0sgR10hJl2C6RiboFMtFlL+kOaS8j3LeApfb9dYdh9DAEwZEY+KxSvMAcIpD1XwqNx816C
sov64K50GmzXPhmsrd86/z9uOZPpHvc6XHHPueV40tRRwPaSCMXdIEgU79NdP5SKQIhR4il856jz
Rv1hW3s3GKxxZuJ390MIJ58tHGO2y9Dy44e4MoZ0ziybZUzfdurX4SX2bxqTIBrZ3maoamqPsrM7
IS0I5xtxD+XmnsghcjTOCP6N8QxV2bH5kGhA8cPNNln1peWuaxHJ/ixN02F72GT4dDEkE1HfYuTu
gwDZ2Mwh9ZISm7SyTX+RSRHEssWjrGgGZqY1A1tzGkp4e/SMOdiqT4OM+SAobNgfZPwk1MPqUswl
+PU0p2XK66xK7bg7FAtk3i36WRrCf3vhl7uE/qt8q31tCM+CWbns+xOZPHwkPfKCtbCoZOch2gZ0
WYtZeFn1hngnVqtYdu+nn67xzuOvmhGZ39QPGe6D30xIQlU4T/K4BdEpxm3xN8Vd1FuJl/bfKiaP
TDfKggkOSE1a/Xm3Bg7DatrQgMYMsmjbkV1bBwszGJfgmCBRH5T91Ezqt9K3XGSwxp+zvTvuxRzo
O/zqY+kbWAkfJmD7G9px5ln9giuL/MqS2NzQ6FqxgVstWHH0k+PRdL0SrYDVksygeSop3NyOCOcG
e2gW+hOg1YaUjzzbpHqUlNet2tmWQy0jJSQX0XjslhdX06MvxquZ/s5kPBl99Z9QykYtOCFQ5Czn
vFyO/2SmYG+MTYp68yfFLCBhJsTDIP4uXtICx8at41W6CEAiybDYYJN4DhWvek7qgQiwOHhWxZTQ
4jnNsiyJkkWtK1BTKj6iTRxPWYdnuNKvAP8RMeMXlZHZKGMjXtGOBKBMqNO6nYc5xAVAOmckck9f
gqckzdDg7LsvM/KKVzQ/h+W9rIUFkZ3ENuUdnlVxyOP1oupxbkLU2Hw6HPnADjFk/akasMQeNRnF
xuBIGSFSJaXB59tw1Xfju6+Qv0U+geCmXPgSmrrAvo/skr9Ze2vqhdAZuAignmNH/3LZQ1qWQG2w
C0Yd0gZxQjRh6eQnFIXlre5x4KAukYBgaO4Tedo7scfhovqlaPVqRlM9UABjLWmCtaxD96ojRVt4
HIzcsmcgDUAH+1HUtDLvS7KEMIyiv81D1b68GCZkm33NqazTdjObG/4LDYnjJvZ4SXHko5fazgHA
ueomEwDapOFE9yyoE1StzI9UECG0EV9n/ezatk88KitGzaP70eM4fLDMXQmf+IVxitJY8x7Gcm32
6vWJl+Jr7/YEVN/kLkWFFKuMRx72XI+5Sszl6K0y+wVF4t6FSo2c2Ydx8naKZhSK64Y2X4MiOrqQ
b53UN89RFHzesoJHxp19MtCSW6q4Fq+ftGCNivqQ/U6Mjc7ZcxuOR6PssnB6BqnBLB6wj87g7/8p
tkUuUhUzWsEOT6Wnz+b1z8U7wHa5jLyjLGqKYuS7bvveJiZBvxdIvqoA72zIBmsRPXJoDJ2k/IRw
Nw7Wqh1VlzztaRu5DnYiRHgNfaSZPPC6VVWJZz63IpwKHEMm91Wev4KZUssb3OeXpqvY08sMWA3S
82NPY+kxpmhq+y/W1/sO5LsM8eGzZjRX94T0N4EvclXJEkqN912HZU0lnTxxsI8tlnWendEFVbVl
Wq8ieIltAr3yYUfpD0lIPxYcYxf/MHfSiqPg70sL7mF45NQ9CTE0oc4j2+8oeV7j8n/l3U33cZsn
5sJDA4BkHguKCP7Y5E/MjH/d0BVrZCXBHQdeBseDRu+nOUT9AHytMMHSL3fC9PjVb+HX0CxX43z+
wKXyOU0uNFScw0fblljmOxOZvrXdUmn+TV5NWXOtW3/R4iPmhUtL07zfmE37QQCy/kQuOIXVx1a2
U03wCseWtOChyFpa/i7PdtTKKR0See+xNFiqvOjXQIcmBIup2EMF1Awa/1pnLuOllmi4nn+vOn+s
GnMoJARsHN8OQqyoN7Luk8MmMvBDQV0+jEMD3fC5NRwQnWvVMHk6XnwXMfr/WIFaaGqkgGfNEa9k
dt9ZxCgJDt5tPd8OIV1FzgmL9YqBjDulCsuGQHVTU53tWBIWqSp7y0lTHkxqOTK2yXdcUmyKwGq7
YzX7kNuvYqGLsIvmnLE671Ds4AHgRYb+vRP9BTkpruFwZXybjzCUIv2RpgC7iWiyU4gM+a5ZGUB/
9lXvprbjZiDTzjFKfBW96hBQLmRyaVBW15CVNYrs+WGB3zw3vCISks6Wx35XLrsM6u9TA9cwpihV
FUQEPjOtNvewP9CeNa5DXGQ9EI1OBHiUv8g4G2zfMgov9aXgedoheCQDq8RILGp6eOGe1aVXv0rY
H/YB1Lr6LBwPcje379T3Xi/AYhim/SwWzgildOVY514kjEp5Meq/+nzUdMQHRJBeW63TfkARzici
PF3NykbMewm2DpGJcXgVV73kwQv/VlUkjkw3gNyjAprzW5sRCKTLnOpRKHcGXHjoffAwfxViG7C4
T7tmBeDWyN+sLC/WdH72ESqlvPMR5f+m7imiBbUS8vU2e/2+OAWeOTjK48SDqCbxAqXTjj2eSWgF
/NaFRGOZVVozvounIyyh07wQ3nqa0i2sNIOSPazOovp1UFSnLZPiYSAjvQtZlm69yDgKgoKq+mij
OieJn1ITe3S0DLLe8xAw7ftZpeRRlH0Gi0KN74orwmozOFRgUNo8FjMryDtejbw9HvyFQQJgm6PF
XGJ6B0u2xPOU/uRByZA3UlNb0CQ2IqRi4I87bUnKA0J0ItC45gRezQETgv1N436v06Lkv7p79MtG
iZ0mOOm59MYGQeCA5N6fh9WrYsshzG1mGiiBwJZrieIZQV7k60KNdh3rRT30SdWRpMC4QZoqE3HL
ttQVinxVKlFxGLOAQ1+McfsghpB6WBz5nHxyjmk9GaDp7CkmxbaXeYngABE2NHb1pjXVWFV2u9N0
kEO78GYvklW4vAOyV3px52gahRJ783fxa3jiOL3X6vXpxtpy6V3u7cMuJEgKd6roOcLqYE983W0V
JQv1v8r+iUuUbjuWxaqEv2Mtf0JbjWYG5OBV8myO85ZZapXThUGNYYQ31tQ6EXnxpXT9Ht/5o9EU
vMhA5n2fqiUXto7m/Gdgm3hbb8l6jtP0uOvi4Ui2twXfgpFGTT8xR7pSrSU/gNgDyRxi3gMKXRdq
eRCG1l35eMiYlfNIQDt74pnGeRSapO0zSK3imH/oKmgmUOYMO5+CXwkDHXtA9ZcfFYp0Z7R3XWj3
kcboHZz5gNpYRk0r7lvUlGTwz/cpgLxpsGYhA0SZVIrywdilWwDJ095NxnKwmxtIFWXIFuRMJESo
Pg1156J9dDFKvDVWpgiEwYZg+M91LJ3flPBnyVa8HcBx0I6qsY2WFsLfH0b9MTKwraQ2Wzl1vjkC
Vxx5ilUt/i07YU4sE6PKUVFO7F78dNnbqS8qpSEAsA3vVZihC18HmNsbuaCiXehFQKOY5njMZaiZ
KfV581x3V7GlQc9/sAdVBPmvyxCWo2tCrPnZ3uFXnohT4pDSJSSVAADk9FmWzLybIKi2H1prsJng
n0uVeVE+nKUPdOzYQLu2thEZ7CcmBSc7An3gY3jJR6cMNq4/9ohOGGGrFmjFr1Ksvq758sft0Qso
FkwuwFf9ao4z8a3Q2PivRSwAyYylBHoGdUZdbAP36iDo0OsRBuZ+ktr0Buu7UjCFh7wQJxvUkyAd
UV+t7VElyvcS3NWYG9fg4P7oRreqUV8pfvP+pA8jJlYPHhwRH7md05jvm5o++MJZcGasSoIodF/G
KOGshaCJ8jLzUQiNrhRfA0pb/NBHFFacJRg4pSIDKy70nOnIsvKw7y+BQAH0i8q6JKknrgr3OBf4
KcTypmCjm9PH0WIpVmlTKEaHLKzS8bIqFv2lV1f+/3FiKAUZrR76jtSci9+fzvw5LGSNDlsIfWdL
Nr2DRlnB0vm0TCLgZxRh5MneO2GLYpiHnd1c7NDTAsf2cczj4P0cp5OvNGXHoCJTKXOQlMJ9GeQ+
bPw/uhefP46FMGTSu1jDRCSQUYUc536kstHfmyG7Ororh0g6bVzB8vIloP9err7ZjI5y3JnkpPJz
MPs/tCbapGXxhpayXdF1K/82wEqzCDZ0wWiaTMUkRS6FARSeyC+WIQZXC9i0SYhdy2vnLA7+bNJs
2Ibd+tYnnJHpO0MrxSS4c5ivODEUnlYE55Ty5qA/E0Zhh28AC5O4aflpqpoQWU87oDbzScyXRjDl
NuKquyzlpfH/g9NhCYqyMUAjddnIPs4Ld6mKVxsGbdf+EqYGXU37gyVw52anFQNklGtG031+2Uc1
L1V2pyQRDQ8/lU+tCyWW1bUGjb6ESlF0Pp2K/WeyVoUbKBPZ/TpAL1JiC+XUuaqaTEIlqGCYlLWm
nbYZT0y1pA+wVjiteqZ60crLK15BkFc99MIZ9rsyeEbog2poX/3FYMUHrYHlse2ilkmA6ROZnj3Q
zJtCxLFM3WCOWGxEGRfKbYCnnyl9Z3UQgtHPu7pjza0LTLWrYHjhZ5qOw+IZku1bosh3SLBVlef1
noMpTrmrd7QHYGhg6PrUwlkyI9C1l9ALeFaGqIad0KbnjRleDAdeqDlKKbS8blWx57cPGoBXwAnG
7RmteL0RdcIFiM1yNrnKoHYEPbZjTAJ3kcYAPra9t+1q9k7j/UusWuYdPXLJE1TIAgpwWrdN+kpK
YBvZzKfy+gPZkb7s52Bh0PSsxkAFTf5nyeYEVxst5n68wolqp5qgNjZqCiPMn0A3lkL2XafsFoq7
o2ENTfo27gUyMPXGxz0YoozLmyEso+ZFn9hhNs0mbxQHMFDlY5YB9bSjwPDugU24XfpaD2pc0xfm
cxVkt3IRwxq0ojnlslHKHNKevnakr3IYKvziTTyGJz5o3rQszDWnwqiep6FUHc+efBXYrAafMLbU
v9wNfrTZFfwZ8X+yme3ztQ25VJT+c7pkvvYBaVv2RJOMBBXH7vqwmc1vW0gom+1FgA9C0lNFJrNB
8zTimBta+mnChEo9619bAZuVr9ilcAkh0cIJSkl8reUo96oSWNBm6ogqJjPpoKWa+C6C+PouZbUE
HQuwyZqN1qW14nTDP1v+SOgldpYL5FVnu1wOGGfwgQRXy3wpOrOGIQDF+zpdg0rLWUEn7HbxMR/K
b8qGi/+dRktw+RGClU0NL8V4ZzLK/Pbxt8mmIM3Awtza/B76NnEumiHp2ZrM6Zig+I+1IdJF3SAj
wtF5+CdprlHvS0JHB29TCo83wYsGLgjjZl9e6kCu/ElhIWJSBB/r8l/FpY4zpSZcsgDbcDJUTyXo
JG1x+7eCWvV3u8WWtqMgvPgUxBnyyfDJCZoip7xYf/FBAzajVYFBKhDizEXVC22doJ850+h8Ueu9
tK9COT3HYX42eTXw0HsZyLTBevjiZVPnQvxLVlQ2LHKKCqMYrAIbf4iPzhJwYThjwhKsQKABb5lJ
kWsK1UJPFN05NubCX9kx5hv2yMW7buFlPG/O8I0W0UYfwsjiLUZXK1Jjtr7KSMTL/2wfkWUozNAp
0/yFAVddnDeDLwC/0Vuwkkx0lK6rHHV6mf5mrxIfrb618Hn3qq3wxxRbY7rDgX4SyjVKLj1K+eBy
auZxcTo/451Tnd5fsUc+NeKxG10yKlmOmp2JrMESOmYQFAM+6qgRRLXjjYDv51HLvLgugN6URa6n
11H544tORA06jhFar7O40SewH9bAOMljxV/zPOUnVQep5LLVj7z9tMKV99A1k5LeysYCmX49pF+q
SfqzkezPKlfg8Y9rHNUA5FZFNuSOUqNo88gUH7Qi5TqMwm9V6xtza4G+zNbpRyIMsL8UZsWhs77N
1fRsnGgW2Pope1nA4yJ6zSv80pY5wOKsCtDNGyh6bLkDResZjOEkPm6QwpC/GA7so3gNqIuT91s+
zWDDdTYfHY07Tj2rcHFrsLGJ+WWc4sfpX4wVzXsB1oEQHflL9z3c5taHWrj5+5cyNGjptit72y3m
GgWFHCkuCLkP3HTYq2QeibBabF6Gu3rZbDwE0M1pSfWkBC4AvGlaYclQY6kEjJQVTkaAV1+AuhHR
b1rP6MOfG3UP1QoqeAxNso7/lN8bQPBYadXL/8+RVmt+RMpoPJ0FQl4NSgeOO0o56xNbG7T0smv2
e79AScy3ys+lOh/Btb/YOrCAmA+CTwWd+bzF+r8ko8liUlJRnZ5m3Mdi1q5ENLDKJ7a2wfZdxXfg
nopKH5LZhAN6HjyXpH5ngdXJ3bmv9gVJrmPUe3w3vWZ8odZI2aZbfdA6yE3ashdt4Cwums9+QNB3
uzzfnIODq5+GR8EitO0tur2w49eSB56R/SwpSRnhmjzniBdMiGG/EhPH33o3NM1UMTGF4obrXByR
EVGxzbHgQkzer8nPnX3xpEwXDNrRxJEMappFNJludqT306uCmNfBMxvgiKcyDu0pqFpSST2EDvRR
KqUZQm0IRQvw3nSIhDl5tBh1KNs32nQUwyMRbbYr8sl8Ka0HF+mEQ38HQ5K2DeIqQfTsDuHuBzF5
fBYaIlpzHMh0a8CzQvUp7EMfelUrS7hnSTzbaNAoCocgId+pabyx9U94IdElKY8c3U6POtIorWQy
YvIu1VHfMwYyh6gFaf2gjibB5N+fWC5RRMSC0Q1UbuOROOGe/OCCF9J7x4lThb3vvz+67AIIruuK
Uh1HmdDD4O0dtgDifmnz0WdWTjaJhxRBd/HPOiEyJYeRU8oC60NC8B4kIoE21MeLO04VJr8czmi6
O8PWqOczfpQ5RXLAPNHM2AQIHrVGveeZYmkZVW6UQRe4epcZk+r6h0IHX1Hj5V5xCuIccseYSmRl
0iPbIDXQKUpmeIongI5S7++LNJBceB6WU+Rz5v/pHPppKdpJh8ap/NfpwsgGvRc5OD+Dd6zrKw0H
x2uKve/bJ8AkfWUb73FkAxe03ueIYGKUOhHOmNMhUbBit3veM+MHB7bmhZkqudIG6pMa8daJzeqR
2iw/uoz0S2DubCp3B6uhOaZc5YUzMffuoGRW1+JrLTQO0GKQdm3VxiX9+fdRphUjCfaRWaa7WJpQ
krfWwEKiSIGqk+VkuBp8O9b/2ViaLwGMQZ0BInHX0C/GsfNy6ICZ0Spw7I8xRu++GKhl5krW5i1g
TI5tAvIlJ59ShrlnKMXlQPWQqz07GmSHb3gIAmiUuT6vXlet9ynSYYoA8urnX4vcs+ylEH72nhEi
XTjgM7BKziDY+DBN4zu30EzVNqQu/SOvd0jVyEE8nW9phaVXpSSS3I6joGBx9e9562z7K1sBVxg/
o0J+lPvefvrzjrZmKCmEx48Vc38pVYQspj378uw6ro+nXPlpEkX3A9JYZ2JtRxdmVMflurC+rO0T
+AkFRVbqslowXOqA8AjnjfCudDY4LP9+de5ZpG2x08WhKtnbdtTAkb1Cd/MSjwPYQ88yeeSDiDCH
eB1SNLvDHfhcjbW2mjEfdHlFXG85U3xFSCBE0ZyFU+jbcQ9WROCcTKI7Bu4aTvgm1XEbvePKOorP
pKri6XDJulNtsQfjs9TX/Vf79Yerv8PcyCaUYD/IT5rMMBxgsd/abZnmQMZYZHKyt16oa74SfMVY
aiIvwVHRFEo7P2+b+6mXqZTDKz3i/ulyh9xur6D6qn2gwxRfWniosXUYet0jS0+D+MI3KkKILLN1
bJk3/LqMIpBpq5x/bMREOzuERJe45Oz5T5mWuwx/fVNTEKvZEjuRz00qJIceg3FMJtlYzmLpp8zF
BPRhIMY0CVTfwxJiI/zCV1oln4RdvuJsNtoZQQStqUFkxTs+0jyWAZo2ZzRSs+hg4fSEEj0Q0U1v
4sxJsgLQ1brPX3NF8HalUojuWZbKCL7sLkwZaoAkYEpb0y5ZT/C2HEy7lyPO/WeWosik0AXqqSJK
Z3xxtJYg6QaxT9lNIGEPyNVk4mCgyiYilHo++1Fqtmn2lRvmgUJ0gyO8HVvu7ugQL3HQYHOKh5Hl
th9BDIa1G6fkc2qCSEcVy6g7Xq4wkqmjWx+0JNBoSkbupd1nibOfNn4Nm/uwXr3E2XKjaX1UAnfX
IBe6BVT9eCbRX1M+5e7bwA8NyAgfO8b9ViCmr3K0qC0/nnvusUpAv00CyNsaRE3o/mPz4mECegAr
aeWjHWYJ1NnqCtM3Ewe3mRX6hPWxjt1u09Em0RKA5so+xFXjs54OHI8qY85w4hyf7UPY5TfJ9BT8
YwCTTVW2eH3KuvJ5wyoPrbY7XZ6gpDFdKPJoVqHIXHhWyFhDZo+MzPfM0RKh5Exd1+tmQmTfjbNR
K4UGvPSfdizdQNTPjaXn6WJKQZyO93+SdG1pZWM2ki+gPoQqeWHGigR/Sygs1urEwp2vRMteiLw6
v7tG4nyoyPAoONzSTltuGceOvqKSnQOmD4E+3A+dCBUDHcLn2KWZFMFKecdUnDQQbX2fNhDGKyRe
kjQ8kGNwMaPaPXw8lnKphfzb4dl0XjgZ+uC0CvMECLGwAORfEl+b/d9pFiab7f9ekrQwpT7c1CrU
1UTRqYi1nY0S5E00zEPmE55SX1Ud/Fy17JbMjVYZ5mArhRamkXPmWvUKSmhGR4vYWmsSqfEiKJB5
5ajdmeCmcNFKDAqqmCEuimvqqSmZvJgKXaexe++adczSoljyUf+GVFGSG4FsfNz/oWKknRV2fd+D
VeGd0pJ+8b1H43In6roNTL2WHoAuhhTrmjPwW+ENhyJx6jfxgRirbaBRsueU+ImgVW7i6ZFuDfPf
mM90qS/ITB+41cyyVtQwaxQ62vPXooyBKez2OEgn2SQyNhVOtnqFOW2qm1tQCyMfx8R1NYgLvT6q
kaTLTTndrcLGLvhdpD4HIcPS22t7W8IwBQX5FsTqqXA0mGf33dSsNqwObojPKYTAQqjLWejDl+N0
xPYSmONRhpc6zEReKA+xLN634+SC0Qvz7YCNCfiiQpu9zrpAdwarbaRLyEJHc0bIZ3xu5IxceVY9
7Y1BdXrUg+OLIAVihEI8t0GPQ6EJ7A7CrpbuSCseMDbTDbdDU3p1ry93OlpXNUMf4glG8Jn9Rg/Z
MjVX1W6GCq1VzIfc21fNNeGrwbqyNaMyBXgvfmx5UaKFMNNmefE/aDGgGVfkhlfXF95HG+a1/a2E
CQoeI+QngFY4IRhfv8e64ak8s4wt4CtHGVVbN1QYIOX25NyL5VvZk921go40jqm4UmADfSSZqMQC
3ITYGkPJynk9LDA2iVISfkaaT3CxavJRUokYqpGb4ud0d5IQyfEc/dl/kPkaFjja9mNzqg+UjOU6
/0+o/R17OLUmi/IkmJZQSnUD4sXxrau8WJGZfSe1V5Q7tC1Czy/gQEUuVI1uofiT4RgMrpo0wRxt
BZ0sGhszUPDEgBnHUjVzRN3knIAjKHJzLTc4oQKLsSONzrMAhjQ17aMu1m2XnzesaEQCRmA9jbfK
APYnN08t3sUwLw3Ryb9Sg2TV6/eirKwT7QB3v1UXfANKi2pTiRv+Wv4jJxAH7kDOTgUk/9ZyHtvl
gR9ArAnjCjUltUqvy7dkxz+2U2EvN4tFiNQyCoVC+lfLLzwWjCKxCcnbFy1i6fEoPqsMsNOOvhTX
lMy7sU3P8lY75k+r1TnX4os0oZ4f9X3yI3D0wGpo7vU+gy4b2L06YtCyxIQzPNqPoNeSYra/rouA
XYGABiE0/W3aQlvn5gVjRpNn8MwzMFwRw58EX86XsW3rkClwMQnmgq87YmzYnKcv6XxI7BkGCxKf
ZUGhPk+Yqfj5hoaZCSh3OOAml5Ws1EPj7KmzA8j9GzzMRo+8k9iDdN3H/uUu1DVWEGzSSdnv5pKO
OVGJqDGjQ74h5WzZDoR042riZp/74Y9iTfpPfHPrZrgtIFFwGwk/4lG8V9QS0A+HTZhSRrnMXhXh
Ml30m3FdAn1xC7f6F4ecLDK/DyrIqpKs++PckNHE0VRoW14kIyN4H2DVsTx6WMEB/AfxxxYPYjGB
5Oh/VEsSUBIOZYvKm2L3otFQnV5fI9dBknD5xncqZcfBuzT0vz3DhUA/GY4mRO1QdpgrQQnUQZTy
YC927rP22OwDcWEYi/nznk6Kuqrq/tTXK0KYt4c5ho7rU9cqmjo/MsV8xl80OZvqqrQFlUal33Zx
3/GJFhgDidX1YrLLjAJIxcdYMnVSdXGO8m1KNJqD7wETjrJhF8XWLdoZMgS/Z8J1rZLJ0BN6l9Q3
jyRk7S1qkTvUNk6Y7ywxsWBV85U3zQtl9nogsfcD3LcOEq6zkApBHuW6sM8zLYwEwv3vGlvxIDl0
y9x9u8vGI2gAbqnII9e7VPq+He6x6OxrhTshFDRNZ397XHl5YHrqIi8nFxyApOmRnAhNMxMIX7PQ
ybxtDJ1uSOBDz8RFHAVzuvMRPoqBB4PdrB6HzNrZZzYJ70kthTFpdhyJmVNjaE/BmLpZrDmh/1HA
e7MnNgvDBeqFjiG/yfg7rMZjbp86oAPFJ4D47GMUVbgnsmZpig9Ov2CTwa3ch+OXDhqSRxgucBFC
LaCY6D+d5/kWJBP0XZu8NCCnUOZ96lHFR6i9odzWn8UVQSO3Wg8ZTTu0r3fJCd7xd2GLh1F6QKOR
p3k6QmE+Z6bH8FYguOC9VNyxsAKMtcZLVyoMNm2mq5C0kXeGhp+MtonzX2aXCQbYiT42XNv+bkzr
KBO8GSHWlczoi7ItL3AHkcVgFGfsNNy2HzLrrrZy73Jual9eqi2gd5KfRKXsthvNtRc4VqF5KG+G
e0MQyFR+IIxITB7/8EkGWsmTfU4bcd4DPKocqhoweknZChwVsRwj91Iy1q3tBKCvg5A+4p4r9FNw
TMz5t/WHfHa8lRbMYfXhRdKOp+V3eU8jCVgQFyWr6eQ2JxUeVCqo6fSLZqDV0FK/vIiBNFVhKUOq
+W8boTR4KGJI9FisCphOS73AihZmxslPhBUBKzUHV6HKMJcVtWaaotDECMz++DjwQOzL39ATpkaH
iYCkigFMZORyJwi+pk5EWeTPxWbQfAed6y69fRXny0iEF2sE0ZWWgWbp3GCTvAAKVJZwRNKUi5vo
L3HDbM3UBrSVz72G1EYCwMblmm00vQS6hyjx0ag6PH8Cv6HrehJcBnb/MEPVUINcXKkp0bmctwV7
bsmOWoo7uVrUNGTA29iZa9BilzOsfhCwly9oHkh+x2b2oaOJquUzYesgNH32bLg9rLeWLeqdEozh
GbozQ4hvVMBxYGsdtxQdP+wci/8OatIUwMiz1T9oZC5SmPWeYPoMY/lwDXLnhNdrKRN/Ge6zgpBi
87AKx5gaemBH1Rq7eXbJ8wY0bUAI5doUTse0xLQrVPbLaY7DsKXxR8vhijQ6zEMt/oM5UiZEnNTJ
xF6/6PRH2pddMwrvC3BOnzbfQwQ3IAg6CygGmkyRFY+6FY91n9JNIYi1xFD90YtiB/1cZcYjMxys
mj1f1OWBNJSxYrUI2qeI+T7NtoSZdOlhECauMOuPvGVIBVQk+bavZMfz3EPUoAfTiyUyh6CVpIzi
P++ETIOdaYA3pQIAXUZkPd76em6DMFz6/QsKMSjbsoAno8MEBvQSMNnDvXXZnESarWY7aQtq0Rz4
Xd8cf7TNN89oxOB2Ft1D30p9O4DIGhTJ2G9GW+1wjzNPygW30yhlnwJCUqs3ixH4kqLdfags5t0e
PfNu1Cl9gIj9XrWsuwG0u2UWx+xBl65N5voLwxdbDy3qpxt7Ro2AfRZkKkPGTY6YzP4QcCVQ4R4Z
qsC5nlxzR1gIpvqFrufA25m1607F7Yg7ivWsOKKYqmDqcZOw3kKj6l1LgJvdMVypzFD+blxz+RIT
1mHOrIPARm7YL/0pFNgP/jclmi+XiI1ROkz3IRRpw7nlRVvwBsIim9QSLbw2ircbU9Wv+F6p6pxt
s3Wj/pprAWHyiwFLhtJhVbEKgibsmtyyVkEkJd13VKdtPYHw/BUfamOn4lSACjc0jaZl6UOMtiZ4
YO0aHiR6twQpbuRDmocigNm8Oce3WgrJDoCWEGh3rsx4m384pvA4UGpfQQapAMDLWqx764mErBv5
u3xGv8x567t7F1KV5XUvlSoSF8E4E6DK/v9p+I+YB0fRL/5ryu6tmlYsQW/Gb9DBMgyQIMKnd3rL
uc2uXm8j9yYYCfWU02ONTzyTcwJBwmIYXrqjkawj5JtITQm9dNd6vW1WJulxlgfWwgInE8F0REjz
xCePWQvaMcq/zRNk82XnrJPs+fgGIr6A0u+b4DYZaKyTXsfe9itDT5YoLyXr+Zs4nNbIsNk42g12
s4aIpj7UMqBKaDilGI4QevA0rxX0g5sTrG60cKHst25hqV70IhaLXM9dYwSMQqG85mEwkRv4ZFxZ
VCswv91Ig6llVWOWul7Uzt/BeQfKA2N4KFWRdAn42TNcOj8mzKen2LwuGhA6BbKou2zQPDnUy3fA
QuzfhSiKnx3b0ZpJPRhGft4+LWoR2aE0NI4+LOA0CezLZQanW0X8+CdFIHo0Eqg/VjPt7daGMHFe
NdlsyUXifFb6S6ChCHKfeulrfyrVIPBvxeQ7jxGshheBKluDzLPzL4e59es/fqTBhGjl3Wmwyixh
8FC4zi6JFflstxHoS9kmnBYtYD1WS5oI023PxOQ8lW0i+cbvUlQZDA1i/GzWDAc/V8+XD4sk8RId
WQPXM1+suS8SHe1qM7UilRP0oqdGdJ4X7n9V8D5FUFFC25zqB+wYzcIfkGRUD4jGdtuPElhMgtqQ
PgaRo0aMj+OOhaMExWtZeDCznkj2zIFlx/4RGBKV9Ln3E+K7kF4fHk3SOzcgbja26IpD6+Pj26lU
RAasesX533Rek9gsiiiNQi00AyCa9nQk6yz/+ZOQnX+jdXpDjFiKk5Bx5g/+oeOjONy72u61dmib
TggQoVS5RbAXnOuajJVUEOEEx7oegFVKKFxfCPDBUc49LVRm0aQ30GX0uwgoZEljm9kJHVEvb9I9
3kxXWbl3LUyK0yw5skpM/G/lOWVKdsTodKlgVsDY02mzPKJAdMJEvGn3s/pWsKItCX2I1yPnp3Wl
GNv8L1kBVb8FvujDythb24aU5Oc3K/0TXpGcKNhMRe8RS2TU5fBqKWtYsengyBMUyd4GA9e0+kVP
SsCvtpJrjshS6aWTUUvjfG5rXCvgCBXUyn6MRX2hQFmKIdqcZktw0A3EI5TmTCSxSXnemnx/Vv4u
s9qyjiLWoRjvmOXgfmLP/pImIJa/J2C6onSPgO+SjH4Oov0mT+E2yo3XGOCFx2GrpH/tX+FKX0x2
/cjf4oPZOZ3CQX9CU2XY4VXMZ8i3bQxNunXvOmdxf9Agi0MK1l90w2lw2Wvio+ax6XcozKM0qxUz
IvL3nudgL3PuTzrEeBXU1uLx0YuMVK4hoDVcqaJxIO2ItLdywbouK+pCSJ1/6MKT82L2KaRmxxhB
+rpLLTY3Q8xb/3yqlcTOgCVX9Y6WHkZ9rdCNLtMgLLzU7snPq1N7i3YQHoDBywbptrzm6F6uMHKA
txLj7bFNSuASrLCU47l1cmrS6EDT8ANz78hgkB77/4OwizyzdyS1OntwYBgwqSVzIpbTd46+2rWS
h6caLUs7+4iQ5fBLTVjr166EqPL+u5PrKFf47GnbJfMdtKBbec3hLDuVQ2hOuGsZQRtcSDY6aCEs
z3nPmMs1phV5ighMhz2Y7PF4CIfjOOrGOhV8jy1Qmc+lq/yosXPYFY+H6zgBhuIkpsj+CJvARGZI
QkWG4ZSnHsA+bvNOkH2pLlF0ypBLFl0jSN7F9mYed2uWdqgQJIFCDzeorVcMkRmbt7csyzu2C2AP
HsgzodwmkPpOUhZAmEWOKwwxcIBz+oKVP1miwEvJ/7+DZ+94p5UhL2Q+LFpibnxksVZ2YOUbvro7
zECqxuF+8iANlqNWV8c2n7q5pLbPrYok5xkwHhfFoAhelVXvbQHPOQy1V9qV8SL4OHJIg4pYCr4m
VCrfFseiVaQ0stmkZlya4Ls+r8RhDGLB4qvgD6lVB8ToBdA7ualZzcU3eNpjc3FWvEXm2SK5oQws
g4avPC4RE6OKEcNAHTb2qkTT3t0lTIJJ4veiOTgRaWl+tO1iEdE+hq+MSRLiy/hh53eGRpIC4TD7
7+Yp2ti5ZquU1riiY6bTlC70PASgEo/ipsoZawyE9OlyBXxo+6T4UBkpvFctWks6nh+Izpda9FpB
UuddSyJzFHJYH6OUv/2YUsW8glYl3652XzktLEwkYjdzJrrCOXv61OuMXR3iW9I37m7rdBF9MSQm
vPEN5z/WF2j6wbwTAVvG6enxYuRBOnVJ2aGakvpgZ2CghDjwHIISEFHPwK096mu4ssdhQISBtqpv
3MyTdDT6h9tu3hMkJkCpcJUbslWFQmXR1wh1HGCilYQlNMoIxT3O2YgJK3yL+I6rYtcVff83mWag
RPknPPI5sp8L8d/tBMGruWUzZS6WGY460Q2ZK6TfWWF/smQpzPdVL+vLGT4fTj+vAJ8dovBzb0o2
TLqsTtdMJmBZjf8HWVsA3CogyHp7Fbx+IG/BL1vFW8MWNpzZV20ouCRGh4bMQatxaSYYKrgNzTcB
1+qMH6ibG4C0fZTKGAyDfGgSq2hWkm3Pe1cf/TeEBCkgW3g+kkS7i3BBAYT24K5Q0+k6JCkbkHDf
ss7dx06EunSeeJHUdGCWdxZrMDAwBHWpguezSLhBPkkxWvbRx22EvBdBJk5ZZP/kGgQe7LXOHU+U
KI6BbS29gNDRo7vyQMkesAdosmMEOYd/8aLspqFA2o1afSaquQYB9zcqkA5Q2mNIOZlDQSIG0ZPI
RzMQNbuA3ZoMgS2JQUa8ESSAijqBH6t+jHc1LCAWehFCtSzcCxp7inYMBGyJCHmK4/2o22fq4zHA
saEg/hHHzax6iTwl3XX572d/ViWKMXo4vZv62bsowh8rRZs9M527PrS62fHGx9P32IbmXBsxfaEs
Ee9emkRtT04+ibpN2CYIVRq5RICzHQqb1PXX3WJfnFBMNMqXF5ANNa4lULdmQDx9QIdv7p3L2J3M
pEJIKOcyeNKE8zDzMQQHW3uaOQ8XMWPzdyb5N/bXn+RcAhQ8NNPoHJwJ6a29SfQK50zH2hDXyYmQ
I4zrQRHrNcB3R34MIpv3HiU3oO89+0fw5gehn40gr27epLag+gGTAFqdnIGBzPeP2/qPQFY2O5rd
IYqZjWCA+ZaRZSjmMYEcOIFZ4EqrZ5AkWSF1NL+yNy3mMCVnrPJ0rxG5xharUEOS+ytvCykbM8MK
72da6kqcwo16Lbn052OMT5V2vw/iKAULTcm4dcdgB3TndJdQHLFk4QK53MXq76/qBsjWDZ6e97e5
/QjSxotHO3nbQQRMKi/4reSr1OlduEDQ/XhsLiiZNIbbnq49RL+EpTou/Wol+ULSeflEhhcN9rFO
tDdSQ09W322f84CZuANDjMqiSv/fPuFeEK+d6unsWqZ41vB+iOzNeZ5jVrT89xdJt2he5mcF6jMm
7xiCTHIlXlXZ4udqIlt0kHC7SVEUCEKZV2Po/CR7jXmGxM1UFq4DAgJYT53WjH6T9jg5APWQbaVM
sbuegjmcEkRDs3sC1QG0A6zyz/ZUNkFxanx5cmuER/qPzHKjtlOzT5+CMglgWgJPzlWo/1Ou1YHB
EumRS+qBXewtLeDVI1vejMoTE4/cig+UMEOCOXJmqgbOkmpU5tZae3VT6G5xylls0IvzZ5+MtEVP
9yh5IZWPHcllzPqpnQFr/uHbNaR1/fLpYWbIsrEoHXlUrA1fIPosJjUU2bzu1UnyBlMp9iB8PUwZ
ekKnp+k+w9cRXUo3EL9wi8Z1UV7d/Q2iHh1LBmI0d1NADkfm7tXZlAuAWxGXi0r6Fy/TxBpWxM3F
jrf2MkAs7gWrGVAScppe3MGukyvCGdvzkQbvcGtr9Pasxfyt6NOjCmy1JdKOn1uqyd0ioYgJ21Q1
e2hUanJPw+4HJgrf5gJ4DB6ISvkRAe7W9KOqZdDKheeOJu3r1JJe8AbOLOrBDnRPidXXtwK2zyqm
G+3B0VpQk+du+70tvmzStFWhl0/M3R3XfTSz8Rz4Dgf6AiloA9qaDF8yIbF9l8255WNksTYiN49Z
kfKkvRbNYPwvh7BUjBBj6vzs5v2gfBGzEgNIyEHgXWyT/jVfbqeFQG0TtDtyZGMWwAe1JC6XEn/G
0ftW2uW1l8eQ289knymwxOZwHr7zcwIm3J6YNb4yiM/P1UTm0Pg8XuC35huW3TpfHDDlWWmaUTgz
5eRQWiVe87/9dqyptyPZTWE+r16abt4HMdbnfOcdfMb4xq1Qn6ZHVAmX2n3o4elc7N68wsfB0I33
HtgH10TGJ/r5UcEelc+LBVF6VXJ7fAMwjPd2wMVucjN9TX0wVGrdtzlfs6zUQbvIpIv3HwYKeuhe
91o+Avkpj2cjrgFzGIEdA3qaXmq67CU8AG1undxIf2Q1UhSH2Ef31hRXmAwxL3pIKCNHaGZNaqks
/lPvta00RjO7S5Sd5dqSJyB9ZSMQiWHZw/sfw2gqoO67eS2AArSJXj10xl4E/bkvPpJhDSYDjgLz
lssIC4eVW2O6+jXTKTB5jg1z2RvWRWnQnUIIajJpMAObuN14Fde8CZ6o7s/7Zki+J+QYSiXztLvk
ZPWitjh/e7wzfR8bTlA51Ph0Kp+1fozdwTatLk0bAi3PGWX1pwi4e8pFgZ7IDVKrhlKwYlOXQyx2
TB0lvW1uf3hkxHuCMDsmi8bEOwgqH+0DLfeeS1ocE1ogJbsDtaBH9qlhpCOBz6kXoAPRFaXwPi8u
R4uva4bvkZp0j6QAQd5lu9peWmchOSkmdCF4A8pl6VblbzpgxDBYFkFnuGZYm7JNYac1vN6J7n3A
uw0CTSHCRBZh/u7ZcG5KSb/hIxXyNEZ7Iz8knL9SfrWR3i/EdC0Ald6ocVJjg3ou83o40/r88FBm
YuBhhHAQyMrNOeQKFFokcrJd86tyD9pcegJqDOEckKqQ03C40HuDH2+AvJNeY/+D93+ZF/mWxg5F
ogN/1NOWH37GSM7mjrrL+33ysG7efB4jnXrn0mnZxEVVduo4V+tK4AEm8vs/k55cOROs/OpggoyR
8CDuCFh/NNqVD/bZhIHv1c3k+T2+76Vh2dZjTJoXMN5VzJhA4RF+RsQA24KRLU5MWdt2f7r80dgc
GTu6araXtvLuUa+qPmO+2Mo2pMllseikMFO5qrrqdGtjtkifQuM6bOt6ZJHncOpE7Hla45cxOKQx
k7CfoB9FGZCImNWWPWC9QrBpArQMuEtEiXPjN4muUwzM2fDYM24p61FWWieWii9Pvj7LrsXmD6hK
bUnXE1XEhKk7zvx/yl6m+Z0rVM9gefVu9ccH7MBLe6VMtEidaVUKT8UWL3tbIr1c7OBIK9WBPKzA
MbL7Y5DkOlfSCnRepiB6b/7x/+ioKFXvN+sijy8SBA0W/zESIqnnoWkMeMTHpZLGWl5L8dNJWMP4
MSGD2vajKcGyesZFdfT2z27RlMRyTXWudi9WEEqDgvB/khxIn5ffeRHIbTjCLesWu16+ETNdXzWc
doUrbmatw7400zUdZ9LQy2QXdMuQVXvy/RjrPvFmUyG5h6q1D0ejaRkO4GogM6sNh5TPwUwBwpaU
ZOBYq31htnOMaVpJi54TcfBGOV9GchM0Xc6aF546YQ5QhljrjKh4szAGatuBH6M1r3Br9UdN4vMz
VCg+lqqyvSwxMVWyBplA2advvuuUmlTYKlR9xlm2PZzjdM9/Up8LLMA4CndEGwpH2pfnDvDJqWSB
uYr2uyhm3+zUSOXZG5tkvayY3lhVKgUFQJNVEE0i9Zv6fegpBz5jytaLFyT2mk4MNtM3ts9iAMBX
dPq7DbZCknXl+4PckNAqU0l+H1KO1gmmJO5LJxKxZRToXuljF/Zj7FxQ+H87NF/OE2KGawBGZx4u
Xq5WmwcBOsJc+EUHmANxTxgcFBuCfBVm/yOCg3rCGHd6srQFJpuksI4Cfc4T8hnJCnvJWYeB3BgB
OAaqRPcXnVbEla+wl8UO0g04Q83NMLKmlpA06/u3xVQw7sitxuh0xnyuiPWK7YH4nyBpolqAYzdC
uIoPh/jpkQlWqdeBpddG0SRJtEt8fZfMXdIXa18CAIbPRpHmCmxu7vr0X6u7c1YG+EJ5JSzMaoc+
VAdIc+wXHIqm3uHf89jjI9TCNQpzWRNCj/FL9xBxn4J/UK2oDeAh77XrBmbKGEzTM/wcGKW2Qv79
URVOwBmfNeZxiD21Cu9yLUCKBHbHziXaD6vxi+jLUpgQEwIQRV7Cw8kzfu5XhI5BirYdUxTo9Q2/
WgE7t5PNPog/4qZ0pS1T0e7b/ybhU3hyI27JiyCOHmggD26stizt6Dk/XLyFVHYat5Uexru1U5su
PwBbqvc9dH3cpLDWqtL9hUvwFQ23Mu6T0z9n2ppS+cU2TWYEfoM4pvXlkzUA4nLg6N+kcD6QSa24
x2gxu1oTTp4zPjgBMN5pQz3RyQmXFNY3SX8AosoZQjuc/3SxuRgxIEuVVZsWCUsvZjg7oCtcHcCn
7mFhZgO3+uB9UhkK+X4YvR+CKpBBGp4EXFYf+gZCrmNUyYul8HAIGnJGSykHkLSuVdvkSqnqcJ6M
yWr46JUyMWyVjZvC0jCiBEOmPFgRJfCEKIvlrDce5cqqgVdkgMHhmXoZNhhAKdOUbDIUb1HjmF+2
PHOzPMCYUyn3orsDqNQss/buIOj3O9pH54fE2C4uRMC1f4VXTRquxKSBZkEgn6SOHbfZOHGCLA3Y
tCO8zDha/F1KX19NPY0k355FYh3yWXRgzoN9Me4cQnJdlIHtZF34CDoJ6aAidvSsnLnu1uz7pjSO
MBSBL+GZ4otngyoo1psTiod5uaBzhw5X5VuVI7+l74Inw+OsKd0zfdKxRqyT0Y4XfDEpsJb9AqDE
gT/JZRnF7XWMFMgUDwnSzYyklJmhvH7h2R49dTGB5xaLC0pih1lLFs9Tus7p6ajqGMjGTQTgkNMU
5d6Uo7vSFQ2e5xd5+L1q9tWw4RuqPQeAuCdHu4gL2uUqUgORQWVtIlY3+DuSl0EL1EheOKs7kDDh
v+AsZLmEdSQMd7C0er27OdeRJyMKLgUyJeMQxE25yPiXTTcAHJ/7jfKd9wCwoZZove2nmRp+g6ir
SiQ+CaCkAyxBvYUwI5wd17QXpzi1ZF2lVA2WlJ3yE6pK4b6VXKlxy9oZWUm9BUH1Iu9maNwjPuSg
qkR1xL/P+0O89tx0IoLGJOjQ9G5Oy2zdfV2al/DxFR15jImN/GGxL9iU+ALtjtxft1b0GKb7xzbE
VsCL93k5ZsRjNxLpLprOeE3Q5ztXuVtax5EoWqRaEK8oEYo9Jv8AMsxNI8hn23b0lbrpBHU39m31
lcjeYGVKLWtUGEddEnSiX+9zbI1ufjeyhQvkFFSlNegjDrIWyT+wjuM27lTBNaNm0n5cmo0FR80x
DULe/z8ofkLRxd8fIswP6bsjVe4nU2KYUez7zPUZ7cYDtBi/vKH8hD4Y9HHUm7JHqmLZQ5t+OPyD
DlPEsKC1ffYm8uoiaYxRL+SH1DyS4NTtuIPmNafPgPdgr2Rn58wrfScWpS+DXLZIU1mqJViNutWp
kkcGyrMXO4u8/arZmRTABbcc00a7e8ca5ny6o1RvkEfzLIS2lHOzLS5G8/JC7vptKqrC47is/Cvg
m9ampQbcrWG/lhSNb3fFQNUONTLi+74AOGZFhCrf1fkWORZBAmnJp78SQVV+waR4mfD/SzUZ+m4c
d//7Gj3S8RiPsM5y2+nFDju7zcp+OJQs1Zn+Bf7AKzrIQXSEUmifDe/D7twZ72y4GWUoI7nDqmmM
9y8Tn8JLmjPbBjmVnbFjoTBeQmyy5Fy64L/bAcUX4f9UQ4m3iS/xIJbl0fDsEFt1YgU5fehbJERg
h0Adusngu9gTVqzdsuewvrSLOs9+Y1cpM9HxBsMrszJmI8YKEjjpkcSM75FqJ7+pAl74CxxVO+E3
/tevEQRNvWJ9uQWQgmhtFRnHWaWTIigfBj4g0o0jGBekR1cZp+v9TgTTtJJaag2sbdut3D+U/crJ
t8bxJup3y2vqNrBzUoYww0pZFyUURz7xMp2pS/3PdqWYvlzT2rOkSUHletmhEytSSvi7hTCB5xjJ
rspazlLysvNKCAaSAZmBIVCLy8dZNentLdPBoPE4wNqEr9XByd2NkFUP1a38W0nvk1GNtfW3ubFp
DIFLCoeEm7YhaU0Obdg71fnM9WJl1z5P5DLXf+4Ic/aaFVmyHMP8f2lZQSrjw3pgfMcBiDpbkVtK
6DIOwh66Lvlv+MorIaEmjVB8f32KcyQgnJ17pDvgnIVPaV76fIXrVTL/siBq/DPWOTUf8PUXMjsp
8yCEALSaBcmxClm/e2lUhjnV1wiFPSUZmADd47YconPRopnUImPTeHtQJMx4GttDM3la0iFiBr6Y
8jwpiC0CY7wbLl1VTyp9q4BiVX4EeK0D/lvV/UDYcoUfvaATdunWBQMZVjR/Ux8oZCJk/xoKmLDZ
lFBT64ADyol7udJNjPpGG8wuxp8ahajvyO2gvupSPMJGsBaApeyWxayqSW/mq7wfgSNOduK5kDdj
FoZhfguWV4/DExVy6sTRV7jDZX3Yk763TOQddGnbIIrPddjrI2STiJNfZ2hYKZzCToStu4gPAzBP
ZABXl4/2sYabWQGA/BbStl/SgfmSeNMh9YYSC75FGOoHort/yerJXPA7XQZ3csjRctaiFEAs53yr
dgZIpkBGkJny9HgdXH31zUd/S2a9EBeZTU5QdbB1oLAg4EI/E2vuhxvGMYOVAJIsCYiz+T7ONvyb
QpGD10iLKqw+/PdWOk36oykWQVt1tKuYwEnQ5K/8DJY9uO9PxOGJwzMDXStevDqSoveNmkZvYV+b
fTd0W3XyFev+bFxPkyx54bz6TCprnSsmFqc7sJzT/Sh2o3L8tFmpJxrjexBtrfd6IuqtcLSd7mzB
kINJtGNjF8QplU0j3YsCP0LwRaOlRyzPQLarAoeMuAQyDNXIr0SVCfa5yDXZzJGashfzvTrCcECW
2DKgHBF8l9s2qqdnVyWYxGhMSkLYZEFWj9iF7Rjbj56XfVwDDh8UGveM7nZWPx9jJvfFg1sU5iYS
eCI8RMb07eW8YQ5silgqqqXDVn4UcuMEn3Cwxwz4EJDGD5QL/ggYa7blkhDXTqj+SFgYrHBM1vPl
hJC/PIFZ7eX83kEd+KhCU4NRc+gjaTJjKbioE2jWbVs/2apePvG6f4CCJspeu0steWdCQQLLUier
vETFrKEZ+BxsL/duuWYdDd6+ZfDIZPfRT9UkEmpfTHxsoHjXn3F5dT4vIh3Vyqr5fF6cm3K7V8Qo
6ZasQ06RP+03YLsXeALLsBAxLmcTNjHakR0gjhN0G3ShQIHemjk0jU+QoZBrtXerXQZxodZdLrn3
YJuDrOKAvQENiUqqkmGNaJ1OV6aSZb9oVoWKQTRZb/T6nnI00LX3Qh5rM98ICyGPp56Nvz2tU/T0
xTA6txTAY8xlfvw/B6uLPOJxg1EFHLUmW2x5g985lH4ClmxKGmgNN33lvaohfSJIvxeO3lv+3mTn
PRyWptk6G8UvE5uPPpHS2Dk1D2srC/jBZkJmYlxk8rcal26BaO1cJ8/ROoYghswW1bzzlO2qeGpM
iqGq5vzx2MH8xce319BxcdxD7ictJ0SCQbGp2bCobiWaCulAkgd+1psKw3sD1Ljde7l3g1nFKJQ6
1eh722VTBjcYDnEaj3WF8QznWd8pZavVP6LfqmIskw4fVs7VYGowWaE6Z5GJ6BH21RdSbnCb3M3Q
uSQ/0Vj+d0Y54ILCOYvRbjERyAYTBYyH0fz5HsTuJi93d4lRTrAaDa5SpKbGzj1iv1Nu4vKOfWt/
g5bs/dXVJ5iqCoUsyTbLfMQ2PooJGYJl0t9ZZMV3m86VrQraVO3VWpkv5Cu9rW0mNfFdj6NkI3uB
JXdrCnLiPUzoWi99Q8rkcewu6FyF19S9+zkfeOGXjFpeQbLzV7AooqYapdAa0R1rHldEIb9sYuHQ
VVl3JLLIbD4DYBXpqR4I8I4fXfw/qDvi+muDEhKc68sy6WZW2ErJYfR6BfOCOa5OLMM4PbCQsVJK
F/LDIDNZ79fX6zTj3JXFwxuV4w0UcNgQEnZFJRQ1FMbWLS8r6Z4ZolAdiJcIO0dygHN466jBLAru
OuSrS7srVgNh6WggpYfsDpKU7wvAoI2PX7q4fDc3EL7xFKV/YNzaSQ9xCibduLCjU1fNPyK5bqic
OaeF2uXKnUkLqDda1a2bWwYBuZ0Swc5YLNbBo5xz2o9Z0ExpPdiPyshrhWXYzlusYRvy6wfCP4VP
ASAKKtRKjsEU2AdZMSRYOVTfgqo4LadHY/H97zZGeI1dzJ4u88nas9D1qoo/BDFBsgCYn9JlE+45
01ThfT+Fps4ncykgpRfvZYEE9ygdA2njgn3hnM36d/4v8yxDOoYCvKrjYmM1BJPvmCNCWoQs/0ve
x+GaSEyGa84lC91sQtLkpR0Uo97j0R8xhYvS4KIeATEb7aDrgV2MvRU4rERSGLlKRiF0xMI9bcdx
wQ77/q9pLh1ce493FIoemjXtsiYPbt6V194vK8M17nlrBBLEl9Sd+/rQCtPxLIkmGnnM4qUbdJf7
6kF6NlOSWxr0zjdOqJug4oH/bQBBpxTKHZnHyV25vraGh4EY2if+Yk9UwBucZWTNmWnFr7FjfFbT
axGpOX9tPRqTV/8g5gGzbUmO9/+BaU36mZib3E5MTPNG0AcZFjm4pNU30wfZR0iqlcyPOm6QfslR
g4qBQy4Ddu863ukICHMTlTbXSG35KSnV4JQVb9i5OvmRF2ehBt/QEF5R48VjUG/Wb6z4s+xSG1Bu
3OR+0Hx8Mqh3oVQvWOuwLCefMIK3QXxV27AIyyZT+vSZ5IN5CpN0zCdR93m6Ww6zY1LXLmInPSKo
CDUyiMQZS0BFTT2+03v6qv2P5xba8djLPUETRblV0E/OeqTkoVFnptIr0f9CijwckDUUMYfwcGn9
d9l+STBqgiQ3owhDXJoqBUZkpz8pazthnH82ZKnIlVAZIixlUoLU64pdCl59UF/0QVpmN7fD0KwU
XcAt7U6qLZY5cwXRLQ5jIVf4543/ZmAAyM3wAUtONnhwAUAU4Ub160g2/z4kgUXEW3brSpiS0p+6
7pntjF2LZIO8LyawDcN6kt0dpEA9yKR8fmyESzk73weuxgQ4FTAnmKj3/huPn5fBcIyLzF18OuPX
7QxqYMrbH2BMZssyCLxyS3Pm3TY+5sz7VgtxSvLTlWBH90AQSdclJO8orcsGdXDNEVG8boJ7O8nO
rVBxzhdX1X/WzzyYgepmwkSoJEIOKyDfVikopgchKSI4jblIw4nS8hyt9qn8yqiVrF7aBD8w7aXg
aZQzrNkxVaZDHxfrDr+RtgEnCCfvCI9XCyE7/k+5GvIVDfSDeiVW3odtdbAlE3YcJ4VxVvt3nU83
33Ama1Ka2pa3e4NmctrORN5VN/1BbherKsuk5w7/EkJnQA91POFmGqeSLcgrlZQG43JyGS46WG8l
6+eKkSKZjFHKUxyCFT1CYkDzenMy1aL3K+j7Y184dsQqarcDCU1VQTYlA6/gS7UYyWfVPPZgALH4
BZozusidTYTgjdT0zayyLa8lrjplwkvvBaKBsNWTRga51nAr+b4tMQA5RcGtvMx9uN5tFT0P1VNf
c30gFvf8x0BDNQC5EA6l11Dnbx/7VaEaTUQkBJHuOmPTPwg+MjDoxRY1v5s9NQRT+RGh2/7nYlJr
wS/rX2SRYnE0D1jb5jCgJUP2G0kQ0nCn8pmuYvBrcLuCKBxUNA4YeMcFZjaiBM6TUALK0Iv9WF2A
34dzej3GlRLpiR6rv3GUehUbAEbUIdYlY6zpGs92wwAHkJ27dxit1D9mWomfeL3PovRf2clI3zRa
NbSDtsnT6P7orAHPuRzk34k+QVvN4S4Hpzm8074D2qJK82E/GB2lbiJnjXhrfSvfCmO8OOvbseE2
MRFtnmL0ReAJH2F0Shwzhsk7uT6iZufv7Y8UFCieA4tmITELsfkbozFx0jpqfv9nuYMiOF2naQek
KuZ3jXt34CSy9xTdwjBX6Vj64oxjfcLQOVhzUqolqPtC+9u2/crzcMrpFHTNROKAP5LA2nORDyFf
A1styTwIg2PujJVBkOr7jbebljDIUPQxg4NQxvzY6Hbcy+zY+8bRkcgoZj/3uweE5T8IU99w1jpJ
7Su9a/Ta244vsJq60VoIeDoOye6oW8jY1YXQxnmXQOWjpx9FL5+Mx1fVqgDwWKoRqmMGxkwMM2xq
EkzmSR1RXj0aVxY1iLL/NI7uvA+yXM1pvRfKQkmRQUOMxr3gqqJ+9zQ5SmjO/AZUePiD5U6NMM9m
JO4xXUsI1ajJfRh2XY0e60/3XORvleKGqdsYhoAk0Qrn9gto7mdMvczJBlnPM+fQkdetEkj8cj8v
OOqBnk6GXzBxD+ESguk6uuky77unl505JkEd/c4U7/HJZyWaaG4cz9FUa9gTCTTG4NUPCsXY3Xya
Ikf5/zaZEWt/Qfbaodv5vsIw9cKi6JqtpURTmQTOpdmScl4816I7uPUHAYfudIb+9wEqla9qlI7H
K89E8GuvT9FQGlujH0hQqopiHV32IHHwhDvcyhdQze9yCrcdVi323sZuev1rNCuIkCxU39jdFMj6
9avQWjGcfmrWWObWu5VouRun+RSeKwyB5CpAQ4YoAIHsX6gG5ykBNPoO2GglFzvooHxnKxlcCCbT
amon/pq0GKVz1Chh0nIuxOcEwG8cyGYPC4C5Fg9V+m9Wf1zz2L+wBbPmdr7EjRxvTF6veeEXZlYH
HmW4ibiNFXXsvm04k7ox5f96XX/g2i6H6NIudPsLRNceBNAFcCgouv1HBs4kpwsetiO0rdUxsNoX
iZ/7ftlEDEl12LcAZHJXT2TR8Tbwxl7TiYAkuvwBRoXeKs00SfyZMIyzGD68dSnSmOisd4atBy3Y
GrY3w3rkQ1HAKgm37t/2pYCc6khDHbEUZtgKfjJiY2+vbV86tm1PW/Zzs5MwptGGvsiGqRIVaKdX
Vc6bZN3Mm8Nm0J5Nf6xAJNCU426r1wFE11+CLTow7NUDnApaF3OUoijDO163AkjPbMNqn6172Bxq
5pJr1+Rwmvseo+EH8lvSATgVxF5sb/xX7TsLd1KNdRlPQ1H0btB2J6r2G7kMkX7CerpERHZTYuy3
JRG+NMrEJLNhOrlCMvG6bIA5SIzR56uSbEykWLlZfd621x0sMo7Ss3Etx5Tnym8iwk+lC84GxJC3
Cb2UQrpnJXXvuJ/g9QLjryIhsbpR2Mk0h+Gn3KMXCJGyxRCIMRsi6p/XXfPBaOWqTABLjWxKAwe/
yWgEDwHdx0uwe/4oCdubXIvXFuWRECwwAKwKxr4uBlSimObmeXVw8L11lGWzfDa7TvKKoy/ejp9U
CaM9HJad8NZvF5fkQHJbHfVNWT8tbWHxLkMb5s6bmHyPvPrS66rAGc7aRt6MNd+SSMYA58WUn77F
8uCJ/TRpaoE0mPod6+VDS2+X+r40rej7+Cy9RJFAilt6CeqzvpfVNRLjFI9sXtVq/qDkE2MkSM57
ISdKEyxoNrIXDyGxUk1G1MZ3AVgKSzMgX5W3xG2Qu1+auNiN10JwBl6l57fh2oCCPkswTT9DZYJN
QYIA/wRs7mNpXN6cQQZKPJ8sGG5+LnOks0ZIKs3dXYMRojSpMYzvTlqz4ewCKjCrZNGVZqI4u0Ph
Ln7wphs83m/Y2Lz2pbsWMtu1TnPYG5TxtOTwz7duR0SnbnKirmhs5YhCHUZw5KIXOhUmcdFR6TJh
Mxq7tTBTzLGrNjmRF+cP15mEJ3OIHB/nPkz9yGW6R4fCEpeaO4TuaPWqfTC03OJYdb2A4TLHX4hO
QwvNxJ2LcPPYF//Bpvul7OQYtz19vROIK33iUtkifJDrGNhVATsJ8ijCaMabcKvChR726zXreHNJ
CTbHBmsvj6LO9nFSXYYHx5l2q0gucMWma2XPRxYJyuk1xb/CM14JL/MmoKWL0RVpwrlR8SmAg6R7
BjO0Ks/X4fVQ6GaV6QfGAED5vxO8vtdvyv3Jm9m9b72gjYiucLvi0+GY4PFgEMD/LNWwnvtQMqaT
/GzmwD4DIty0+R4Z9UKInXdKFvfVobRtHJCsGXMPnbdB47vJ9ny5KTBKSBYDvaxKkebdUIoRrgFW
X0uUfu8tzoVksx7f2jkey4uEbVAm/AstZnHl55cKk4cygSF5urr0bMdum/F2u8VVeLCYqQwXrsxx
IHu4J7GS3YsGzqr702DjGYsm//AbAwfaU3qP4ukl5gESbT7VsLWtMeh1xYylTAxUcbvQtEpykk6F
HmKpAVbEz9/a8O5laY6RxPf8Uk2kED71SsJWe5qV2P5ihScpd/ZBkry+/ecNGCTdaBLVvaxdu8Bv
GaP0UO6SSZ+FlVcw8ULKYfWwREj98h8cl5FEX2JVshQSg6SHYCdGT967/WJqo8h2MYCtLoIRhLqy
OuKyG68OK+zrmengpZyLPGe4GcDIk2P3pgF4SNujZykbfGfkA8a63z8M/WvRiUiPp4bJOK/yO12C
ep/neR5WW3IP3XlnzoWiIPMllc6UbKthxOL2dstwE6/STlFIlPCwEGCxr2S5AwS6Ubo8IR9DRukE
oEkwLzbXxDnkAmLTJH0yIxvzbCvoA6We1682NKUWdYsnKWB4UzHc5zacMYKENa9r0s9HN5Mvgc6r
9Zaac9pHKF6pqHTbxqjnNPAo6eDZfyMRsUr+InrdiJOjf6zFyxx85xG7VQjGyyQcQvgij636DR0H
/yx2HNtVURkUTTkPazqSD4hn+L5wPVY0pR9yZfdgTPPD7Y/rtLOeDguMFinL496uZtsusY9ZCBjG
lX4B5GbhNFRgJBQ3wy7cA6B6BW6tJb5Bg7jUEQlIWNC5JpgXg39uxm73HkHEgXI+xbtH//+08UxI
dxIxX7tQXZjjALdOzft5dOpf9mLYvxc9XdpQOXqLpOxDM2oYoaIZgYFhKqhqoTC0N9Cpfl4lMgSa
ug/HUnmQRMgoFYeAkSEDEUNb8VAkTOjc1OyFpf6SJztTOIoopJ6gHctIC5PX1ssRDXXTzEjACL2C
1WiPnMhdK5bB7JPvQzd3suIy1/8eyNAS3HJCgphk+vxmWx1Xr78O9pcFIZiSlroX0tP8wb8D7BRl
WD19a/r58VjNxwq1W61fH1sJd7oQQq30TczdaCX7kZOBAbp+jmZwddbUIeRiS3rrUkhRJoRuktgi
Gm+rP2R5RaRFLtupl4ucIu5Ojn3prSypF8Ylrofcvs9Kk/LTdH2QgNgXjPdd6FoGOR32wHI6ogdT
aVYY3BXGu+/f6kNvw3GbaEjgkIHuWC3PZFii+GMlk4Wl6CS2A21sTMym44ZmBpy4CIHd4JLvjY8v
xkdpH9CsyDs2q58lS5W0bJIXRHYoY6M7w3KuirnysrjcwFMwLZIO7gKsRVOmB5q1gYLqWnvB3ZH8
9lWkTkktihq5g1nyePs5QpHAzM7oHKUvyH5hYz5cRB/hpUOEJyOjggSjyDIpksYIYtEQ0zBtpt3G
1bqkw4VZukgNA0dGi4bTyuvkLAx61V90JGC/qCXX1KbTOfbM4ltnclCZ7k9b1wCVVO0pSDTIUiGE
urf6dguAE0ZBhpAljxKsUgc12uSSaTPtzzQJPczje/pl4cHLAjI9jSe9GxbGdMMYc1qdIorZRzag
MOeJS89RuYFzfESlGwahOXp/gh1dRsJmLTXS5dAbK2uWmGfQYGqd9BNXX8dvYfbJn0fWFhHFmWR7
/Prnbv3Jks/ksO2t+8Qu9HKzPA1zyu+/r7BXO8q3dh5+UOUKdZ3dwdL4ltmkBFX9NU5Oleehr4BJ
C/li+HXyMfYbqf3WdloJ81kWrcsh9BqrInPt4mq+MtqAsaw7Z/Bx9w+EzSahS7IA7BSxw62mLUsK
EmGb3KFt0Hy37JcAMuHmvja2K/nqX58+vFYvmPdx4bCYgfKDfSZI5n6Wmqh2abWzmvMVNZ/rvlnf
Nr9qB1Ily5LtMktizPDRdj5da2UUACJdZM6nddmWNm1GOeK8bahl8DTXn57UTgCyeSlN8rxOy4mk
Lu6uo48aq0kJ1oW3uDVUV8s+2uV25XyGQBe2JtHwuV+eZZj5PBEIMFrK/u75J4CBGJXrmRxnV/cR
jsTgr6UPypmeZtc6Tnl3XLO4lN4peMRlMrxoXg0575nnMR+23qdOL/orfBkhJj/NPUgQ21fJD9yu
DRDeJcMujr7KhHyPNFneulCv4IP42ZIvvcTX4KBTW2PuScJ+tJ1cyEiNPiJC25k+BzfU6viKMFQt
smCdxLafs9D0pfiLTZlhNOg80IJxOkfCLUfeNbFH4+kmjyAc/IyAn7Dd5UqX1gcQynRDs1RRjh35
p9hvJeTIPGGAAF00qbOGElRLe7vHb43aj6fMruJ6yvP/3RugTQ4uG33dvme7otW3wLkDs2rXw7po
cTep6W+wxnmRVbu8pvabvfFdoAH1XKKXKHFSPPRORwUuwPYXcIB11R0iZF5aBLwf+yskHlY7vO3p
lkNfVdZD7JMzfkAX/lihkA+m1N+czEwUOPbHc83EHUVyq4C94lgWnqLb6+MeB4/C9QEfUhfOrsNf
W/5fKn4BWXKFK/US8kQojUTy90OF0WGUtdzWV0CWpTuI3xMSkIrR8HfBUW5xAGDSAifkFYki2RpY
Np6TOsNXxQo52MEcbX22UKHU2y7PYwwflRRsCEPhS0jpvAbimxqNqsG937zNgB+kscVs1veElIaB
7re/MRRncdZhYOlaLk7S5ZZyeyWbIvXl4LbVCQ4v182wSdDkPfW53ikQiIs6bnnBedSor5IY61m4
4PaYwt2GtA3sexKnH1YZDlBCAAiAptv09uYYLfcb7HLcKZNQN3ih2ifV3Xfd7ob8lXmdZLr3BrIi
h6BfK+RK9OWsBLhrZtaMVKgsaTpFehg1eJP/EWeQQI65sbjhhptiWjeoQfajYY9DR14w43luIkCf
sPP7PGVLvPUr9/gOk1I9ppFLhrf6t3mFuphoJTtXr4EwN9RvF0RP7jklGBV4gYD17Hh1Fx2lIDDw
bn3ralnQ0UPIekc75CP6n9xcidFfgsUg9L3eXiWvrBMbsOhqXWIa//aCV4zUhVpVB8LRsBx5in8g
+58Vu96a2sbQTUwUuG/VFRbW2gYKiT4JuKKSeGi2Fr1L1y3ot/7LcFH60uYcyC+SAxLDxHnkVW55
9u39wpe24Lw+LcZKH9mKmjI6yMhPk1FzZaCqnsFi6IyvQJCiOz+U59fy6YOVvSFfb4LE5UH9ONYl
NOJkHftXHt7DJ77ugOsM8FxdlWkrOzx6zaWCZc6thr71bURd6qUhH9LxDi3ea2My6Qj3rylm3Va+
iRGdmjwlKVhIv5OPSCxuOq6kQV9yZbDbnM/X2BBO7FByM8EPWqW6r6qpUmB0hIZ1Bl4ZQ1m/gw0J
PNcCbu0Suv4/QOlWrUHWTETWBNOYgNp4VyFPghMwYMQAYDjP7GgXTJ0rzdxMu+YV6S6XvcxLZWF2
kaz93iCCunFfZsHfPuOgUPJ6Yz1XmG3aP6PIcy/RR1Njp13oYURGUna0ant2mjuDt1QiFq+qjwXc
5pHvSiiLtxZdxoNjklXOO8YkzQDSGdb7/1guUhqdrSlMnghN8mPLflB3NqiLUc4mA64fm37YQ1U9
x0ELOUvi3gq6DJ4EvtwGf8SykpmbECszK0uzyPSEJ/Gm/vYwcN/T42TLXv4AC4dmrqdtRJrvs7BF
sTV8Dcpw5k7Y8wPp1zz+JVq+QVfklWPoOG6Y5CLYbciQuk5qpQNQx91v9XacB5wl1f/eSLW/Y8S+
S8vuLPEQD266olEemc2sTufLpmP3Fv5v0DEuGv9uyNAUwhmMXSfFPbd2SEN/MKK26c7MYY1xukkm
O3EU+PgQcFtPHvIt4ZoofPN5+47Dd341LDvAQge7+yLTZkAlg8LgeuU/Wc2x9gH3Qjbt/dLOb4Bj
cYpOY7IDM1gHea9ieo6rLygBmZPmRcelPpNoOmZEH29RRimmkOGEMguRX5cTR9uwCIclVoDdliJu
EBWHDUIRyk0oc7A6jdXHrF0cnrTpRPzcg/P1E+CP/qHLuimx/6RNNwf3g9Hai8hGQPNNMV0HSEaw
TMFpA990i74eT2NTQ+vM51CFCxmOr4Qm04lD6BUjKBWPldeL09W1f91MO2Pg6mUTpz4yt4jYQfpz
bSu19Ed1kt+QNJU6gm03s+2r8MZDfnuhh0rVU/fitdCUdE8NP6jMDbi1Ed4d644ZTypleyaLIKDF
WpPxk2oqG4Ua5W5yYeX5sFdEVbnoWN2pImGt1FbyH2Rc+YKH9xdl07xyv4TumStRhvFM2lS6qDAH
rJZq/WOT8twgwOZTXI0lRQESw7FcUxk4w5oIx/6xkSiP6Lh8b7ST6r2cn2MFlxrKWCvbmU+VjA3C
kBWWu6Ywf4hyzWL6ZajmwxA4pNk9VZvyOsfqt8Zc60xCtPgaCDjTRS4/a/Un1XNfffyEls5qsjjM
n7wSrzkMWKTlYi6+YgS/Wp28txZtcW+yo23MvemlwJatk7LGdCT4rBHYiKsa+uiLcnoYYTHGXIT4
R2BJarxtTMneQ+jcz5y3fsHVcFeM6oHuSwj3Yd1IB+EnWRRgjonwrd75swjHCp5NiBGx+MLp5IWK
A2D5s/KDQY9+Weq0MR/FknyQn+NNr1jhvbiHYnjfWvz0Kv1g2kqh2XbTZ1mdfBdRY9Fz3PW/dOGm
VGM56Y+5ISFl85h9yf/s55C1WShdo+5gUfxfnn+XAbuaU1HSW5jhnbQ4WJpv6pQtL06A5ElhXmc5
F1bvlq8K3eSLxSoeyyLG5e7cRV89BWGW6yhp9aAtr8Ge6PGKih/xs2OJZHHi/g+Q36eNMonTfoUF
2yhTa4ZZdicCeKDCjjYlMLDfEZePz5KgkxSlbj7PGAPMoQ8+PCso6HZOXQjZ9KXYjfDEnPL/YjkO
YSfiGwsqB8XnOb3qJCsAYrf/uw2JiOrUcRaTQvx/x4EPhd6Dce4/xXA/mxQX4U9tL5ralQqGAzQ/
h05z67elOSWecZ5f4VFx47qEPauPqBy/lBN8l/p/XvLCg1ogMnZRwBPtLRsID/B/ZCz0vqCYOZ/o
Me20fllaJw4hZyepHaQmXbT2SS/Fv3jpj6yal/sxxSTjELNeTP/VsmZ6au+jht+b45prKAAeaN/h
NECFoBE2kxFLoR3kU0yRaIx55ZRWxkZF3JWCdkIN1z2P8IcEyvzqS2VolD9A/88/e+60md/Wxg9X
S5zQH9nsQhKeeu2JwB+1EZO58w7fVlN5BUFu5isft98xkHK/TbkZka5len2kEWsuFZlHvAs7ejBh
01sWc0N6s5v25bn0uXE98MD1kAbC+B1gpu7mrgxiy8AQKF87hG3BtPOCT/sQHLHf3+XMgBtifZB9
i5AOYpvG6yvMRZvNl/i0Oe9V6GdVGi87QibEhvhpwKzEQYnq6+v3i9p902bMoC0GWekfd+mcyTkg
9xBvhVbQkHi08+NeZs6RJwBhN6HVJ9o/1l/lckRY28jYkJjBlOUH2n/5ke3mRsPbFQIT25B+2yIN
WeAqzj4Tflfi7VqOju7sdvfCiFP/Lg2J5kC22PnokccaidUGYOJm0usxBLYrAb68TK2wL4gTexuw
SweD4RmwchZHL7UHSF2gdfrTcwSxTtCS5NYb0Cg2zO2sm2SNXIGyDNpxA/k8d2HymvS3I39vmxQG
FyOyDPbnJ+t69r/3qPZvgukfEwRrGTJhzpkvOFiDcFywqGGxq8KPF0mMJITg+rLmGOd6agUSae8W
SSa23pngShARnvqbj5Oce+/zCYXS77t5D6n7TWZGk6vTvFn7VfCuquCsCW7lQxVq3Dq0g9JVFyK3
SKDne85L7aFw/mdQ8XLSjn4kn/B35T2mTMOKxINSPcayBl0f3WeTIB+l2Rk0tGGLSk/TYGhASpOj
0FyavaUwqouDrX/PhEApVx+TpP14TJGQCVMJGI6FVR+OFc9C5UQs2c60L5i4VVH+8bmzyOIsfTTP
5tc632tSxvQwYqkqDX9Z1HSRrNcrzVcTS/iPLszlSTt2IeRZFpywQvONUkvEMrUYWdx8hHvEO/Gp
UKdHKrWr69PWpGmPaXOp+Nq2K7EXmHG8aCNN+dhuHBedK2N3ldIQepdO3c09azdbn/0ggcbd4N6H
KVuGyCchl467XCWncbjBnEEtA8BwGV5OqP1bABVPcZZi0XRVmVWhUhfXzxa/ckSL2MzYtel+2NDI
DkUZjvqjVP0QCkx7rCLGRb58jwcU2yBBMuvbTlu72xZ8UCt4nfgh5QIaXbS/vADe+eRg/QwrUlKh
OVSeOWwRgElUop9Cn3cFWdOrZekz+ghBIhMMqXZQkvRBUZQ4XTosBGm3RnkjQDM26LasJtryrWAY
etabwsldj7+3Y5y+NSLavoAtltm2u9RB8Rckyy4F3y/xgWoWORngKgIQGTitR2QO/HXnonZgjmm0
vlHNyb3nthJha5tGi1xrNQNjFCb/N4GYdlTm5dgCDfKIIEcrxs7/0OF+6JHjkLAaVWCD1gHeCvIr
B8nEM51HvAn/wtbPx1Ax4gqLbTbjG5KcXC6a2xikS1vYpDRpprQvdJC7xmKhQ1XdU9OTSmzuEGWR
wwaqL7GAhUeFZdmvFlQkpP17z8PwGB2Gm3ktcRW99bYWwRiqnUywqLI8kG7wWe+UnmxGWmd9STdb
j3SuUMoP3sBVGwr3tUHu41cfcluyczuiAXgkSaj6/1unRJOuh+sWpCI5mLGqG+e217b94FmZiOk8
V91yV/rvMU7rKWE+cUxM7vljPDZwdMCqsZFmwyPEghIaze6jukchrxrWyIP9hCGEZJW6ijgMJrpW
sUF6/DMAm3eYhESvKq3W8wGNsQmmFxksVIOE/lxP/8ET9gAI/2K8h9Rea+HXjO4vIF0E9ZyuYQdd
6s+mIKAvoS5MSuw9DX8zQ5OmFPA/2VchjSuENyrgNoPdDemcnoppTfCDf3QKIMS/8GP048BQLz4o
IqMlEE2ARxXnaqUt4nvvdPjB/OVDCMdlfXKWN+1paEHJ9OJ0lVvEPPtPuwxVsvTGZEUdwBvcKmXX
TM7Iira9cw5CbNvnPBh+Bd9rYcrMmqTGOBFeYkijL25i1DzYRnHE5abeMNTslrJf0Zxd0Vg2Jr+G
+cE0Djl6+1TOPnzCsqAcG4K0JBAtnYVorRNTan3NhzyWfwLyMflb/JmZl7QWt8MnWeh4KHdm6EsA
47lvEc7dvefj9E0hTilKJbIeSnmRhojUF0By08q9d561xTrJ8I135wMhIbR+edEwG7CpD1M9vtdq
xFb2phW7xQtCmmgYC+0RBBKULwH7nzcCGEOisFAAR3RTl3lCxlZAMOOsTZnq0wpx6FOhG0rV6hto
xujwOZryQP+hbwINDl4emco6THEYi6jqxT4x0iDeQlbbdCpQ5DOfLLcbfk6objsvJoIrcV4Le/79
yqcbI97QVzRf3GcT4cVjTjYHwQC1NFjbzJ/VCccEaBywjJ4hU4wLyiwfdJFjiGZbLnr3ygWE0ixK
EgOHZjUWrEYUn+ZgzlnocP+/8q6Ikq0D1PIBBdtoZDHvwQICjeJM+VCuyA1aX0m3e25pqN6YLKTr
JYofoAX3U4I499dtvOzuzqONQ0ZFMNEtqAV6toJMwfpyeium9EX5VpPjFFs29cn4ttudf/0j8Uuv
bj1dbu595svrxbjKzuzIW/fJTLRpj6KO+Z8dHgZKg53F1LI+hfOjDO68q6bL8fAt6TeKFqRAAStn
ZS/7bWnI7qmbSaFE/XVvIMgGxBe3akpP2TUEI/YkAjruPksmdfdaXTWEiIpkf7pdWsjg1KNY6Omr
aq1JIK6BWh/UA/edDI1y+QbEQPEglW3/vRwaqYW9akMSe7uj9zTI+SZIu94j9ZwQmklTdvFfxqzH
wmq1a7HsOiyXcA75j3+dD5lMJ5FcTgBoaQn4QoNzUzH5CYmY820qkzwDAm1eEcXyefX1JBvzz1gW
ym8OHt3KcY8hCIOgKi3gPtMpjvI4rIWV0hGk4jKB0Cec2r+R9P+TMtaA8MMe4xlDK3uDHU4zYk5H
qTq4aBqpddgpOWtx5DjoJQNuymatauA06ftXhks2ulPTPmVNIcJPFCR1EgCCHWUvhqO27FTtJLdd
uZDR75xjXXa5juwNTGyJtWg99jM4Qfu5slGTp5P4slnP7YaLXTeYdXG4AlIDe+ibyALJ8Jo9hRAY
6bcaUrYrJLiobEEHSpf1sIpXr59ccd+Cg4Xoar55NTYykBdXENhhxCwb0RQNMBpKWDfzt3G7jttp
BX+DK9IXyuPP18cEsGEHdzMyoI/NK1LKwOVDvRpeVvClrGNIgwAWzhdeuLfyOD9mELK3xLvvdBOv
KXPB3Eh1KaGPe7yoRbHxmzj5ZsbE1SJg/W+oSA43eBTLKKi6ydS/yobnZ7q8ZnDVsRQu7dpD9zcW
ZAwzBIh6X5jEhg56CQXg9jmMllYV2O/+X3Q3pmG3jcKSNPPzXErCxssYPgaoJ9qm16VSUEafGKBT
7Cl9w1i2W416i8ymk8J2SvJ/sbp9P0c3vUrQj1AOk7pZyy+a81+7rLXkyn4A3DtjjfORK/BEOWJd
ub0MflPg/wcpML/m/eCBas6r6oZGvzY6X6nFyaBMJNgP9akSswhOTswHqb+gOWPLcanNisfJ+QF/
s+jZjkaoSHAZH0FH7zx2q0ktsGX94NaUHwBcPwgDRdwldv/tYd3whpe5wthitfdGd5XrWg0L1YvN
IDX/zQksnHQvSZfRcfiHVCnqg8XL05PzCrGmrHMKeHfEE9PkBntDVamHUyCBfRWjDo8O66bN50bc
059F87asPLagk5szyMpULE99Oc5yED8YOlhWT/J9T9Sd5pdxsDpw2wSEK49bXax79jN3sd62FJMS
hc5iWxaK8GC0mTsnX/ceZ/opMFrnbfAEuU1mWNEIPyk1qTQsjf9v12bOb85mb7AIu9q0JXwFof4/
J98ZNWGEKzCC79Iwn5Fca1bnkoh4LKlTnwO8Hgd4GN2sJnxJvMqe24ALiq9ol9QPCMGyGM7T7cuD
KDCyEoq5MjkucJGYT9Egpw6a8ufgbDOEpg6PxZDQGGcbZ2GlaaQN4rXI0lrv4v8Z5Oz3mcOmrb71
z41g7go1K+Q2rNXKGgiKNsvFPjCnzXKaEmyR264fD51sRdsn0GWyqOAeuFTzWuYX3OhWoXAL46Hi
cdKr8oao1BtM5h671mzm7NotAPQdacFX401L3isNAR0orf148Td6pVjgsuqlfWn8WWo2pN55cEy1
waePjdWpWEi8BipGAmIyLZfNiS1dr9aHTdMbjgNhyUq9B6WLTo9HcWyXDPayROpYG++5inNj+YdH
HYl4jreq0qHH+RfQAnYbMHEpeQ0ZtGPQWz3pyj//Am7p2pJlEUjMJW4Ykh5qI2x+qqFeLFKGMi0/
uKYAyloC9Ixc1WWed6bfloNXCF26YijMkWD+mm68AXESMoUeZ2T/c8uXIysGmSPGfvZeZkeyusUJ
+Sv2y3uk6oG0cvw5dTPB9pXdZun8jiyqbxUPmORr7/KKeooNo3LfrSJM1oiFPjT4vcD9IqR9kR4N
iA3hPJnBB2fKYsdpcQxKaqQvhB6vyBlIJEh1PhztTg6mwAE2ijKcZgXwU21tpJoZQECtdeNJ2Vys
2CQNtYB7vmVxaX9xFHmD788Klvoy6E2QUfy+Lvfr5G9CQYaSzfmnEqWARWuM1zEDiN0H86WOu6jC
m1RUAXXRdD/PRpSYZhJ19BJ6YZZMRBDBWvnaPKRMuAovFlRtUE1sZOzTQSZKxif77ZR1HKi0secd
qVlbhpemHsYQnKIG8MGR/aeYvxeJ1YuO7vQdEPSw7wAJ3e941ghIob/k5VloZBj8OndIR01hhl4s
eR854Mw10ngroGmNS6wpvI3aeMIDOs8VO67EllOKMfen27JmYqtc9qaFv16+xl7MuYwovTWFensF
j2ZVDK11wDCD6lHBu93/TT6x1Hwv+rcX8+ETZsKtgFeT83OpMR6DqjQKz2faU7/t/H4sbRN7JBUd
+BcJuoKtFF4aUr2M4yRmXyxz86rD7gcqWYaaTtqS+Xuk7jMZ6XAXQg6hPpDk83L15Sec6FhSz4Sy
y+rIBd68qhgX5zntIn14AawG1mWSYcO1ANiD+bikHw32qbPpd6OMdW/MMc4fSdISJZhxSgE2bDfo
55tBtOoc/CjG4siz1bwceFBcL8U7Lmpl7QqEOoLoUOpsf4a7S0Exp1CqR8syWVGjRt2ftx7ESwj6
vsbXX7pPV/o7KvWJOgiHDhHBYy9yNGFA1KUtLl00//yOwIZSBut5cNpBnJvYsqDZsCtILBQQNA5q
NCASy6N6mjJGn6OYLJZlpSahz2FXD+QYk1eNdjnnc7/NX8+EtYvANtSGUSC5W/+ewZV1BQv6JYbF
K7SNbViuLErYjVNSvQn7xHOJnusGj5flS8Rblh9wkEOcaTHZAiMft5szai1IbN+drz1684S5FW3G
X+DQZv5fPBh1oGK9EoLmwDUV8112RRdR1oZSEMopdLfKABajAuzpOAabEVYyrYozEgU+I+iIf9he
OEpwW0UcbA/DQ4yh42owrSN1OBveUtzdoMiHqqc4xXf+WMWOqxi0FUq8l9Uy0UM7iUs8cAgwox41
xMfufjuUJTvmhc/8eKwY98PAvwsONBulqU/amHZqXUyGpcNMR1peROelWe3mi2uzZm/qhpVLHWVe
M5Wsun7C7hrPE90Dfdawi4MugnT2KRaRJZF85CoWwvL16H3rqkavAiez0P5fWYXF8cMhI5RKZvaY
jFCloth5xxFx3lU06q7CaDnFE4od7R/m/1PioaiBSFc+FKI51HxOBP0Ss2a7TYPg0G3HqIjNmU6Y
v+pi9KEJ25iaOeVrgd/3lU0GY+Ta5rUsOzlr9q5nadZvBgU1obUolUupD7tk4VeTaHfloZpyZ+s4
W7Hqpk4v6UutTlQ7q1pbtKbV3yBLWQ2SAdvXCCpLatHVFWjV9Cr5UfAtig0mMYaBppTlzJ2B/Hwi
ywhmOHMjRAFryE5LvdLqqeKJ7LPB9rCWklrhka06Zl9UrM+U6SQBJDKB63WJzwS4wW3C5Y12O89M
UxXJzOYv/ORrpsx98r62O2zC99wuiAjTenX4bQWPFKUCcEnALlBUM/MIUcFRsFajwWWrtbal/4A6
P/wxKA89Zy8j7y8UpQ8A6/KBuuaeDznPPveX7BqPQVdFe9qLu8LxLMlm6einXt5w2SdgAPJJ8YSK
vpoFLcf5H5bmbAKF4djQylzwi8Q77S39JyjKJeve0B7dkRkvI72ke2YvktudV0PsLlYDXA/STnqd
FHKxEUylQFJ3AdRmzmcL+dGYGepLVl6HFo8zN/BnnJfE4qWPVwI4Mm2ikbbscZNMYnch3SlQ/s0v
J1UmxZYRmlZdw8HwaCynZBE0jW1QVzcFBSRqA/DHM4/2Se5pX8JUMRdVULtrEI5YdyRHeBLJxS/X
i6tWZh5EEZZquEao8oAgh+Ev+SZYgxK616nmK2W74AbjAPcb8gv41bOpkhGQ3VVvxtrVIfrUvB+5
cifu0uyDNZr2ccEuT8kr3scoxMa3FFLTzRkBFwTv05Xz/iFyPKW1mgUEUJXn4iwFvN1cPBA2v/BX
a9lZmTTecz5BemKMELabmhd6CW+kIwXOejQfJwvL54Mf2GzWW/HlmdSYr6hGV/B1rSAqvF4ySRiM
ubnCk9o+rfeEwq/oMLJGwJ7blaxpvq7GTncsvyPoEk7atFGkTn+Jfyxs6AqSDbc6s+7wlsyhI54C
V8kZcOiaDbxenG88sBVXFHsxgggarnvg4JTfvU2N+dz4TakDULO3NMeLXFSKn297fGlI7HmHTi15
EvciFkTtZzafczf27tGBbvt+7cwlCPHz+VjxoMkd9J1Ace1aExQ63p5+OqXl1QLJ6XXgdDjiSiMP
1J6UmliqpnptQ78jMU6EGc8GfLAxXdoyQBiCG+vPwlILdxIJsefRQixe0ptqkd78jxf4vdq4rMuM
RXeHeDynrAUlgk03nNs607kcx2LmLX+i8JQDcNUTcPwwKepwHCi4RSFXhsn8yh6skJof0RA3GJc8
OJRmJPDIllMiwlBvOKAsRtBw3GIQSsoLcIU2BK+J3Tn47B0EppmXrR2H27Gchp0/bQ3byjiuclLT
SMmGdZfN/ihue1AjDDOsoUhH5Tfo7sYJjLpTstzKVuFNIWB5r7sb5tBSfRmRvNg3mBCkthqXlXhb
fuaEh/AEKrAuEW6ro1xj9zuiehWGCXGPdYIkigeHLmwiBs9Yu4V7W2GIw8i5Yw8lLUZitzVpUT+g
w20Es0Ftt+8u3eXVuGiIbpxOW6yGX4bX92ypPC5wLVqvvv2mph3aUxa0uVlZItYL6iDJFiHQzSrQ
uFOwgjvF+RAhKGVdI6e6zeZ6kgfwcad5WfvXug/esUGmNqKA4FZ92qQIrBf50G+DhH/i925LRTys
8yrlsdQ+cTErgPtv4c0nP2jR40U4bKP87SBZcqmyTSwseeq4OzbmPl3xYbU7W4sgZC9v1kcT0TQg
BXCtlQb2aM+bKnqSXUqfkDqFOXBb2TYDy2MGSwEQ3bYHNjyIQ5OcZ1CH++jCeXkQxjZ4ZhzYtnjQ
zWgyx/+O8HU+CP4Fx79kHuJo1hMDSW57hHVkbzn7ksta9DshsAuXuQBMICydYKQxXqe9DJGmZjY1
QTfP1YLOA5p+JO9Or4ZzILyVXEUy1IDfeGD5Gpt5tHIXfZfVMeSkPnnVQywI5F28sJ9imjEmcneg
/kCEEHCaLGexpMu2+37pAM2OdafDurs50aC/bW3mtiOyl0qltZGERX6ZXZykCI333o49zPm7g01G
BpbkPKFMplei2JxO+NUs0Us5jFUillarud0C3E0lyQrMzPM01l70rMP3/az5YeH0XcxhTTw4xMb7
1NfHTRbZJOTPgwhJjPab34Z3eQ4JOkGKKbn0yMVf1mhO09jNuruYhA1ZJ6knONUj1aJmdcSupiu9
i05XtErKS0DTAvuxvgOq5rY0En2HyRqzjMY3ddFgihr17QxMD7uu+DjxdzH6OGTrAp4uKuVKfJD6
ukx52Oyg+Z49Dcvi926JaomwhY+WcrlMymfIeGgjy6jtBcoO70sqUgBdguue19n/52v9IJml1fmP
+F89Jh0pFz6kFdvwgY0D04CXMgId/mOHj96gZfFNvAk5ki24X3OPLbUYK7oKJDj4lSf+HOEj+Apz
B3SZAs8KASsEkbxJZuvxvJ9JlMrnx4y5Gamgm41Lp8kbzlpQfIWJ4R8ldAHTqdCqOMlqvoIFXYFy
kVnCBk0jVy8NdwEinJq7Z4slrIirxmJkyVPtw43WkZ4PVrwDdlLO//lJERkrXFTcxGgOJRJ+ae09
t//tcmXIE2ZS33Ksw9NSDUQIfbm9G/ZEn2zKKqPgOoeKg9dXQEnxYiFvjHZeGHdDZVrMPg1fQNFc
G2sKtk9EX5MwS/y1IhlomgRlQ1CLe4Y5262BlTDPjx6sLxjlMh7E23d9OxxsFNwUTty/0ffWfq/7
XjsUJPK4+DSjnEDPaeQshAuvytgV+XxnuXLO9VKfpCGh1fdoVynr0bDUjqTRVuCQLg75Kh9Bm7Tn
lZBEvFs28dQ1QW24ELnNUCakA+UAWND1rMKWN7wmbUyoRMufUIjA4k3hVNT1DnT75mBtTTaTdmPG
iwjOENRvrNFoZQ6XD/1ziAkyzU6ANLoR7fYWjjRcVKIQR0RlKektj2f7G9gfSV3PHO4tiGArQfDj
kzwgIifHyYcJicxvY8FcLDtuCkvsLcqzNw2deo8GajZYzOdGCauXpG4hH+lN9kJt12+Qkf06g9zn
aay5OqLybbnoMC0XSxK8YJkJ8fkB2qk9issTQB4Y+hvYahq+4RfGNjKmV1kFeerfF5gnKata59Ug
pIMcAYt8REDB6+hFc9p8X/qVaT/uMYgiClaN/U1w7vNDUKUappklYT6hJ6dwLw7hLzQ7INRiOY1E
40l6apT6FZYEXPWDpZKz2xHVic9QOlx5rb8SlEVL25O23SMyY/uVYeL+HJSObJ/CVoRB2usy/wrQ
fy01roAJ1SI8+1gC0hrIxviBl2QCB13JUb1T7CU4ylDna8O2XUNySNwCX49NGX+T+e3O8zpcjIAB
gtjbnbMUL5farc/vjLoEWN859DpWweqQz7Lia7qe59e58x2DojYoRE1+RbD2AQSJNqy8PD+kgTWl
7GENSQ8yNwtSLARwBJq71x6WnTMacD8+oWpfhAV8JAYILHEXX+rYXM15BRC4MQ1gRd71n7zOJZ4N
foWfEtjWs73EjDCk/MsRWHcHPrh479kH3piAmthfuQjyGe0JwHARZUO/5m8w2ufokvi9gGq9+kga
RNN/DZi5PhSObHs3YdSRsi0t5B3RAbt/dZlY5y+lKmKzONgco2gANF5efulVta9/3sB/0pWcwzin
ZC4RECrNe/vN6+GXMj2EBGjcG1jpQB0YhrLZaEJSb+Aq7cW8jSAWB/TsNGhv4G7drEgSe3cNK8EU
nEAMiil0IEdIU4lO74IUNm7emt/ygO0oZzeGI30nkrjujomEvwc/Ok9Pa/uoxsSpRVb8ouY1FmXT
USSX9knH8QnxaNMZHGLOHalQxcwUbMeZteWtekXN1cFh0L5i3LsQ+n09T9CshroGFMMbt0vtxUqH
jFeYWikKLIw4aPzJ5iIRk+73bfvOUt8nEamrPIfYOOozitgMgFbGwHCw8muWIO4zOi87f5s6qHBn
U7p6FlQ2H9DdqQVYTF4uPOffGWRyyTxG1Hco6EbdCsT6TYwybXZoWZU/CG+tMjiPk671I7aBA7tL
ZqG/hAu6SVquk8b6UDkmOUHjwG1xAFU33aE85hj1S+t3EOyjRQ4BmzpJtP6MDA0aU6ZsK0bq3Dpd
+PUnVEne3Ont2WM6WxgKSkqQR9dSjx6cAYHjJnhGZ5cLAUTw57Tu6is7RsVTWKB0sE+ScalfCwLq
Fy8n8uLaC4VrBSGxXvvRyE8DOJA0JncaIvrJBkGD4Si1nlUsnXqMXs7Rf+TEbA81vGDhfOHsha5N
XrMCEMSkFuHMvFYlZIgB4PVxwsxW2VJFnV+uxDMURffW/byUS84T6ltLFKGrW5MF2X8+YiEbWk4v
2NHXIUqoh2T8MOxQWeFbdghSUT5bX++odX5mHXBBiDuzuSV1bswNU2YyLBSPugCn7BC9NK1SzGdI
9wc7XqE7jXBK9pMkrb9H9Hb6r/8j9hh5T+nlx+yffMzEcv+Yilp3wADc6crP3FhpZ3qPv6c9x7vO
3DmyH+LTZAGd1jGxo0r6CQZcVvNtO7eP0Y5zNczrbSEIAxqBPmd6xrBNRBjh7k8VZhbEmekixZME
CQSoAxKXTZsCPAKHxmvF7cjkVgm6nq5tSy3neIwKW3W6q9Ztth1JkTQab8jfq1PS4vSuE8F9Nshl
riap4vDQU4TinYbpS/pFe4ZvVC0XYy8TaTInoZynxqHAYMdrLnJa2AetH58rjqEo7rT8flU7QzRk
3htjucVjto4k5unLTz3bWVN0/W0PsE2tsWUUT/GlKPHCcJdq/FAkfqZDtsI0LuSWeZuxyQpNQcYs
88V5SU7YjeXvEJoEo4bg5+XJrI4w2pXu7oH1xQHBaX0pDln53qa4+n6qPBCMiGIeezrRnvbivop4
36D3fMMV2vEyIXpBCD6S9P9zHiIxuh25hE+YTS7yftX5RCEzlW+lM4E+OHKbIxEZf9V9sYAnSTYj
EQfOA6VVCKVp9TYAGPQt4OMGWbphGl3WAgKdXP6b3jDk032sC7/Ls0QXe2Ns6ZNmBAal4NHvw+yB
6FQnbhTd8fTgtmpCeV524vvf4/E/2f+DIldePMn1KD0ZMqjhk7uuiXG4Kgk75CD9TEKhKjctM86d
gFdhITNaoDfKtMle7Obs8jpOJmOT+va6uYsJqcNgpvq8xpQv31qut2QMpgL2GK5qSI8wH7UcrASV
uu15Dykj+qwsbv/iqPN54s250mFpBZ90FkBSCnwZ7O4NDIY3KwqB8IUodNIjAtfplv2smAI7sYXH
6hK3/axJ1SyyKIRkrlT2T61xtAGAs0yFokILOpsTJEunsSj00ZMpxd0rpHg8Rs6/iVD/FBEqFlsC
SEmGMQwo/XvmkWKZCb27re6d+h5kABJcf/Mu1c/SOsvZVQ+gNc9xz5neTiOuDbfcTVkpI09GVsk4
9LNRoi1X3IX1x/h8sZWB1MVviGeoA60m12IfrXhuzhPYROiR44UxZElzYkZBIO87yyq6DdSz1hn+
OInjhDKZXzNxWxcM5vLtPXWrluuuCaSHiABnZER50oQkaS3RAld2p/J4U8/D7GbbA3hEUDbnXZL4
l9jfwvyZRRMibFNHTo52kiBKoPgPZtCa58D4onQEki0Opuc5O2ELqxycDG8WMeXdcTxO2fw+MMgN
KaN18RTND5ygG71adz4GZD4sgi984a/CzaZMe/2mG4UcRLBz9q5q6dm4dtQVm/NWa+EmTRB1p6Sn
MlKz2kRAi78m7X8xFxWB2oKDbf4kPUfpVkqgJMq73YVxz4KzmYvcZAqyHq4z5RnFpIZ1/RgsZGnq
OSFI4i0/kQzk3XupXDJwtiMe4JKaQWiAv9WuY16WNMSBGYxgfC3VKfk6+H7V+h5ryzyie+CWkRnr
prhd1slpuO2nBndYA7rKux2HgfURw1nQxUy2CMV17CeVxnQ/hpEhQxNKYp1Fdt8ze9JvFJVij0JM
p2wSxX9d/iX8BH7H1l/GL/zUr7J7aGf0XFgOFRr/3fiiDtgz/PLrfUvYdUON4GQald+CrFzZpa0I
iHl7DWdclgySZIhYVgnuEaEVLdmWkHO9KlRcQyXI/BTwWKPGwgHgPJESgNmWcAoTPS4Vk+ssazbT
D2OflU+uJxVpgi1DU/kGiHMM58uaclUFuOjE1a8FgOrx9V4LXb/F+hasOc1KsmwbT5giEYRUQ10y
7haQguMTutnBSl8TxBDaj8GF5c3XbXZdiCcoFVQJ0/RJqYPlcDvM4R34pLqBElzH7V1MwxnLDJUz
afwB8Std7ISPVCHiYDjaUmBuq8l/WYluJHiMrEIaifQgk229HQyrEMlyksTpORzxBlMZ516nIyJz
vPuoY225VNO+e3ol36E/wmFzWCsJaFFr/lZhhS6phj2No3nyW3wrbHFABBS2OC2b97K5cSfzAn83
exCJ9f2ZY/EA0oSg8BU9i3mp49mv0hdstyPA2CPrXb/IMsOkzMHlNagj06VlYBvvtQz9ksdiP2LL
7tREYSY4B/r2dwn6LCzaLAGh83P8hOndUK4vnPATGzm6hAogOoBmZZXSUD9krS38wUtsd/RfCusZ
PtqPYQn+q0kLMHra1WjOI82C6sYbqt+tFzjMpkxIyKzVY3RfNUAcZaQCfDYeB1+NrCmHB6Vv2Zat
m4nbi5uDZlR0KCD32kuG/KmbzXaZcOMI8RZHpp3+GodFG8EsQycKXwJ1p4JeRVvLYQPv+WWeX9uF
nRkg8aJkiMZcjVpNIpYnjewjUpVefe4GUIHuYrBSNgIJlN8nu8eFHVqCFAhmbYTtdI3Jv1UW6/vy
QOMCry4huiIRjR8Ht2ctZ4o151AZwViLjOrjHbUKvPsVc2f9MV49PocPQmGJ7TTyuXR2E+QAOVbr
oiZUsHT/+fYMNJJQr3LkIKHXkt0sRtsogD0ejbBmrHEmpK/EdYkPn9WjznJ7r/wQlrWtIxQ6AI7j
UcE5Ua2QtgaV4fpSMAEaZBHmQ8zgRZwhuDctBAtvz3+KFo2TjMOpuTB/cou/pvqHVfBiF7gGB0cy
om983Ch4M3plK6i4IJRBpyo6PQDngTb0kELGOQlr7xBi8FMh3H8Yj9ate7cDJs1a3ulonebi1hl+
ZFyOtuNr4Cj7o5n4j7txdqpQ/LJ2IEIXHJljdToe9+LlgFKcKQ5JGwC506btEYu28TZKGzXiVY5H
PMcvPiytTea6t04l/4QXhyRwIjZ0b+77UqK5XbsdxdBfLOuz3085uNgTIbkye7dZ2tR+UN2Kz2tf
FAYE6pAe+Q5qS9Rl3aaMG0x1WScJ1wAKR8fW1vYmyltpcfhOp41FrNTHsz0gkuAiOPj5n99rnSx+
jt3rnoXXfWhRDoAzR3CqJOKaS4LCktARFdbT6az2iM2B/ZGvgEqtGiXPSDwK/ys2aQlBzdDu4LPx
xSKGlwHAT23ym12G1sQ48zeQr5YWqgetEVu8VHDbH6C9tlf+up7PlBhbqfuRxY7+EMtnwYz7XpV3
AD1lUmxv4dI9QL4Dl38NqfdyZXU1IXe1hpOfXP3cmFoOl8c6Hjwabtld4sDBW7Ijm/k5tQ5CdsUT
TJkslG8+ptVMUFn+pFm/sgjpPWrn0PjdRHtQBrYbeCtE/QuVU7KRL7jUAk5KeDJ+D1eb6KWWX0hT
tbyI9AFbn6j9tN72BhAaPy2nQ3K6F48eZpzI3aT31ATvT8g3VfbW5GjS7rZ9OLvwBkkXWazUF44b
sWdyn7aEFRP4EXDnO4KKZs14xsF+hLTD7D8UjwbUIqH9KSutYjf/tm5t2FCxmwpSG8C0YZ9LqUXC
CVP+kryOQXATGv6mLVf95pBAtLyYqw76mnUMec2XPwdK0frwECZOCgnIgBCz1FykT3OrzX0pYuHb
Yo1otZmN+porWVxA7lx+fp4g8FFY/qmiGrA9sOoE2/b79yjN3B9mo4fc7IekM8n1t1qA/7rM6Q9j
l741PoVmWHF+RN1LSooXZF3WTp+xquqhR2U992hcQkhWrjoMqu5L+EBVibR0VaU0pyok4AqIfDNv
0a9AETsGEigtgXDm7lrAm8QUkB2LXqyCLJAHWgT7F146nWv+Cd3y4J+Xan2/dNCl7d/oAvKHz9i+
IS1AAowQupwndZQcNdZ58oUMlNIe+p9m+3mAs/Av4V4ng5QoTVUoSet6SIRmJAzIL2/rKRaKKf+U
p2pLB3J7TXBmBprRdg6xkYiGJHKIY5sOgNaETw6iJREPiumMdnzmUEvI5W8OJifWOIgfYotNZr8i
OABp/PO8SOPe9C/92Kj2aLEnigfnTOhXuJ0NBHw1SFbXbNaU5PvBX47ZaEqVNn0YaCwv1/jgiSMi
DIgZmQlrlgnAi/QQl3HsbzRpoOc9+SHPXK9OCttHq2KLgpRrRNPtaBpNBexvGIooJ/9uReYluKxV
uksbyFrMXXpURjQzKIuCHGdPCu6eUp9zTKZkumCtM4WVdzAGomiBjzxf4eIYG0p40r2IFjLpk+2c
/VuiE1os3I+wnqha5WDBfmuTAf72w6ttny8yLRb++PwmXQfiq5MspuzjaInuiAZH48hucHXetMCl
zTSnvub/iVRQ1GYPGiMgA6IbQ6PhotNnkhzORS4VqGpwewaSZi8eVg8r7UAOrJRnA0iq7Wnhr6IN
tj+IS8lwg69X06xDslup7NXGEE2vTIEVbrACeo3E2//Y4jPFnDYWIjlOs/DxXVQRj7mO/AQc0wp6
iyf5ol2YrQ8DdnLh0EqPVuyTPr+6vq9AYYnRjprttZ/R/L/yiQT97fMjPwW+N9NzCmVQ7b4C+UW5
YlvQkwpH3DF0GJzvAwlNM2Hry3VTKGFRchgMqicMV8jMx1baVx6yPF89qB9SSPPCwBM3u+YqMlho
V8o0AJkahCgknQHOCTTh3Nxwnmo12rNrd6z0sy0LtX/YoLLDQCmTi6fplQH5sLJ2p3prfqUhrLzy
BrW/7O9Udm4LBbrLhboSGhEc/vuylw5fM5P0+Bf1K/iQIr2itxoBeck8M2C7mj4s1LkRKx/bza6I
2Jyu+pESJ40E0iPLzbj1F+IT6rKAJ9QO/8kzP2ltD6QIRgdr5LftqegpMBodCxWI6V5OgUxcXqEd
1bR0r5AI/MwuLK57o08ky3R44w5unLT8Asq1stgnyRShbyXFdtd1Tpnz5lkECQg3KcBab3rmHgr4
l+dP9uOgbA9iFXQCBnIi8pZpfhBiegRdXVExtnW0eRqNQqgEr4Rstm9rhwF4FLA2EEQlR3fs8L9L
cdI3hEoEhKvjy4RBdblQqx6OK8cF2L3g7o4rqSoCwV1qWMJwZbhZfzBkwoOwNcezJwOmwC6VAUp+
DpRx7EFhPClyQ5ck0nF+8nsOlKZaH5mo6Dd6exnPgiqW8punILjMqz7kPGLOH8Dg2sPZXsdDavdB
ap7Nfiee6viCdF+Cvwh2F2xGW+fqpjE+/ANXIn8ewQfn9igTymtu4Q6LI23pN4xD/CikVSd/hLmf
4CCMoNnwikDpueJbxsenS7mR3bsqnicKpT81WIlE/fiNlhu5aK19ndxiKyy7IUcgeyHc+hr2lrFN
1k+b2bGWzd/vr2/KgeXn0XCSFDOkpJe8AVUihtqz8kHAoSSlic5nYYqaSwt22EVi3kQpw6bfaGDU
Uef0aCFQI9xvLZZof+wpTrgSaIOgL4gVPyN2iAvRppwd7HnLUBHePHbxj74IMJh7C7KZFBYiPSkw
jF5RwEW8ulcAtTWgx1lb/2Br9eFJBEzknEqMUl5ol6sYxht8kuKIc5kFDvlTvZUfy47baHM7IFiI
WsJKqssdQPWbMVgvq+fA92syZj1AUdl7vu2UoNt+e/F1l6MaoZqVML3XoeLbDoxMWQrlKjXT5GPJ
Hmq8aRlZDjYPFf+fQlhlKDRZKfYYPg6rbwV7FFlY83P/T9OTaEplg36wZBl5OGU1KP1atH4XcHKl
PgSnR3asGpRuZ28VGpN9Ny9U2uDcEuaoZNMpuNH63eJW6n35uGLKItuP9SgwKDM2njn9iNb9kBIV
UFAu4vauQpmZAMZZRZDU+/3kJlSHh6qFMf6zw0+1yAwtAp/Hbrt6CNVLc5Tidl1Pp6JdqkT4qYtA
sP3+eTygh0wTo8V5Kg3TOx+X/hsHKOFHkCuiyC/xCEhpCA5EMdquXH7MFhmSrVbP2XseFefZMDrX
7slr/Ycd00lF3MC+DCz8Kwt5nUsdFigRQuFpdpdhCgJCh0ntPq0DElg27yUtRBEz/BAzJweyrFzI
5u4sDMY8OcpArmFz9lUVWaopvNDeENUTUfUbMW0bez89kyGbp7/0XURVflPI4vYtE7MccpS0NAWF
6k0Fzm6xvyXcsXschT/J5AWDDgn6bjmoXsyHrxMCUJxkfHqWAiIVTuXcBvwd41IKeORiOdFU89PG
rp2LRbFNmVS1aEDM+bC1K4d4q1gN9VoO7LU+zj0pYZAc2qLB3vOuP8oCo6u2RFUDpc6Q3Z8MkpgE
+DynzYkfvbPSsv5ug6aMa1AbldbHYOJN4R+1vQdglV2uXAqsRMMdBHIW6+sbbF9LPD9W+5UblQGN
NwBCKHABW4K+zOQQs3w42u2oyLAoB+1SZ4FSOsxwb+OLmu7Nqyxima1IhQknNrfgQg0d0Va3orZQ
MJf8k6uw5rRbMRWrRByLIvXBX5LmWBEiEC+S0HqnZfwmzeWENYmpJL7TEh+E2R78fy+AblBASbch
Ogf/LWf9zH2BUsfhMbMubs3WZPtI3xLbMrqpUoMopplR8Del6OrdCibcUcPyU1DR8ZSTlZ6aM2lr
3HE+xHpvxIsxiVXa7Sh80r/Xw9RIy7v8Fm5MLKl/zfxb5Wb2dF37UqFZpX5sNBMSMWWZ+MteeFfy
9jvpE5A74XlojSiXDJ5MNb7TdBnYuHoPVwQfpm7WjQS0FY0Nm7GBkhhPlZ1JJtVhFrtUgMvyEAUC
VspyCGd1B3GTFc4GR2xA2FV8nqHIg7TGFR8y/4zEUumtKwNqsB/m+wAXhBxgb5hc9Pqn5iIg+Qfz
k7lSYU6+SUckD3qT8xJyqrJ4EWoAPCMH+eWyd7Mx0F74EKi6UnQokjZH4sdkdy8xrYvKenLvpXvb
MOyNfSS3U6eby9bTOyCfb3G9AuvLu8ZB1hpSMvS7Mm/vnNCMHjx9UNEplIcoRh9fLJlm9zVPY7c6
KY58z0GYvSGIkifKdj0Z4X2+qCS99hKmWRsy4ImPepcXZ4xCVlzOA6T8T5CPDQ+i4z2jAFiL8DTV
f2Hne8Hh4rB2b21IoQJ+MpS5FWJRHns37AtXAf6YxUCS1T/skhM8dUh/YDrwRSgqE5NQM//2+A/D
mOFtWAuNNHbjq1s0Y/gasjdGLFFshfqQ9z9uEbMI4ezt0OEv/KJbooi2qQi8iauO9dmhLYEHAXQ1
Ta035qhAUV/cBDOd6kGeD+Pg8z6+jNYUsXMwo5Dn8+C9etBy4kwCZddxKZD+kPwltYjrqylykbWD
KgTq/GN3iY2+nBKIIjN32x58ZyJ/UNgTesyEYw3hSqCH1JTUoLKgap/WBLc0Y0pnCRYBgpfiuAmD
NAvZ/gWKuZxHwVPcGux4hFlPiK+/3pESOBVwqHcxcpqIbApOGJ3mWxAzn+gsIaTIRPC4o196/Ty9
nypolVWE+3fKymYjAGe4sV/ONwXv1BtlDs+ltJFa5OxsA4tZolCgfKpyrYeB2nSXJOpzB5imTsCG
zcsG0KDpIeUzv2OEy03gXqFu8uIxXnHmfgHn8B9FtdoYhLWQaXRabWoCPNpRcHfBhWuvK6iQTtry
PjqkMDIB/dIaF3cT5LsiTaHZJc7OrfvfLZU+XYijayU53eWRbOTJhPi5JzBl+LWdD6gs4Oq0omAj
2m315f8HRcarPHrHve32KVheUo1W8aQXRj7bQ2dVJbPDuIgEqmXgCNgKzIfX13jKV4l0GOZACE2s
mHVNpOj0W2RBG9BM1Gc1W1jZP+x7nLKaCmBp2C0Ocx2nGXN4VgriZq5xpbVXYQsCzREAOnj4pb3o
umS389OAOks3iw1BRqpvcc+WzOkDK+/MMqPP6usK5iGwgIouXzK8XPM5n/+YBiEKZMWNO8RTQuHX
ur4xDu5B4GYcfBGvXgyTRLguHA7bzLAH2errE+CbHPV5Nh9Wv2WwCu99jL0UpUvI7o0N7I8sLkkS
wGZ3CvYfUsXWm67lAUSrUEll3DUR3mlxsVu+HL3sEfLpqgSC+tyZXhWkqh8ERJkBfUPgqUHAauIK
g0mKll3b4gLBPYANHZeXgWhrsh13OQSiuJEMd/q/N/oBB1MkBBxwcaueyXnAhCEIooHunjRHZOtq
yctk89AndYrvkpIMb+PhICF1FocCXffJpRbiizrnTsWEXlUFYqhLwDywLMLq6gjZUIa6H//zcI4T
z519n74x2raVjGtbixJNGS0Vki1GWsQucZoFnzXXw8P4uaVPoKwEm5b52JfAZbqvNWhm7iYw/+EZ
gosJQpUCAVTIceV3gZlR45vtdWmSvPLRB1rjd3Ru7gf1rSTWIqBIzx1PKKjyI9c8/mX+rP535W3p
c1mr06E7UqD7bY6M1tFUx4KptmYcbpgua13SKOvW2SEBatQ7ylfSf7oYJq0b69B4H62veQwZR0xu
yYb96+28l9pHcA0mCyKpfBQmkLhwQc9cRtT7N70g5/+oeyMWArRjmXdntGbSnMNLJaF7Mpm1CZef
soZLdKJ9pyTC9YR7FaFWtIExQwbSt9OhjfkujrD2mn7Eb3WA1iNQSOH035wk1h0Gz/fWj2b4tYrm
taxQZ+beWDPvxLvl+GHjgphfVhl5taRt1BzAoo1H8UR9VPC+0pM4Hs70SmdbYANoFHpuCRQgUJ3R
xFrFhRrwCrEn9qtHQ7JQxEENxVweAXg3r3JswGnu/NKwNagbGCNNI39RJNXIKAD2xUwjvfhdFh7y
3B0qUzMe+7T1l4uDCI+on3/1gD0n6OevNNhLbWaJPOolB9wh6YJfB1bFuV/BoWsDTTbM8xOKnAkG
EKDVO6st5eIcH+S+IaP68jybMOYQ0e15tG+sfWxfNmuVae52eo27rN89hPMN09yRFWYKveequ6pB
r8dUiacwb5qaKkzZaGEj9FQEnXX6U81/YlUAubnSctC9XxWnhZ9zV59A8y42vUAZWMsmjfdNFBWM
h5Rjt/icQr09UuuKEN9MYeCv8KnC310NVNpRGMaMh98XP4LiYwDJgVqVXxKoa1WjOVXYdlH9Yn9p
1mfZqPtg4RthId/RhAtvK0XTOYxFr3j9sL3fhU3g412MLTnyhWFE52/dMRJj8HUJQOo+UwAEH8Q3
NBa7Jm4zLcI7GVARpJbM5Ye0j7jFqBdFzMfC7daeUNMZSEIyv8uqtPfsivlIBINLC4xnnpBfgglY
+i90qx7upA4cgwrjKAOndg6H2fDPZpgsqAGQV+CzF+0xAlk+twpDf8mVDAKrlv/JTYmCkLMgEwy7
XCimcR/Z8HJz/iBD2P1C/poECvtYfipoLxGd3ecfHRTyPWshCODDyUC4kF3oWveb4tmS6+m7tPMW
Hw7Tt5L5i4GMuUZAl1Z28OoFTHdubSh+YbBwcIUOEOkfkViIilwyHCeA4m3a/nCercvoGEbH/hBH
8HblYl268adO9ZX8VzThTXSX8X7cyje8Z71uyIMVkXl3eDskt6F5WXXx6vwsx383sR5irBw3gh1T
mM8KRjj+kfm02HkD22WX0JqI7dR/I9ny7ktc0D6hH+9G7HaiiqAgOeAM6nnDjj8125MQ0+kB3+0U
4+IhH36O1A//bGcFNPoj3IYtUJddy4yy0dKTwRdIyUmyYVMaxk6ztHBMgosXKgzpK7/2kcL6NOI+
xYh+qTmYFSfN2GzId50cRNRsMiuGlpGNYiDjOjQDlQZfVss9cGceQw+BlKhrbI+/uIRqe3uwuyLL
mKlVH7BMcxuUofrk8DdxEBlNViycHZrz/rgk1OuIviZmmE2rvzN/m/58QsSjC5GCDDC2qPsIYAl5
+JX5m7vEaKFY7WZTUDqAgOK11ndyLXs5qVmswz9iBzYEB8PH0AKfnGqUHXg+Zl3PKy8qQBmDWEph
pQNlZ/IER8nY8c3ovIwXmfv4Fja1OyyFra8D4wm5APaQUy89+4qnW/UIxtgv9ePzHeQY+NaMIFSm
hpb8IEttPCuOQZpCk7EGivrYYmjVYGSleGL3gRYm9jGwFxiatQvhb0dtjCyiI7s6BnkVsZWWWQ2G
eGpC1QiZNlcU8CFauSVKGNa8THeJHdF0IxwRADk62RkDUp2vn4KJ7HZX7UhGGPtxxUhK26rl0/Wo
1Zk83owTGWj7yCFw/I+E5Jdh0qdzT2FB2PKVF0Es/lhPKRa92HMyoVCOA3XpaxwYwHJ8CwSNbZ39
XSMvgx7OW2pRxeMIOY/NsdLA/y3uKdWHFKWHrRPxwx4ZIGddE0qGJBkMkKm0NMabchJHFwp6Yn5b
wjlpknPFZmO4xTc8jB2VSe4lbR3Zhb7eZVnjGhSW43nTLmIiMuhAcvlN9lHZlydF3VyQOULjLAUv
Bv3kLrBnVPuEq2AgpxRRoifvqjsQUQ/QmpSlxOxco4NZYAudVKxVL3lTyvTEHCxw8Xvifzp6cVmB
35mFN5c/1d7sQv+A+UiVCTbgSnpX6X1hPiyFCosbVVX4PlyJRlKUGLL87RfHqlMnRtZkCXtSFm/t
m2zuh2IknDZv82xE2U1Q9YlVekmw1EBg4c71jXml8YCgr+xroSkX1C6+m6Hbk2oEm9D9MjFvUyuu
mofTsX2Y1wPVoesrRCuZCZuRBUkG59gF4vhlJAYVMaM4ThCD4NWLHdEjGti+v5gsn+ReqBLamsYK
Z1Nx/As/KVjLJXuZCu27S1fTvLPZWO4hKOD04BKlj8gMZ6TJo3Ag34kAmkHZMImY9RucGoU9Shpb
17i8UNmC2BEWlMm64f3LgPatn39ZDuQvnX1IQA3Qw9kxZqDJFA5lOYro6+hgYEeHyDvvUpXMGyx1
cqkrYkhvD9WdBBjswjsWuiIHNWbojzHJ8sivJCS/GE7Gu4oXL3JEYyiQMLVMyQcNG4K5tVd4Ug/m
Yts/3OjB+EXJtC15NwJC6CGPqJ1w9uIH4wHGFAwAjran5q3qIoWF9lNcvFKsHu6XTF3o6q3VIG79
ib4yNS8qgDi6Ttc3Wu6lYcrMUBIeL54e+ccX7EGzT3JCNMg33dR48cmSUtr8F6alPFO/bSU+1waR
aqWRjfI14Skqp7oo/4e9HYVdl7ybAq4JIJadVWXWvpGj6PC5LYM+rOow6uVwKVvdr2bAm+F+WOt/
ph5U/fiBORTorz+cGA9e+bgz1a/1GD+01ai0uJlID6YKbB3L5DSt47AI5WCCcDE1UbFNERtS/J9i
2v2C61tRXUS1MEtGgWwzBxNogo78iZQRBYjAIOpAHITElS9au4dzns5A1iKE3BsHAVYeHeve61Wl
ZUJtzZLms3P1/56P+P3JwJvYYDJICnDNd8QolfgNVecuavDSaVe/Ph8chlFH9q2TtQbpQy7KKEnS
frvRH0GR7WhhJr52S+VVc3mOfiNubza8nvK7NgfGjpqHYhGcxNx/Roriilq1g0qaZNNgobV1PEDw
jd2PPj1mVmNefXNld24NIOwL0J0Lq/loYlpUenTxesOhmjqHVjpu1/5lLsjnVyAsD7B0c+uAtniB
SDmZZWaRSLTPH2bTEcnqp9u1ao9y+TFwUYuquwV3BpDJMiEVzSiWWd83rlbvW/apon/wKGIoGG+D
snGGG/1lNXx4xdF5IRkkCZsiozkmjD/a3YdUm16fiTTJuEOHq8b6Rxw0HvNsg+rxtFpK6yKxcb+e
El4/xENMbKmo9sCktFUXZVAq6chyjonoKNkQl8zGSYCiiJHY4msKdJHFQtH7cq/o6OcMHDJrAiBJ
CiRVWTzZd09Yz/F5sBs1bTsKj3VxGE8qq9yZp7KS1hgna/4vWz4AuQ1Ghw0EclXh0FrYMNVw8GVw
6f+fjvmZCU2ClXUEs8Rrk9JQPkSpTwo6Cm0mi+6i+pZDIIKn8zjaae0kx1759jwB/7wNaERSZtY5
ajFp/wzJlvDRhYRjNfW5+tXjVzHfbyXjYQ6dyTwuPeO2qegq5rfcNZOnTXQ8+E7ynd7Y+6znkmIb
5gM8+6L/x1Ytk0x22IW+8Ecc3sprXbooizA+wRXiJprjM6AWTeU+imbQ+MmAyHImqKC1YXYVJVHR
VvOH56TUwNeWKT8cBNuHXz7YgdnaHBaFsPXktHcfKVw4XzTmKZOK1Vlysg2SHqdX1Ngm4xIOwCbX
S83WdSzRW21Zub3pxQBfaZuHrM/Pgk8y66qrzn9wtGG8ZMlYG3v1gVPul8T+2NETxq2vEz5a/taK
5+lrTQPUNWjfENd/K00YWhxiXb3amuSxHioo5uQT/ij6NXbkRO/VgjNV1LtmMcGSWoN59QEW2kQ1
AhFZR46l2PCExIqes9W4TiGzVzAm5kdWTitnMvlo1KtNy2/G6TxddBCXyWLV5cIgbzP6q5QJmYr0
89IYxXIBeQZWlvaANdBaW07aB9L5/iSn9QT5xH/gWqoNHwQFLpBBS0arLmU027UW1uEgg7ypOsjB
hpPp0Wgnlbj7g+3WNR8CpROlkrHVBmuOgHWLIdyR738sZ62w396PovYt+DJqrWEKAAJepDRstDtj
JCHRVFo3tC/aRsVwom+wnPy1WtBzt/KN66lLWmS+ywnNrrLr+Ko2xAOuh+HcIYr5FTPex7wjhqzb
1VT5rUyYxQAfmJeLLKlW91tY6OZq3MdXmoEf/+lxBZUluwjCWVxJgVGbm7coh0ZfMdIcRIZnqvYU
7mZv/ZS1CBAYrbAkgd83MJPHCVpC/k8os9MacZe332EqHLCGCmuriGOxzMf2S5Yi2sy1PnVg6z5u
fXuTM8PYAmVTuHyi8bkGFMGU1iKCRF6Sa15TIrW+l5dPBk9iqa4jxrT4D1/P3OqarmVPnXCjUFf3
EcMBUJX1CKMvW8+aaKCY28n+Ic/aoogWMeMFmX/+459gqohbJd/ya6H5/idOZbTXWrnZqI6SsJxP
lnKTjGAS0ii8OOWIm8Ak/j5JQiup69HGvuQvh/82D69HRFctgio0FYBacRVon2nRLxcCDirAbFVk
Aj3bhYy4P1qlT/x3mYzR1GZ6rGbWkvsq3mj4jKpxw4ETLpDoHn6grj8K/37gZNamGUEowfCwcwgV
V6h5Pxa8GMU9ZqiFKrfJyvsAaaks3x6QvJJWnfjS1mWcxXTudvolO5of/8TyojTwr/Fz5Wt0KA6X
nS6nUjWhOLpYkK0Yts/iew4oPFc0G1rGiZHGsyk8tEjosBYmc/qwCz6/WG9Ty+WLQHfa1QyubxRx
AFFwcuRyHYjRyrJfhpBnDMDfzCN1g0/R2TbLRDV81MdLink3I2F2fXULYZXM6fAudWz1gzq+JCMm
PC8PAVEXnX21Fi+81xWAllYQmZB+2tj/lCAD0yE6FiPqYEpCcMcghQYR098btz+zKTzcOtxeRVCW
9dWqAlgXKqJb0VQ474suC3kxUwKTjMnXhcxA/WVv4SP2PvF0zHqVSUa3y8h6AJ0y55wdPx91ZCI0
i85qGaY6n6danI8iQWlNwJmsz/bmiXUS+/13Y/Fe+6o/yNb3s+DMttjZiR5F1d+RgFJX0i+0Dsl1
K+/lbz/Y/sy4fkZWeFZIo1TfxQ3EVodzZW3RVcmP/XPQB/mELvrNI6njjontOO6akdlVaZJJW2Cq
QgjUCvA9aY8BWOjDMDX3lq7L1OPYvwOQ/5eKK0Xx/jA70zyVkUKVkrczjW2bwbJR6lsddffEec21
8p7s5Ems+dFM4gL+38d4XILM3Evbll/GW6RYAKN4gNOrzd0uxr7fAG8I7Wte4XyjkYbVrsVN9e6b
inZwolFsjtaAcxnVH+hRvNlCiQ/5DnuHdZ/7Fgypj4SCuAeh4itPFZIlY/jy14FcJfuvEqZveJ0o
Q9W2Foam+AV24QHkAIbracQQtA7z1rm71uk/t0Cez1PEXLqROIVcSIhb5Mj3IOf1e7bzYYkCT8NE
Irf421HnNwlQSNII6JQiA88cdcpiL0kWJr7dJeyM8PTO4DzaCoydExRpPRd6un6dEMhVYQMnj65g
XgZ67bm90/Ehh+hk/PjQzOt3hazSefgG5OVy/7kM7pThU9l5f+bkJwLzpzMMgIrVH9DWaaTeiPUi
VZHAjoLFKFEQGAg79u2U0DCJWl0aKcH+25SUHJDa2rqxXh9jxkoHRVKswbuqJ/urZjnizUQK2Do3
GMbbV8AkmX13QSIV4TSMzM0y0eXaFgiQpK6Ai930RePYl3xnb47vYn/yXDXq2XE5mrSN6E+AlTFh
ylOjH60fAMTCAdXFq9/12qNdrBVz12a4oX8gqWkrGWieMc2Uf4NPPewknLQcyBvmUdFvbklmILy7
lW93R2CVLvYYcxFw/BpklgpOkUBu4OSawW5euQclvti/HsRTEWd2f4KUWud0Nj4dGrKEaMLRZvUu
oxjTONKthijXtK38ve0AjY6V4TGPinCSoysWvhWAe1XVFRHgh4HRLjr7Y7mUljocIBwb6U1o0wSA
JPmk7SIrJrJFFAVbUKLMxngnDjkOb+gE/uEg6GImwDWc+DnZeM2AB8qdpCQ4peVfEvXeV0zewwOT
g0gRHcQw8GXpreTBJcVeRlzRPZ3jXMHjZq0G2lnQ7jx+enbO4ucq9isgX3YLVOu3G+wKSTXl9VmS
MwpcOSm0k8n4FZegcKbehkn991NHHRu0Ty8QX/dCBTTRJiJX1X1TPcuXeQZk5feCikFVc6Ub++J6
L6mJxme4WPBnBySYh+beLNv+PvGeiNOHaDhdBYdjasdbwNTTCdhKCiPYCbB8OBgY58wHQw8XZqvf
nXH4R+60YDWH61JeXtI5CzoSKBDadXbp8wS5Q6s1VBd7sYJ8UH7In+4YFz2JWChf4BkzLiaU8f8g
A5HrTSd1tFFwAXeBbI3iq3Bcln8/Gn4Ps9MeJ/L9QpFuGHMNbBTUKo/Mg1VlphouAI+dqbf7gznN
+DUSnUOHJuCGVmczlU9gMaq0GvT4mQoHMoR6VuYY8trfbZ00lRWS5jou/3RhAE0nxYn3z0gBLnzi
kOlHposI8+R/dQGzazFS06bvs7I+DyllrrM5/I8TLWfoO6DaBGgdlOFZUf2OE5x3nhUtimPNyex5
+sMkkK/RR2JO2A6+Kame6MeT+X1Tudy5nzLWsOE+5Ikz5icRN/WxBia+w0SR3N69jz3a9hM1rVDA
7xiWayZp2x4Acapj1VKdxmUar44egaYPAJ1dJTpjY6ywEUEeMmvDR8Cp9BbFQMUMOEsZH3pkqk0B
mQVNbFierDZPfiZPMwecdB4rd/PnRhQOV203IHqnBKWxof1ZJM87bJGg2cw7jujpDEnPDCTHWRxC
T9iD4f0dNMA1SlTF3NMbr+8LpGJmBOXebRNNLOyZnsVOKG6yE04nX4kFhA8lvdtXB7hJPFvF2i8c
Q6+9QrmP81QF/8oR9jev+vOURtbo4/9+6xp9zMEfxTN8gnW2FcCSfVh/dg+b+OJ+nJ1/0TO+Y7Zr
aXcM17NkQDOplZ5jjp4lJcD3hvluPRgv8IJ+rb8y2Z/VjXTwlKNJr7WZkb1RUbjEI6j00h3ltlwn
mY7kX2hoJNUar3vuBQUk2wxUYmuOPyiFhp/GTb1Z0n83PpbUFCYkBtqROhNuG3GUNElKgSYgmUDi
aU+mB8hCTyXkcQOWQBzZwqp/470WRyJR6iM2YVWte+uXTobyFDaBfKr1FYwy6zINaOzMRJ7d+tna
ob+oolZEBrer+bFDrGOMhbPXeP2rsrpQT9BUN7BRCpk8867agJF8mgrnPqeplP7In9A6OpaVQVA2
tH3bMzKD9/jyW26Ypdm9Ih3SGOP1m9uIINPbuVvbZ8ZAiGmK45BZ8bNYEXikeg8ZQ/WDdAYxj9z0
ZQHTdC3aJzNENHh9OWQzLsrFNR6CVztb4T26MDllHMf/69Ft0+N8Ox/x2FDr/3c3zJZz0Ugn+BwV
dQWbq7S66rgg9XooMWdNAwi+CqZCXL/Cb7NcX8jij82J+fpVACtucHVUqC9/V3CbchSQK2FDbt5G
ttcSnQ6jJ8BIDrgTDdVOHkaAT1T9r0YrerbcF/Hm9k6wjKilhE1sNFIdiI4h7jA+NImOoq4mVxoy
7IJLgMgjl96xczFJMM1mi4yjslh4nCiIrniug7YhzCehYtSZFTFQyonq0ztdBIvFLtS69PCG+qQ/
N6ImD/FH0bOucgw8v7LVRFycNb1paeSQIG1Fmn3Q1ohHpumtlRGOF8wT+gk5mtx/GrAhyglk6sV+
lZs3RLncgNqDUmtB3r+ijyDGa1tRj6ZAgJ9+RdQROJQeuax8Jic8U/ubNjQSA25Vm9drjdktIKjb
++zMw0+eN4eQ/cI3oMeCtxAjxEYl5vq59M5inIQuJdv0PFriTJCL6to1ddZn/8BuEeVDVZZ9UkQr
WRKrFbHxLLQxw13N4g7mMxR0rui3GuT0ZeH26a7SpXSBPKQ852ByU5YKiiNbMgaOwJqfTr9LJv/u
4OYOtswCJetvXO1w359Jf6G16TCn8hA6NgJcTPg6s5g42clk4oE93Y8lC2Xqgi+tuT3WKHmQJj/K
vU1CukOMNzEYB5h0XkeWoNS1pGW7rkhxQm3uQbuTJ/z3JJC4awnH19qCf5x0VnSvhdJasnxYdSs6
gniu00JbHNQ882X2X1jMHaC6NoeNYNVm/pMaeBLcgwdJOkVL75DUS4W19gkjQOX3h5IrWkODzzvA
P+qRPIY3kJVNhi5NaFMdISL90oJSpCD6L/YIdalZkPU0FI/F6uHgXNMs8Rx1B3WBHl/GnKXKVjkM
iDtVYsYiz03B0hGpvPIF+DWgqKZ0lw4aFQ/dY3EwYgZVV6/Dh/FB0cu0F0ehZfNfNUFuFrlVD1ti
YC17ZYauvppIPNPpfnAwm0AYGvhhYlemmXG80j2/JxHt2lo9FvtNta6wB4a3BkZA9wKh910wES0S
JBtjarI44R2ki3KskxwAMGfu4vDXbyJM2jAcT01f9Cg7Jc3fOQrI9AX/7fpadj4zyyqLfcpVC+hF
gF5n5RrM0MtxcoDRPaj2W1Bve3sdtxH3gSxsyZZpn9UUScPWI99DnuEgK+eQzny8CiaMl/dMniBZ
nrDvIbvcHN8kzRbcUb1GDsfOP9yN3BOtzgnDHr77sWvyFKc19ew3tBsd6APDYnD0YZo9HGIfmmmS
C6VlTr60ZrxDWqjj0+0XusVJHMJu0pq77YJAHUFdLPqqv5l/CW9HAGJfBqEcyhgknsPINooAkwDU
spPSY30f15FA6k8dZoRFB72czmhZA0gxxhtPx9+ew3fmYBMWBw86Tq9pgDu3+JOyEXaVcPiAG95q
FOjC95bQRRZaZkFXQB2I/3lDrosbKpnLbIVh4qqAUhuBgQkMGjcj/qtSB0bRIRg7PuPeHich9a+6
C8wIonjj+Q1KMPnvf5bvrBChQkRqvsTGtHB8SQSf4HeP3dXWl9949AjkyZa8cGYcJLml4BZsKgPL
X64OTDeCkKQ6ja+GrjVk+3QSxD09edUx0vtMCLgfyifsW3LlKlxMWWvCFBWiJlGHu972nrflO66F
WDOkx7XGOB7DNJEhZdUvyNvxYtaZMsBFr/65eRBECa9x+wn/PoQ7BUFE86nL8P/DD+kCle0CSMAT
dCvu8lt98fB59tCO9SFtcIG8+gZ97eOeOD6aiWoo/q5dAwKoSRVPzSsC5BqICMYSnZiUqkUYj3uL
Y9MZ3CemNk7L6cf+gGSXrCYiaADuCA38oAPE0DuYBDlqwt4qpTrvgJCfqYIl7vA6rVOOaiMmRYS7
lmjWCvMeQ2BWvKllwafiSQJYFNMDceK9pPaD/KWq6JvJ5D1OSo/ZC96912gm/YVXbY8KF+/RzHT+
8OpSxayOUoLQ20FMdme/thq+LbcS5UB0G/Y7uaU/C/YCwl0S7/9hVWPjLYf54YNyF5zCXX4Z9vYK
DrQqs3n0X/0zv1hAsWZ0cKbMD9jyeIAJgP7qTyk9wlj6fYKk07fLLgxPN8IkPOtqJU/JFPVUdKvg
ZZyqXohCcnCW3I136YiCdUAyp+CGxk4ma150WfGpq1FHiuCTqJFQMt/AG9l1d8Y9C3ADy6dbLEwn
nPWlZ1oSCKCZbeBKKGqsVHYWQWXh1qvnHa8IHx9q6t2lbn8x/d6BMnzvnVuTjaevAHQ9CAlIpmJZ
ECMmR1c6B/HE7C1uYoBMdYCCLJRb2b1A8rWPksTPQbPgeV9tuVfQWjt9BBTzNVLoD1I+f/2JnU5W
411U7i+plBbstlWe7+QfbZBlE+I78anEM30UplzUbt0GA1Tx0dAkPwej0XXogwgLyU2SP1eMfLms
yZYwlgv81uwyWMfK8z8BCzlfEtzkSYk1lgmydUC7Lk/xVpobMWBZ353/9oi8/W4VVE5nU4NjMv0A
ZhC3Sr0s5fPam9Y7Ib8azJk0PaoICUQqz2NAyqnO5A31BQ8Y9LN59H3UFamkKvR203pZGJuYfQAT
2Vugt6OaJe0NoXiRa9iEmraGS1tHIjYmpdljkBTZ13vrKjNVc7yCYIisIDguY1P9pDoDui2frA1X
fQa9yKWPFe0to0Uacbbv2Gu7bV9bruXhNk5nNI81Frs2DlGbsavqXzjtXdFNunL3k4REz/c6ivtV
yzFhNKycvGzm1Axbtfn58APzin5tarQaYTcqqApI0FY0QYAyqzwmKQmPg2IdeyHXQav6Jk0tWaCv
TjJvEMkbpeh3oae0sboaI4IVu1S7PIHhaizWtCEX2QZ1uMCcwBWEXiZ05M4zO9sV2KUlO2l2AGv5
HLpzJmY1n5eoHxk+equ1kqDVGHgKNiJcJGjZ1n9ZbyBvCYoGBXt/0uqjAw04FhfjfX97kX3uPMrz
2MkSp68i2Db9EpfrcYkCyE71HQzqFkai7lT5D5e0gK66nemCpKFj8UJPWm60qmhVFAbww4IR//16
P27+xTkHG5Dmg57b9qkDOmMp+a8jonhpVnjBJKAzn/EpperucV1QoB3IJd+AvyIRAxSE3qZXMbz2
pS3V3Y4TLNqXxmxEOwKTKz/Tm+WuprjnbYifIeb5QnN0KQg+/6k/DQusUwXfTDQh8cEWvAMc5oJF
FkOVLIQDaTisB/ubhWfcnIWm95pZSGjXDKQUxCdywx54Rrkbpkc3MXOWupJxGhOcdlQXUQoJiclN
907pjkmfOqangERFlJhuOb7HPKfn3RBHsezPPTyTdv/WyMBsBoDDbo+qKFYVze287ZmGr4wzQ2Ey
ad2t/8OdezhgHFwm9VEo3YBDfzFCSFc8zznS5tx5ZYUX7HZWYFnUvW0+q35+l9Ttk42MARsMcgAE
4Po/dbA0UIVHCR0cIeYlyc9/G5Y0aEfsGaRY+LrgYJOG/JYJoWesiHAYOwEwkSmqs5plKOTUhhVa
3J7vkuEjrHZ0yNNlGAN74av+V4mX5PkHGVRLRMU+ANoNW7zgn8iYSAzwcH/XDRj6YHEbt2PyQ4Ja
70+a+DDLq9oKzs1EUwp06WEv+CZpGw2mPzXWE0T6NgDf6/zyD5nla0oGUyvCUsQxxsk/w6XS4DO6
X1v67Z3xdJ4s4H066UgJ2ASeDa/cjMUDj99Pjxi6aqwmJRiA4fhs0dOBjHSYpC5HI/gh83tPtIjF
VMJnjcJtNTGqqVsm/jOpLmNlFPDhjHYfW1sPH+45ck06H9Er048SdopsQhqg0VjGScf9C5+2gg4M
YfES9T4RTxVQYMKCtNrjti3S3ZOw7Y7IaTLGjXgZhJl4XPFChEUFvDytFuOD92TNvKgd2aNO+7NS
HOfeWKQLkuNLUnaHangV+uR0wYV4ODRwtrsSFKyzXWb2aW5bMlNfYwKpwKnmfcVtBuMKqYGz0ciE
Pa6q0KgqANWRi+BXuAv/lFr6DQVllF09Oqhx2jmZnCyD3ZmI80p5xfNh1Yh+jv9FztQS0lD9SKsK
jqc6Xr0eOF89Xu9jON8fEBae1EPzyKsIaPT5XiQQcYLgMDY4ClOQLG/+3DjhDQk4PDagfsezC8Oa
BQob2QHLdUfFqChMirzZo/cqnxcQawdlkEhjIfdosRORc2kDB+9pT4Nn+huxgGMMA2ZS+R/Tb2hK
Rfy4bm8uB/yi8E/kUbuFfwmQjCNPOS1GcjwCD1AJVJhvB6YIFaySSaTJnKY+7RbPQpdOeM35axdf
RHiFKhQ+gDUwXeh2gZYLbb1dnaHKDxITJO6Rk129bIMlXs2V6gaXqEPa91yjg4BSZQE8LmEprgt/
1z68aGlCv4gyJi0nxPM5jaffJ4pfR+3LiaY9Ur+f0xTIRxGdRHa35Ov89J5chcXlsz1Fk5baoJbh
tYdtm8HOMrmvupdret+8JSH/5FEYJkJ3knQC7wL+Xn0sYh/N3XKkG7JSk7KenXOhcvuUKPB7Qcty
i7Kh5wJI+dQTVV26/P0LORBEtpytMPA/ZaMsvQl/fvMpdbWjOt46y8tW/7Fbbs30XZtQwfhOXqNb
dXZcHFZuaAjsIsijTIk5Gmu2D5SlHqbM5H56wBx5L6wLYelpVFo96XRdeoQwWqkv3bFXz+Uhscaa
mSUZ+2ufOiT7dd3mK7j6gGSs7COeK3Vv8c93nztOQR7vWtFBDVislWI7HKCKFS6qtDl4NMt2YLrS
FwzTA25Ce6ePYM4/h6wF5DbmpBpUATGN4YGgfD/VSMGbxPq7XzJObp3mLpkuhtvJmylA6sZEbBnf
YaM9MGLQlSzMBGFxbeGmBMiA6P3TekDmaLyLgYV0YArXv4G35eHN23lDI0dZqzws61BqU01piv3r
HX+TD99E0z57IXuz0rsk/Wtsfxb8/QWAIMtXRQ7Y7dFimL0qHZGmkdzGqwIblNcY7iIuF4Bwb0Xu
UbFbCSvMJgE4R/CSijAKpw25J22slQ5Z03uxJSFPU8Xs/Kf7Dwl+fuScFjYb6VJm2G2eS1dc9Mu6
dQsIqJA2V3/karZAkYaCt5DNxIqFqctahbk8AwsvwiU1Xv5UMwFbHrXMJld8yZv9JP6T27ERdfMq
zjGBWmfduUA2zCvcDVL3AaD5Km6oeinWe0hjdh6vETGq501kqRcCbKB3sHzgvNvC6E3k4KzK/gW4
4uhYrEMkEsJ0AY66i+s4i5bvK1/K8075fYXcEFSkzYrI95/8XeLmXZyldeO56KgWCtRdCwlmfGyJ
gcbevdIPk7/SzgZZeoVXJrk0gUacXvBzw7hrYPsZoHnr846pFnq7uNTBkZCt3j/4qpqe0Jd+bpua
th8hprtFG4cEgSibkWhVLoaEmMNdEYT7lVerQhF3rPwSzyniYE6oWVoqhFNSJHHv5bh62EZVzZGg
mDh5+jwlZgM5fw00mxXfwUDY56Y+lVYuHfpyl2s7h3jtzRsRl2/MrUK76blRR87NFfu69Bhg1sbh
mKMsoNhxTCNarDJ0Hi07KbwauS94XuvEZtC2qECiz9ozq4AsZB+slelDjkJ+6LyuGbZozyixCEvF
OyPIvtcdWlgg8kPQBF5T95I1fjuXdOXkUrMyHHZJRYm55k3ZSImgBA+82T7vDOH1Iv11cAFluTmM
lSjO2CyBJ23zMXjfheo0aQuE14Egw7/admGuhG2mN3H3o6Vj1RHpa53fN3/YdlAqJSJNQM0rXCaR
jlwWgyGxy0AQuAGSYZgZgEv1d0+t1M2kHzKgBMxAYNBkcGxMhmgtUtdPi5of0j0etGXUwjEDd0GX
9Apn9xPA3X9215w5sU/uu6uFIWUzyuNoDTxFlkdIU/wSr7ix+iKMkXI/PCvMMq0lH86AGCoiNfih
uEHSKIFMZGidxcSecxl+ZDN1PD190gie2BHe/XsbYsSs6AexvGjBZk2cpLgSwxjDFzHv/JAztLbZ
AgzJjMIOoPL6CME17tdY5nb6N2/vKOdjwPKChTi+qv4O21U3qRVT0ln5oZhIJ8Udhf9joVaR9kkl
DWstqgLn9PZs4FINISiHoX3uDlZqV+j20gemp0pneYE5uiW5QA3EMQYI66WB8e+WVvrCSniGvUtj
6tuZcbymZGwjT8TA2yYq4RROwakfta+aFiEdqOlR5Am46TeI+xbPnsxyEmAEwSF9KEGoUWFPKp5U
bIGoKFcBvfSTA2zvQhi26HuAyXb+iEATH5ZsbU0Ih58+ZQvfsT5QNdnJpX6HAeogM+s7wk9EhkDp
XXMXatDc+ReNt7AgV5KAKop8uARdAwzMknXmYWg8ND0VbIk45NrEnKrWmjeRT2O+ATjQ4LO7D2TZ
ixI5HCTX8J3wKHpXZcFOwFtkyBjQWYj2ilVGTAJFXfo/AGpIcXSkaPmTl0ZNuAjTQBtVNwK6VetN
gvO5SF28wOXLNHsOHxHIO2H3pW1KejYBeUk6QJ4ELRNLrzUdDLYtN1xsDRpLp4F3xuKkfy7RARM9
Ng7uZ/IoUDKo1EtK7LDh+da42D8f+k6jetybzF4CzhN8aCh9YQGtpuYqOJlHTf6YLq3BN2GMQgR/
jud8TtCEe+bowHwNzNYk2Uts3PYdjhzHCirNu6Cm6LBbCgH2+yjc+Azr4UDRkznVxCjrNDFIobPK
FMDjlFO3y1+ZCQeSoe3lCxMnV2jWkE+nVwLB1e8Hj+r4RiZVH/cn571uAvXaGq5VBiVmJPuW9Ezr
zVdZLEThSM7Br8s3pNJ/n7HPy5Fwep9Ptu8T39/ugxVJjjgRWh4lxobxD6kDBPdGfVy7WSvo0t93
8GMigLUUPyc44me23NSDdQjhwFbxXCH4GmEflhK0kN90aaVWCUZoffmQsWSTW1QtGGPv2K8NQTC1
AE+vaqzNAT+OxhQ3KOwT1ZTLAJ1EWcFlHJ67ZLG4dwIIezL7ezZWKxHGUfj8SmNMFRD/31F39aH0
llGEJwqzQyfypxJ7jLDysJ2iZ81PK3/495oznzOgNwNKIp46h8/ktPXEDn3Sm5uvMz6Ow/2ie+WH
c8bHE9EUq7Jtyy86hQTqHdCZI1BoWG9DlbCLWY8kdIV1KvDD5Yghv6nRPfS+SXnd0wjFFaKnqsGB
i2MTQYLkDrDDJ53DzU1PMSwPf02S29Ezm/GSiXE4ZSPhK0KaZBNfzKO1pF9HGKa0YqLlVxFe1+FG
68A1c2tJaitgPeGnzRnbVbR1zLbPqmsA9mRB4RMI4r4Cit2VLd4BWcHCGm723ipLYsKaakrrxhp4
1m9XZ52zA1jf5hIq/O6t4RE4V4u78OM9Pepdc+CI9gga35UnlSmevYOiWJkSHomLHbEJRGmZqVfJ
K7NhRCstmzSGSCFSezbBu8xCOVkUVoe4NHUTf7KZcCMBDY23MRmP4hmR9YYtuK7pWpB7ka5DIqze
wjKgptvJ0nGQS/MndlaowE6dlMAQAhqyU3q1o3YGKyfKcgnOzQjHAsp0oX+k+cbFb+QzGuPtue/N
OxQM5wQ/ZMQ2BNZwNvj15+C4930imsPUIv2qQnTEU6B3hG2w0WLj1xGcyxKXUJ2BTcMa+RLWNu1I
zncGdsDav2jI1whg8LbvbM+Ku7+7H6cdK8L5+9pGNRT+CozWAS3PlqjVytPQwaf4vouPShQ/wvFA
Hb2EymB4EapT6gHdNWBTyHmaGV76LHcV3G9/NII/AnogHjuVNAJa0l36/paDyyeorxOTf5FFczcM
lQHRZ3irHl7SEz3kETbAg+1X9scmwkc96JYfYEyvL2pu6hWFgPMgVmAKUT20adsWjX62tf+g7fw8
V6Nqrd3cITlLdJGBsBL0EyCdvNZAfJFQu+Vd7EDV6baJ3CWUznfLgMpM0cYskiJpsCF9bnJSoG0V
439DHkhxdv2BF4+x2s3iA2p0DQEl0qqUbodmsNYGJmZd9e7iyf3xj+fL8LBC6WkTDoiduI09nbbe
ENENq510r3Wtbk/1oubrVksEiE3EgWnElBrQ9S4xEXvxB1vMvRAlZ7HAQfrcALp3f1bNmXRFXt+V
szlXWbOp1SsSj4/GOopb5pppCv8g/vG/ZTVjkpeLEifWqptFeNT7nV7vZXrM2StaJycsRYxImigc
k1OGIY7eZqOxn2raCp0iYznlo5jBUwZlH5mOkdPAcVvDIU9ifhkZzjMOvsX7Ei/cqk12SvkWyTvD
QxKYn3Ho8T4I7qh7KBR6TxoMgWEton5GT+bGN7tj78rIWAnwK2q/7f6ecXgexYuRPvs0XUOyoo7W
JsZ1qi+CUIwugGoarpHI2wvBcxDio6E8N+x2T0TVPSmHX9VOA/5ymCVropOesf8B6d+GJOGL3N9C
ZquAj3ia/bCIUH5br58B4t3M9C0LJuCLpjGvnqL52hkJQofDu5qMUyPG0PDwp8oW6N1JMexa/13q
0i9sEZE1c059TYWw19Z21EZ1TErD8ZgAjX/J+NG2Ucezc/qk7eEFyXCLVnzzOWpb164OfSD5Cu93
JBJcbcnBw0/dcrAZqiTAaWHW8F7XjiDVnkEjDkBfcvL+fBVJScIONWzrzzxQjJxwsZ8PUiXWPBYX
okC07tXxPhjtT+N4TTtwqVOUcTqlysu7kJ5tKQxI7/OjRdL7NzDUcdIFB8CaVauVcawnod80AhwS
mi/DJkzDwLw2ybIPDFWj5uB4QIvIg2fFEFLW1/RiBlpejfVTNsOP3dXFTpSiGkLbitfIRn+nG37d
6K/c2EktwpsdPakS93xfwYEAjDZPpAvIaxhNIz8Z6tep5ozVKouIFlOICEjWvb6J9/nrdDayCVGR
sJuirdZUPhPT25GsbEfn3V25eZVvu1LlmkRVFzYeHl6hNY2gLejNJFBnmukwJDfzZ7ttZjxzmjYi
4mmNcURBXQrVCkqNKoDwIqDoV+ZrGh4sRo/+7Xh4TTLsAmhiTE8C+xsIgcIDR9q43Ca7oG7ABjR/
rJvwgZmWfsK+kEcRoF3R/ECOEbCAiLaTmwSkuNfCj1EDHjiL1Zhd9enVAEiP/6k9Xq3wNlwPBZ6/
2o3RJMNMEA5d/XfqXgN9flRJhSbhW8q5inJH1nQT6NSHqDyVpTBkhJGyVm1g97TNuyvcFw5hPNYN
IxOsh6hi9s3UwmGwU6ul4vlF00mUAmrxVSnPAy+mCKYKnsTvwza3keR6XcCEf2RBA+Mtpv4u8SNl
UMCIvGRY2EgWw7f4HPrOsN/2mEl6MG4NExXzZhYnCUtBNIH9BGyCZ3YFG98Mi3828egNBdSQfi1P
TOZEx5nFLo4umO/rJSfegMyWkCGO0hGcUbIAoSeHszVB3Nc0/uQ/6t5ayk9yemINSdtipaTiEiD7
IU9yL/6ekhmIqpucIjw1woD1dZXoZ7CnKMIo/qrOVOOYsWpZzOLY/QyaVa8Z7AGYh7z7ol4KV2iv
hHFbLeezlh/Z8iG0fY93BN4MILnX+1O9+KweXTOtUG8OkeO30E2FOGnegdJUJJxNu+svYmH7shFV
SslSpTaHDUsdjxhquY4OcdbOpsFfH2+4Iimm/8tEO/x98lM0VJrFd2qnHcm7u7vJls0NtOViqY4W
6PE/k0LO65dBRDnnqp0+0GqadTWuzJLFOIYWmqbtoEgKLSFv1ilVzxJ3Ov8PCwfB/iZM3Ag1AvF0
ltSep9c16bulZVNsc3+jy6cZWIMYG4GPNHGPRQwfRShIzNRs3w8qEk7KqoxCUt4xq9CUFaAIlED+
IDgRSnEaoDmpE4N+w2n/alegBmgjdIRWFW47iSPL0eqJG5R0DfD0LfRDxBLPtYJ4kHgVV3kH+XEO
WaulayFib7x8ClNdODG3nmEqyXBB5xAu9q2jQtWsoUL3MZ3GfHbfpZR7WgZH3IS/XFfOHhWL76j3
WAdMxHy1bL3SGWqbwyr8E5q1dTq2zVxvr/FQtmuf1QzwfWWVxiTyhb76H9ZqKxNomADiSoK1bSfo
MPeJ+UK5yqWO+RNAoYh9ohcQSgjCmapOy8MpGmUXNZ+xsNSjiC6e+ixUe+IUMRYWEqaoS3uETD6l
cegpJEt18QpvO3jINss3PrVnjjQ7BkmSJK9BlKdXLa1P22WqbB3sfd/Px6caZSrD31O5Yqq3Zh0D
gnuvm5cY3oQL/i6z8otGasa1lweKh0j8/MTfxtq0xfntNeaIm2S6IMx/Pevq9+M9zR3Dl0lM2pHj
5aHyS0CMQAHlGFqlE0FOmvLTAl0bn2EtN4uVOe0a1SVIAuZKnULw8UZHxPo9jTbm/W6jkFVnsr8Y
4QZfIEhRaFEzmve6fYR0UPhk4EwpFHNaVgk/RyBVejRQUP0R+aco10Y5UCck3hPyJCLWMjnFFwa6
NQBkogeg7p3ozU5YB89+dj8wkuEpd9+mq/1u8xuKnTs+JdAfVXTTe0AzoA0Q/LZmrbMXrZcXUpBN
ACFOPPHg8JzpbddIGhJVwJpYO5J5poWZxncYJuUBosEplIKs5bdPs+UP/fFObcAYiiWei/dNGtF/
38XFG6vZtBDzm9DAcdn315YL+wVosgo/lCek99HIEdGsrGWffX+X1N/SK3DSmAtR7E/wPO3AJJoz
f47xddiuDy9lw4uikm1kQTSx0g53BuC4WXstBG4gkipfAi2E0Rvrxhuvbl8jtY5UeSGOSjUOELFe
lsj7URZutKDXMetHVHeRnzJ8Tmn95FY4L4ODfMIYkesW5otgFkzeIcYspEXY2oBrA/ffNL0gjztW
EG+ML0CwDL9QasMlRqsHAx0YLSZ7YLx8gwX/zcqhqC7lfzcacay44u1bc/RRHUHUf5hm4srIuifL
v+onaRIFChIPjRokD28h7UMkQhD7VFckTU+qCbFNPPEnSHE+TQqSYwqGzc+3RxuAqgT9q58OQQcZ
iY5oPhHgChoZwHn8UdZctenaIIf/bVCR1tuyzZFezODg17BWrYYKDjSj98DAKh1cnQwBoUkx/tGv
7XubisX36RJLF8v5dmx9dYRqjBS31FHLmkLp9l4lajllsusjh/ZzkZf+Ht8jLSjwH2NLn2iwg7o6
uVL0zKFegDSO8b81jlVAVlanEZPgnx2CeMdOVTptlz5M6kq0bLmyQecxMFJ+h1NGN7sztTWN3CdN
0gJwT1xq3MTabV/LPQAJ7HZRWazKTbciPKLZ4MEICOjKdiA09aBmBD7fTynOiOEqY1OfbldYqzzw
JaRl/jHw9Er96m/wuyQYpTNFhHJvVfe4qIY3T2wWqNHSb5C2gTlt8kWZIccc/yxY7RQPuMBQFZYw
cGBbsIESrIySh/UbwtjGOq0yHV+6ANT31aSogCywyrydieINos75hKnu0jgoMbyDMAi9j0C5zIUy
x0j2ZwguW7R7If0V+DqQ2xJjVilrwr5u8dg8sOy5T4hgorzH6XUcXZBaagIEnKkMGJLHlsxo6e8T
YzD0VVunGKQJBpjRQT/PjJBjhD4VyRjk6h5T4B4z0wXi6BBmjStY9+6Q0JX5zx3BJ/OMei2K39Cp
f6sgXDpXcwcyznHFKtRze9mUGvV3nMIiMO0mT66kvDxvERJL9Aw8hwvAytxcwWG2zaM1wsFCTiD5
8aLCyfNhvb+qageo1ckK4Ty19rjZnvR35drBiRjmTVp7HQFfDCGA/wKB3w7gI4vPgR+0dN3TLL3R
8NFYhCZvrnfQ0hLeFenYGJhA9sBQ1f/My8J9gqgexkgSu0mnxdJJCPsbGRmVJkM9P4YAoJOO1jL9
azagO/dV5sB18tL4imk139JWWp5mYKGLSUCZwKdNcFC2sn+RtOEi1MBpUVIA2FnrbwYgYnOFJBoJ
tkD++2jUpkxWGWsx/6s2egomoxsC0mqCpyR20x4dXcxjNM0Y+ys8zeXIz72vOtAt7bVYHIRDtVeM
0/4/FtuOEWeWLe22gC3Zzyhg+VoMwG2JvaxXpZBOjmv9Rladtdr6mieVMg6TOWQOQ6xNFahTKBri
Y9ADueRwl7PYJoVab6ZMi//cuqYsmVTmRGoNVv3pyilYlwfRUNxZfTMhD3v7ekedSpmrYCXgEYX4
thX4vFCUdV16XbGWVMigIAaEXwHZPHZiOgfu2tGUmuDVaTvVAZB726L0mJeGXE+iqOV82fje+svN
9Mz+NFJOQH1Ap4LVgdrBYQNH/nFCKWEnXbKiDEU4usA4Hr9W6gnLLv1lm79bLUt/hCl1/lwER6qA
B4GcFC7Ql7Xs9HvJgmjTOs1D0lgDuVD/Hdh7OoHz8yAzbLzoPt244JcVhC2E6PTvJtjc5gwyqwC+
iLJdbiP/s06R254d2ReOx2gmZuFPqwu4JChDFk+wZdyhowGCF8fw1yuK3TG2lKcZwSkunwvEW9bd
/Zqvr/P8PPydJCXkrVRv2tnWcBBRKr9SpnNoLGHDrqokfkJJEPRqiZnaB9MVSjefZWNrcvHmlXVg
83TVudK/GatLbOQc98MCpvnTCWYrA0kAMYNMSwarcWuhT2LNNBHNwTJIFGkubghV9ZFl0xXrCRGJ
BCnBqnGTqzMfZqLvsc75u9p4vfckI0vxf8WoamUMV/Qq7q5XiBBJSuy8RIo8JJK3vDxXi0OItXrJ
/xgi9+Zg3QPoXLB3gg2Cf6pH+XSO7WHlxAX8l9qNERyakaF3EqySDmBVbnvdflfvYplYZRDautyg
iSMH22IPCfITOsfgRwyxWj4NGOF3r9KimXVbXMbEJUePgUO2UXl5RrfX/5FDAnh/YWpuFhmQXeFa
TXenA0D5QiU61+89h+hmjjQywOgi6A1yNP8waRj1gD+y5fRoW36ZwMTpvYefBzobkWjj5//XwCGZ
P8DttLn2T8Qe+RPkk/fS8AmgJG+pj9lSYA3eLSbG8ne9kw4dMoe8yvDhgG5Lty7ZYkAjtDcix2Rk
rFCbOy9mi519IA5fO/toJG7U5qXqbmFVEfBVdISOCpYtUtPhJ0kkkDL27ZDSBh4FTKzqgV2iWtnh
Q0RyHiA4okZUcvnbEfDIqmakEITZ1yr8WtGgv4JblV9frPUVYU9QqzVIwW9uSFpId5VHa4G4PKut
h18Ll9f8S2kYEYEU4hihgegD+O68aVXO9ku+trmYdAE895ZthRjAKi996pRjUYW4xwIG19zYmULw
ecYZVLBZtfFXE3Q+QwcLguylUd7PYJxfpXWrqd/1P3HmFIPq+T0bLi80z2KjvT3gTVM75g2LAfJ8
R+tmBW0iJyVKcayjcyGbZBGV7d3aPhljcJ5cLhSaclTMnG+K4dKnoecTqsA6H5otTJQtkn15bUhe
QZV4GX3ynA4nz3qNnA73A4AvrKk66pQdsiqbtoZU7B9MrdzTsmH13ij+0JUd7BqE+XdQ1QqKzZJs
hB4FS7zskrkFFZx8i/SUJe63OYJEXnlgw5dQ3FO8hrccdMHeQ0vMuaIThoETkfDsCsYDemSNc76v
UmlCjnQ22CcP1CqQgJTQ4nSrAgc/Xcbv8TSDNG3LfzRo/sd9zGR5azl2geDLsdAQdnB69PLEiIYU
jgfKFlEfqL7kpiS7EQt8WsUn4NqI/WBZdqNuzBH3hf4oBI6Vt+S8T3ZyQhoPKUvKDG4SjSCyuGbK
qEma5n7VTnUOUwCQag2ftlTk/dv8oV3usjd6GjPeLvZanuwyKjstAwTMSHOyh1XbsleJmf/Y9Lbk
BZZDT4FaKo6vHdtJ4sTo6xZ2VJ3SHiqy1banRQBme0r4yUev9p7M0cRCd4T9qOw0+Dr08l7SI0jb
8NyfVeR4YeJXpkosvj21a3eMTJjlr49J2j63Om58ye/kId2cX3uxfdy5kDJyy1I//Q+1fmpevYew
OnVjpuxB0XgWBXAzqdPmiFMRhCgEIzgCEiBUStRUmmuINfUcPt9vaCRBOUaAaINvqUF3uIVpabZR
wzZTDiB5Q/jep7Dk1WYD1wF59mKuiJIKaZ+atIiSNIjYco20uAvWXt5HpnCCeE+awhPi8tivBzjM
GbHymEWl8BGtzFdHTgDimcrFlkH3aBq66HNjgtwTXardB9+ADoeccz0w2VthPGXeFh217NK1lwxg
y4rsJFpCdsXvc+M+blPRJoCmlkQoJ18TOsAwnAJPCLLoEPoGxnfSTcqa1MZOl2GfiW+61MY3BUdJ
03KNOfmj14QjwZYh9rJzX7G2wkdOaCauv1QQ+7jvXX9FVMu7KNXeXpp2zUTV/dvtPP4TgBE9GA0K
IWcdOBQddq21o5qnbR/uVToZfcK6tQQ0yFq3JMa+PTqK4rHD20wDZoWLMKW/vppPFJTjK0oB8WY/
yd1anyc/EX0WUfI6kPr1+uACdvDwl33TE3zbMpjF7xVBMazSEgtlyeu3/cjnZ4thUyZyyNuCTVhk
5bAKujTasRsDSRcoUGyvh3uBCfjISUixTd5CJ4ReGZZtxrhXoi/+LFHGO72iEcbtGQO3QoDY7ifQ
l0DUktCVlMT/lhFJRanXIz8o+8Chu4++Ce694x1kqUUhG/j04rqqrFbxqWeoMAUp5lPzAPlJot8T
Kq0Kmj2/ESGiSqIzDZUTyKK6AX0cCG4vz2s1QSzIo2c1C8spkN0k4U133MWGx36cxVQGIR4UpHn7
GStJawJcOAMF7YIIPSehuwuk2GrElCsTkCHg9L3ofSNKlWGRBxHqS4IGKjsM22Lum7WD1EMeOTwA
DER8y1mj1yh6lhTPijAW6pCW4M/QsGAXKYfzpimSqqnhXAgdRDenEgEqXw+pV3jRpyVZlHmXmpVT
t+jq/gCdv+wFPdPqRX51gjo555kIqihVj3e1k3Y44HpntpRzFl8a74dRHOMtMLZxEHxz/2uP/3VY
6G3enoyoCHGX64cRFeh49tOWnAWUH+CRCAZDE0J7gmaFays547tJh1yvhJzS6hsg10Ajavx5dlE4
1wZscBDtdyoQkM1o2UXpNa/PCl1ZrqFiURAwGtGkicts7ltKo3WjlB8HQtGOK0HhgM+Yz1L7YUZa
sGSY0McWAv/mIVXQMbBgQ4qyiqzbJCOxyVr0K69TMCN78G4les+2l4zrea5VKYALrxKduQqw2XZ8
xeiN+e9flzalgq7s76GqLNrTiyhdvSr96F1r7T1b6C1D3kNc+UHjQcnr9m2bgCiO96nwGhXEccci
zbj8m1cVgJ8HFHxekzsfgkfwuWxqgZqrKlOWe5wS47+Q+/xmSn18GNqXNl8pkbBOYKLx/jbZ5VPP
c+5mpAmiwh2mGkmT/IV6qfWvP1hYaLatLdwDVcJA/QSXtzuClpEzGw+nikfgiIuDv2sYdUv0z0Hc
nUbUmMGjkBp79kWYWqrxq7lRKBHwY2Fc/zA2J3tw1blgblekQOytbZciEHEh7yuDP4FflfRBNRhp
yJphOFSlr39qPJqtTKRX2u9cAlax8gA6jXf0dCY4ok/reWFZ2p29twsvL3M4eo/ju0QiYMaFI6in
UA3ybv6X10yaglEThSjTY7nsMdt73ekDJ3rive9YylVkLTVyq0xao37frz258LFdTPk6Bl8eXXfr
BzJLavGic+QT8AdxgnO8CDMNFCyIj+XTlBiey8ylMqz+17WvOGGS1NQ/LMxd2M+YwtrmLBWRUzRP
voJEh/2rzErfejhiShskF0hUQnPKvT6Rz8U2H4f16zsz09+iN9jlfxZJjHsTPW3jFsyOBlxvIJkv
LnseLx/9H9b9RLTt1wdmgn1xJWQq20S086H1WeJmhVGyyuCBH7/1ki16qDdNcbXkA13ipmnsMQ62
rhspGKp36mCvo2M94zsqVfASurByQpOFYZKJmOUZtN0lp4n93B7WgwXmPHfEPdTI2GUJ6HIvXsIC
uwTyzFKaeV+GVF9Y/BkOVUSeWdeB+0Z8hJjQgU22ESuy9H4j6PpAyNp9OFvkJClHv6JPu5oVExOl
RvMbKWlb64shs8jRKjG4e0K4xZ76AcDxcgNA0iYz2fRNxgxa7R8u8GV50FJy3favKAnYTYRQ8DsX
Tk/MQB3lV2KZ73dV+xKoiI+d7Czkdd1fpbpz17/DOzY1+bh34Cb1NADMxJVkW9NGXLP9wfmOEZuK
lMsBVZxzu6vpg3TQdo3ZYRtCVPtV6ClMBida3GYvAae1lxKQdqgg8LsuOd193A/6klUdKuwKNAWA
oKw+j59IvcUN23DQAnAxoDxHSodXl4Ekyg2TAoqXHN4UXozAdNg+lVOzNB5ejByAhRmnPnPH5hvu
iPbyQpQuhZzxDCK2B+Pn7rSm3vb6N1PnrrEiiHc31dEG81SwpuLEKTGcoLiCDF+D8w2Hq9kEBbfA
stpGYJYEgUPAwq7mT1xPTdHUv5QZp6yFPNQf2qiQyzFeNeyr6qLqbQIjwwy1HnOo6h07fD5wzMz4
3ZxkUc3BNdVHzVsak4C6KCtQhhlO2AS+c3HCIJTeeuZF5DAFG73CZ1JTOTJoDjWmsu96fHDncLic
lET0obPk6DA1RD6Le1Dkj96AWJfieX0t1ZsRRWmE/Wq2Bu81mWTnD6EgUXQwsAM+uUeNi+mdziN9
QDNEEPHoO2k4IzkrU5QdcEDY3Kwi15Gf/jAvC3W/lpJ27yOymEDAOZgthyBmMl7K3jZc3CdBY+8n
jnFuY7F5OVPKox2XffGu21CW3y+y2OLr5mmWsGHUxriBiu45QBdUqh+7ua4JsbP4ZD78/U1X/lCf
etEEEnY87pbjXKjHC6lX0OmJSpjpNFLgU7M4iaRe2CNV5KhU4dH+TvwKpnF8S/361VjKs2+FUrgY
wQeQ+p+MatxmmYrFq7i40V4cxTts6FFI6yThSNh8EVvPlGqfer7uQyracHAI6cVOHZMKaYnxHnCe
YiOKJg3Tj01KnozizidWNQ4+NhC4Y4xcUzNYIrGY0+eTqMjHOSbJVQ9kqmAeoHQXEQwHViZcZw9+
GOApfAI8l81wTOwBPCNY9fqlbQeRwuFiNEcNOyAi/9Nc0i217l9otCkWk1smiToe+RJZJEPmWPyC
0hFPZlbWyoaL/7Xw9o9ENH/1/03oVMToFjlPNkLiME2YewBCJV9PCazHxS1QqNAkUJso/pHwdjRs
9V5hcY75lKF2p88WFmVXSP9CSh2u8/whD1neaPT3dBMMgYTmTSHqsYqsuiSeIlKkZ/IgaSm94u/C
CRMwl+yiTAXEmz/LQk73VgUarx5UghPO2tLJOu01KsVDyzIGqrxkmeJzjc4YgtvS2Uy0wDXCt6tk
1YwbfHFpK3Nze9oXGpx9+fJA00qHX6Vn67Dxya1dDmAq8bNoan6WkMAoAdwEkid6iFG0JQpQT+aJ
NM7z7vJ8OIVqON7NVrGBEGG0fe9GBeTx9IQSQ43RjbgqiymvKm9xslmcaKJ0iA0YqGrwIsDEdQ8t
Xrx8mD+n/KrBK4hDLeuR0Tcj9HW1hlZxaZfjDkB5v/Cs7yY2fpPupt+hAT0DsuE/FAZKuo0/Nr30
7C+O5tlVTqS1TT5Ot7j5UEqLDKOlP2o7G2jI9xmqYQPrVJf07XKksiFHIJktfkOitpK0tFo1MKnb
wYBE66RsmOcs1/wxFTBRsQoFkwknWIO7wfNcY+gzeMUd6Z0fGXNqMXDKZZXjZIeN99ttki3gCFoO
qK4F7d98bYnr3mLwiIyoXqxbkBzvybU4Gk5lDWjiIf2d1ttlAxQOSgXICoW9z2Tn9+ZEoB5XHk9t
Ie5Fc3sULzOS9IkM1WhX055mrNNuRp8qQ61cfKsQpvguDlMoXfSRJPeq9NDuoNRxhJEWmcRKXYHm
KeVlu0HrPRpNVVfGFb2dQdIxpawh21LREdeMVqrxOvhFtKXAT6Sv3kZ6wNtnQPNI3S073XjOcD/Q
tSCBbiT6T9fprX/e3hIF124mFa4IBYD6MiPXruoupbFZsd7AYg+un3IF4driRZtVLoLBycrRfart
w+7Jj7YuFLcQYJMtl7Ho6Bl10TwBTt3owvBFrKWxN876igo8kff29jVcTCHDD0/X1JmCf9LJvtLt
zfURgBOXnSsPGrxwjgdYOF1nWtyCyzALD4WVPmTNmMUuSkKHtD+rfOiZCgblDscghJAvYPF/rjXE
8NfTYi3dE83Pe3R0dRluDt/EKn590mbZihVLRWQyIFmvGCYf/9BNiErHexk9HQZ/ftXksjmt8gH9
X4ZY9GRPendGC3f/ho3BwVxFoZjL5/3jOcjVq3EYGQojhRIHghhtYNNkbWpoygOWBbzywaNNyLxw
GjPb21qWzbAbkdvSSVLT2XC2x0UknROwZh+mB85/2SRsBYUGk7P1pBbpATRtwfFFtjsMIXnnNcO7
EZkZ2T41AS0vl4BlxOtIXo+WHwinFJ3keKK+lLII14b6iKSf1hBqLG3AJoiICWMjQo94FcMb0Ysr
wyckRlIaqyruOF814I7ZF6cQ5v9nA/CyLpy9qQNelvASOFqbFBDcGaMARLzwUXP0dYTLF37v2CT5
StdOld5Jwp3RPGqoh/Q1hacjhvJPX3uP2dJKMV9fiTR9tws76j7nHN/4e56g2biaBjvrte+QUIAD
L2O3BsKz1U1jbiu/pvxNoWfPHn6lVBbUB4s7mi5CHToGNz/1BKLU77vDHxwIBO6FcDKhNwqWl2vc
8Z/x9PC4Qu4J+2hEc+PJpPAdugIW/NNwFWAQ3Jq1lWITzjVruQi/bdsnt2JktQgKG3xCyrmf8nDu
hh4h2Zzggov+6aFKrqzEiGJisfnWwu740LO8EaIuDi9Yo4SHTSvCgQbJCKniZAr0auS3Bthj6EiJ
AFWNXey77x3P9HZtK5QG+AEjCxlt5PtV1euZCkBE42uo0vrRPui7CVzi6v7nGkk0eD0dzyDOQOm2
Eugc+Zkq2RThChamngQz7TOfcv5049UV4iOTZ8Ji3v21G7C16UnMQynsAurTCBgk9i/2/cvWrYZe
mtp8rAi19saj+3OuT8fhlhpSIH6ueLxuEOquRlHZqmUDCnyvxhqrxp8PNCq9q5RKSwRBYWZwS4Z9
B6WG30a0fqAEHGGizloBk9Gf51/WyxxJeeiuo8v1LGO/p2S/a2tzmtzNoBgtl0hoffVEaQwmmw0j
PeuqwysMrRINtRFKCAniYvKbfn2WgHKw4/MKdO7vsbHvJtO9Od81kIg2fXbxycOBTheExEDMu6X5
8VwEc7B+lSkYBCYkkQvduyLXa9KpEElqLwN+Mx0gQgjr00yPwR+ZZwUD2V/c1YmMv4YSYwL9ziIh
cHxVYLOXZ+SnDQUh6MuJpdhMA+VBCWtY9HM5vL6CJNpYDumdARTP8crq7EBOAmBOhYs2bCDeC7co
y7+SSSEbkWPV5mF1A4tU+49zcjlMuGgSEyb4/u7gjsMNHPG5N3+QtHq4g2ZzQG2Wu9vVj2CRzRlk
Yc8wdzZpXmdOiK74eE2wJKQTv4rx3pViH+aNBLQVcoDajP49t9FXyzJg8dax2+R6v66JL+UgEVps
oLsb/jdx9TG58pEPnu6jQq87PkCdsKZoqrJCefFoZa8JmM/Zy6NoDUdKgZ3yQYpZziWEg8l2iRVO
Ebmq9vhtA0aE83At+ZBwERO12chk8EC3WjjNl5ezvfyQ67VfijtR44iiCe7K0MuHAMuXEl5+tc6J
O6ZRsDQpAHTjx8Ub9cTyc3pFBgJRPnTA5Hip9OrM2xJO0JDT+VQtC4qgDIb4/tvf3LZkq7V0iRZb
v2W4W2RhkmqIx/WojN0h0w+SG9OIOAT5xGNjAFK/2EM3O4GdxHQz9zopLyj9blxA2nN/7J+g2kai
2rQTX63m5zcUXmY0yXx91+4P36dpKklPVvRqqX5JwT7LoTrokiZ+hby2jEy/EQGViF5WgOb7VIrA
2xUodZz7z2GbSRcwl3gqi9k3Jg5fWNp7bLCW2JklnveCFpqGiyoMjhBYSWUWnQ6pc1i7Srnr65uH
dfXkglPRBmFhgf4GJiIEAHViYbbptqW3qYEkaUXluFJT4QW9wpLyHAqjS2ne+PKIgjGPuO8Mya1+
ZUU81rVTTzfx2RmpfGlrIF6ZenWsGJp72pOpyqAqfXArKnao5fVlgyKbbq+oUwpNf+AayNnJ2og2
/jremXL94gO+HT63ZwmkSf1Usr5NATsNy22XIgM+FD0l7aYZrKgX+iOion4SBDXYYygEhuagiJVN
NHAkPvJqL3si5m28arHu7exTG0dNUrKNYX27nsjBoKUZ3IvpKKBI3FjXJMUWU2sYE28tqVbvN/98
1oajhv0mQUZ1MNUE//mzEVjbzwtR+KSII2fT7Cyvru1b6kxbs/EpmeU3ySRjI0P4eh9HCGywwZ+I
Bfp/HOkFhMFT8dUMPf85G5nSv0PzaiGkJiK/caxUsw17JtkMaVwLdgcCzzvXZ5/qjFub13jpuCUv
GOHr7F335BzvAkFwkjbuzNVJcrC6Htsv51Q5z4B5TsmAyquQmqlZ1zT8GWceanUJW0a8A9bCc6Wm
R7+XGvelN4B7yyvq3m9EYVkurzh4suIecAolJrPcuroTosFdmsl/8TvIE4HT6bpG+eiBmRlgk23j
cDQN13B8375W87Tc2sDw69B4yB/pQfXAF8M7UAmBsZVOcHEGDHss7D6lHlDygXI3NrKQ6hPNGoyy
ftnV2hyTbPpgj+uMUVoU69Pfkekq9YdcK6yuTAQRyqHcE3zm4gXidgRDMIUxbm+OMyUbEz1buAtp
qZuD9iq4Lgjrb7hYB8MEeR2VQs/74qeWkK0b35MCF2XhmL3DT+ZTv2QF7d1f4li3XzlaAsIQJ3X0
4kwfV5MwPl08jfnH/tk20ZCTfGmN2AbUup1n0cwxAr2uLHuZ3UF3if6rNnUW227fgrOdq/7kAfNm
B2VOIqLK+QtfNPzFzXeOzonA/28zhI9/oHPsqn14TFgwEjLnVgbqolv8g+6C95Khf+LarfUbE1zS
t5IEtj64OkFvsYL0vHmsKf9kmDifxMMgUoiIn+bhfnyz/iWCTrpOk5Px2P8sz8przgfUcR4gsmlG
BLO5K32+3OmYrRt1rKhV9DIPdIlYgqH4tP6P7NDA8UjkT2nBMy1rgVnxUfGiwrpOkKatlMUSJYgB
Q7O7hVWvbhKm7G+eOzirWe7nOrxnlFp2KStyP9DqEe0t3RCELkjYA1I6IFl6W6QI0k8mB+zaR4J1
mwLdBVrvWCCW3+uivZ2Th6tSvqqnLzx/LoVPBYjMGog8a53+yr1CLm48WgbNRKq2/9iKLRPMpml8
0GtvEoQh5rczLKPPdP4tvQYdpDBhD4Lfma4HrXFb8Nzf/wjJ3fEK7Ow31Rtj29foaTWXwTPkboHt
I+R7t4XObWKZiVCJ4uYc6EhpyfDEG7kAVzymB+lKP0aQBj4XfU+wO9p8MiCox1sMfAWR5ZiQTI5I
XaJIL5VvKyi1zGBx3jYJCRV8qUUtilZnm7VsBs4RsCsksBOZrGEqk5IbRxKuIV+RMBClG0YLSirq
L1Cqkv2aEBtDgFZCQKkDmoeC/dUFTHM0CCGAeP+wUVyMYaRKc6kwrr7XM0W/2MYe+1HtIy2TpNOS
gStfbVB4Uf94+kGbrQ/OVvvVv0DofLkEixtdRtjyACmIf2o9IGS9ReiPYpPRfhJHrBWxKFYS5AMM
CWmBGKqn1S4ClURyc4hdwAkz6DAFzO+qjv2xjxHHJEOfgERai44yqkIhdC6sGVBDETd6eRRRS2fp
hJaklvYr6mIbIQ+qWkznBmVIhdO53JdbJvxwrng5ZbQi/sSW1qgSvTdj44oW7fFRzUXFDz/k8yit
gFcZbO/D2KFi1Ft+bQc4kJtQOyEnL5ol3cYDrJhpUJpP4wozD9qYM+JlthG8V0DfZjyods+pegVd
hsgKVHPcp1yzJGXfOxm4JQwK6mjQwWn9XD6RhJipHFd3t0Uel6OBmrsrJtgLU9MR/ebMvmCTVxg1
w6e7EjU6jLGAxynsNrI3lro3TKeckqnk3FrSeyJPFRwi/LYhperUE/17COLOQt8aIGOBItEnCQGV
nMOhj6U6Ez+H0y4i/+ZlftM1rmpBAhL3fQr72lj7l3zbdmPkGqisvb2ruKd5vHr/Hv25UPS7yCuO
V+1/4aKXCrLQOa7rFw2p6Xb4GWBDc+AW5OI2I54G+C17JUFXfqW3VXQ1DoX5EHKsLvIzgTPWQYI3
XSKtLwpk/W0+lfhWzrt0CNAJAe6u/Y3PmzqTucs7VQIWfIFEJ28UY/gRUUfqshVhnzjvZcTrDq9e
7uh1NHTVIKRf90r39dpF7qId9YaeLTFiTdQ6YQersuUvOjKGXg6x7cD+1rSFZF/GkpjHxVTQGkSB
JcivplOaU/7203OYTariqCOYv49K4VufacAV/4wsXj7Wj0MrUJUh9jdeZOpf0Q07buCg3cq9rBeg
X/zAaW8zuebCP3H1fafYKMEEnihhzthb0u+SnkZ6bqfZtrhj+KthHam02SmWaqAyGfpMCq2Nok8F
DoZkHNq8l5DniuEk88eZWx8YIK0caq4Jo6lRE4fn1VYosFERJDCq1Am6GYXBv9A5NPkY+Oe7FNhP
bzTVUZXrC+CH+dVcZ/LRSJv6HG2UMg1ZWYYTTTyO0/fK5XYNtUwgUb+hJNBrNzzAAVKfWsd/SAyr
bH80i8y9XHlHerkwIpWYIj/dJ7KJ2UpX928MC+q7sjq05KfY+tuR+mJ3V2BfNVtbKdB/DNG7SYNZ
jAJDAjBWX4wS1pvjCQlB8JPQL+CLGz6woTq5z2roDg6eREKP9pO5zdxZ+datI+fCeUg19C8m25Mz
/rzL6JZ4MMxfAnd7Q8NPbT/x+2OU0x3wddbMH/WaJYsPKDwb20O+WcZYMggKwTsyH/yQIGLNH/kW
6P8gwiVDXYTiukN7H4394c5srhjyaq5cZfhov+XMKVbmEHAuVVo5lqNT67k8MFt3rXW1QLAr+ENq
+xymuaDZOQLDL8l0LRj14CKGppWLcCBUjVTD06wLCThtNz/u/yS/CQzhx0EGIYFP2iIHd3pHrkmN
QtiNf3vJ+dYXek+zv9HrICBHB5G35YImfUoch3egKiXpJDPmtAmhToEZkVSWFKuSeu8RxV7fbVd/
KhU1tFHvYZXH25+YccIIX0wLOtTiarFKj/ejc49hM4RNTBZWOU96f/HcD+2xDDy9pQ5cPK9FhzcH
UHRzn38xSuozBoNoYTSkEh/gIyNLqseCPDJGMQL8yktrY4JefNtxgVEpNPfci4yQz7XN6+uJNCh2
bKAildWfnjoflgQHQI7hFJ9C5wiAjGX1i/rp7L+vKV4rWYSUiY41h6LVpaNyLMc9EjgLNNH9f3ZY
zuzC0yZqGpr+ODgQWDsS2p1WPEujLXjJXHXucIOCZUXwGltU/E4JZmYtBNqcE4+XqHT/Ln+2uYpW
4b2HXwAvsMNyHvgKtyt4dLA+HX+XYb99V7CzPeW3UyUURCDN/KdmmiUCWBDOvYrcHwP+Ph1KyEie
1Ece8zktch2wIo32zM5Mmklzl2GZqtARCSpd4ttuW02XjHuQocUDo/54tyi2SYWPBmqB4Zz4WB8h
GHZucnjaFEd+ppYkMSbqw9uASjL9PxBf3kAqQ1RKWa6yK4xvQkVk+mvxvI6E8EC4GYEfAVN37KdR
AFchXhOWwjPMs1/Gf/ClmRc0TmC4zP4jEuGxKetW6K0jGEq/ukZ3HUfARjotpOgymS7CXdiBymGh
Xu1b6/oB1LhVh78gKUb0lpfVJC9DVj2sXm1a7wFKWcg1LvKmsiQxGhEwc12Y1fUIdktXuqvILM85
BuGNiLrvYcD79EJBa1Ed0f10yuP6g5NPDMkobTM5bQsPVSJyZcOGl52vW8fSGZtfRob5BcoEzb0q
8pGuWVjTTiccCN3eCGGS+E3wG6zaNtyJTN50bD+3S7rF6lDI7OA561TZLecdk1ffuCi/gtuGd4et
g2P/2cd+3hjmwHpg6KN1kV8R8EbhQ70/bTyPMLf1J/Z0WqV/Qxd/IIp9g8WPHAJo87XNhxsPWBnz
G/c4KvHJcbNiuyogprm2Tc7EBauJV162Cb5ZaLKxj21wjDC235ZvRvzOjzMqBHkGBuq5Ojswhg9K
ofJyu3JSs6PuzO+k/A++KOKkIP49zH/CkkP4KvBmHoaD9MRj990LERvR/joysk4OazR+Jz4dyyJW
wjthXETlYJH3zU7O7ltpQv+Bbh4rry+aEM6wBIqVpvBnAkZvaKuTOiA5/IV0CiLUrpiNjfp9w3iE
31xsdls29N6fxRGaCnJa/+/3CYhIJTzwY5QXJdf9tcSsLPHTWFQqwxfxElHqqen72ifZf62CQd5v
XWRF3hEmQgF0MJMlNwhWLOjYUip4xnxo/VXl8uLumWQ/E4fOLfgsfgebInmBVH22piTL4J27Z2+n
v6JV0N8pnqgouo8QPETboRSNE8tMpkKeNXk9G8p6UpbBc/2c6UA6NdR7lWxCCZr9QtsBb+lHmLUc
zXTJEUdwqTcBK4fr3MRIAHYFPISmi0V3oR0kVvJoxHiXhyEDMKu6snzdUFU5090f4F8ky2XT2Pir
YMUsUfGkWaY1CVCgEWUTK93bCj6bVG+nErUHKTpT/UNifyRNqYcYkx5V7CZmwCOh4ilZLencCgE6
5tNisbuyMAV3P4anJRHEBpPNXKk9QLxjs1pLnRtmV+qIxf4gqX9BMeJ1I3WcJMaeVvshAT7EQaqk
snLk4CpHr013ctbmIOncwlJfvVhmLyluZhDif/fIjNuZuPv+eB7oZEr3Ehpent8aTT98trFzSxvh
MJ18nD6uQULZqyJ8jh3cOhc83voShAmUgz5sNuXBbUMWfJOuLTl4ZSE6rcdPisRoIXH032VsRWf2
LUbE+o44mJG1MfTGX0tIY+I+K4QKQ71/fFFo+6dZ7vJSV7j5/f92s/K+7SSi0f4uavKqCDGUoubx
/X5UypN8OTfACnyfKi2EFu8FRET3blWsYGvaEdEUX/2ndsYNNVrGyJJ9I+EjYCcUgKur1OqF9rDN
ln5xyI/Ezz/PHFzPLbZIoFG1IppBq4kD/Yfluy72I/0Kt2ayS3hUxTjxJBz9bz0UEAqKYGyLHPFX
Gu4PuP7jgCt0axomm87drbUpMxhY9tu303vqv3fm7SGsbvBiY4330vJngSD031NpYQSNJUo6//W9
ndmGHdOgf82xCAVLb6fmFIIgNDU5GgPvvlJy40s2rMIyLQEGq/cmInP/CnEkEQVD8CHEvlcE7KRK
/9VfAFULwajyPqxbtSZJixoGzno7zt7ujIEXzl3qxiswLdByVD3NmlvSpR7R/n7vyakB2xEhrRIj
ZP8CnbOKqt1SWYHk85J7mqEbheRa/GY0IX9zZ1HHC3EAN9RN0J3CMPnhMa5ZJemG12MMZ5sm1f44
vdylR7+b3neQhCyq7oGTAuepn+BCitvHAxZ/tgzdBg8w0vwdDTHEkgDUKB+I+gIS0WjnhQER/z06
p75RMX6+JJV/8ifAMtyPOIbTTh+sUsvFLWHRsshhJKKi7hUEHT1MxhtC+XcVIRA3/UA+D6VGNopq
gwxnOlV8iQhO4szWI9dj0/0SQfpjSMlFTN/V+Ma7r+GYfpaP2VXNCJmr1te2VmJAlGzaQWYser8n
HaNJWz631igQvRb3i8lfGBRd6NcP9TxGBI0Ys44E8X6p/CZCgHB6Q/n9lIVO/FNa1FXHS/0HqwMr
SDkrMLJJUxbA/MT20ldW8UNFVgD7zQDGlzSSp/57sIAqzqK68AJzRgbAtefKSZR3CGaQQ35+Al5o
Kx450PyacGvGE2pplTIl711F9loW3tMfNopq1c/yG2Y2IxCj/lcOJdWzntcUiLqm4H9qyVAW+z9v
Wsv0A37sQf34z9KvUIb6fYCPpI5CuIzfzO4TNwpim4UDdzUe7Em3L29xqmP/ZR636Ex+wf2TjxyR
mthd1SEg+T2G8sXE+fafIKR5VW9CykjyqvNAjKhfo9LqpaXnQ3XfQpv3Vym18ktI1VnTpI3FUZNa
8Bx5GGvlp5HG1vf9cGGELFLc22AeUzhF6cNHM/GO8F13W/EW9UXpP8ON0qj2kPCrsE/qNdvvvR/c
xOWtiIRA2m37CqHD6q4CxmqAbUhT+6+L3q/U67MDbmT8lcTqK2Cz0I6CEdQR9QH8M0zZkcF1DfxU
cPBAED2Vhspq2RXoUwhSp3127zh0wTqPfxUebMy2ZKns+xC4RxpAs/8SILIIwK1mbSD2TcicnKGZ
B1z2/lR9pMZALtvTDNjNvXQC43HYi81ZWGSS2Jq2K7Ar0a2jv4pmuKMBjCWroaeFyowgi/pbsY1m
UHcFSBtKswX6DhHcyxiqBTejMSpo6hWC54HLpsHNjl+1PdrsO7rkRWZq3k3M/spQEXxXMHoLmnYQ
5Fh+8D9iJk2kyBFy/8qBnwUETYZwP4EPha2oHPLZIlICG63n/VBoo0e5vzZcqbV0h39KOc1aUe6S
CmjsULdyzNAXX2n537G0sk5nJU57LgXkW7htW74clbbm5KlBTPu7m12G9hp9wY071phQVZTHiAfK
/5XR654dRYdaXwAm9O519amyjt4J/uhmIpBHrL77GfC17Lun7GcKfa4KZZNjcDAhJK0KjlewD2kY
nq/CTUOuRbDEJUJRBPHzqhKTcjxMprk3g6gibzdZZDfY4PzMtG2F5buc0VPZiQocBtXsCrVHBpJa
rwrTQaxO5VVMSJmZfriEQXrvGIIU7/HMLyUK/6oUJ4amXYEjA+hO03HXqrF330pBULXC5wnm5Q0i
v98fx9E8V7316UsYUtMlh6kxUn8tNxZVFCXh2jYvlIBgd4U1AiUe2FqBcToqyt5hyfqFbCV0yJcJ
RhBOsa/Rvjl2/QS9HeeDDI7rDUrUrXfz3FpQ4OEnX5l9ZhJpReVqiokiE6rU7e0dc0Zf4S17YDUP
80XSgVtE/KGntyG4NPWkTxmi9rOYxzPhdoiMxKB84euRxcIHaKaLKj7kBwscAeJqa3Z2N+GIKinT
wuwIcsGxeWsRU2852rcp6djUkdqNPcM0POmHJBx6qxz/0VYHIe+FD8CUCbuRk9J2Cw9HptDjL2A/
rTyJx69L+xb8N/dXD207Sl8LlKNBbPTNJBLGsMXKO085WD+cdTGs6ejVR1VNV0W9B5ktjEbg22Ll
zgh4+sya8U4H9bjeWdQzQCkXGofyaJE3KpNF0uvRR8EERjTs7xJgDnxsek9P43cjqRvEyQKmoT76
zci0ooAQxo7phcOP2CZ/31QAgY1iPWJleI1FG5PxEr6kL+vHUXI9pV735aNjotcjiDaRNwZh3sM9
usMeu+tGzyMXdGRIk0itzwlvzCn1FfcYD8Rt0BcesCt5tDAVifg2Vl6trWLo3TjVrHhm/zMgp/Ac
z4COTTFWya9vDT/5PBipfWSetlxRIk/AQS16JW4uhfXOHolMV0I5Qhfj8EWZrYZx4Kuzw4+rZyDK
nV3NAWg+Pc+kS0sVa44M18UM8rVW9DVfTYVFQTEXwrzF6myL7X1mIYYPHryGSfUpz15UbRqKIQC5
b4M6hNegG3GFn2tijceoJ8LQwzdnBUcBAFbFIA61B6mesQXDfw8NwTmy0ExzgTJ60GWQqv1JKAGp
CZKm79/wZJQlX206h+IVHRCLQzcpwBnHI6nwdQSjci93d8uNVTy/MB9Mn18H+1HYh9P86sCgYkeu
eKIW4nCp1IvT3eo69NACohjtM9QGxk+nNhhVLC7Yj/Dt5nmH91O+/JREN6YsAWQSm9zxmCKvzmiu
ugwSPoN/lS3eQLg1+4trfZ/zYDKqM1Uc15cSOTXUUGxPpxiX0bCXQxbZz43G7StbHmGjZB/rWzh6
APkKanHe0EoXxMkL4tZScImaGxgRAK6mu0+vWQaSS37dL9gJsxe4oASFQ19pyXei4JDVpm8aD4So
KkeCGzrzLSnvp84pZ14XF8b61WFETV++I0q7CiQESa+IFURjAETew/kjMChokD05OmYCTSlYg0vB
UBr1SqXsErDLDuvZhlDkGEiRwq5/+OJMOpriB5puTqexdIRldDspOeRNb8kgElLjhHxeRxDI8uPh
wezsZrsAWrK8Br8aux5l7z+Rdz+Z9XF2FchKfH2pL0RBK/TgGcyWYVxzFLdvbyIoqz3S61hkI57z
Asm7KWtqYx9CRPmKk+guQoS7ZJjfjb7DS8KQooOgJvhev2wx37NFI2cNqNnhuXhMPz9v8cTlDPNK
VspGV/G4t7WtsGVlqmqKx5zWurY2rCH3DggDqr5gdPbgk/EEGteI93u+1vOQJxjKy3KYx1ulGxQC
CXAfXU0IaTbrZq80TLao5Ne05BSYAWy5WpqIfknm4CUSXmOD6FH69vdBOR1nQVxqyeL+YmAyiiE1
NT4MaiPQHTYNbZ1YEk63Vk77VK38aW5on71L4i2nXpi98Vd0MpytV0aWJsyfNkukpY3l4Jxo/8ZI
BGe0JxA69ZBHGIbRtoJR7Ysat+DUAJMRXhhOSCT6yZFlrdpdXrYzYOoM9RrsvHR2kEPUhr5j0hkY
f/uIX02Ot09gWVFjMMu+u+6+mnYobEVMtBpCQ+eeZ1LOxsiaelrPGLlMY0iYFfH09NvOP+KwoY9B
swxl4hMfpTvy8Cbk9BwzLlHHpR7FLxIgy2oDtXZNK9r51YROHX2qkBvqrTTKXZMtc0OK2ZqXmlMG
PrpcoFM1dzN2MILDrJmYsBP3UieRVxUMu+6yCHUBM88mwUKyP34tyPbEW3XdpCActq4NN30jr6Hc
ScFcs6jPyvmsy4Gt5IlOvSAQkVMHp2pQWMWxWbcBJoLb2Q5Vb+pzC0Gi0jmmaucbDOVEyZ4LIAXB
QEm7khHSsMZJszBSU5HPCwpcvBshvBRZPp5n6r8xUav28aQ4KT+AuNrZPjYq7YbrXepgVfWZdQCm
vPDLt5q+5bx9r60lDhDqkqCUnImPAgpmyZ1vvMega57y/U1jYQF6xrBOWtlL17mTVcvJZeu7do40
p2Y4rT44wSwVpMpOhF1Ks4w3eDKvsCV1WbkPvIvMxYTSHgjVEF9SU11SllybBGhQ4Pf3kkmABdsL
hbYuw6o80g7Xg7SUKnWJsrGslDm4RxZVAwMWAOG6qDUJW8AVfq9/dE/++6llqCcX89zGNK75vbnc
tUCF0dhY7Id15B7KJgJ5htU5REB5UnGmv5JDqcX3bFlwugfAY7DfeUIaU8r9SuEA8QDVlviIXk8u
EE/owU/z+/zdUW18bVgoDHj5HTYze4qYbo0+k+wzEJmn4HpRNS/Rzcqdu4IbKe44/alG74EjSAGA
ZaehKAXR1l2Y7JZluajGUyJt9FBBvDdOcR/3ar4bXe104SjdydJ5z02VK4Atm5ywQ81gokfsZvJh
g+/sdNGXCKteB6E8co5lKcqLiD/uUeB3GWQoWlkt/xpDRTsv3Xivih0u1hEgw8v83tnjngbncfFb
iW8ufhv6U+MHfZVua8VMUaxRAIlcCRbkf+HTZMX/etxtxX2qWSqZyjbJ6SptP0zZ2Elqj2cOoD4D
AmUPaDdBONaxgb5ytq3ElE4Ge75gAy2Buf+As6f5G7v6JBzU8ou+cY/tKxoKsqJuOCpgkBzOVabs
WBrx1MlwNFPjuGxhGYe5T8j3h+YFzoeYlEHb7IR/8f2cIbm88Zy6MpwZ9CpPNHEnyRRzbrbPUPae
2+laMhrUjNPPUaDzbzhBUBGaD8ypT7rSHTiojrOzdSiNwqeC3hIQBT/ZY2dQVDpq0FMayTf0cfd/
9Wit28LrgeEQ45EmcpyJLVv08qbL1lY+KzEtnDIj+GG+/KD7zflsO6Vkl4r+ij4jrvf1exmki80w
JIY5u2kQW9IePmJff1wNicbtiEmR8b6vRjOg2+gCBPGnc26rPw1JziiworqSDZPlUCwWTarEnEoB
hba/W8CUYQWscrTxms1g29QyqD+y3MurO8v0cIPXOkr/mRgPB/wow5F58fIegj8OyWGcT7klHGuE
G0IYm6uOooqQ8AHq0sABLy5jiIVYdBOqIisZJM6+idRypwf8MoGP6kxxVXuDTIF3xAGi5EgIKLyX
IvTvlslSm1ReMlxG6EeQMSkccYs48klfL//ZYS+LjCEt/Y7LTTIz5WpRDjWHnJIyfkW3H0Db7GA1
UghJbc/Os4A/ks7HmIDIsWO/hvJ2qXcHcQrPj0OsSStL1xb32GCITUw0+uLhRCLmSX8WjpKBpmso
4I0tqW8TP8QfrmToq1EimsnP1KLklLhGi6d133CNIHK/d3og7JRGHqbVPswviwYUqKitCcPFvPy3
/Vv8zJO/T1zpvLrLA4/wUl/3IBHF2aE9+lUx/VrwkxbOYq+spMKBY5Ehq/HGtFrVXk7vxemvlgwb
gk2x0kiHiIHmedKGtkVg142xLh9g407bZP1WfZz4dS4EthXpVQxpXsgo6hHWXZO606PoGt9jtLdz
3wD7wryCTkIWoHLmv3nz+MpF58qys7I6GdpgGoVZqSUEM0jFeTDZoNBiBvntHyH76g9h6TghtgQe
XvE1zx2RQdT2pqRuxHlCvc9EzmSBaF6NrxcNwaB8t3VIq4WcQtfS7mtv7tIJ8OXl/JzOE+9rQ4up
0imrt8okmGaGn1y8CXrjeEEzKSwxCzUyrOEN4M0DJfLLySkZCAK2gHJSA0xKfXQy9We+UvT1cNUj
uNrbHIBQeWw9pm4Jryp6/NfSopeKZ5L/VQBBp1X/plQv3bvWUNfaWZJpmA0YtWZyulDQxKahTvhu
eFU2KBxY4ckWOkF1JnLKSkhgkF0om7hLnqCyuOonT8QkpjpZhclcyEAC9sJzR2L0yMvsqtmXlh0W
g9wC2uCH5HWIZgKQxx6IKzWMIgGfy4ZFSgjtfJpoGC+qnxgrhVH36Q0drly/gaeIZp5NbfVH/Bqw
wvSVfLsZgGG38hE+N4u+oKXbw7I4M6vD20BYZ8INcuTjJzBwMEHktVzXoTcgA4OX344jpiK36aY1
iMarvk9ikDiKGXVKNW2HQp/6I3OangVUxa8HnioWgDQJlKj4Y6whEd5xrzor1MU1uspLqsCgXnDN
uNPHP21ez6ky1lNc6WKoqgEDs0EZ68xmQq7AbkUJ1gUnDFIC6EZecX11HVevQw65H53ceVwur7Pz
/bygU08omZVy44Zm5IBeBLcdP9I7Y/lRTMwKt7IWWY+iBOE6HZV4RdBA7LEz5iMRqJhEO2OSpGpn
js+OkalQ34m6Q6NGcFLC29chKBrQ7cBiZin4kriRVMRnC4lEO0i0PXjaNEKSQ4ea/BlpEt0gbg3K
nKIcmJ2zDzZVcopI9Y9XVFCHs9qL9PPcfWjAW+iabX8UNwledcNanRPFtVBWOCeMUQsXFXjQvqwn
G8nI8uKsjZqsM0MCvgP4xByR5DnD2jPOMlu2rPsbAy1OBpRvMUlg4aFiTRsyXSsd2gzTPI5E1SoW
kE+RfmndnZdaJ0y4EZkPeJDgqo2diej+xXABCAstzezWvj+ro99A6m/XKz1eUBFv3K8uhvGn7m50
BDLt5LnrfYIlAMuEecaxOXLijA/dlpafQXZpBtiFezrees/m1EJZPdErGwSadQhWmZ4PO1FlBoGm
UbTirsdH1vhimSh2XoqO+HREcaJFLJTspk4be8cPKkdUpIbzgRX5L1g39Pt9OBvhFawvjTSStfrp
zmpX3CRyXtblVnY1C0Wsuf832/Od6me84IwdNp3gjatp3y1ZubefGj8gxakz5d6OU4P30UmJO1TW
G0Vubyn/8xv6kFYQJh6mR7uKS6dT2xvUCo1oYxCPi2ksayVlZHuHxZc5I5K5OvZWIOmc1m/O8YU9
P7O1ci8mm6sVkETkUq4J8RvFvO1ecPRWEvQQbYBbYe9WRtN8OE4GTHIPgzbkK4M7Fosd+DM+ewqA
dvRJPkrerfkCQHFj4vSv6OoV9sVrClddvzrkmtc+YuezYbYO5hMVwwzP2Q7Ih1xz7HLSHyCHztsU
e84ak55PyIC+Cw2eAiHKW/+qWoItfwZ1TdEpZMhREPMVSGSZ6x1qt61T47/El2TGrw3yoI8EhqHI
QJb0x3FnNyHwr3PxSpg/FsbZIzg4whR9IxBhB5OaT65cdJ4L9Wsapu+t7klNgf1/x/JL03g22puH
/+fglNvktCMs/ZlXaojzqnuxXqCJW2r58IRmbNUM0IUlGm7H+9fMYkj/kie08LyQ8lpH/qlYiu1J
uOWFcZuYpQF07wvzSU/c4XYriiSsgzjo9PNYKrQiF5e/fRzyRgo4Wq0XMyeksS7nEf7nnaUig11h
sZ1s/RKCwZMOzc7wC16tNj5txGAQEhgR1Jk0KL2zIikoyRhMxmh6hvMmntwYXDLYKzomikzMhsto
9F1gwiJe9Vf46BUSj6KvDgf2mxmRQ76eaPovoT4HJLrEWtLe5/d7e8lETbtk/g7ec5Caz/JFVWr9
laDBg/Ju0aExo0DlfnWAxJ4Mk/UEL4CwZe6XOPW1trFbkQt3Gc+vxuS4iSwZCMS6F6KCe4xdFwcu
HzYYItDaJsNkfqSUPVMyg5/ZdX3yqlA96xfDhva3a66p4mn11iqFCdVoORvHOGhMuRMDJ8p4lsy4
V86a9L0zKKEeFWjxYwtGyW+b5/lCPsZ3TZYq+Pm3Zpfxw2qI8GQZYxxhq/HlfNyMIWCKXS1UiEa6
sHfCpTmvgwrgPkNECiCfjago69HRGzHx9pmCUC0+A+VJ/nrhiTAtvzbe2M2Aw1pholVQb5QMTo15
gMUV4MXFURtdTLiUOVtMzt14W0P7aWTO3ow5tx9k9H2PVSi/OcxwGQ0oxMUK2tuxOu+nCIYOrRcm
58Qeg3DyTr8/QZP4ibaYkr0uhiHeySeCKdZV6bw4h/at59LtXCGcicKNIFqvxdNUI9t0S28u9lMg
/W1qSWSnVzykbAsKP0hqdEIHNTFsunmJUN/bS+bOAK58OQWdXTc8R+FxEl2TBLpabPK7UFmsPaj1
PMVIjO5pF5fQVbMaq7hq7UAYGcqN6NYCJq1tzMQWrgD3cDlUDcX0LUPlylRwiBaoDyVDUXMKrZ9a
cdjPkQMAxJzYvQGkniBYOAgRLN1++BVZcRYYjx8gn/EXf9NhBXtMmSYOoNgAxqmN9Bfa35oXtpz+
uZrQKB3Hs8qo9Nga5whuZw1i3ZbqeaIZ6LodGDZvW8TfN41Be8I1KvHbDsNIT3YD+xGpRtTb+Rjq
xSZ5gnlgLQK8/Vt/5+T1WAdTOpJcFR7Hii2+1EjmLKNEHgZDiCANx81Y9lnHUtpGufP1BXe5nHAc
1TuDzy/BVt2+vxyD9U2dGiUnph2krFrPbiBunT0XnQgU+et0sqV7+fH0R3iaZekUz4G+clFdJgd3
aQQofY2q3pERO1ur9nAqZ+4vcs4vk6nXZtAsZGDYF65N1B0ngXe2rwCN4U5DhSAHxhR+VJEE6h6s
cWSOFeB2r5ipz+Jelw8B8u2M3mKeTLZ1ADCoFmYO0LX0pQkDSmdYvmp73uP6XF5tfVqopiMeYrRP
As/JWpANfMOxeaZZnk90OON42vKdqj3lznHZpDjz8+YemJOw29Hf6TI4C6YLZWiaK2L04j+vMd1y
rAB0QfuaEQ88fJGTcg2nShZxKDpXohIOPmCeqIy6GHf2htK4N3x2WDXEdKF5uVWwUq76GOmKsc6G
JNjy9o2nGhFY4mOy774hwItxRyVzPscgKRcAOfvshtAPDRAJzEvrCNHjY5zYikDCTgvujNxLl4Tj
n46Qy1IwNz183d+HYrAva6Gt6bWQ93BckIW6IIE/aLiN76lQm6FjWW0WZ96pkDucurIZ7WnILP/b
F4j9Bo943qdVmxb+JsYkp/Wai/ndhvNuUIXQHQiLPHbv1gYf2f7Erqcp/WId+/T7EzkDUBM1xYDh
ijU9/8su6dWV6Pa0S1rVE3YuHZrFDTvkcYzlzKAG0apsVuS32S42Gwt5ZARXjpWtl7IkY2SJZoBR
8ZxoOOZ2G23xbsSTro/ZR6fqsOC2t+a1HVrLPTVl6rWq3L3XhKuvj4+rilTdbN4KQPNdxTRvzW6K
AgdLmEPXaQWbYnDicHb9S+LfUj7ewxB+NKerGS5RarspbbJh6Ube88Sr3mBGgUYHGDB4Ovi3t3W5
PaIyBrwJbt2GZzmfM6++Swy5WKp7YXIGKxhHpqN2noDq6ys2VgfObUfZu8rjPm9ngmYbuWJEj7GC
KGB9efRXM7OpT3sEBJDZDxF6NJ8ageQyB/rOPrCp+N1WKTN0WVjJki8XSEOZl4xjeJ9vuBN2P76T
c2GIvK9KKrxFVe/0Pf27hMcIeoCCfchU/w7bMN9VV7UPjl4QTMHYIjebqUil3aVVOG7u4ofR6Rzz
hbm2or3m3/3QLxWGxirkEazUS+5Xnn1xqZaH+rYVjuJtQm783HkD4lxIEJlYhnze4V4Ry0ioyp4f
zCxnGTVyqogILVURrZcIgbHC4zHy+JjhCdgGOyba+UKn/bAeQmLExGPLUkFQa0vPynzdkshQBU+W
jxwMcWQGvEqVA5lFcrHJ9ixjpA2/lJhAXU7fRk8ksF5JePmftZbAIF8CwK8APAZZokY4vCsnCQiY
CV9Qua2XWaA1hhP76YM+C+sOTAiVpO7rltGZLTZW6FTTcGRvVzqcXswAagHEzVxxS7xbdR3q4tL4
I1E/9jjvlGSbol1Ush8xEHoP0nAzUrswv+QpnibP9+5Z5BQSzGLIGpsiPbGyLZTvn4rz7k6lxUEQ
hWXp8yKmjV/ud3dpy0St4ROjzKNZtJVTVdD5bYfeVpP9ORjCPCcvsqc0165JvN5G67P8tf1osypE
aAJhmQNLnbmFk60yQMIkjNcbOlppemRJIhhyr582wh/A7F0QykzwN6/T/lmLuR2b5Pe8kWUb4XO8
/DlYIYSk84uuh3LcnkjPpjObHohJyHGUirPDU2BmfVdqza/4xbqvN0LNYM9sRrGfTro8Gt0mXrCN
7dbi3KLvV1Hl2YTGn8n49jfRHq7EAeDXhWfW/oxsRUE3M7dFg+ONwKmvZhwpYJcodZBio69eCl5u
y5KR0ZgW1goKdx0A2akZw03jHctdY/jR6v6sjxnL1jzP7WcqyRAZKDYNc0eAtBRJxNJoizMN/cyW
JhNBRojdpFXlcZtmK6OqpAMpPpR0ZkV3W5naLsnOeRLe7j6/SGL1F5MFu02eWg6vI5Vi6iwQqsRo
6oOEo3uBADY5WFTnmve2s/nUIFuJ8XaverUQlZWAaOClRtr6mECOTtgeW6y7SWcipESmeiqASJmi
KK/DE4crp71zRsBvEADUTzJAgJk0hUDee2DR5V7CgOi7VIjdKRZZTORZgUnvFOPBK6ujF7+kdZ3k
FlpzUiIuRpZ/6yi7AGopJgRGmWIGl3HG6QejSRA/wpopFR2WzUTQxYc1QKzPPL0Me0yPz6Tcm8k6
/34gKURFy5Fdr/jO1CchEOnnur6PYrK9Rx45ilZDQPrjOsXIdwK8XT0XE+1OQg1Xg2YQufRHsZ/G
w8lhQDVqNPQEA0tT0L8KL7m0ycIZfEv++HT9pPpe/jIqlERS86gvMWhqToZWbzaOpu8VKz1YCv4Y
bYACxsDhjtmxQkupsOG61Jns3HSnLK0Aqc71MODjEWz0fHWF20aO7mPzrPdG7ZOB9ZkphQWsjHfN
ByA8/1EDFere6uXBLfaQSXScTjO+Caw0+Fnh0GiO3JkN+zevx/U4zL1kSGIJeeRYP4J8qovNk2BO
ALkRH5z+eErqbghPRqYJvjU131FbyUghUZqqsglxTUWnSfpr/Sc0BZ9RQ2Q91rdIOHrkLjjfIayi
oo39LBLqMDPLCHsavS1zASUKbuazWWHQkFRs5u2fbT2gEEKJT6IUm7dnLwiJLjf9cp1rIWDSeTaK
40iTBihYPdLAQPSFPTe+xhbxc+Hz0fNZaytKSOd5zz7H5104EFRaM0CcdWEeC6NH+GwY3AENwlON
CZZ2MjlNMxit91PUZkHziy0GYC48wkiqbIJfNyc+vI3tOz6AkObJgf3ZxoKYI6yuVMzTgottcmjh
jeRYfb9Wa16wFMgDHuSpTGqaqq3JOyptkWooBM4v6ppk53YmUsfCChYBDe+VAh/O4UZv/pAhdJjH
TRuGT6xgEiiv7Wultr7vaN3VZplkKH14I4v01aQQyZdLb2VjWCwu37W+WO1RZNHrwNc2e69vKVmL
6u90E6HsgKL/jZ/dQ0E1Ku74uvjS8vWuV04ZJ7DSspBC2x7GFLqRD1VWzoOICKz9Xc56o1Xkg2RU
K0a3aDFsgsvXvLiMZB6VEzXe5Lt4hWgGq6W4uAShRTJz1YLZBvZALV0sqclobUW1JeIF7zX4+Nsl
W+8VoilmW2tpvVczsB2StjDgJgJVOBFV814a40u2Pi6iDV2dWBHB6/AVePT8j2GXQZ1vP4LEk9ql
WfbrIWUgChblnO+RAoRQICt1peDdMr5cJYvcEMMpwjg3Z51OKxr8/BmaLCNYai2BKXIqKBuPC4+h
oyBIheO2/VcckWPm3D8OXhyODmEgQSTqfFTTwNmC5qslePwgk7jNEaqYunXMqdeWl72s1zuujiYh
QyEuqH9dTbgbDcU95q26fkdbZ8iL+zF/VqoMkh0it6WHgG6oxV3LZgMxWhnMOu/MVLBMux6c0Xv9
Zc3/QloM+H1vo2xWcpdYYCif8C+E4hcAXPpReOtiWD3AQ+Kx84D3yAKLa0OfGdSPkOOu2RmZx1S+
COyaeb+SQfg1+FCs/dwcEZidNPK4kshArcPRC/5NOUNvpYnRCxS2xS+G9tkgSarZeSjzFDXzG3/i
amihNwwdmkP7yDv0MBG+FaIYMzLKDaYfptEejpnnGqyR2tXDdLV96+k8Hqri0f7bAFvRHcAP15p4
l0T3fmfb21bffLMvvjoF6PuIBI+0weK3ksrpsKwBBUDamQqrseKl3xguSbSFXffNlvTP/sGJctQZ
xfjvHbWmkHQq2qc9MOdp2NWJWc8diEMLD3Qbx8ZE1yV7LFfoyiQLDZDn/++hg7cYPxCltn/tlP2c
7O4RLmoL3Ny1TIMOQgfbPHOn2r9SFBwpc+Si1LLD6mdx15ColKB3cIJRu8vMcBOvheOz7912W826
qh77DfSo6HdAkOaVjBB4xV6N/hHybiMeiApY/cdSSxuagdhRzlFS857WFvwW7eRVePTYjWN8Dm4s
2rfFjGJOzu9UvHY2DniCDilEZaNK3EEn2rsG++jztD7s3LdGsz+MHKhrCxS3pVH+ayKbPxcbNsw2
FblAvZvmZg9rDhB60mqLbEFnnjYfuocO552ZM4JJO8cPSSuJgS+lUcNKG8Q2mOoBNnCDDSHR5257
JH2wUe/Eta8Gm77In7weE6/qvVaZ33+mDGFU+EjVCubfo0RKOtX0TlgZ59jN7c7XXj4HUR8g2t0R
U6QRZ+5LjjBUAUgtOgBrBGk1R1hdAk2pFTJM03g4rCI/IjA8zu84lVnOe8agR2Ey9dJJXAzCFJCZ
bleiS/CKBgPx5K3Vdeb1I4LWUrF7sXKiCJQ9kKj6KvWDpTxM9E2Xh4ZGHgx0r2JuYt2cqVHzwDuj
ySYrsaMYd/H6+36ujvinOblvvdISMU5Kp4B4ZoEV4wnKKvCs4DT3Bn98N0zWb6xsfyRGEPcTBg8P
JoPTxxkOIMW107ExmBz8VyzW4t/ZTeCCG1REvDNNHsqqyoYpmITUlWjsKbYjx/nSeuoUtKn78xTx
Lq/oezUaOa1vvAuWE/2AggnfmcgqEiYZlagVjKyCLcCO85DYukj2VRSEY8RCVodAI7+W5k9ThGSH
OqDjPf/KH0wRZvlw6P45orwKvVw80R4q3BzIvg0d4EDogmnVeI3ZXB7wcQOr4Z5hY6d0Y7ZOHl3m
peACJTZOwWK6+sPXlwnih1WXw5Oy+F7KdtGLibXmq/6I16EbQyk9nLop76clyJ/0SC8zJs3VlBvZ
sMWkw7Sf0jCUH0D0WY2Lme/MFEtyXEMwzRuetS5nZOvXkp7infD0P60jv9blMW1n51o0m/dgckep
xKy1UjSlZHMCIM44WdxWWTGdQvNvJN5E9BJhOmhAhKf3NmwILQjlY/+UyA4eZq5VfN+KmV+GDWgG
xgmG0M6PYHm7lDK/wkkvwuFWiMZD0hFN3g8SIWhDbaH4cESwDduoqa010guWxnCbPqh1rVQaSg9i
GzNk/Zh+FB4xjJOJOEtAV3yaWMP7T03dBSsV2UUEv7HwSpGkDEq8UAPGpiCMHvDMlPgNR+sIR4N2
0oGNsBG+swL/QnuPWcvoMRmzeb5grdHbusTAH5nIReOiyhpk5DOKhdUUOV4oIZSng4w2rlSP9ttR
+F02nfvgjOkdylWCac7QLvV/e8j3x3pjiiGqDQMB55vQQjT7RBhBHbCvlFbeajT34m8qqWiWg51R
TLvkbRL49yZcwR1OWnJ3TnNKzfWjDbFtX2UeAGIoQ+AL/FM3rjZJPBpPBn1vdH1vxKT3Fy7oqC5z
PD+elZgD1Ma2MKGo4nFFQoEPiNKFm6/Bhu7DbKiMl0zeIZV0whJqbMnl9P1h/5RCR/rBKRgZ9zZn
2bn55MI0aRL0JWv8nBqYNscvEg0F1rnv8GzY68dpQsWzrWfryJmbuQHYizg8E1ZqE1HyFBiFjR6k
+M1J1Ov2eK4xXz30RvRhaRhyQRn/94t93Bh1rsMkDy8/7T0fW+0MxzjDZKeDGwhQE7QCw8w2aKOl
3MMkNZUBMLD2Yv/ddwCQzz490E+NeMQbjA70Nmp0u9z7qf3mLG6OhISLiS/cRmLY/Z2bwIrwQIGr
axA0CP+mCLr3CP7on0mzhDXsllnxno3PsJF/JS9tNosC4p5cgORJFcy5Om22zu9Rch1yV8TiFgfn
MOH4oXN4wM+MCQk2/HrUkeqm6x2ANYlFv0za76OfJ8sCtm7iDrp+k239qvk8jQqsJ5uz+szUdRqg
3q5o3zoY+n9es/e7Ppfdrr6wIcB+ncVkxwFGfu/26HGjtfUcUhdU+tQ3MAw9POxKAFOuPEB0OS/e
rZfDf0ttYic7lnCx87W1xIDI9oO4P43GRf3RJGRc+QL9GXi3zZ5uLJgvkkvpfC3pl7wxXNe85SvM
np7TriW3DbsJTkctzdcA1X4j69oSjXk5ADyGgtM3GU2+E5AG1He5xKP6VadeWNPsvhAadHveK5Ra
oXUxPvS5EuKiwbOIz+9zYCcsFc/owdvNstEGYm/n7GxduXCK063NJg0FT5cG06CvOvzvEZ57cG1/
WRZwVjXPh17ZhZZIgfZBJeJ70x4iB9Wip6jO30fvnkGVtS57GpgzGBL4QdUrhg9+Sr3Hrmuf8ZUB
1FqjZqzM8s7tYTtZEB63cAIb3Tk0oABMkItfuIj2HB7PKfoWdEHZ0oLS8LAzMqLCFD36X6Z5FF9v
rxFPAk+Z1sDhGUtLQH3+fkq5H0U+QoKfwVRItXh+46KKf85+umFb773tp0k+2mdILNk2kefLTh0b
QZIyq2SyxBALuYgUy8Z/nn6hCkdY/5ym7Fwq7fm82WM84R4J/FX3gQ9H3N5gyP0jfFQt4qLVEA8X
ih2z7JYw0SApQp1PJQTv4/RapGltbEe9sL4OsgtWQ2bn4HWDHCJ33wUOatoKtJ6RUYcsEV8RIl8t
56veHDROTl+5ZvDhArUiL9WwUc7aO5jYKj/SKajkctRYBntFGgxItmKjXOJsHEbxEMWvJSCHEwPX
4HJ9okqoZD57XDNeoTUJaIhljgd8u4LfmnMqW6iwQ3g98/hNrABAFMj8S3or8SIhs4yL9cLKBXM0
QevaEsc1JzWfp9nJKyeSU9v2GmxH5CJRuGcXvfQnPncOTEaW4PWumnH9VqNtPU9Cf63ezeMtI8Td
IhzFbjGoFXBXIjfFHerVHJ6V5qwNE9xqlz+zwxWLBrV5Cx33TuSmU2KAlgQSXIPP+xLnUdzMMsms
UxSDdZxK+npyUf64F/HAGhk415Ex9ISXY+qPni93tGV63rO9de7oHmjgafMMgaKJ2DsQM8AOGrza
/M4trjNC9Kh6EtlX4dxa5rhmZCuzjP4Nkp9y/MFAde1jM0kxxuPPGL5j7WbgFG/yY5lzCUIxwJ4h
5cQRTRkW8M7vIxPZqlFGDLbUEKQLtvNfaqwM7h8af55BhMgZy70/5nN3nLPJJI2b5wHgmI5kd5aQ
RAevrjYGIUwstQAHaieElJlfkx0qgE7S1VFTvPa/Z+jJRWDHSYNPxxZqjJRXJolMhytof4fC1zbm
acYQ5ONRB3mMl1i07syrZrnnCx1JzH2FXK5CT5ZNi+e3jauQssBQeTfUqqy3JacEajdAhTUBGWl6
+YRYSCcbh/94NBTg24q8nzazHhWXy6+FD+KLkGRiT6qES27IjNTc16AB9ZqK9o0XEDjmWZ8QOlfS
EmpYJM0+7Pf2KoLFn8PfGlXSa4qcN4Ilfj5mubIZnBy/FaFOQOk/hRH49bB3gAA4og3rNvTFjhQE
2paOHu5F2HiOCx+YN8bo2jauBAbE5D45FqQKz+vvN/8dcW9hra7Z2B8dIlXh4ffYcsKgblQNO462
6JWs5up0tQIy4K8ljhg3acGBWuWyhcObU2mTw/LFDVw+xJ202oJpdsRvznyY8UldYjB0oCVnrBK6
XJ9uQZR4s3dvVCSb1WZ6rL/beq3y9fDKpBb6nxFO56rQbqsa0zH0//2xHrffhNJVXnbthvi6REJm
HdIjLEZM4KLlWwBxId+vdzE5jr699IpQ941Xe3YpmYhLfMr0f+0p2emd5JL/T0PEiJDpm46o0I7v
Xn/KvTJ2J80tJcc8GdvrENIwhnd5PLYVNC7FoVqout8X0t8RgOIdbRtzNAIKiJ+p9oKocfymdDUa
xq+4oGnyvVbwLcTzclG18qOZs7Wnlrc74rVOAg68gVGus2uuwqYKVm6GKCZ1zbQx2FplPvKGy0zA
ts4lUPB4770l0LWhMJdaKvBM2UCk5R+j+wisVF9aNoa+ivYm3OlVYid+M95D5eQyBN9K/f3SMAgD
jCzDtxZn21OXObZ4/OA8p+ZnQ3cw5JkuI97XR500xPSzYl/myc/yEj7ZD0x+XS5veGUacmn0S+Gp
BgiU+/+clWBnUSBPFxPcUmFcduWd58lDeFWOPqbkFSZIBFplkh9ho7FO2wLrInwEXnE8aruXZMaJ
8SMvMQZtjpVvhSWpSRZ1oMN81xogHfV+WD6SDuUJKY8/lhYmgWq2WIn37cbHEtaynXrgqbnIn7Dn
nvbVDIhmiv1FzOgsXykiYBwkTYnkSpYf5l0j2tA1V9IMK1fGE+isDgYInWH+dcDUwzE0QQZ8S38j
IVYRR/efTc7Q2KH3bWFCld9nKr1NNgMlrtVm/a2e/HRzSBIR1MJmNWtzNQ2gQpoQz1Rj25N4xWDV
Nxu5qPhCSriqYxPJmZX2sO7TiiC9y/EivQEha2xD4RkcWsrR/fMMKIwGUd51lIpRSnVql0dLW8WM
BPjKUyrev6RjZ5hSkrovK8SO/MJCLhgI6zO1lb0gVPaj4iqMrEytlOcUBz5jE/vanz2X9ACZ+yO+
BqfJ6vXLLH1Nl+uaIZIbAn2D7lADZTN+lGR1FFDTnTkWKRDo8nJyduuBVLVoFJbSwi6StgFOOnAn
aEEXrpDKrMi7MWalvsmoDH++zSS8VtLKUEX2bJicowJDLbyTGAc72Tiz9UYuYWZSv67lArAhfcqA
85vPFfkTR9LzoWKY7VsgOD7SkHZPcAwpQNspj9wOTpGrRfCOo3abGHUrWAE7bsrodXSGoaI5JtCM
jNFy4vu83qk6bhDSE43PjuTWdny/PeTrcAWHV92kTZ2fEd+2fwN/Q8ML36UmC2x47sMi/tiiwBHG
3ylgvcRUQdJ0eTUzG7ZGDE2CxQWq0CPOOhivkeEKxBMrO8W5utBeQ4ljbmDur29GRihotT4S/tOP
4J5ZTKJoUT36eeU9dLcxVldaMeQgW0b10mm0RQ7MnnFQaX1iO0dpn9PoHAJw3totD6mdGkRvUz1q
YyQZe8rt0I5MnnS96zAiBkNmAj264Iangh+z6rLfGNacW+igsxFOEcHdjFcpKwHoLhwDOQXoR2jL
H/knYO1uaT5KOQoR413DNdiE2ipPSZ6f0W5SuV8i2q7cjZYOkjIGLgaayD3LbiB8b2rPv3rrIJYt
YKjUEaaqNNK/dQAiC60VXh3f9GZiLldfFxem2f9ArGQX8UCN7jFJFtgyilg/xX+gBsF05kt0nzre
IysJGGSD0uGV4VoHxJY51VozJvaJrV6OQmjE/afJ6wqAv2cMnK1C2em3/v3UM2FrImmU5IiCDZP+
7vzyJo/XpauHPAeCXD2g4rZPPzQTsrLYCAca3hPFJMeXIL3WqTPzChOmGNwcGql0BVP48YPcXgsh
as3Jr1JmuhsbbszNSy8KUPBnnN6BwI6a0Fz8qAs0SOZolXzUaJC4/fW67rOaY4LT0LSZuw4LddnK
ZpqWnxlr0raicGiAn2/kRmjYyR4wgRvYKc5hD8nkElTqj1Q083yeSzy5T26tG4gsRweWVSWaHBfN
q4fUHgRGqeLVRq7pYk5bV7of3N9+qlYrqfxnaTkbeZK/kiCHcwC5lt+uh+wgbx1d06spSC9kyT1g
TnZyHNJyZQaXbDnkTxuQMqlzY03zEGJQkbMta6Bom8eryqrHanDgRLez+93s5rTJ182X2yz4sOsZ
j5ISK4+0/VhGAUL06aq47xQV6y9x0auSSb6aGR8pJqRssiZmxW6GmsL9vFR+5iabs4g7hOhFhyLo
n5SnigLEJSr/ysrXljsiLMMDf7sheu71LzUBxd7YZT2g6mkwC80CcTs0roeDHPnHr4qr2FsueJz7
lPNFPoN54ADeHzqL29yBrOr51hlxmFnPfbP9qJKJ/bNs3+t7P7J94j9Vi1qbSPBwr9XOzuEQuBXg
1a6eLca5Lin8oi/2fUCE90TkL7lTYu4anTu+filF4HDaGG7qqOi0B9/yFdU2xARPbXB3Epdm6m6p
GyR5z5FxwaBEFbAK/msH+P4ezM0d2yaeme0L+/pLOQzTBNQKhnEXpIAhiplcco+Zng3AhuKmkjbo
lM8ug1bbVBXqy7ymmCa4/DlLZflk0lewDFBUyza4OrLwT4kr5oaqy3zkJDrs8fX9FOrqr1+SDYYx
hsWq7vkx6QuQ3rggwD27IzNZT+DaZ/FBnSda8pAd0a7FHTBTml4WlQa+cfJPgudIZY6GfeVWSytt
nWxSiSsdwWtaNw4p06O2//tCEqZUlHReGJ3413hdnUO9neuRwKh1GB3ewJjH5dTMjbCMalU3+bYY
AzOvkpt/EtmXW3P6MRHYgV27j4Nj/ooC9Gal6V4mj4dcfwoKYfCVenThe9vhrJJ6khbKH8wH/YxM
dwBlGR85LEBjy2V1Zji1xnMV2Gw+PQ384iM5wNPA0KuRYXyuhi2iVB0xDly95ItwZLnrsvElrzN/
Jxi+TjEOhqOJRBM/gCO66QbUT/YoMJZPADYiYMTcb19KU0ozgG0E75EfxwQnWv5DdIp4DbX1OowJ
8DHtTcMyEmyJVz6jIdNKZvR4uxWnx2xSIwRemITyfQQ5P6XwM7ioYH9Y2Ac+8zS//RlZFkztvp4T
dJ1NkCm4KuBBTM1BUSnvICpD/eE53cU3Cv896Jt/mJIJqz2K3s1T83CVS9EsKiVU9Km2eLPyTFCG
sorlPZYRpKrlzx5M0hGXgT0Xj2a6x4LYYaNyWSSOmH7LTwlHuO01/+C+himZIQJ+6pYCV2xC4m05
1iV6L38iZ5QkBsvbQp42Zn+xdQX1mFIgGwQQXramkakLs5/d/bjOW3sq/lZxhYHhMgyA99xcGEaG
ikZm06FhHpnzO7FPeQzsBEp1k3IuPxyNb47qGvFQt3PABJd6HuDWgrrKFe14VtGfZi4xaUGbXEBJ
nQS6ZN9dyT273tCLs4PKHxhp7yZrgr2APJ3soeDBDMYZxTSvP0SpXh0QTmcWDGx3tme3aJo7Iwps
lcqmatBC2TrpLetMdYl+5NauPqWw/xvdzc3m8ii+uS5svFnHU13/zgCKbEEJuHt1aMEt3WTcaw1C
De/YONg6YS4Hf7BmWK2Ndm3pwU3xpHpyD/Ex+KIqUxir/xOudNYOpeZOi7CnknRdDuhS8EOZlJ3M
YUgoTtIrYtBXVfsLBzI3R1x+qdsh+WMcDAPURvb8cKrIIDkZuUvMCHrasK09ud46911PKJGUVtZ6
q+/PLf9B9ASRe/IFnjf4IZRj4gV6Q8xXuixya+enlUHLlohuJCjh7HqeiSyUHQJKA4BSPFtIyY2D
8+eFrk61/NQCSODOPqMja4IN4s6d/vIxMm3Em3WwMNOh0bdK945uJyhmq9KX0j33TTdXpwtwCBiN
VKcfkSDZvbrKmnzcVS9nv1NVZ69LBNe2SZeIUlk4GkMqMFMqQwc58RvHs5/Yq7jdB+YDKxeejt/G
tuI18zaKox2xxb92zeluQRhTGkFHFgkSjPW7cbhU/H6jv8n41da8Gwrhi+O5Kr9X6TFuEiBd8paG
rz37kQFEc5SPINssq94jooenO6mhvf+36GI8oNTZuGfSjPqTkE/NiHj17yL4QaPF8YBofIzyS53u
cCJLr97eHlk2Pq9VEy/YybJqhCYGZd0virztj0mWANkbUEbFvasrUuq9d3oZyaVC5A8eROOt0QPu
ID6SSFOPUmcos/3HvbJHCrxlBbxY46TCAv6tB3i6VfoLeh2iR1RQzbagrf1dn7DObsCu5BrVm78O
TZbP5jfKno5vNRphi1zx1ISIx+SehkIWoP+POys4bXhdsyZryUup8QXV258SmWP+6qrcCMiMyVqP
SX8UhWa3Ezbb5sTgadUO3Pb93OgnXIKCQTh5Y/wH+8YiVZjpnUIhevLky+vNxwvLCQLeitrOXq4j
0eGeoWmLtRem5/r0u/lmbvX7QMREjx7tAKJP8gWDHVEDBwvszBpDTf4HrTAqZcuSqXpuKEFqxX2G
u1LPK8VkV264sTpKqY3czpn2s/3VKFMe13l/zaGwIDdknPt/CvjOAJYCIkhzUVkD/sPc9UALgUU8
gJIcrH7lp3ZRAGfRmkc/d7AqbrS+BYWrS3P3Gg5OQeRJwk01mUXECkeuzK5eFpli7IjFoWMfduTB
kOvm4I7K5c6fF4KlL7J21RskJMsb2EMYe5oxbsq9GwW/6clMNIR7sx25SOfJt51j3ZZjg0LUsfji
wLIB8FEahBmzLDv2DADFFu3ut0U19S5OWiL1l0XcIXMkiAmky43DRXkRX0x1BGqvA/Q96uLTk3bD
wncLXdfCbNFaKnNrEmp/K0QNKoWEe2sLYhl80nebD3EsHaZOUy8gowu7vlSinOLeiY9DwZhPHiha
siJqKsjy0CeuaTCh2TXCpuIoZcp0K5G8yoklQ19VYiAaiPMPaG3wHyxT23XdMfGRU06GZVmN9UwH
oW1NDkPsKQtE9XHjsP12xvDNiTIfkZCXGem0bpUFWgnzOhLclrKt/qoRMPl/99vj/wXL9upWuOBd
1Oai0Gg/Ik3avTHUwDgvDujUJ7PKFhRcW3hBW9KQdXZzto4CD2i9yclcbipMwRa2LVyO50VP+mkB
Qv6HWu9OnRUnUZFq/zOdKMUS/GcQgaApqWU2ymU4BOEuyuAvZF0SsUNFtu2lV4v/Z5+lITfrJh9v
02LqU3vgu7731UV4tuHYWS5S/3BTudhu6puWgnO+Hvej+B2Sa8S/i+I5glxgqaVp5lUkwe53n8MQ
G7OgPhCu3GxzYIynpa7D7BUPei/m6ZEdmZ3Ogmk0Xe02FHG5S2YlDHbqoObvXuxIRKa05jwas0lJ
sL/sRUia2zCe1EsbqmS6t2ufjCR1wSTX86aa1ZvaxisyzvjyL86hG9iR30ITW122202JxsilgbvH
doh1IjWVbH+zpufUmBebpHmWmXcEyTFdadVaS6HYFLHprePiclojMWoE6OErxwpak7nF9simYv57
TPYFqu8QSRgdvh9eMVhJbGkWD+HMMpNehPHzZMyer+KGJsdS34hCsjpCZCnpDzG4uVtIaYvn/ih5
rwy6qvo/3/eT2UcJUeGcMKxQU+/bJahCUdYstfF5Skjo5aD0Pi1HreWX1pxF3PwFfrPh+OmYXYSX
b1YrK9wh1ter8AUFT3UKWYnfLfOC0XFPpljXFcUT0exrLyIx1qTMi+RSOAVVY3iLnAb0/Awpxraz
hSgBkcKeFfgOab1zXNVKwxgl6AZNdSHDcgqsJqIYhqiQQR/0zXLYj3qLbuA88R6nhy8OZjhLK1fG
d+GfZUs6ZkDdauvmbiidDAaCCf9q7ue04R0zPNLJXVe817SvN3pJdXq9AoZ60dMvPYnfqquPEmr1
7urSgbLm3S39s7dQkyclZVFqkKsp9lGv2wrD4h9sgPXYEkb1JWaDfUhqrVv3xcM8Lq/gXzww9Ajf
0BOk4QdeJYDD/GUPdkuRuV+unwXXqHL1EBoe93GLR6BtAG58DVaMDYZ4pZs7JOBs0RadZZ6GLKvs
XW0gbvvXCBznQvGYqeJgD1GOMORyJXgsLx7PR/a4W9YZlEzEClTRGf2wTPPpa3DF93nS94mxn3Kp
n1vs+m7GCM1tXwiHuFpxosMvU2a0XikzH/Rlhmf+O3TZQSLyVRnZSASK7IlenUsFaVkgTLDfoDH5
EdytxBOV2c5twsL6Rcp2liHvF1HjG7HrwpnHRC7uq3epMEd4gnYuc2ZV8yj0oMl9Dt05mD6JR15J
u+keXVx+eQA2oqSDN8SxXSznZwx0vtSFD6+XroZ6oOCpVMQd5UZjyrmAxaK9Xj/Pr+sSgZoJ/H8o
guKo/5VxmGoTmGu09Gmrwuef75NzYzqT4vqgTddZoN8dSEvP2fgdBEW1SmpNIdQDIRXCb/OJQy7m
y4cWu3AB7jljNIAmx0T/qk/QK6vM928dkkIzrsLrIkQlie5fWDLkaxltJ04yjpkTUaS/XS1gBGLX
LN/SY+SRg4qoIecM0Skd5igH52P0xWWWXkYtnzc/zIiZQSxo8WLyXaEt9Ii5/Eh2QmbXLFJhqG/5
17VkOfVX1F4eQ4TNrXlU65e7WfcSjhA349JIJGmcyQ1uLmffdV+n2reUKfEL95cl0llUFxpO7d0b
YJXDI30ekVPAxOdZR4BySk/kOapLBii+RsLmOM+h6VUb0Gmsu80vwNKPi3JU8h8rK/+G/B2doxYG
+Wrmm0LdtftSgt/EBY6cxQBg7or9u6KnXbeQ9fJVmEBjEIdu0zwTSK9VWCwSRlwieoaDrPBYqJXU
aub2Xi1zyGagqc4xzkOLrGlSBICFm5yzAI0Knh1jEipoVDcTju1d1wcsdNcUJYlKFvkjV+xlmPFA
YJKcKWvxAU4Dvgr3hb6JDho1Pmm8yA50kiOfLEh3qOsUSfA0SQV+FV4Os+oDHXjrdbtpLis665bi
xcJQF0ju9DfDAzDufmLTXvOgqmfSNKCM2LNoYBdKqQ3cRA9s8ErRiEsiiuXQ5psBOxp5/NsRjt4i
ph/tHvt4XSU2MYD9vol6qonFPqe4O95X2mPCNpvr8LcJsL1h9m4VUTNxrBhPa73z8bNVHyul6t/N
iPhcVC6N2fdiLxWXZrF/D9HOdWtzBP89O6fqCE1nxTKFK8AVvI+cm1V977pIzK0+6UpQg/nOeOjA
/5SrMI/RKv1x07i8L5gmXZcJeVd+4Bl1y80Nv2DTdXSbJtJegOBWTQeoWHJTG2AsEfq+IeDQd19m
N9IeNfbwdJvbOVLHlYGDSa4tC7NGH/VxOzTQdIG3tDw+0qSlmp64H/5Voz2ygPy0aet7n8kVGrF5
193fd//dnK+ImFATF4rDDLY2BmH0LqIOeGFKVPANoOO4gyAtbuQsTuweyOtff7qblMoOM3zntErp
5y5Hb1Rq2K4vqMgw4iAaRJVINZndJ6oPRtToAFR/U5qVl1/07I3ybdYJhClDBVx05NBVagOqI5ox
C1uXKL8h1VVuYRl65kSWSRPcMOCO/duEYsnp20jhrhhiKY2OtoOFqW0i8I5yoVd/b3WQJl4Ec3ID
HuJutwu28MR7/hP4pQQzWpkFLr2HuJPzuXp1mzEoc7AopPtBXd7ApAGpggOgSn/e2QO7GwzRwgu8
QBidCM9Fu62hOBsRfiTiNssdsXHk5/0MetMIvOhtX+rXE+fHKJp+2M8KKYv+hgB0aZXhUHNF8A3t
pumLc7L4O+XlkGSzNc4IpuBg/0nYi7dcvvf8Ct0LGjup1dFYpoMac3JeQ/pEexdqSoDEdvWGc6Rb
wCodjnMYykBAi+G4IC0vFD+U3taTvnu9oFeTBYFrxfPOORmxXogE3Kfwyt5sQqkwhOFtz/+smh9z
VyRG/1vPzG7PoLsDHIQdNn4vCgHFRR6+4U/42+ERgma9f2vHWzWQ/uuQTc3urP0nS7PDzAixMHlK
Cx8Df48MMAav2wfEVMQkkhgMoxlazQnEjAksllnEtmvBzQciP9s54H3LO+mgtPtBmNRQ5yU5R5zh
/1cSdVk8BAZlaDO+5WJ55O3KxDnMWND9J0nA0GqXPg9mGPAccjmKp4hOGo7mUETzq758rkQXY14k
+rHNdE5hKRH1gfH3zla1MlLldtYy/r5veO+1xc9sNGaFMaE9BX235XYZ2BFyhvGLpnLLMZReZEoX
XOIPlG2Bh5Sx2KhMG05e5w3CJ66fBW6Om2tKxCVth+IZkw+wnhRBTZlO83BSIIjNi24xz+onK77p
YintcztAMxfpcwE965z+rmYBmPxsDjZMXU9TW7vXmx3XnSPMz0WjQHDgtUSIZ/gxlKWgqtBSoUGx
6LplSrSCO6H4gNtM0pKORNfvtQW5wDGnZON8xKHWKoUbSae8B6Ktqrqp8qjUPOyeeBN12n9GCDSc
8rbBxqKmDDF27uQEkU+QNlpDbJ7M/vdh86RJiJdaHwYdpbNAV2rZ9VqVePFPd7jn4iGWGYdQ+o1U
K6dY6cOWGSjRWys06f8key6euCH1jByOjFVBp8bgEFOFYpLbHVFECpkwySCApv3ek0ke3aBLYaES
xcoPQfvIf2owQnqToo8NHIx6u9rXUOK2XW8LtuMOVuRpFIU/YGi1lZv6t1TGfgSEMu2D8kqb31Gv
0kG3UO1kXzaUMyf6JwabBaiJ75KrbF8A5Ud+4o0a6RpHCHynUBKFItI+m8BUi4EyPQWoBjLlgSlG
nYriUjQbVKx7jIIl3r3HuvYkKj0ytc21wYkJ5YLTv/nUpXyc5mIgEvaDawdOb8oaxePiW41EZErb
Ao7xkkLg0TLmcXIFlnDTRtJX+R9bNYUDIsErO0pIzpUawTbe3Mov5vZNF9MWSjdK2nTsG2br3JJz
dHpw/KREhlpUqg4HL56PauUldzbI8wsgjXsY7SExYeVkf+SFbum1da+a2wusvd/kFDHu3uLuSDB3
JoF+Yz9CiO4C2BDFhkiYQz996BshFaMKukep0m6XLVHgjZe3elSpE/VLPAJ9dDQQmVrrAdP4UUj6
66m0NSt8G+8Co3tIy9RdR46WeD3DXG5lAecrFj4JLFZZsw78BiZpwCLoHyON04Uf4FQu7BrEMC5z
JtrJ4bWJ2mSeRfi4NYhduF6cvrVLpEDIjxOYfTsDo0TH9+DOGXxFMbF/Tn/umdNTwPOHd4pgUZnl
NVwuz33oDYuX934ymRHyIGAWmIip5Bqjh6NqErgInDqPoaJbxBe2h+RpE65GIDvN/Q+UDMlEWJdm
FV3SdoGpJdTfQjwllKW+WoUoqmmUnQelslnYZx+SDsRG5nhBiT7+CIAo9/lRg9nS9sTW/Mnc3t2Y
taiKQDkePy7RZsAKkydfkF1Ee94EcFkc6tohz9hVCEAAe4FjijsJ//C+kH7rAQ9bkhuOzyyHkntk
VHYwpt4seLNXfoAe3M42Cj41IREw1bX5RiYy/3EMFnj6QuN0pzm/Sa6VnJdHLb0Z3nM6GLdTy6X2
sJYFMRFPgEOfx3klXM3kp2l6gq7ES8lP8ls7seLcusN1pI536zYryfnbQRD2d2SkIh9awdG/l21o
xwl1aaG/q9VYmIkr5puA0xIXpcBqeyZTShSHUdFYQjnaXHZXSxqB8yU0Uh27SEIy+mohUwPrNEfd
bTkvOPV9yJOZdBhyD4b1Ijl3pXcZq8pXFTM05rzqwbFwt4JxdQzA4J37hr8c3JJgS/Sm6VHqVZRy
colp3sXRBwQInAubF5XqlRyZ35+jGYsrfyC4PXtxpCMhQsZV+yKzxUzxHqZT1mxRPQSuf47CIfKa
5uRf7F9fQQpa63FmLDnrBZnwxKFraMHgDdqA5I/W/q056ocsRufMm/K8aQQ/dZrbM813TCVba1l9
CDc8OiFlYramVxJmjDdczRMUaMYKSLXThOwUdJ8LPdkpwrBzr3I7Ac9WLQfXwIfIkYgcUVlc/3ut
b5PfuORDyMXARyzbHgMsfgEk8WR7qlU8acHEGUM4Xl8Ou6rSpep5s5HTIfmdixX8I6itZxUHcoNR
B8JGbeypBM37XFksZgoAXPKcbmPbCLMpE+BT4VZOdtIkMvxR4UlOd4+H+CvthlknpyAczAEhaRSR
gqNMWizpgMTxLMDb6L3sOG4TNJUR8Zq8kMQUug9e+p/gf6O9XX5rQ0Lqh3dVWl8xtHCP1tnSugjA
3LFHMvxqCEQ93paZOTd876YJ2jIAvU5HwfD2V8lsQcFkt7XPXPQQd4V9WZQLbVcj7U8lxSd9+ETz
nmpflg4C273Ud5EImyMv+JKN+TIjvMNbdS8vSdR1Giq7lGSeaXXdrSjKamQK+0Mx1ox7clHsXR9X
ZBDHGI4+0gEBrOX85YyAg87McmskavMosOduKYiQ9+cAoC4xGV4hJqZKfUp/YDdx71C+hnljBo74
FdNu4n8beXnR3YbIBlg3WR+J/RTERg78diBmI2Cp0k3V/RLfts6JOfEXuHcsJ2pb1dtuPYftewiJ
0EEqeDs4pj0Jaj15961pSGoCnTptWQIg+UaqWqAZM6+FhPmgcqDHXkORxRJ0UNJkhCGDDjPNYCOC
DowY80VNZU9weKkbSF7sZcmiI/bAo9B0IUDuuPlqTaMHeNwQkCCQ95d8G1CmGbgE+9ibWNV0+2JP
5/wayRcadtaLoARsUPhlTvKQEfqDAibLkcwqGTkL7dD3EG+NNjG8QN6fZH93plV+OgF0S/M9efGT
N5hRxrFdgW4ptadSoU9sJu+35Zn8aHEqOs1LBYn+CS9PlB30IvvKTSl9FfB0d9D/UY7luV/LstYu
qU1TNuDKQdQ47KlwxQIyIKU77sryUlRlb78EYskSqQb/q6W1mIQArFIn3EwY5FpEX21YztIqWUEa
Z+6dYacU9dkKn1Jh2a4JWXkJIfTkMbT4iG4ZvQ7mftXUzFSPokIRelBlyekoDc5usBhyBvaMXtTc
fiGLyKKaWpE1oQBf+BL42AsWZ8m5VT96Xz+ubnUedvyeCgtudoxageaQilVbPQoYDuIDNlaF3FBn
rPMGuC6W6OkFlTajWs9f6bBPju1SVZLhE+21slFbg4GJwZgFksYrxFibzuQiGMQ0/u3BpmKKiVxk
iz1s9ykMrzgiTX34P+KEBI2QoFKs+FjpBBJUlunnWtLi8Cfrzw9a2FOCFRwf/JA6qKoSE3KZjXmJ
g9bI6jBLNe55uUvFSz9vcBgjN7cmCAcCjDWIlPCOoVfsYCuZF0eZdfmrHvDBdArpNe7aNm2AUBZn
EaJYDmAlxJJPXbZ8ul1lWFUCYU8ZdcyT0XKWkjfATIVma1m0WqjyM44q3dAnbBCqUtv2nG0SbMJK
NLrKhpqtd0lvQuRybrwGKmoS5sl3133JeuNWzx8af6Ovd8H75uc1GkwoM/mkjOrY18GZHSG81dmm
nNnGF4JcY3v5ImYAVGst/UYYH0LO5dW//rzo3olyEpn+2pGwlVpFgE7NrQAu11fNeha5tgpHyqYW
RhVH4YwFMDAaGqSHYTDLawDEl/7BTYo7QU3qAJ7/I7P8ND56JWW17x5rE0Hoc3AOkAO+oUbb5KKb
f95zVW9bZMmBxAt71LPFgRm1PUqVax2GtKag3PL9t3bNHQ/9tPZf0INjoadKQX8Xf4eOesozCGkr
duOwzCdtRGyuajHG5UwQ4/0CYjupXxsJ9CiX8x1EEAXancuXfjiHdrSsrKLP+eoi9FKVkoyPrAAg
Y+mg0IlLQLwH0LvdDA/OGL1mvCtD3bzjiAUrYNiBQADmQZFJbYpgLae/riBsVCsTM5oWOH9mm5w+
T8a0V2HPG7x6BdqRIGyjhRg116e/XEToTV6/fSEVZabs19EIXKgVjFnv7sWuFyOOVRBbjm/5QnaK
qJwVXrFciodjfeMWHnZmjHi/ThiWfwXBL2bpp/yhO4eWWtQbYrl8Skz73y7vwn/KRlbcYv6wNQ6a
oUpqoQWA53xHw5nW/WwVR+4g98Qof3HJ0URlbd2plaJ51AbDK8q6u/9zNoc6to5qCId3gbbMyJe4
37mkaocgWU4XNgZ6PlToK+B3qBq3UEn0ItAwFIPIyYCpFlO1NDKjWoPnEe8eO3c5AnbT/94fCfbf
rG8+29xuc3fPDTDVcEo/3/lfsxDJdJCkc2OJ1W+QFcYcylU87hRUUJWRuWE+6W+K+5SbUSOlMohM
eVdghb7pqlwEWMjN3GDGNCcB3xdb2CLCQMovrkZH7AdzkfHWtr9S96DLpMAyHS6srWigJPUeovQ4
MnwoSR0n46OGW47r3CivGGy8cED3ADxIu5orLa6BHKAqVPwGH9YLXI+j94a8MRrfeLHkmGBNHEJp
qMG2jQKhFUpXEaHNcGM+WWmqEJxOuxnJjkYj/543Gw07eAVCVWOATaObeAfRxsDFctxBqNQ3Boc8
iAZ4F0vv/eWwFkqT+XiKDb7QWhdybCZHVgDhasOPp03B8R3xm1NCDkuIV4tb+oqSvYkVHs6vkOmi
lKT8yL9nq69ESLTApS1yCeRXpt8HmMFPj4pmxBCWXoXW9c/lA5rXOhLIpJji2WDKpJOfkEmdbY98
FSUe7H2aBjJNXtag0s+OudoOdYQo+c9gErn/M+DpLrH+GmdH4EfhCNw/QP8nK+xSdS2WncQF7nLY
TGhAchHXDJ0v4XfPYDDjiNu9Z4UZ4+CEfYA2AEeGpc/jOIKZifObc2jLMuI6+iD3Jrc8sYAhcnLa
A1zsolAPwxCdnuzinHH7wO0hEbTRmJWQU/LLuzBFRB61hG36YbzC8KWWgcQ+rzQsi90zaiT/oOQp
wcPnjh6j9RsE51TbCfE3/a9YAYYDgrl2WQYer/j6vrjQVGpaBgNDsZxcI15Ir+sv4t5Nmu1tu9ae
OzK8q86HNutNZw0gYTbsWg65129gRTn57BR4EYlsfMToH7Fv0Vr47Z/lhHbBC2V6MNmCJ8vbwjeP
bMi5adVnoX2h//nT7JHcHuUM5uaxyoXQLUwiZUvp/NmnGIaOkc152DX+BdPgZhgMBN7vBDwPdCfk
X07eg3P6uDtolvjapW+31JydwrXC0nVxPcsejhCZ+ZBVI1tsSg/8UwvPv0jlygEl0RhmC2FF/LrN
PAN9kF89EYvR5w+GE/t0ACDwSPFLXytVJO1R9pqKINJRHUtWIdTziaMIj5X6wQTWRNEcWyNfMQYF
0e1EGT4JKWIRWzKtwfl6JwuNXlZd7DUB17b4gjDvCtON8QppzIuOXcpeuGnbpceic6IRFVscmj0t
72xvpsls4FxzV2Ni0k0gGpUSkM+b+vSvMaOBFwOKXyDBCyWirIFBu9DFsfno/WY1unLZhVSjZEcI
dd2VIzsMP5nRuOmO/xZtsrAH+CzS56ztwfjNAgudN0gsnuEnR6LNb3bHR7WKHsWBsbsb+pDEcIHr
39C30LRZej8qpbI/kqOVio+Rjqrec0FSSP5wl8I66TzpGGTzGSgg+xKV903hL7ROqmRVPGHfrBKv
b2TSoijyo5r55Lh6uV0CufI3OR+OFtbMqSsLZXBxQk+RNOusppNF3c+QuPdtgUlrlkt3v1tmxrlG
KnVsGtTbLrMx7o7lZJSBYfJK4rSv8TOZeMhrKr4woARLjEQU+pQLsaNtROEGyf+pL92a7aooYZoF
37g4BmPqWQQ0MKQaj1jzik25eLrVPgS1ONqxNEqR5+9X/zjJAONY2gOcAcDxz5pqY/58lvgD6uDB
/4OQmjllKepsxvVa4EMspXQA5iqDvyqbSCT2Vd1gsFCAEtQVaM2leCstGwGKn8XEPrsgbBB9eEx8
A/+Ce/3FwjeCwM7083KbO9MPmD4FH6h1Mf6MqSpm0CoKidQJTql9D/kXxyk+gWwqzKLfPQYiYmQ/
w7giOIBSfjnhyj1sD7niW14vl9LEkkKRGibL+Jowd5oZ20BkNkiBfDtA1MdYoCog4GI6CitsygTM
BWul5LNTtzHaRoKvQlDGyAEorJMedqpOApgQYAqh/UYZ23rjfdsJM8MLMh8cDLKqFx37EO86dVxH
mniot2C2zqb/rQnzPkSNf1MN0B2ewLapeeM8mn1kkzU3Y3ikQuDAn+f1XBSofS7pTAKhSM32OzCG
bFAU6Q0Lqe+Ps+ulb7LTTgIJnAnV6pfRihdRVxnIWE1zBnfrw/fyQMR6iSHFcr88cr44L/VBpsQ8
KNzrDiprFtlAcX8tjh54V1py2NYYO6qQRdVOXVuSOtKjnSUMzZMRqAMoDPfl34ULRkOUlOMUYQrU
Kv2Q8VOCfmY+Drv3UlE3U8BZaA50B8sc21vZdFw913ovMiXPL6YcL3zdiJ5egsYxpq6JYKkqUSZJ
A37cfncF9aBuPQ1Oz23V/3o1izSBe0h1Y1kLlCdML/qpD+Bh9+2A5X4tW/vPeNe2J8IwZUMBWYFR
7Z7ptV2rvh73BE+FOvenip91DDCfnavIAATrPbMxCmgCfI2DaytMR1IXKGb5tJNZjffMxFJ8n2Uu
JMwyrL3Kp76BI65xnZYe77HNyvYkifCbJBeqxaJxILCr6Hc1O2zozIfdkQ4FdvX5R6CEcL0iliyq
qAQG9JHT5u/vqJuWTTT7pRuKN3uEMzpvv4ScMhN8fwu2oNUxW27Ac3QwyPHAlSvA/LRVIVhj35Zz
uL93iQvg0jlFbFPpZBHl2MloqPkrunk8U/JbEBD9xFbatI8Po6RySE2OOesrwAvKljmKMsK5AbG2
X6ZGkJvORRNuGODlX4idmBUrmSsQBD5bfezDMrV5lkFNtzMMWs2hKDsABnDel3dbSQp2vk6IZy9Q
d1pVR8TxUgjSSnJ6Bb6PSGsLvV/Zxo6qZ6a/cbE96kN5hcUo0mIchPUIf58d+kdSCnIQZUAHxEta
IhUfftKX4t5TWPomCRUs1VpiV2ozEcOz2lDqtIWE70FnMJE98BBGpDxXwV3JcdNPr0BGYun462z1
h/4/TLboqvt426J9w5Kfoc/JXI+ZDk97v+G0HRe9PtTmjnrixyRCH/u1RiERD+gyr9M7KLlOPYZb
zBVM7sCAgXPZzDNa2Sqgx7OPrbJt6kEfsZkDSofhEonO91hnIMJp5XxNNA7ZUOSbIFFhZfvMfYZ5
ZD7Rfjmg4c75kOFSGvY9KNc653RP3LS778bBqllpHan7cgYqhlFtyOb+E+h3eGSAcceM8QBytQLo
U3FIIX7+sB1/m79oIAGLgW667ksfKR5+MqQ5iFfEiUCq7kx3vYhCaACytDBHfra4iYt8pik4m88G
bI3kyYsTYmklDgcrqk2kH0JHntsyH3JO38pUOmy8NR+mOQQR3rDF3ufC35LQieSc8VFUFTSoYNIR
v9UnMXqWnPxnysA61cOWiKJ82NL4el13kx3KJ8Ey/nsOVqC/07FVaPXbwCKjwu2mfiCymItAGZ6q
SUP4sxzgLMV6tm3O1evQNrekTteN62lvXVCgzrvS88vCUYsGlWmjVs2XSYhIdmw6sNniFow5ToKZ
JmBBHodXK6BSzz/l8QDk4zz612tOEUz21eLYTlA07upi/+0Jtpj1bL4QNHmhcKjiL/TuR2O8twAh
1jWnxn9unfH3y/YpMEfaAb4yzDPSQpx3llbQcxRZSv0eXqVwFhuO2moh9RaP8dTPGox5+UMUfoS0
/QlmbQ5Ww1mezlRMNEMB4N1Mh5ovKqSBNLZIi4Fd1pBu6gCyhS1al0ljoEZVwIOq843xOGkFgHKt
Fb7FqhoK63xllBspW+LV/+6b60pvcUQLNSiLbHZ18uAvxROcnQziyYxzhJlnNXHkIwvSOof26cSV
Wnf3XJOL22N7buT4iEp5oiWSBmYY7JP9O4bURzjmxHViZk70bl2LjfMYlgSR6TI2MOEC0XNLi2tg
NGv8IUm0Pg79xu/+M2QygGFVWHx+3KzZpgnmPtnpciTHQIGD+vGafXwDAp2b57pc0epbE8Vcrr/K
6yQQ3HcEKXJwYLZ/qCGTfZqjUOdTL0XwdA98mzrqyeTHxHXOT2jKibMsejDeQ6tHHGwpX0LiYBJF
zf6Llutb1pvtZ6ugVmcFuImqtq/UJuwSEXxmUPQoS/3nXITufmG23kHGX70/5MlHijOV9fRCRa5v
1lhcwQJ43qpKGJg8zBI/bk76Riq3sbjxRMs23rZQuk1SjaUZxOw8ijBlLIZTbIJPWlAlSoTmxLDJ
tUVvVrGhl2k5/14CcLMLF9JBTY+0/YS53KyZWpIN5YFZPTFnmHm6OxdRzdsIKi5TM5biNoirZkWK
r3ZIILLEeVgAQ1Ql/PDleFHz0xz/x8J7K3Y8C8X5Xzj8JFInV/huM+WQwIDjO7AizHsXYeI/kdAB
d6IM6VfHVCtC7XJj9a8ZsjX1rc4MbrgmeVamo1QtEPgUaxFqrpBRuruha4BSt3sihx6kf59osGzI
L8upmkpjtOaK+sL4fiXXVbKwBZ5KMworVR5SmSbIAuJzvN7IYN+XI/bdlg78/3l+6cWJXDc76KmI
vtr8VqKvg8tDlHKeQwDYF1oX0TU3lFzGxoy02n46v3+Ii70iW5qSartve+MRQHr+/LxSKPsOBVnr
tqyHViLNuSc9Cnl5oHIVNx3HDXGp3PrxvdKd9pc2OKL2KvgKXvIVnvC/PKgaUCegHSGy8PsXibi7
WNqBs7a7bU8MiPdVnsKjNkaBcLvxJPY4687Xc516KmZpwQAypUipPA4McImIifngOzQbXd4pvJPa
k7RGaf4AgdevnYrWr9rl30PclrabqhB6r3vubIDPfvUfGGHK9+hM3AZPcW+2DjYpB80hLyZjNbQ1
osfOUGi1OfXizqrkS+171o//RtbQGeR2aDGrn+trWLjP0i/FZlD1lCQLKZ/BWK5uPYNUo+9LBp67
DRx+4Fqv22sDAX1fPQXS+42KjkLRwOs5ySu/CBk/mHxw9iIU1Et8SzBX5pgvsjXyPWPCiYriBNK5
En5dV6FshV81KCx/7ayDJyFmR161PB71XqH8e4NFln5O4P+ghdvQHmdXKGpDzoWs42N+EmnFgMA6
U53el24930FdWP+oNI7Ze+oeXFG6u4KTabytHRz78lnlhilXo2K6duFWSTXe4WEVhLFsAusTdsma
E5+NiB4q467zaRn6rMaUg4qwgIXe2xlFk+8AFfIXydTQ2ucVrbcmOTVI4W5Oa8BtyLghZMcXjUkg
Y425BPkU1rTUc4JBswGM05++XNO2WuRIWI4yY5z7l8RKYCfNDzCV1CHvXIUn5HgzyvOnrJXYV/hk
GibYxOX5/BNqwWAyQai2pSCyu8Qach7sRN9+ZbdakU+AIM1oS2qBaaXUgHLFHd22t7M/4GEmCLt1
KIjuhs0PhiCCRK3tbo0pzonEPQeLOVpHf0Qa+zx/PbG2Zs+hccw9zsNjgRhJ7Axda7N7MJBLntFj
eibufqUIwy3ZYJfVQ7lId+l+eKfHh7xRNjw39+PTjpMCcf0D1Mce3laLM5jMYkyduqaiLTc8qtjX
D+whi6xJDRdT1g+oRmgzLu7Cp2vYMoqJ6LWTUaewl9imd7X5Hwcy3+xrh0qZGNYITS4uwCpb7/Xa
XiNQMxTZ6m08FwKHS/7VclzOIpY+xMe3jcyuBiVzDqWudjKagnDuTE+jJpBdl9RMzmV7HvssFRGf
J1m0qDD/YVcmhrJJP4ha78agGKFWYe2fr6+bj44soBC+Op9d8cAevoA1j3xF1JzSlg0z0woGWclp
mOPjM0sJ6H8Cu0fmgZTR3XABOPi/DYzCPSddqa5TOyW0+NDcWHPVwJVHxRxFOnb5V+j5oUZpzBqs
oFM7fxNf21qcKulhJiRb8RTbhQAzgPq9Eox31NEmHQoYnkONPYqkAYDEtLhk2ndS5mA9a4OSFbzf
elR5SU0Rbpo1HF78/6b/uldLNbpvFYFVUiHMO6ZacMvemt+ATpMQhRIEIMVBEWDUl5Zfh+zQCyJw
dcDfsVnjkW1nj3SK14FYM95UbewQUPxdx5aoh8UtYpL1OqHTvR85prnCl41bXMcxqQRy6lrTaXHo
S2Qsba/HZbAWAeFgBouSbCjDT45FZkftK2OQbz/y7Sgi5zVj8vzHWS1Vr1wO86Z6bDBwUtN7t9W6
YFKhNhR+mL+iPl7qSWZs9dEmOiU4eeolDe87vymZTcJpUtYQ7d59no11i5Mf95GOuzNR1xYeyqrD
lpKTn6ml1Qie3plcVSUMR1ncewqWd0Q4X3faOZO0s89LlLZR818OUaGiY7wvmoPesUQnGmt+ppbj
aZdPu91VKSIrDv5txPeoliqKkpf7vzY2zgQF1aXelMKpoi/iw13zkQPnrt/I/5pVdrW8pFTJsU7N
ArtsQ/4fz2An/7wyCm3QqYkwSYS9xeMGjz9rsEwEwZkYPIArxdBpL9u+mogNydoOMbp3cDkF0zri
Jj9Bcrd/Utaeg9yJL/t+PQosPjyAPUYRNtpvfo4xZyA3xxE4LoZaDBUzp1Lz4rSJHuK4A1S6OKcb
wRO9jj4lzg3ht8vEJb8YXBJwR/Pdh6aRZVfhSunuZx/GCqCjw9KW7wjaapYItveHVcQkhFoDOl4O
77C1l44koR26frkrXdgehQ6RDHUiouEtKTVrY69IgzeZDBFYyvfw+YV76d8+pzE9UCOrmoZeMHpO
75JuMc+n3gE/ckJW6qISTyzsROQOCW8EzOCYFzt7SYJf6t+z3MqDxK5tJXlH/m2yWu/v1E8rTub1
ZWMdAnDDwSFmaKovfINvjqRJBIGdDHfzsNdcT8P9oFHj1Lel8fKy8yicc94s3khx/iLs+f4W8CAn
mANeN/hWsokbvzwzSG3wq7vuUhlg369dZzNf4e74JE8RtHRJ7xbIqt0fFMu8M0xFoy/QXXHRfBgl
JnmvPzbdhtuu7wbv2f0tTZ50o9GkBIPI7dVIWMwTbp89tve2gI5kdP/Mol4JXu+jZn41Bolj1koM
ftpUpdtjIwf49WcGHWyYwkftD+Fe7nzsozJTvdXRHjyjdxib0dWJEFssvqt82B03kGvtXkQ37euF
hpVOMMsWbca4gqZwHQ2jBumsp8pe/fyZ6ryaQY95B+igY0kK5T0IECJiepXuXzVXnX9HFViqLM94
3NrCAYbr1rB5LZlKHjjplO+KorahGje0PRb0uIPJPM8vUNbey5+G9nJvfgifaZqs3wWJVMr8Hwq4
PqqC5uz3Kqnh3HT7Rkf+DhMwE0EGtYcbTFk11Oct2wqjTUQX/8Cdav2PWXMqn7LUiwYDuZwLJ3e1
XublIC1biA0ec+WxVpgMIAlykvjXclxYUguDeY6zUg8KEIuqFpA46DzvoYUEB2ptAo7S4DCvRX8+
A6vqb1UTEXmt1+wvdsfiXvTQHnUhkhwPC0Bd21D7cmU0B2Gd3GjsdxKnQG4lzr+03LzxdC74MHu1
U0cS2+Sy0S5sC3VgXW5FTd6yyKBrGc/q1AeyRD1hoSPYcOsJ8HLdWVEqho4YuhBAM8ckDIjI8Ixu
m5gW2UAW2Swf1NMR6fTM8MiDBxBTkcSSxEeAIpU5H0xyMm/n0nqvdmjYgiMwRHoGwh5FPZ5A43oL
ur0VKPDyQMyhBI+4qCM+Hx5PtLDSzelV4TrrUuJ1gTAgS7INo8gFkVonIMW8hE3tQzSlQVK4Jsv+
vsyRSdh7yUkNR29ig5cNqxJyggPJvKLXKKln1nphR1c7JehMQSzsQ3CBLFEm+/R60cguIhm7hdr3
SYLVhZiFvwIKTNH9tio6ub5nXvJbnmvxfO8P7bf9286doIwg6jbtET35VruDXqLC4F3bYsnwrx8H
hUkZjSdiFkZ1SK9z22ckHTLIxYQ62QiBMFfgNsUebFZO8dg2edIa2mn5n9Ldjprrt5KKJk+KsYcD
e9RuQSveUmkW8d0Oh7kwHSLPTBZj6k0cFRiAPxqNhtZ537xGN6YNCHGFfAQvcbDGXCQ2b8Km7TNF
UdRVR5MhBF7LcXGLM/PFUi8eV6TwzYOxSJI5zPjWGZew6zrFtuRv+ARjXEONeuU0iP5Yi/m8MFuW
v7OdHKA2PZSDU7Azo1IwIsTIJFOES4dFxsw23UF4SAu37JiXUzqXjj5SFOBJS+ZXdqQ0c8PTJ4my
6/42yjlHm7KVxAiTmsCGByhPTePssRQsirvthZcwQup3mzO0NWKF3YC//igXZJro8+M5lVIFGs+w
en37cTMJzo6Wh5PqIciP0LCryjzVosAqjwc7+e7QoDln7aTegm/PPJClkdrzEDXM6H76sU1esnLY
1++kchk1sxTRrL/Eu7t9XtXzs9FVcddd7D8i5r/JJp2Ejc63Or2QxpzkAojAxTbhPDV8GmJ3rzYy
Md1W6byjjf94blQeMyLhArO8t+QXKWZzfVYWTae6ufmSIjECY2XR6n4ET873WFdfUveQdNIUUFKZ
C37rbTpt2Hzcfi1t04wsNlT7rCoXNernXPiud4nX/iIgm2pfdse9x2rzL8xbNUJyLws6xYao05gF
irZxspBkwFxg7yjBYH9GLmeeW9wmkNz3iJAgageTzQxoeSXkrNNqH069gF8Om5UQVi7av6lLTfWD
8QbHQ+nK1jJm4b3Pj312O7539H1cpjKH+diUui4bG02lIEjqrASXak7l1WjqSfcffq3+9opvX06D
X+EWZfTvZYiuW5ZXTPQZ1ITJPrTle6zoXZ0op2qDJtrL8Vyj/zTAf2Da9NQkKqylI79QXB9x5laF
OQthZII0tOCzokBRi1sOmMayJHofYNlwHejd45blmYb85kb2BM+2c87wUzQgZOeUHWMJ1Q7M0ooX
5RXp5DgWag8PoWB0oL3+vZ9Pt5t71onQ3TiTmwy8+0qimRXs7FyZHlxhnr6YItviWSat9JIoWXLC
TEGdhyNJQHxlR2GE2iDFuI2bqrqIYQeSU1gLAnwleTbtDFaQK9cnmlspDwz2TV8tn5pyq7qflpHM
OtiWPCsH+KUv6rVxMVggc41p7lNTH2A2E+e8/8b1nMWSH9zBWP0LjAGvvY1ujfadfAAt3Z+igxh6
OfPfDfOCXCxCpzCCV2BBjXL6nAi0sHSrNnBYYuw7Uq1bXoUZXToZztrJfeprPDaWAfSioFSPXn7N
Cx/RqYpE/sHfeKJvlZ7qOP6tnV7ny6+R525O9g3HqoP9mdfSYF87e5jvWm6BGyzZk5kA/t6qabNY
35rZ8KF6S+NlHvktrhDGHi3HNimL4/lh7RnEjAWDVjb1ta3NLboqwagC2bttaSoSV38E2L3dLSFW
XDi9H1Px78/xjn/L02g+n6/+YMcofpWxJdjzfIdY6HRF5R/H67hcx8m3dpjRMPytrt8o0yF8/oo/
+lQAgYpEbX3WlKBhITI4cgpZEXME7RBGi5vOug1T+STyDPnGL/ncIFGK0R+NJr0v0luOsP9c0+Ix
IW8NhoaSRVkGX0W1THuSrmkDZrIDYj8uIRz4Xv7h3T7MyMkszkYAeJsWaCXpY1CghMvVYW/mMiEr
YuZUxa/uQln0tsMDvr+d3HhvbQWeIaMj1xMj+A43Jo2lClchF+5niBumbQrAH27654ZnlAqFW1hs
Zi7qOzKqnM76suH2z/gRx4Q2dENKb9UPN0jzRdEHjZJeD22ihWik/Q3f7Qt1rN0OFxZTgVoxvP2E
3uj5eKzSVS6p5yKm17C825uBiK/ayH9ep/A5yTZZDT/faQE707zrHtkvMs3crZmfuXRKFZg7Uu9B
bGQBeKUTcTiKbUX3VxmRwBWX6c4eZ01euXYp3af/D6YAzvp05Unt1UzqtFtnfYyyTmVcEG1yGuFX
oKHq3PdA9azDfZN1vpaCeoMNUOlaIPtl/3J2F+U3HH+qDoNGQZ1JH+GH1+ZU8gnyGTu/VOngb7c0
ExXxsEH4P/YzYbsk2jewhn7ZfQFQqkudFPn3incAatvtHKq+Cl5fMw/QF4BWOEaBu/EPE7DXiYWF
qMfD76WNaeLk9Aym1PHK3rTqVfbClO1EBqysWawI9ACSM1R3YOKYbOHhz8JsS0vmUjxAQQPI7ziZ
5O9dPMu9GzezyAgQVuLqhig2r2UxWsKIyDn3aWnFmcKWoyEB1kcRgzYGGHWPuKZB70aTQPiP8M7C
bPvBpbLJQKj4TOkefzC80U7irA+++M7e9zoQ35W0w60CQAYcHz/nIG5q18R6JD/bcuerFmdfyr/n
BIcYhTluL6bHncnCbrVfQs91j8VytD10kg1YBLjoqhXpJf1B3amkuwMQAgUQfc3CswXVMmWSZfZC
pTk686Qvb8JeHRs4cTBnRq1dPtPlDXVA/VF6yDFy4HSS2FkqcFkLLrF3bfIzI6HHm/0s/OPgaKWI
fPXza7suNLejzNLZ31RcJq1q9sOhHRwYf5RklsdLU5TfqLZP7HWi4xsKmou2eLsSXLpULKh9hFUZ
iwsmJciff2GrAd/rLxXjQK8Pihzwn19BRWmSEdZ6nJd+bpckCmT6RT8/5ofhdjccs2qDvDvcVnw1
QaffZYBFKdOTkrbzYLDQWWZTLgg8NiG5Jwi3lu5EK5xh/HSADhDXGDz0HP0xNYOfG38GiN1Rpw23
Ce9ZTAz3HsqEpaTqekO3rm1gQhy1jlXfM6wTg9h5SxMfjM+DO/iLAkBZiJ9YnnCQO2OXxoP2fAM0
3YI/jlwWXB5iGK1uTdd3U2Amuxkm31oJ9/k3wpo9Dqjd+MH7cfmYcZl2OyB49JFY15uTQUCOxRLg
C3ieVWgVCLJZgCzbcPLtnP+ZH+5JaaJKWGX17nRPX9gcIAzg7jKryfyWvgG/eVSSM8fpd/sec8di
nMmORP+SsaER4EzswDdR4LfUfwv7whdOgD545zM7DNjDfAnD6kwdFHlSXkUCVcd8be0ctbpPbUAB
ZvbeMaF9QCrZ6Bs5dlMUtTY8wmCIn1JqKVpxcHJA1mU4R5bj5fGDhksL4m5y0ZrxLTNZTFea6rxZ
a2MVWJUUKACu31EHaAjAyfkgAV+D2N351zMCnaxZurbf/ODUyQi/K+vSA7YD4dWd8/UTddgX5GbD
kOriPZhlFTJHwNhCYd6etK6p4J5cBfjV/kvC3Nv6z/KCJmWdPy0AQWXbeTGTaJOTtVSBLjDUT/zX
okDB7AvT634epz33eLE7sFn27t7QBMKY+6++/5/6Q3GuBj59xil49awf7dsu3mBnxnJyPows2+8t
PBRHtWPbFGD65ZIZKA2c0CqYgqPrk8kpGcqxW36TbelmoUwqnmRMQWNiQFkgjT9NjiBmjuWB/MFp
CRxtUzrsLSPk74GYzihoCpCLQYi8tucA+MnC94cmoMStLZpJ/p8iShAafgnzlitMY96G39KAgngX
+hnIn9w72zczM/a3JCCSACeQFqMR3S4nphmfA+PqdFf7w8xxMHBS+VvJZ1m6SBgzp+eICxxqCd5B
zGtm+NZaoMeV8MUDZvc4CBPbDF/ZFuHh51k7eiXU7ZA+MBah+U1usS0cPPdXf7ULh64KpchEdADF
XNmkX3a4nKzyOnTXiimMFALS9zuI4I2mAHzlCREpQOGrRPqriSb6hUmVQlLW+lV/ShtmVqb3KPzd
V4qCLJVRh6KCXlBXhzCcXMgjfPSqcZMS6JRLQ+Sa7Ww08qoXpqVHFdlTM5iVthw/GwprreyE5Bzw
x3TephAcq2XirJe6f+iFHuu5CvEdRx7rXpFshH5EoIncc+/ZoBZjEqDvIKY6W1kM6Gu8CkshSsOz
ePPyZysroGmzxbNhMGfi3y4rRSD0yx42cxqcyTvuIQujOncLjubY4+gh7wuH4ag9cCA4F9jSlNk0
wJ6ztp5k8ZUw258EZbexfvhWVAGJw52Z4RbxR0ejVkBCKmaOJwsj62zhTRA6FDhH5kfcSueMhuXj
vYP73asX72mHAVuYEG/kg6rQGx+cFS2kL/tMo3ryhX12PE/Rd1L4JrNLkp2iKOpE86Tqe7wMLv4+
el2zukJnyANK4480nfE53D69vITXqkZw/M6Q9YfhFHfWjKMi2weWoKVIRrfF1eBGbFHLgAyAkSwg
B4WgCTcy8OFgJvTI0YlH0zxkqo7ebOp+ffWLsNMpGX9u98/a9Cn2GdUumNzXRw68XY3hYVp3/qtS
ibMPa2lvzx0DDK1X2K2rTsVVW2f/girhRD0nPQO3v1oy9EU/GOvlAhavSyWNyzFmLU/P2cThsI8f
DVz+MvXU8Iodpkm1Z/I5hKtXg5nIX67WKTD/fe4/schyGyEu2AAO1tJSQTJI27AI5TQvHKSjZXfH
rBJFX0W9bsDMKeGqxcIuP5XSEgUCBe0qAAXPCjJUxVZFYybCdTq4lxVixeJHWPkTbmmnKLSEzew7
i7hGnrBgH5scpFuo+mQzjN3JjfZ2tvrp11peZSkYyrL/4smYlX61JUH4LhFh1Ff+5beYuSYIt3c4
egzRokw3Fs40S2J4SBuWLK/JZ2pwzZ7S5aW8u7tnGx2vc3loc1rjMprHQUc8jSpErK85257ra1JW
8Geo/4ywBufKubO62qkznX1tRsuNJFfeqwKAN6MCo1whHJmcuAUtwpf+j2d0ztV2Y4KjAJlA6efQ
714pV2vKzKO3u1utMjNvSPKu3MMEIeEWItyXzh/L4wNAdDEByYR6tlzsfjdUOszwJXNxymrTiqXh
OpJJ9M1IPFTeL0Ej5LZu5SSDbHDfkJLfBceuF5HGJLqyKydqbZbrg08xCgdpl6O0FgwcJYJ+ZPJW
3R9ktsml+uFZtrOD663y0/0/SjD/GiYZvEgETwciCVJrgW8grm9lEp8Ej1jeBoPeCBK0kgeoFgqh
GCIhGgvTa3sT3jlMHBo/LZScmkF/uGhdlkW7pnO388gwlkxQvrbVSmMFgkJFtrXzkvQptj+awgUY
WdwzGFzuKWvUeYLIQtqihvqQenq3jx6hwMxc1zzFqY8BKXvYKTpkJ9SfUQ+FBXDEz8miGbO+/WQE
u00U2N7efzywwvfwEXtHVXi+ixN5bP84rySnSrc9hRPgEx0TIJ+JQAbL1lm8Psns066uiLLU2mCV
GL/9mdP5jpl0eTUVx/J16+jo8BAMufns/BjGVbokz9XZJVcXc9tP/BvnCjVmb55ZBzqHrs1u3cMd
b9vnRIu3/mYeMFyQ/dUjA/gCfxKIT5z4ScDCVSH3SdGx0SIZH/N4nIFnBQRmGjQYAEJ1bbe7Ncoh
28F2NxH+mz6dbYJEaa3j9WRmfitvuqHkR3KjY6x7lcc0iLq8kYCUHRBhg/7LhwYe3c1uSZtcxvOn
DVLS0YYRmgTqd3GzD0FDkD1D8UW6KUbKerRapMAkUvxNpqGGUyNZAix2GLxoJcolZEfcEJJdE/qu
wtco2a8wFwfGzG69JYCMMmQs+Rp7sBxZsiG5YGOYLtTetIaLsUK5kHhRZVzEu7JaMvdrUO5cUgtR
xHanaWtp+jeKOmRnLfA5+sX28drsqJunVOYRPllyFrLP4aiQbOt9R9HoG/aclzdX/cQMCyHFBEim
W89gxQefifirk4xJlNfli5IZRD5J8HL0u7cYSCcDUCE/07wn5jCg4rYpQi9UxSr98JZkR9JGK/pg
APk85Xw26GykyYLyYWiwqPBAEpEVhOkovYcJz2X6CTeU6z45yllsCoZbcay37JzS6xIVBkR10qhl
K+qu4nks7ahP0P5dFZZhmz2sCa2OWpFuZJ8o+sjbEnuajMvqdjaV+2hO32TyK3yU9EVrC8rmqEBL
l/xfGcLS7pVIvuovqMhe1+x7hgRDYgxf1UuG8PCNOFzmiMqXVWEOFjoUKNJ0QSG080vbWG5XeR4H
OnL+QOJPY2f4GlTlfEfZ0rH2MgFwgwX2nkC7fVy2eIcU1LzdQbe1ZmpgDb6ERU3Wbn7EvR4//cpk
TB626nEj4IKdSCGs0GfEVqYvBo051iE1Yi2D50TX5pARHViTDe9GvEV7RqFN6W5QtaLbwvKIi1jr
TiLogEdAhY0nCY2VAHbdok3z2/+semFDHPiuQ3Qxfx9rJhNbpQf2qpFPzR1uFbtcrk5qe+lkAgXF
QOhO8C/Vl15jlPYMI3kRI7CIby51CK1q/jTPQZCU+mXQwZPkzGgwjCGqPBd0YsATw+Will3FNt0O
qv5bOq4mX1+uW5JGsXeOECVko/X5WeWznuQOo3NVNI3giSg/g45kkvtRd6G/nXgfe2yeEB4YNUrX
g+Mtrf6rnfSAgUZrLvkSUvlQz4BQTc7w1eFnlq3hWUyP5MzuBm/4hpq2ya7qC8rNCWu0aPAL9eSC
13zIksyeaQuiDLy9c3iUkoA2YlZzKK5/2oRXFst70TDVYFxKF+DjGG9CkcPgMfpxhCgSzoAMeLRX
SRxU5Uw/wyCXIrK1LusgL/V0Nzki31w0CPPpFYnT+f6NT+Bx4ROPZTlAHV9oRbERSDgOST89YZ/t
Cpbp/+DcfANolsSq3Ldxi5DvLpNUxkQRupqeUNhuXaNxfwWlKEj++0ClvN/loMxDDFnTT1yvAB8k
aBHQOHbu+HKW3Tfj5vI3b4BZlKSkag0UzLE4ZzQ7f5WcIyh7YqqxuEIOAuZpLFp49zs3yyr9+0kG
yvmnlguplm2EaFhdrtpuWwy4xWM93h9waJcR5JYMwu5a5aoWdBtCc25yBLzKYhOVJWtolctczMCu
eaJ6GIg/TEPwKGqI8rS2YA8IRj/1Dh05rIDDDTDW98wlbNL9sisdjo9GCuYkIKjAH0VTPY6jnOxD
cYvtTAR2Pr52cE8d/uq7aO5Yvg4YD02BnGP2I3Xal8OSZrK/KDXi0lyCtfPj+5H9wBrY0ag9fpAm
M3VX80gd8z96w8g7bpmvJ2u58DVlrjtjqnvP9tTq7lFx36IjUlEANysFR/lscuGzzXEa3Zuam2cx
VrMybPTNHLLut1UCK34oMg/me15Bf1nDqc+BMiorU1XXhoQHoxvdhMNigiPnhwg3geLkfVSrgoP1
KRjfmTZSatfdZ+mc1g2dlde7mvFrKYjxQGXfswgPyXbA+D/aPZTXDH+zo57f/6u+ymneAO3M7qZY
FVDqtrNsn0Xw4RJH1lcd6aP+pDFJnjKrF8+a8WG7xo1kxPcfTg+heod0c34F4PiBX3J9AN3HN15m
/fcxIjtrzBs7i1fvqn5gpdu8AihHJmnZfcLLPPgrwr0tpvZdmXEFI1FyGKADpEe11zBN34aAxk6b
MHiIM+YbefytUlUom78yRixmc3eMff/u7rA9h3hivAu66Aia4QV7PwFEbkkg2hzbZ0qW5rBqK19F
nus+2gwEt9RDcYd7B6wR276AhMw9j75gQGD//7z8w4zCF3qz5s9egNdL5SwmUokzHT8obySElGtA
Kli0O7cB3f9aBp7TI87aaSkPFy/DiBmUvCv3R6W4T8ZihLM+90ojXMhYTPfz0j3RJRsxeYAFi45j
R1mUJVr2cgOjkT92F++JG2+QkP4/sDbNRGCeARphQOVWR+NY/7R6asU5fzLxmwJaGeks7W2jevjY
b/Euq+o6Wy6qyEBjOFCjgn/usHJSrVP1Z9Z3stTtFM+D1M0fLOzMYGo9jZ+c0g8MvNyPMG+v/SIP
FlfZF0SPO3ps9lWaEjZMoRy6uvClJ4mdlAnghBk6IWPdWhcyj4xrlGspx/TISHCOgOMvhW1Cqthk
nOXISMLbVK+mZtEkUfthuQ184oxmkYxJn4/vNryCcxmyaEYcbHjxB60jKAdGgvAOp7RCHNaj2K1l
IqbN1p/mNIK/CQmIqHROEJDlScfyuhBREJvHPIGi0x7MeJheaWwoNB31K8Jk4cDhhC3i6KTJsG2n
a9T07sL3pUKn6nLpOX10IZUrBrT3S5zq4qcNK/rXDJrnyluFFTcM3IAV/1HBf7yTeO5J3zu43x+n
EQ6u+/Nu+IDzj2k9wRbNos+kyhgExSJaCTfYXHwr7b2GIfZpfMYgwP41oYA4y+CCM4tBpvo2wiA3
dh3N9zzrFttACrX3qgVCWd+doToeF6ZK6fATy07FqZlnt/xstwmyRxbV1YqWo/v+RfWsQP1w+ZEu
i+mCUdZUPN+Qp7PQ4rKsRsYUxXYMcvF6ZWPTWGgkxyVKMdKd809XMryRazdQZUj0Il5ht69/e2iY
28+1Hr1gqf2ToKfk6D9CrAL0pVcJuT6ioEBiwC3vFN6Lc2aXIrTzpUalJITOQqRUwNn4ms2Qz9j4
Qyd+i6yH4AnEfednbj7xrW+m9V+jD9WSJ9TPsMUsuVLGOKAbHRsDBUSIb6o+nXWvsn8RovH8uvQQ
iF+dGxJV4OoFdT0lJEuKvgo02tlh1+nhCJYWBlRDQduYAWMgcxldM7czEzGqOH5tKFUnY9R/nA5z
xLcX2/ivX9fO3RS2N8mV/4IrD8z0xTjr7DeLy0S2HNVt+bAY1aB8Ef6dn2sv99M2nZZs0BYrsNkq
0yJSY7Amt0X37OrT5CTwlcmdfiiKa1l56QoLVDxqyQFRusIFD5WXlgJsrdnVFzYVTlsBi+jywfPY
PvCmIscuOpJIfcXvT1sCMIbj6EE8H4wE27frV5SXqEvAK9RzVQJtSLo76z9LiBe/Ja1F4hKBsw0u
s26khzCqmV5h0DhH7L7lc8zoKFUMAVgFbDo8cTl1Pr0e0CHIy/wJkfiJ/dEk2kqSQYh6kvXgKTWB
5JBOj9j+34vsF9gB7wIVWpt/ni/L7yB1UYlSS9n6C4BCcGNpmk8V46J4TEPfwaz5ggJnbXzhd2EX
SrgtNtPBbEoIzP+9e488jArZvC0L1UFmPmuQ6JoAoFOi2GCeTxPjfsPyuio2HAiFbHa4bEBKB1Y1
lYRHGFFFzZ/+nnYlOuNz8CE6+r5TwV5l+6quM0upD1JDYnaK0Cf6lZvR/x16Z7pPq5Us3zcCLxnA
x3QM7Em3kYcEdoPVf8OujuoDkdlySrc7h0ForuLwlKuUZYFA3H+lkl8JjCRtAxcFDL2KUd+5jrX2
bzUGBgvjk1IWkphnL9BltTxRDMGz7lG8RI7uhwgYoE1KZ6uoFheQ/nTyCTQlYwhXqTdjLmlMvx6t
pxpnNSS4du8m+Y6sbSiEvcFH+wxcE9t7Z9mwp8pJXzKy6z+m5KBM1kX9IkNJkTIzVG2hdZJbtPcA
df3UXY/FY7JV/Vp76lj0sTQb/ghRI9ARLfLgjwdaHH/Y9AJQL3x2Q5sEy+tIjtRPl7OIk3WaQrnt
YHQMh/5E/zPX1Nr3vYPjcL+DLkZ/2Dj4Juer9azgpU1j/Dnu41qpG3oFgxSP8FVxGO5hwntvmpsN
Cf8kTO0owQ7I4RBztLn1EuJpXt8jjc+hfqbd8tvF6cYiixMARTSlSEos435frCbCvZfKXeKd5k7z
EnCipYU2ZPj+vy5/oSk+XFE4iXUbbTyikwGyHTa8bteHUOzjWyw7G8/RnDoNAtNf6pp3bhJaJAN1
RhQ+sDSSGCHJeLIusFeY2JX0kFbXqB73PUhyZDqV9s4DnyX9EUTa3aVD0wN0rzU07c1NcFgCu8YM
cyFKrlkk9S0zjWra4hKO2qUEoByBAWfvD/qRsNw1jBkC/oblDTfKnVK1UIH2XcGkTeDHSblQqLn4
T7Qo50WBNwnLIvl3ddAAntzFylWR9Q9NAXe1sHBvbGInfZ+CY+ly/8d4V0n43qKYml1MLPQOT2MV
yotXR4D700lErIjIkdrDr0GpzD3WalpWCLVKqNs6SbRv7DX28FubMD8e+fW58fN0aVkG7kx6/XrS
TE6Qbs5MmNEuCnGgkkWRW8etKQpMUHG+RJnNSLPfqMA5QREt871E0VNaTj+VyZ58094INfg6xZRy
oGGhKsJXmJ1zNtXvGDZlswulsTvlsSP/4ijPjsFqo/yZ46FKpH75WbRerzaDJBgs1FS9PxWYC4Em
APy/506pwanS3EAx+EufRE+LOUdtHeIKu22PnRg8WL0EstaDTXLvc5OxXDRTjsd/sR8iC7k0LGz+
ywt9dFHYaAvhOu/I2ecja8UgBXU8qv/T2D+US7b5pZQ5VFcNSO9b67AwdLrymx2mByWasU8kvNRs
ojQJAKO6S/nFW0j5YbUZEL2UmQs+KyrvxZzQfgaY0GaTkmNBil/tz/pONDubQRrRAd0LQbwdtvgT
N06XBvJGeZMMwED/yJRN1R6wjObksTqt7sg5pOod33FoTVXGzah9tdAg9v5hYOAoRS3dpzo04yXI
SlZK2Y8yEqv+jw5fY/may2Q0wsWQHSAsRSf7HzAZ1G+xWo6MLiCg6akh79KZvovBbhZ85bGYnIyd
C8hzXGlrTfqrQ/l5STzwlk8YeS7ATax4eO5MEET0uuzjWZ3XGheDTxwcvOHU+depHlnOGpE00cAk
qCY1lrPLRQIYhrXMjJtifAOcbWXXyejOn2O8j0uhXALYo4bmQvJARTP8rsev9s+4vrnV9mOnCUTb
MsOPzIAof38SnmYXjRNmQHbC6QqcfjNZghmavZUG7/gyv3VCouTxzBbRGo1+gq1zvgdFl8lspKLL
xdJQzaPL+BKA5kYU33u6yAbedFO3f8N7AFlEV4LhDzmOwwU4AAt7edCkAlAd07jFGKOvtGixhBwX
LtSA4FsL7OgOr/z5RWaJAjRIVJTGIPJ70v5Z69nCv+DftoCbgB2cAwNz4lH7kxfwBCHxGuueqfJ7
swbw9LB18NRJHM2k5XSJJ3OovJh7muv33rx6KFXv5Mdt11nE0fvrwl7bBKKiM4YNwHWVkUgQIWe4
hvw53AKzI2LVVKLT6CarWoUy8Sp+OSM0ghdh+8ejUWpZ8jVrmMXaYokOS2jfAnE98SrRVFZ8pMd7
OOh632AoVzclyJwzfzN4RLsyzUiwdBlSmRNXuEVAeujkCBsxZODk06FGvIu59JRUHI/4+jS0c7fY
wTfKbVMejJMEgEPPqyVvl4rV9A8SzEfLKzOnmg1qPqChy+zL2ZAUtqp0gLz23+DiQb6RNKutW+VV
+ZAAQwq+F4ze7jmj+uM0ig7a20hvIV0r+RrZrMLfQUvgmyC4mHRVMyRdN1OUslnCear+0tgfvLF4
rG0EMSTWdSsaG5b6niWuw39OPwVgyAUPekPnr0WnWRELA1GQWyOU3N6WZjm7MATdrNXPy9Ops5Ut
4VPK4FJbVx0m8e7Nwk2mnVRRSv+1Y2rzZii+rg+0Q5SLgV9g4ITh9SxigAeU6IpGIoDcaga9t0H/
xg+MDMDNC1qQDf6YX+5oeD1TFBNi+erycFnp6YlDBsomgcZYR0OXUZWWo61KwEJqvUO+lyONqOJl
ZBYg0QXpTwSwBE4iOu3bLqtcdfyHse07E72KMsZ34tN4eYnbBzqM2eXGhq8oPVn9AsWKJiRv97BR
hhbkI/mLhWaSm52XIvkLGv2P1I/8T0IDsKthy0zmSFhxAtQwmJ7ptu1EUZtiJvAngfxAFigq0NjP
vvoFVxEcfYLJMokUzCETnKaxkSu0hyamU9LJ6sLliD/Fk/8g01qjwmxtk4YvnGxbEQqePkRooNWT
b2LVJw/2VevCmonMHrLM8Tg0lhFMpm38N2yI/J6wu/xW5JKH0sBArxpaCzESSIhDbpAu/mLluPYy
qso388uG3+koF2e4ExkO2b0vbKj9b8vAj9IIzQOkZyNQmlHajDxHrbB1JaTzwVPrnJQbtqIU16CG
PgfpNI1NwD6lljNL+B9YAvtWt+zHkBBx+9PkTR5AVx/xfILtHcIN3t5czuC5+TjQV+PzfBwJ31lj
luTK3+wBUmiByXkGZNV7CUuUx1jpuOsEUoufqu6D8GjUYWtAG7nv2yRALzV7Za1cD2UZeDdjMhYB
28plJ21fKwDg9h8LKBAl9D7jHl11DDuwkgPv031zbdNsx+9NxA0CanW7pe0WA5ZjKZRrTUEtmkFk
q3NxzHKVfAsV81Vd6RpyXvynJ0ME96n9vaMKZTcS60VtDdKgM660gVimuPaKomiXtzk8qMuzfM7m
Jre4wlpXhvuQLyT8hOj9bXo4oHpFkwMb47dZFaFvbmzvz1hQcgvjVxht2UWKWtN+hAtKnXvKD7i2
jt+y7I9d38sS92Yo3feXVRTtLvZWCmyThCBWVKbQMHWhgeO2poI/6pls7iO1vy4G6LkP1mrOeZhJ
iEqkk1LSbUNzBzq3PnIgA8CIW/SQ7hOfooK1MLIqE3ydPOFHc10+MCnOJKmIR0DRhrItpoA8AEYq
+liQ5XE6xfh5kD8mwwCdxJ2YKpKm/4kKHiaWJTYR0AD+9L+d8Zvhn/XyLsVqmMTX40GYGXNY5O9G
xL/wjQjATlzuFZOjbsIqatgW/kbzFLL7tcGMcTQFzWURYeVM6YUDRUIRopTOez0D22Qpk7yvbK3o
DP8slIEhYTnh7nlRPWDezsz6HSlo6g+ILlZAXlsb6snRL0Yr87vKtcpGbKXmQylZ5+arqtoEcRbq
x43HY+kjIp4HyHo3xCr0Cft0uT9aIq+dhwV6olcIOKth2qxNe+LBO/OQhANkowYj2/EcH0Tjp8sD
h6BX5ltkn7tiYSawh9UHIsb1cjIOH3YcH56Ep4C9G5EzAWlZUf8PZDlE3yL+nnEg5l8EVo6LIQDa
oeorax2Bkt36KV9ePiyI/RtCG39V1WqRhV7VKc2ijM00Wg7WYREUloXGUqctLoy9V+gLt3ennjIO
HrVMpxJHl/KzbNtl9C9tPMVHw0sA1Eo5VPC/CgGiP9Hnjx0FNAn6f6OJxhY4MeqxTluqoMW5VLZH
lfn/Oazs3zBsQpMFsUmazJpEq+7pMGdsG1JCPh1DpfakX/mfQBDIMAexTJgBFdcCs2QstBw2EMmi
lCiTSw6WedJQrnbx5+qeMNq9xkkWT3pcHhlcusRyr0xlXXOQubIpLKQyuLIeobD5YC8ibePye7Rv
8bsK7J+fEEODPSATJWTJeL+rWJmpZspGPlQ5at9hfOV5FIgA+QtvHIdAVBvuVQWeEiU7q+/66CjC
8dPYnFLTu0X2V/nmBxvZP5MugBS6zVtit76FiGSlra4m+MzkRSMCcXmqHQCwbYrZIKNDjfxknkPh
ZoGLqBWbCDDcpmGA5XDYHU5MzfLaqgMTemFqNH94oBG0NGxjVfsfY8Xd5e4cS+ZtWKCvBtMOSOJH
nbJ8LCFD3vzRugBb4pCpn9ylIDoJlBiD2khWL4YYhMNyW7bAfD4j6BvQrlYhGqZ85FIn4ZVVsUDT
ec+w/+NdnsLlPgSIfrROrnSID5+fUgbIIUfY8IaB3SAClOb+aO63YFuWE7ZUuf46xspEzrwjoJaY
o1WLrf2Llszq8ZzWe8VCRpfHVWeElw5GsaBf9DZhEgCiRLbuUPBJh6rCkezpj5YKGbDe+eDuM1PT
9g7MTUJjwLzMc9+SwgMtPfEau0frqdFOV5yCmooU53a+nz1RSppA4ERD8FlzNyJztiSX/8tWE+/g
/H7hT1U2jbjiH5Yd+cmpX0HOHcoyLgC1GlslIw/8a2uhTJzucCMVvKQbcZKzGO9u0QMimOIotK8V
iRydfvt3iSYx/fWb9pbq1VylsFpGKQgZSoYeu7Xg37KeIRwiLgyoJEM6r6gDXBlPqqQwL6CtVxkr
XPdveP55Gts3YhdBA0Jv0jXOCkD5/3QtsupKooDo+hz3SvhQDpCSOPmkiGgfKO1wASrwFT4hx22m
CjX3AMbqimwE7s4Z50Ta5D8QtbEvhxz/+/Ji7JzqE+SxzLDEkVNFjodOXUxYyY02bWY9GtLe2Ij1
19e6UwaT9/c48El6DrGjomUmtRb4vWGfA+ix6cyBRNRdXpm28xEvVvYh0i3RkZ//82BReWWuW/q3
CQp08Yx/5WzRWqXjHHWvVFBvbeENl5wKRAvfFg10hGhHS20WXPDK2t/oGDMa4LQDJ2uXSvLW7t2b
rplzjsEAiyHeF5ygowh/zzOnJkfgkE8C9VZxTMHQNRf3Spiyy37WmTnmamixI24/4yFceazy0Una
oGuLQ1uRxqXjaq0tQSSkNWCbfH/vxYNnMeGEb+MXCFUPCVkH43XyOBuGqBORWNhUv99MZPbFGT+S
0UFd/lwvqExEdI0FXLnh/33+6G/Ss/2W5KgojjjbB7RAII9BGahuXoJ3i8pp0duksatVyd9dcHmm
vHpF2RjAhCuYCfnmW/3MZjTbvIStIjB2fFsje7z8r3o5ETY4YidBUOiEL7+g/On5Iz9gUq7aIzpc
DS4nqUea1Y80rp13faRT5G1tHNoa0tDufYDauxHqa7kjV4OyVlwiWXqoBLqL6dHdmWPqvmpwVOEA
CY4PJKD8ATtH9NlAhyFxxQ7tRsh7s8B+T9HH0MrV9GJRf2a8agn9s/dIHtuWpuLfTrKR6zEuSkMw
Wi1qPwzrQooFlrMvkcOUqBnBjZMwNI72BabA1OybC/iw4pqSFiO+mvq0XgxdYLxbkzQgBEsOqS3O
UOrjsEqbwj7L81Q7i9JoG2qx3rxLdc2pR/RKbNH1IEf+DHyIhKqJcSbUiDBWEDj8QyIM0XWJBJQ9
yPPL3wc3Yz7xAoVejc4FUW0xLzlu6Aywe9WutI/09VeBfk/wy9yGcVz8s5zZ+pXQXFgL0CyN7bQt
4RU83pBJjXjaKQPPDHyBhVd+ONEEoIaOr2ExMKHf3vo+eJ+ToS357Iv/USsLFpLnTjWOpRZ2gNIu
k9ILtw8BsF8aiinS8j6lrPNj9hM1I8n2CKnfNpvhseJlHzYi9G3dZxD+GUv21XzfI69oeOVrQhPi
42N3z48aJWnRYIckDQT8nocX2huJ0Ohi4vF+O1uiZuL1NHOIGwMrvNqj4KiCQMeroQ393GwWCaVN
Kcd6AZOd6EVuzM+Sl6sW0s0G8dtt5vfGJlf4PxGkasogmnwdHN4sH8XDFKKemXAU7zfqY73HEjHk
clxkbv3G/RpVJvq12kmw8vLLSfMKJDFW10G3jmeDW/KAloO8PkQMyYrdvHCjzwtl2NIrnitt3zSw
TMU9VSeGJGzXakr9QQeCdqpKG/Zm1U1tc0Kdebwh8FiXDHnRrUZH84sFkBUbguKCczSd3hVwT1PW
QZuGHEjB1DAY0tNKUV5r8M88feGRkmXaZFWx56P1+pOfu27EaObpLAAMEOlgF9/Yie6sqmhfiLuZ
6veL928RT034g6an1wUuhCr4/HcUbbdhm7ea08fPe1kP7rA4ElNdRZ3nkCzE9+XR391byYkh/AQI
D0swQ2Tf3jKla1Yqaths03zF3DvX2o5bkkO0cGcO6cyN9WxOBLNYF06sO8DU5OOUW1bDLawSID54
xle2vX5HlnYB35KXIaxgGja7E1G7w3DLfZEaKt3qrdnq4jrPUn0OjGCeEnUWBStBL05WNwEjjCTY
DXuAX1/vJVbt2p9m3hgX/xerL/X8UaMBCocc1AiGOtPoHeafoDICZLuqSpyTD6/oS7E65gA9hUcA
desIoZn2YLdsS4ZdPbkJjc3C3yguyHwyJoxiC5AVCfTvTFHCjUeo3AVFO3Ts52XnJh1rAUg7hvG4
TFAvH8jWUepD1fePWnwxJp9Sw9wW8oxWWvvd4oqUnUGK6dtxqwp40v0drIIeHu7BKwdk+iapgh8y
hq77TWag3jUrAIZDrdy8UBzgPxmbGXg/4kUNupxW3QTSR/tDtxHIfJgLU5b5Ges+6u9gN7tbN+RU
bzLBxXidnMZRkPSmat6RcjodE22zZe6//0YDHcp/hdf/BeSNqYvsRi6YyM6/WF/i3rvyPVZgjxfL
U13rbHMRF+5BUjo56Y/2OsuxJqjNmvIDe3tip+4XlGMA36HqFYTf6BcNzghatVJ/RQyrHs3Q1Br5
ZLTDwiPlIasdAAyCadx6NEuof2aOgft/w7/SSYxdwxW+Oyx/mXygMrmOMzeKG8++hFEfC/jdg4h3
iek/yEZRwatGkxk3rxafmijZmyJ4FfpJPDQlZkJTxbkzltdZJJBfgPChv9AinPxGQJKTcy7UhaiW
kUqLcmlzvysBHVlFhmbwPjV7XGvPCBuEfguBTle6TMNxquUECw6+govZIa4g2YckVW/cn3EW8D9t
wxCXpm8EbIiAj+XNl/XcsLhvVx0zXIbqt6Tyd2upOGJvfNB3/53L7TOASk1jGLNZfN7yRWG2F7cH
OP6l+kipZ5GCaWxcvGYXLKQhZlJ41Ru/uOc9dnPQnm4866JlFUYQ+PVyyRf4e7WuCU4w5uZBtv4a
LJEDjuFlqiCRugeI/TZpulCuZPu95xy288rrz6H9i0rjQDpt0jtJ0O1Spd4a/Zqf0ZfbMCMh7iKc
dcGXxZP42Igmr9Q4FtXkJOLj9N/uJjR7F0BRv9fc3V9Hpgte7hYK6qfMDoM7A5+wVf7Mpgvb1Tzd
OLf+YdDcG3UzjN1ekfSZ+ZRNysKLU8jmyZNBVTEjN9ZEjRuG60fewikN2w2L+yben8aaupF1mFXK
uwCu07XouOoLa4MnIRv1ZHSOsQBfbYQIhGLiBXpputMST1tITZyMVn6242d3On38N+MGqEMEBSS0
krs6FupFgGaCfgx0aOzqBVehUsbMpq77QVGPn1tvRgfvFWzHKm0LfXYcfbAqCX0EkV7kPv/LIZ3E
1yr9OqPQ2ULfU2J4U3I3773fH2zn51e+XRIw/LXqnllW1zWkqlE+EP6J2imlYOP3KhIHUWJpLygu
U24aD46T9utz2nyU+r+5Uzy334Z4C7MkE3eaSjemS+CphkxP6Dt3R99BGiiaHubYRKrJ2M1iraiF
W1XNHxd4CFMBIdof7nARIjfLDgrCzK12sfzwzMebJ3waYUqsNBP+QdIZ8+zGcCpDS8Re0j3q529c
BUVz5VWWq2zrzRZR6PXMIScHHRr6Zr2WWOQCAne5DIJwhrPKHyl6qBWoTxtwp09OZKzFj7kzpM9U
9IBu45VbOMoOLZjvwUmTXoD3WKu7Y+JUzUi7UpmCpGzy5Tzb2DM/degNwO8Q6eDy+2JTRnB42cdr
dSRGtvKwA3xudtuzEZdkBjFp+s+5t5y77pgZtlTJS1xWJAop3/mu5ruHUsmSsbpjbf/hEKbBNk3e
OZFtmQEiRbGYM/kFfKFv4WQlZRPwu6SpXYlYfQig0O9Bxztjapo8ZUhlPX99otpSknjR4dR9GmRi
8T/NzbpcajdMd8G5VokQHgpMEdnC4DwPzRMpLbhWN0jT8W06Vpp9K5LpW70a+QV4flsWEvqVq5eA
1wIM/nKBa+oOkq/U1ynKt63rOeTSHoVber3ziCY13MSBaPEb8G1V81YL4qVAsWV68KCmasSLNzEF
z76hiOHIwciBndzTixsnc9Ql4dlgoBF97OSeFXAMgotsLD1aiTgJsRccZuC/G02sDuYj6bCXH/Nk
NYa5VMhBOd4aOIuy/dw+ngicys/qhVBpIyuCpXS8RZEf3RtTur6mmr5jm1bWi1UvVVx/gsWFZLGN
eZuPzv249wnv9825bN6JbW+nNn44QF897/vYR5Fo0q0WmTILITHQENjaKRyyUZTOezxjYMELFhkO
ktGUt59GMxjJLAI0tzqFxA6fEYTD9GMt1pdOnhDdb6oR008xaasyql0V91m+R9t5LtpTLUxBSSAv
nkwbAzIVQtZbfN/s3P/RDSzsTr8ZmDBZBlh/TydMZTGzGaYeSx359EehQ/b3h6D6erzuhe6q5JEp
t2DOIMBGAWofCBLVZVrp3IwZT6+kuvBtKetSSegw+eo+YRf5agYazemlQRXNd35lKFm/qq/cviXm
6ggeImY2PYSUjL36yAtCvJrjthp/POA6+8lLx7hSwMVba5ezGcd3Bmk0M9446jFw22AC5bS5UR6h
plO3UAbaMYL2yjwJKBQqxZdbO0gPDC5NGIuLc5+GHdisPi2d0umixEthjanpIbtFEs+UZkmMCiQ+
5MX1GRioTbJLgvL7D8iHL3EZYffQdrvHkmmqQjl39U7jK4s0XI5y82LuiCrdVjay8mP1X66G/7Fa
tu9zg1QvdtkWwgdj/aoQuZLA4hKn9SnmUYSMqHxtbFkG4sSlM78QrHwQSec1r5aO/lvoU8FyfnUG
DhWbCIiZ0NoG1+EZCt/kAJ4rV8VGAwmvPyx21Y8d/Fv1yRy5MKj/EpErn9jCxyYYVAMxssqDpTAe
w9rP/jbNW0QvEyLeTgszd/cfS0hILMzPaak2IbrL9ju2JMInk4uuw/LZcRZuZ8oRSCjYylnpYVKh
JKqRUhAmw0ItNDAK1MTu1O4rVRJxlFhG1QAjcGzZaM2z5kcZ2i4BZd/WrANjcagcJDCtqGCeWMwJ
1kw8xK6tPC/hm8Czwjc3SCgMFw4sgt60Qqw0HE96UjrfMwsRCz9QBB5puul6sRxo6T6yR4o7D3w0
dyNFgBmxaT1qw95xRjF/oTU71ZdSITwQb2wzN7AMu9o/1x/YaRvzwtIFs40QI1sKB8Wn88py5Q/p
WG6iVPwYqpr96p0Sz4B7AvZ6660sXszJvnRKNzOGHDRP17p0WmFaWuCftUmXAcURFebrmp1NnD0W
MY7TImgmvZHVbqW9fyz8HL0ah/8qVnaF4xFkkqBLCbW/DMpqysiGtiXXOAHxpqkHanoNOKyyHrsg
sakCgrBds6SgNzbub+9jiAPwwKKM2fa8eWrvNELVgGI+LuXYwBwz7R1jNzF6kgB5LzUaTV8w1XAL
bUPIjUJhpnlzClA+4zuPDc0+kGTpL33BeBCCWA4ox+F5Kon3Fu0qjZxq6Q/MlsM9e6Lc1PnLoPgX
lUesxafBWLPbqirJHBEJSKwmyq4tUfiAac4fegunjm7ZW3NwZXc6W4aot25cSgMvye51UsYSvpkF
81TB53ka6K5CuZxhQonSE6XsEPOdGvSWuq7Fs7ZcdLgxqTjKSY3vKETdJu+NI6C6z2qHLc7KZUOr
Q/ieB/KJXBJHWhbndMwH7as9SzgRYwwJC89GvbQV6nyWmlEoSaqObCe4ewqfZt3WEMfILFPd0wiH
AfKaqpmezUvXKlflgdxzeYLToyZXT3CDz4wY91Vf0LhGbRk8Gtd0Z0528UsN3yhEByWzIV/ZvG2/
zgX9kPNDzCn/aF1MyF+h56VN/qcZhK9DqA/m+vdAezGJ9YT2w6N1MiIyW19EgnIE2CPLIX9xXKFy
m3UHduuxihAIltf7zkwLXZFSNNirMO/A/L3HI5xdTlC3p8Bc1rnwlm1Bcp25QubbZmWnQz6Kvw4Y
5DZycehrW6HOFEn72Q/Wa4/A/ZHYuGUnDPispAINPSpcMkyHaM5IOdEgPRaBOH/G64jyrQbfRgaq
Fa062SLgNMm6D5uxQopwrcfjT7VGZK0Lrq6W7NEeLOZGNNPckOrXTCGZ/KMDIpn9DU6oP5g65tLU
pvOk/ChFXSzvpDZx3XlnWKP+39jqlAwZTPcTAE2J1c/swOgtkBUmN4JkM6xDvcBRgc7l2IpneN41
JPQ/lpYA/Y6Gml6orDSqLgNZWh+nio1FoMSV1fDihdLf1c/tqmNaE1iD0i4OR2bteQA1w9jWNbwb
VF4ZXesNdLmJu47MGIYmFsx7kWcZBQxKfva8UK6fy/yjmetC8QYBv9mrO5NRuS2CjPQJhUha2ac6
b95PcagxiU6wSA1oi/uFNKTOrjfyDQC1dC4Kcd4c88xddNxIKKnOATiewPMK0nVP0pBLSWZlfhvF
giGRyuUNI4tWttTkPsIBPLVzDR07M9X1ZT73v7A+zwF54dB8K51qgerzlrTXV0G5qN4qHFFlc42o
UfU4rgnhiZYZbeXraExX3v4JkJJa18G7cgaHcPlNYfdr4XJOMOlTocUM0LZ3cy0r+NZPowXcEEWD
6UO1bjaxNvgITq7LJUeGgec30fTH69gAZ5TMm5a/LTpAFSJO88Z9uc05ydYEd1XTD12eRrYA1NbT
KlQdPM4vrhDqFqpP0uXYIucFMFKrCK6J/Q22QXu5pnkIsOM5iCFTtQD2/Xf3g378wk3F2hgmyHVg
swLUe3Hv0cSSC6FO0VMLX5CebVJ8eiIIEKZ8ldtnxbV5ve0dJLpoz/BXvTk/eLI6j8hJscBdt+nV
Q8MX56BQEzREP/J3w2r2v9hPkMhqi/tkMLJowZjtyw6fbQWnUCPPD/+HI91vv6Fes189LNjj4H3Y
iPJSodCLAAYpeSP4E52WL17wVhBr7r1HXSDLfyYBwJ99wf4izYrlTXjHQzitY0QHhH12yEXiNZeM
JnDSDdp2FRABsYrnZc4UDfqfubyy+2QNC5kfSr2ZqUZ3/S56LUKrts9tK28C+tVp0NJ2elXqE8yC
xB8xpAr6cavoU8WhInx1nvJR31G2bpk7gj+kZOiulsxfFi4CoCuAajNvl5kdL4ZBpKAcECLSbB48
sxNiFgv9UoCvgdvVPdqwTRuAQRdNZOO8f75HirlJXRBXEcj9zJ+SPxchHZd+Kt7pUNtIGSWhkRZh
bWqT7HMBFM4D9k5khwN559yXSYwO4wAHkbHqe+XrXJRguqfQEHaMttG7PmgE5ZuDcCMF6plGPytC
/469HbQ0JDxb/GSlj/Qc0aD0iQVNcb5n25srdhwzMcl+zYh6EmfJ7AyYARkwT72uTy1eRRubJCU6
2n+DImHnfp4i0wHc159nTv+xR1lIBmbv/HSMJNbXovKW67TjCSz9PclSyjjMkpQiYpxEC97fPjyy
u4NSyiuk1ePIMqV7WBhGrbw7OxmHBBb4YKWSBEun5KVQ4wtyFyDf5/NDjJ/ZZ478Vd4YeU+aYSr4
SxeID199TMOLpt8Ve6G25hPk5IQTmx86wDhjwQPM7ka3cy7xchHISJGumsX9bQnngk1hWtGu5Trs
MR1O8VFqe0785WqDkL6MP4Rybxz8ZSm7sc9M6prLkPKD1aPBqQaO4Kem6sVPckHi//ASBvIieJ+B
GddwAP9hUZhEMZcdvW7oGqPA/pm01YhP0zQpxAA9fcVON8VLGrmHRj7qI6aIZJRgqEGyu8q1gLt4
ys7YykqxXzrKCzoAKfx1ampDN1WebftMfwBIJpJjzD34ESbcVA1xk5oDBYxOcQreB5wH0vLPwLfC
jLaLh/vFr7Q2F9uHosE5PFVbkrqSDZDO9IR3NuTy1GLbqqH/T2+Fv5u0do6522Dy08TtEi9daBEk
pfAZxJBrKMGGCM0KFHBjNgs/5hZxszLlKIvuw8l8ZF5vwao+PIpHWatMpIVN2Un8okBZdmIJwo3k
Ew5Gqgz92L+OVafZgi5ylIGVR9hS7x113PMyiwz0q/AbR/5+ZTWueFg7WRWW9f3O/7JK0RhbwJBH
DaDett7jmw1mu/wJEtONCK2m2OKZzN/90g86vATY+eHBv/QfSoAh7ckvy/+4VNuqPrgTtTt/VPSE
BW4Ina6tlva3AbSivVnZlCsaYQDhOC0pKU7rWfoFWIB7ggNMg+0eBxW8EgI3O5YhIOz6P5StZ84i
VUuBAHEFSm53VhLwrjF9miiXsqfqyqtkwW18LyyJF/h+Y2KBaugytgsjuY0kPo66wsl704mW0FTy
ZY5fpbrTdOAFTAxZgnNN7heaJTm5nf/wcaaJdiHHCkMiNgyrcI40oHqgjJfxMfLblX6H0lJv9QUr
/f+TR8wpVWVpErTOIDgvNgEDDNxSS+hYQLxFtQPg4evxv1/fnYuwOuti7GgfrBu4hUWxc4uOwO9n
j3qjE72EAg5Ov46T2+/UMVHsx3ejqX08gKVpOWV2r0cq9Hqh/TfXKs5N5wTpHBagUwlnGXYfbnfC
//cSeVJVjridSp0S1rXC36zlIhSRrk0TAPlv+VUxxgTqT+YcsRggBqv29dHYFarhdvzEWLD5l+vb
u6RMVGrTOjmkfaoFOR6sfpyz0lgPXb2xEW2Ufk/bTXAFFIHJCcXl91068TvLF6GYZOtlMdClGB1W
QO9lr38r94pnynmBgape1wePkpoQjNJ0DZ/1/LbSFFW9CHWqBDcQqkxBP3qvvVXm6WMftN/PK1OF
rEIvJi89HbIBX5Bl9nOTDn6ZB5+9aDde0Y8a5KbSNg0EbnbCxpi9JyE7iCRT9A4HAV0yPMVR3c1C
LctBm89eprN/XeitoPoMVtwf7AAh4/JeQBquPL6MiZzAATuMAyttpNyJ9B3Dz7ZbwPJtW1nE7bSk
0fPDvoWlbQVgW9s5zb5aTVCTYuWnrGK9MBktg9+jaiAnYMbFm3sXzZf+HtKhULq8sXvPm7bV7orc
aX1IsGe93Wk1gRr9khgcxTO1PzEWlCK9sRxGUxCpMLUhaUgc33QA7wgBBUrR/+IC6A4hKWc1HLX/
lp3G1gLyPhJ1YkiUHsshWUxhSlttXtAD9jzFmFymqu3/j9G4IdaT1L9F3/2cZ5zOB/lBdSnPTIDE
YO/t3V0OmitpHCCzCGhtr8Q5n2qqqF4UNuZynErJ3hzvNU/QTS8FPH/lhc67dlwqatkFbZ/VmIPX
FJDikYZh7Dq7usp1suE9HLUjs8PHZKJ7a7L0cOEOEkTzxlRedXfyUCj8AyF0L85mR9ecNDeckzC4
nbN+VvamaXCz4sBolKbY8T07nxleopATRLJE12RiuuBeTAsWLp77hKzVtpfSQL73w7vGWD9Xgxgh
mAya4Oxz/6h7v6zEGziXquRNl2KP/SU8ntZCaiRxsK+sP8Ty54F1wu+s+ChAvecCg8gmYayolUNW
1QlE+1hTB9uYx8MPhxOlnzJmjXBkFQIKP1Y5Q1tP0M3uuvK/vd5nWhAxkEsMOjX/XAPq+xhiaLUf
FYj2B/kUM6rwDRmJWnilWednzzwYkCBl//T7094QYmtel4cAKs0j6KUVcQNtx929NLdKWFLkATG2
RVTwiVgX1hSAIzuyC/MS8MSPbDIF1EmM8m+zKWYm1adX1txbpgYtiQP4rR1qMjkiUHFMQjuUgLlS
vA0gyVYol3A+UJcjZxyqNxxsgkFXD0UrEnp4quvBeNQ28fZERISMdxEOfu4ZkSMysT5m2KX01OCY
ufX1/1daOVXj5LJovgfW/3rZPEdYJmon4fyk1N1rLKQhT6qZ2A3dqV0SDUfitaap5BepcSztwy50
7l0lSCTY4PwipsCILjc8N1ERxCekHW3jKCNpBa+QrMF6e+r41cn0ySGzW6J0gMkQja/OnRBfE+VJ
drZZatidV33OBO8aa4pDa/xxVHN/6LvE8h/HQXEstUP4FB/ptIdpn1tNmzU0+/uX3ZvIE+TWymka
sHf1ce8csqOkLt+KpFbn9NKBrU+lr/9/joESwk0vGeJTqipBvuIsl48oiO8lLUYSUWzcBPUmtBKl
UgDnEPH6UWUSKQhyh9glNtflKYh2jeUi4BX7Typ3wozptq5KbuT7EY4DSbpya+GrK8c9AuKBjzGl
Mih4/8rE+9twLob7NH9udZBOHnWNgz33LEmcnPHtzr78gVXrklX+6oDHxT/EFOEKP0916uFu0t98
b9nE4dYY1qpf9LkHHqDaF7cBZjbh9utGQe20WpAhvzAOQl6ySvXxHYIN/7f/LIPQfUM//5JS4SVY
JCtJQ34lri12sW5EgIXr1iTY4r5+0akawb+G26JJxf5I1kcl+aioVRf9WBF1xTbfvKbo6keoz3vw
g2ndZw/tTYn8/2/3TUGqziRr3PWA+Yv4mH6kEkpxf8F4TlKxF5P3my1nTIh5MkHhC4D1hsAG6/Mg
tJu123OWqoi1WlOZXbeCW1RV9T/Tr2TQ6I/ZTrC3ciNdE2fUl/hL6UwERbx+KnQlMDYKE+NbwYbo
NMFTgcM/w/N7GD8qg4h+imYccgDaD/iTPGR0GP21gy1F98QYE33/88Orq1ZlSp+mSiMin6Y3fUDB
/lb+v3qvPcvnlpK4V7vvqhjH28AXIYaRQZEo78vZBAIHxgesltwLxvqyIHrBGY9Btgj+G+XNbLSM
KqWGFWWzH79FNEkMaY2yOoOZtrFGy8ndNxTWQmAupZALU8vJmzfzHsrlX8bpK8PAuRwSaBoZa6Ps
ECNjTm86Rvp6bQ5RKmui16Y2YtrwYLnMQPZfaVfyX9qRFOkQNcEOzJfH7C5FGl1k2yVzfeUfcq0T
sea0nOjGNGU0KqdeUfjm8qzngqPm6CxD8dKPdX30xlhWQHVhUU26ftWXpnm9BDmIapl5QMqFkIn2
hwL0oSkoSSCduGfAlmfzQ2/aONrNxJOYQG0QH4kh/xOWLIZilutVjt3O1e6mdrRkai6htNVfE1DL
ylGGLuLshOCwAH4qplUUOcvU3UgibIwucKLhvx50gLqKxvAvlZzJ37YALsqZ3UPf8Y8WSu9AjI4m
iGEHgqaLU7DcAplO4mn3q/hr+dozq00psf+tPSYhQvkLMHjNQpV8JChnLfMCwyD7/+jwWeU69XqI
gv9WY6J5r36/m70xBMECPqJWAovSZwKq0K/NFqPkizWnF6Xos3pu2xA3nv3wk+cqWNZVitB/TF/j
aXs4S/6ClycZn+VbMC3+Xk62E7NqmZ3zFTexj69fOI29OQAHpgpV9+z0J25YPNkgubfmYqRFN39z
Lj0FlffHzHYH3JJ782SdqNGVMJysQAlecmmfk77EuEfv6wzuN9W4PAlJhNUHl3J8pAZTxKJrxkdl
RWyjgOx2ONpyKP6exR5BgmKRS9qDpgf3xg3cNi97jDySUShA+SRXqdIyV3IQ7ucxrzrUXS8jOFy3
TUq2WOEmzzPKdic9OnaTIPK0XhuJDIlfVNY15g6gLW07VggVxd+tRvMgLJzXNQIdMVfdEyXBgISV
daMriOoVfPXAHxWKjs9u3I27WnlJWBpSh0QgzzDSmwOvupkSAE5dHoz+5j2acbSABiBp47j8g4Q4
A02Zy5be/JRBC+uyM2h4HxCtyCVKDWdUUSMxES2yY3Lnjbr8f52smRQdC61jr3bfz1cVdnlaHe+a
u2mDrIE6F0bavVCI44D3kgY0b8VunnoZE1O4QvxSbyZksFL3WhRaeazqeY4ou+qDKV8/mFPSQf01
hB29XavNir0mXdSdBFojZRzUqKvEez9BGgGe0EP3K5getZmaHPd95bn1k6WbrtrnEzSuCwULlaM5
GqhmU+9fOg4Ocvea1hsK7lAZ1i9P9t3O8jprBNg9+VyDoWCEaKv4uBjWb7ZhZd0OZWjyO7qfROVh
qlDih/DbVGuSpFdDtJyxGpHYqTeJ10CA31bUpIRBzP2wKVARI0TQ58S0fpNuCO7mVw2CN3ZwG7gg
Z395zf4RClZJsOXhuOkzo2yaNm6j7Eb2hq8K4/ENYoQ16c9PBL2IlDTNYOloSbu+ILDJXr0/83la
e2wUQ//aoR7zpVecBpOMDvBLK9XHvQybPXivGowHLVyXhOpAV3xjBVa2wovvJt4SxvjJK4VsDxw3
Inx5qAW9WTOOOqvBZf+EgFUJHU18sYSwBhz5za/YcxDjFiAdBzs7nqmOizBO69uSijQGV9VO8xEr
QKl88JwlqqaD4MX4BhkAY9eRJjJmbEQCMTeev9ofairCPVxD86Vk3pUPa8ABBQjkpMKjEbLDodDA
Ekg4s1/yymI8xZUQIXd1YevO9bu1Awoy63bqA5IQEmplhXRRduw8PRa2/zebj62uEay3EWX1n90b
sJWZyncTlIe2SRQOcGDbDKu/IDvot2+ngQzC7XZiA/XsxIAd1+JlrV5kkVp4Qx79PTA2qA8XdWqt
YMsHGEZbyB2yCVOtyrJ86PU4gWLuLWwrQlclrKbIUsW81zsvJiOWg4PtwxeXj/NV6fR0g0bd7Q5h
/sGrkBIXWr086SUs7QMuF6YgorRAFM35x8lvmcjtPPHnwhU/WwW+VXc6qSe7+a9/GKVJi4Io50J0
0r/uGx/vFahRZaUdTorlx+N67Wjub54H/EKkBewqiIrh8VUtrIvh4BTNCTXcIknYOMcu3WsBA8PT
u5tYHRy9xOw6867Wj4ImEHsrdE1mRNvdmCLmyh793M9rSf7Vfrollid0b+oJHfjo0mp3QgFdCpob
xfkcSUsUHctgqqO6OkvAswjSgmgFk8VI8qUm6OA/o26uqbqhCniy7SD4xK10d/PSN6ZiUyuNBTE9
zZe+xj/lFVS9eqPHA1kHpY0KFTMYSFDVEruk+fTZ46e8x7qHUgu3vyrU1tWdxcCpKtg13+DKUxN5
dVtgBSILFBLE0/SUVSj7/8AFHtNwbpzki3cTZoFGEFGh5NSAr0kl4tJgkbNNaY4I2PQ10VPBbYlr
RkFQWD/XBSGgD1eyl8xoQjCEix2ZS+r7ttP2hQIYGonknB8jKmQ4fr48v74LMgA3TJ21jo34jSeH
sKcj8rGFR2yxuQYaifp5x+9YTBK+kFflEA0UCbfrgYGY5/zfhlPw7YPeFVSyuiRaiyS5lpMf5Ush
9j66ijwvhJwqorv0hQhY2B3AAiFO1+JQzEa80YYhL/JiSDpO+1DQ56wiO0v0eyiIbbotjMau/sRe
E71ueT6CcG9A+klk411ph1wbIP1ygna7AIYl/TWU+/l7grRpkT2WEyEDsU23axPK0m0g3o1gU4tu
qfmgm+bPMdqfC+rS1GjkGAc1CFn1YClBKslt5yvDzdqeKwRgd+hwywVXyXd8VxOjP7nAeq4vtM9M
IUAbnrOcNZqUpkachGFjUhC+SrVpMkOBcqqyZoUwssgElBaXxkM/VrlzSaB8BFFuFbCbYkjkPOxS
6ASQPs0tGr0QZQAk4s/dY17yCtWyZ3CUhLA1F0pAZcJ6OpJXnJB/X1Nx9tp7ZOwb2zcPl9Uf3o9w
COVZau0d9dXX8BpzZOWrjnjyBYrF7Gjt6/chpurSL8rvKZ6ZQOn7tylDL7YECs1yvmIEcIbkobPB
jq08HnvwI2JGZ0BZgJW4HqFriF8kb5aLOeBf5LOJrszic42pQSg1U5rF2rAhVM24ErN2shEgrQPY
tjI4lJjrnfBHCKNA6RSPawLMsmAq5cob4Jm5QdLpPHkomJ1r74Z9mNF9ZjA1dRHfDpkJcJA+kgnJ
MLfCIvuXl2QhPhGXJTYrZGG86pcBOuX2wqhAWnkQhq/uUhp3fOkpOxqzPo/g96UkkzyRRpLhfjDs
I3ybTk55Fp6slbnks99WdWgXk6NQPawAX0S53Kpz9aAreaeQnpNsPb/VEAdIvk2MSBtvIHWzMlQf
pAzOF1XH/oe4A10uqfqhNbeKdSOJ57Os1ub+DmuEPcAEhTIOIrDgp7l9l3ZSTnosXkLHHhyQl3gz
vNYAilJq8o0Ja2bY7TN43zJfv/qXPXDqX7bB7j6DB7XNuQs1VJbPMt7C8sxJ2t9LDXApwtL1WHXj
C2n6E+5fR2Jcg83iZBtAhKjukJ9kQvHa8w14kZwDKZkVWHTYvPpTBa3n9UDqjscPjY0yCWcgUsui
/9mu11C+agDgDtNzZq7+faoWwYQ632IHM835TDvUAwu1zRBU7K/Adn2AwkdPIVbMVs8l1kJwF3be
PLGDddBwePgaOvut9sPTGTEC4/FwCwSfQLNUUwG4zGUOTcTmF+Mjn1Xu46Pi6A80UIIECwgzZVzx
oD7LFUzZAAJJW9ibjOdGbcAvz7chnGpHdeKCoK7231DOQqs5GVywZv1G7TvfND2t7GDX1OY0E2DQ
QzxReHZfl/V5ag/mQdJE00IO2qNXm6Aj1UxgGOT8D6qIG4gZwTTeez4m2Chl1xgglXGfcBzw6pss
izYs7m0wcB3yeJuayme0ZaHZV5o/8J51TSGoU6eW2gKc37AECOls3zGtY84ZDhhi57xU1EMT9XCB
i95lj5fyP04SEJE5EiDYF1too2ypartsyHK2yH1WwNiFA3p8JbDAMUOvRU2faeiz/daikt+cOBmf
K+17Y9+a4EoJpr9/FvsLfGhUHw8rWH0FHOhSQQZ/zsmrNKnaZLFqjMT3kLHDlZGkTI/kGe28mz1y
avVaoSwfzBTn7g/iKhENWHm4UeyqJiC6HPWDcqjKjLzRebAdsTtIhdOKqFqr9wer+ikTf8X5JC2M
dYGWS4GM/9rBXk3TNIvNEuA+DXqZSGgckfmJCgruiTAtG5DmnKEMljbZKaH1cnMMW94UI2lbYsuZ
8csGnfRdT5TyGYQ5fvgR/y7ikdpKcTZt5Aq3FKNTokzyI8ublj/l8+s/vwVrqVys6a7D0nxmX1wN
Xv2p9RZDnhJnSQRuiEKchZEDRSUyR9U3FD6qSCEvDwqKL02pl9USH6w0ShlrLiv+cxxmzZGweaHc
NaHYaBiUS/iOl/5LA/znWKG6k+2wb3xvH/26kv25mPM/AHsVMFjRzYXoUIFCFFjtlP/IPxzrqZY6
+3ROh4/8Evu7YA4jHlmmIx72OmuzSuRNfn8c5XTJUiyI0O2ulzUJ4I8ZYa5WTCGX1i5ElOkS7AnY
FFGQVelO/PtnhrJP7BGFQv2d0zzN9b9N3IeaG33EPqEvOFF5sqPwrzI/TUPzEUc0iVFPRkMRxBxM
vIBOpdO6EodoSJc19bgfxr4K3tqc/HGcY078quoLcw8ntgdtM0pa95SH5JqqAhDDIrj88coskzLJ
kadle3ThKo9pz8OrFeRR93oj1n5Th4X3XxRUFJnaSOjHHXEXJCI4EAGfON4IOwEYynHlDEm4Xcbc
AqMmjYQBh4sJAi6Ts9Gl9+/ydqrrOO4oHvW6FrV8feSpVT8snTtYvDC1mUD4epyaqNLr4EsjlWQd
gxaq0FRR5yvzQG94pi/+d1Hfv1S1KMJZ5s18/LpMz76kLL5XHQdoQWusDTTwHogJg70NWptjUTWC
brl1h22Pl2HBtjJsZydwK93Wf/h18x13IkVdjCLyK4EdeP80CaFuJyJOnIz2HtrVGYuEdvMC53Ny
LOGLCetc9BixXHr5qD3PEW+GVinXx6X0BklT3vKN4V8KX5kCYMEkarzkoX+YwKtgKx0A17mH37PV
1QNmejbrmS3oYJFFjf4Gy3t2NbRshHzXWpoa3B5QkvZYqZ2TWDEmycWWuhYsRoAs+nAnQDKPfwFT
k+3TGd2EuxSfUCVWg4MOXkT5iEC4OAX5ToA6vCD1jtn9+3ThrbJeI5zAJLO/SStk+iX8mTQ1ZWoI
HEY3AFLA+L+FISPmjcUuz9Vk/IMBOUaC4CLI1eUsCwMuUqizf7Q+8aQoUeWSfwxPJvv21Xfuglbr
a4jNpVJgy9EtGTbs1e5LGHbGrWtdRoStUH+n1WCrVzDr3cleTcdz1w28pxqsqybcx4Cz9/6obeEc
n+osJ+pC0EoCU3yONx+3NiG+3khHDpQsuFpul3J8nuZoHDDRRquHdE4eK8uEckX9LNbTAGL6CQuI
98Ipic7jVYhTi4Q77zRqNjya1tJR0ZjLINmWum3uS49RUpw1AEmLB+4bD6VGGHRO7+tYPG0FE8ZY
nYHwtpEhF3yFhrtpvc5DJMeKpvO7CaAfkvzgDi+TQzv9uBRL4nzEantT66KoKtbaqrqNIo/lDmS9
GBCVZG4Mj8gST7ZSrhLuRTQ8xCyzSlHRDD0ZvQHdo2o0fr8Kx5yKAK/5PRAXrZMnQoDwKW1GN6o0
tCPXcmAvIjZtjt3sbtLvDHMPo4o2rcmO0rGjmdEZxOpspUoV/1T+uIoRcEp9tOvjtV/19zjJUhBa
Jb4U8N8GDLlrX5I+dMRkjZG5yZEK+VKUfu680ZX3ZYV0zkU8zqjrq3Zoln/fL0vYq7KNnswft/Du
wmtcNAQA+EVqvSYibsPRtOrq51U8kGtwyuNrOSehwEPFkFPuibSlc+rz6SJq/691AoL39mkEdnZG
kEg0SqE0pooat+9/pSrzuOSibryaH48iseVh/XXEadEXRbPsnv3u90H0nM+YIbpnQ4YgJYwvo6CJ
vCIYQy/fqm1mc1tHxOzk77qzgiKsU8ytrXTutJjnNt1Xv/TfP4/RXMuPLcFl53m75RBI3Xis+9yK
LHCd9WP7PJWbQZ0y5Y1QXFAigRiJAIEvVAntEanXrDJR6+yReQdRZalgKs/sOiXM2zAip6zzk1Vz
ICaVJSvGpnrV/Y8TB32ukTwkWrNh37DBLcESK4DXUr90AMLjCwJqPR2gEspmQ5pNZiqYhTNa8TM8
DLup28GfXBr1i1TSwRczhSS1QavF5YuFYcQSMy5RXr5ss+ciyT1Mi6gO7dbjULpBfhBkeRGIn65H
cuaynkFNF9/WguHZtl2ycZ/0u6yiru+XTZR5IunQ2U1+M1GSwUV8pEDZoGP7VLxhnd9a0gqGfRwi
YGD9cgwM3ySbETcNa28HtRIJYzHqL5BvSSZpETx50NwTl6oDN+BNzUYNtfAInePP5XeK+n2RjirB
j1EhrXhRA22LVHJ1WtX+yOxLc29m5Uxd55zq/ZzCUEJiVEeEBOtb/oZWNVpG/YMY4tXTrzT11E8R
yEtVveejmm+cVjgLnKUG2mtDVWEGhrEgw0/+vWjzL3u3JhEV99lHjAjOBR00a89frpNRn7qoQiXP
5CtQW5gMwBsRLCGxAy1X1RVnkIitd2vbBWFIg4HqMypb9lVRVF7ybyWLh9SP0mrd3jhlAHlAlLiG
UaMuydmyjJ1IZd9lD5c62noIAEOUKRNWh+XkIGa8h/NNGuHx/p3mN9P23/9LeSLo87cS2vchEnnn
V6uE8mb4yQsQknosl1qGYOz5PsIxtYx6UVT9ZDXwus6LKZEr3TVw/vLEMVrtPIPtObOQnlxN1jht
P0rHG2FzrXmW1SN7xG3/hwakXtFOJ8smwC+fIKPC3e6ncRIHtIynQIhreroCSOx7ec87QrtZJKwx
unHK2avG/bVgW4jKs2c9xzXjoy30c/ZXCzhB5T0+KqiPiOLVudFdcaFA89ROkmvnnlxphwco6gXT
S/YMhCGu9PucYT9wMnWZn2Ab+824QapACmglz5eArqnrPudoTeQFXFqQ+uLTk20btns4g7YRaDeq
ZuRFcpHYjcxqtscf0D1Xzb3BjMQALFAwn7pg3HJaWyQEPhZUeMZMUcwFzwaHjwFjDDKvK3LnF6Xn
t/NyCCDHYEFs2cUfsEfjKMZ52E/HvaB/W7NikgBTOKDL3d8/KIbUZDtOtOKB7JhaNX15+rJbHsU1
njSfcgiHcpbYWXwzyb2Xe2VLloArYGozkgI3uSkiZSmECJ0+cG/3/4qpXc45s55affYAgd21pta4
G0+St91TxhkneKPiJZCZkro3es7HoDEQiCpr6tDBTCJp8N+YpIS7i6DUhxtUFWcIsVJ9VZkUGaEJ
+Dw0yAEEeV0JZ3jqeGk+/bplubb1ZUIpQBficFWbGGEAwFqRFhwHLtuVCA21NzYjpA9aK/BwDpcu
ToEgLkTEY7qf1HcGCXwmxN95HCNrSl2F2O+lCIfyhxZh5/w6oScyozV/nPQ/v9CGDq0hOvjWXq41
hW3fFlNJ4aEkJ1qQA+LojKcPYPpB/kZL+F1eBLRT3wH1JUX1uYm5g1OlB/g3mSX3X0DzWXGcdEJw
ijeZhmkIVnhBF0jVTQ6BUrFSXPRlTFdWyU8OdlCm7I4AXj5ptA96PCExbe6K/fU7TUNkCfFdquIS
RnT1LIXIWhC3cqiiWzKkE00hbmq98uh0uNHlGx5lwjIdBo3OzRlO0MJCRlU2FrYzdilgsbYXToIK
U5+dZHwbuNbK433eqEM4rglKAeptOhtZkqsM1oZ7FrKUvwTaPy9PsRsG+tH5ugnZTtpCvIUcJY+m
1j+phKDYWQbfyR9hAGus4Ez7xId7H8gXm+rkeGAunAlil9n+q4ydLn+jPm3yoWf2LqDyfXNGywMo
j/rqQNRTTh36vxcfP6vnRqvMjlUshdQFIw72E5qPJla8pxn9xnIDiKa0P7WmIVeUgnlSfNxYOgF7
O/IPaTFG9ycxGzoiT0FuV7hXfz9x5HqECmTdxVKJcfcPrdR4DAmGKvmjnMsLmalQOSXEb0x+iP2g
difs8JFyOKX/IdPWbLMBu+fGOIvDY8VUD3mHwV4R0nKvCZuKdRGxtS9UUb1oYQ6g0UIUi4LZbyQE
e3qOwmZCk+Ce6E2UXKfC+mKHPwTgowOllYUOf7CWznAI2eBKFnhBxXOdC8/jL+P5DqKcq2cDvU97
JimV4fCpEjIospwgKSY7nATEnIf9g/tG4Y8+bAHroRqug7Da3BZsvNN4fJb3Ddk87utpA/ADD3Mw
4KGX3a5ah1jCYRxg21kCRmmbZZqH5Q1RKnCZkvzU/7K7kVOCv/VR9LfS4t1TB1s9//wdmKotaX40
F2j+gWgobtMHrkvlB/j3q+riR+ZAmY7iWNtcoWJNwh58WvMwMvXmIyvpC+qJ1iN9cBJOk0cwvHwy
ExqX0YeKhebLkoAqWusJWxhmrBLpGZ4mpQBo5jsT38GRtPCqBK9sqylgbDFjkamE8hi7KfxdjOxl
pQ4GPhmOdqPe0T0eCXArKKMLaQQRVJ4eSgGYQEQxaqmSYzt3OPBu50/En6wWDjmCtbzYvFA2v1lZ
V1f8VUHqnMyQEx/vyGWpkhqucRvVljVqaAiHXnwkviEcuRqYmYDHFKksX8YpxeBzmPcwQkYIrbvc
sfNQy+EM179SKpaEwK0ldiuRpV4CEA1buTxwupa03O40wFCSvW2HNqooF9A7zPezvNtlS89lATpF
CZDxwg2xvK11AEdImKhHoeNm9UFxlJVZ12uaqHECGOfgXYMy9ufWwIaKpedBEhPvxlwc8uSCVM12
1S/y6HDYbOL7ahEyyhtVrQL1775vVgOUbRW6amCK8VKAaTBAmAU2TIlTqH4pzfhRg16Amz7TVpbn
28xu1vGLk8wXXbDww7/kHZpix6bwEiMT1Tnj9vIYYXZK1PRqXp+60WRBtSi074yydVOPfyqp2aLF
lcVyi6Ajg+q2PdvqmZxKaHwpoBwJkjvzPlmEO87de5W6sN7D3MobcZjqDdHD3mCf8yEUzWYgYJot
gP7h8evzBO4ddbsrHGqoNQpyQdtJ60BqmakkPYMe7VHpXF3LQnv+wCy6FhWkrkrWSVgmw356TYfK
307bym1N2fgfqL0v8ScToQNEy8ogjBxlOlKOO3gluctpGqOvcP1178JU5YIyTMKaZ7/vVNDBrStX
/OSkrlFjUk8ZEpRenTLjHZpKhyjwL3/hyvQEzOzaHHtMK+A3b6U9NRL7nrNjfNTCu9ypYJu69sAH
vcFexXEIRmUGHhVglnQxq5ClJ8Zn+Ll9DPbZnH4Xq1O7Xu1QxOEBQGFvI2aR5GNfzkd9Wx7tsKch
Xi6579WZVk1XLxC1DJF8LkDynurlsGPW2ku/cSUhhY85q9axbcseeWd3kktuavu6IF+EtKisxQZ8
DFEh3h8zTFtczQjRvYWAEX8TmLTfcruQrbz9Mojuz9ulURd4EuR3D5mVE5Q9+lMh0K2za/UA285Q
R7fkIJqZVGsViQ0Puhg6EpQ4ASeY6OUHbNNljqFJEOFFZ8C3JW2XqwMlikAL/uEI1MneSZEA/uRo
ob5LNqgpBJc0fXmluJWBqDDCdjRbkiNHashYyXz/HwkHUBFDedyDvEJ9kP+Opu/g+b8bdJq/jGJq
wKtEoKzRqqZA+LCcP9BvT+rNIcAOb0csK4h6PQE1EUXhhMx/sr7bpx9xdvEZpEQiRi7IrH6jjjGs
dJM0jIMRyNai+/MLszewZfI0GYG5onDDgVJ5Gjnfc1eOilu2qkDe9o3D4d9hIBDfT3o3UI9rXG6T
8izPbwNX5YGUNsOiP4Kw88JOw8k1nr3RmoUDs7mCzt8iUyPw8C/VZX+RPm0iLkCIRkzCUQsNxZll
UlL/g0gkfLnY8UPYH9mhJBKv647H1eGvQu8jum+JeHgGm7oXp1kGoW01ZvkWd1zG/fiv1JH8hnq+
QduZPpEVYge6u2lUBMm+3C2d3co7G2yYJBq+xm8q4H8HLRm2QsNsuEGNFXBJSeB/Pqwbed0OUzV3
33mIX4bPIxd7NpAjDOwvlVuda7NUxNapVdWseih7zSJpEUgnfl5Fa7BG0EhLjuqv21AY6fJZSCL/
fFmycDT8G6h3HgNClTUygdL6pK89reWTuJtODxCG/a+EDnpSzre45wn+ztl3VPEJd1aJPiB25lSx
v4HbPhbeQtiQbOsiULB0Pm4I2eC7sHPDEjNWV3qkAl/EnkmlM3bqGT3hgHppwkKkfoh/TPrjWDzg
9y+sYOyDvxAmyhCLAcH1NSDptONmKFwIU8wD4oeEPtZK0ahTaI4eZfzjcu5y5wb7v4R09raXTTi/
YSEaug0srKQTaNeMoo1XM+tWKntbn0CZjgt77aWdEN6TDcnJFeA26MLkwT1lJrJN/sgiupc/3oiE
S+dxuEvhfxodksAlzUo7T/SSxhNGYu74IEyHhYPmNNhXWXhgCan9J11jRww8Sx1ehz5LJegOxQ5f
y8rr6EdbA1mtdk2MCfXjdnFMTYq+2Hg5ogBuZCcjcMeASTcXkcY1lfyyuYPS1iyOzPAYMHoz08GL
AinF9FR3CBA+gOXaHxA8cDJrvZlc+XcCmmrjhBCToDuT1WZveOQHvkALhY+2uMZqCE2CoipqOOl8
uRwPNv400RmCBOdObC0mh2Rz0LwaJNstIycn467FuQ9y50CNC8udQpBNLT6kpFHDtJp+cPhBFcLY
bnA3KHEjm7WZZ4CcGIp3L7Y0Y9a9FQgClA9KZ71uWEYNHs6JEaQLUQ/p7hkJOAwM7zDupCzgd9xW
CTeCcXn13lOIdY6Vb2vJYXpe1pUSsGb8bZffMBHTKoHzDVEqsWWSajM9XHCzaidujfqtiI6polWQ
bBMDsIjq88i12gLpBMX8lp5Y7g3/lq/5jH1WF534w5Wck6X9BUJh8oiZ8dup7Q3in+abJfX6XZij
fi99kopFYKWAOtROfqq0E0hoWoPGCEB0fahbFec8Z1fJ+ivKn7MyusEMo2vO5QES94CBbNf4EB0+
peo51FQh7SxkS3C4woKc9X/I8zbure6Mpq01cVZCarxmtJMyTmMtRSq/lXWapPBPv+/M0nhpJIFm
pXIUmbIvXSJmBojjW/K6f4O2rnk8gfpywZ2B0Jpj0ZIvA+ySNx8Fyd92mvZUKibLbaVXzGhY3JDf
okNYnx0Ju/4x2Om89bqi/ssz2d11Uk9bCZ7H7ikDODBKNK2a0sZxQIqTGLw3hVXZrp5A/Oc4qTId
oea7+4r4eDUBHUSU6f8wO5ftDcI/Lw20Ww0LafimWGNl1Ap+8rdeGPJm61AIEiR5vwzhaF0s1OSA
nfcmh0TfPTLzWNd9e7x48G7d1d5gQjK+WguUa2hBklc96q+oFIIu3Ta1+t7QEqzIz/8E/62T/oJs
WIbnE66rMJH3s8RIHFVfCrBifBJATUDVlpLHe48l8fMkxKgUwkVDlTWJHLCpQ6+ir3tbpvz5pEiA
gIfXlsJrQxrBGXyF4/9xBLlv9OVYHMAPNFfkHfd8qtHeyvA+sUF4qDy9ct6APE30moEhPjKAgUTu
4Y1R6JF/vbOcAxMO6rICfksU48q94vAnt8tatID17TN2LqoMPwdS1CPyxgHVGXdb3yqOePYPH460
QYsVM3ZFGUnmhvuiiSGD3oCWpXAF2+YGt6NX5olTemBNVgkrvbe9gKXmpR3q6aF2KhRj9HWzaJm+
wl9AmkKPSBX0bUGjJN/inTJ77aOZ4p5Z9CoSo48HHO8tjcIJ+xGlttJ6WzCderBISvW/Jn6LZZuH
xaS9rhu7Mn3h/3Y6+Q8MeFcHBTfmjJ7WMByTGEAEg3dH2rCDkJkpnwwVQvS6ZlYRQbANkMR1Uy4t
y9LGCfdSNGC1t6nUVkoVLAqW5E0e6Minhm1K8JGUMxBhKxLUAm8al0+sfy06AecMO5maQos/cztB
P3wNto/L0I900lIrPhywQz+EEEKHf+D5Lo8WAZiqYG0/QFg4L/FN00VUDQiB/2D9tQQ6JZHVDDMu
mp3VqOQ+RuWFLvKDngn3ouLG1Icl/ZgRm0QWSZAFR58kEP59sYezS3y4QMcPzl2O6paW5WZn8UwS
dEy7T9HxEXhtnHzxsKhVe0tNWlQUgO7vaoLQrNSm3SN25W2Esj49hMLO7nlaSVYYhRZ0+uEih62Y
+uKcu83ofOn2fVe+sIzlbqN/fbFKvi/PvgAZ/aoLOZDtmgCMK1nqma5Iq2xTMelvKzftDqAl5kHa
a3pEvWMsO27jKetscbo2FgWTmlBoZqZtFPmFWo/aBIlUaF93i+0K/IYz9fkN+yuuieYkvTSLWcik
77e8L7Z010lw5nKs/KanswmzdyDLso8Rw/uegSNxrShHnqJpYzqd6NMBbfVwps56tWkEeNisSAFt
wMMKSn1PYtdxMu25fTVTs39XFP7LxeXwq6NiRkm8eIou75nBgjAtnSoOLEODMkTO2+qNCzMXWHjH
E8rfCAOyKWZPCWhN8PoUqENmO5AhJWGg9L4BiW+sFi6UsHyFJt3XbMpPx+xqc0vydFZNwOK0OMVQ
LlOGuRfxvWHI23cwG3b6ig2N6ozb/CdKehypt3ysUioeqIEUKSOyPcVvg9BKXRU4QupWwubYr0tO
T2ZzPcKtaPHnoE2TD8HKygMVkJwyncDx0uxI4ZdV+TabOml1MYLMM8nNVTmiabM/rFnhywPOn0m4
tKQZqgA8b3xtIPZZ8BAlR30zzQx4+L44Ofbro+oil/5bk0X/LRoXiiZCwUZU03PlzaPZlYFQP6QC
sug9dW5iM3o9yid63hqzJ81M1t+ybAjGdm5181X31/e+QpMpMG4Zui0/XBHEE8EmuRE+B0Bj9ay2
XlA3LJfCILd/5KjHGSR+91ZicgfqncNwKNo3uMTh/XWERYeby6+zl8Vq60fwKkkG1gmibeNl54LT
4e84QyS4g8KWQ5xYzBMXJqSld8qPJc0HbU+iIhcbEmLOpLQw/+7hChS1pjKfiMfZgVsT7nQglX+1
xyy8qksPMAIC+QoIeBSjB/+OQ80k2Qv7oCGzn2+TUM+nIr6XLumCvYq3PoRAPLN20+dPohewV6Me
URIj4kZFGjljhbjGHwBssxpqylcTaoGvPxfcMupatLoMu/r091kJuckHHPb+Gerc93z8/d6SjA0I
71vdw9FNEZU/EQ7ViJHvPBDvPvZZ9R0MsnF5kHemiRZci8RYOky2Lrc25HXksz+PiUSuq6i2yObO
SxlrwqcclUSJIGmYYkGf7HVawxKDlyZfCtrjtTZxHiy1HixhcvsnOFy/WkvXIFuaWCgH09dfEDfn
TmlfoVLCfWFzrDQEvXcuc7xSd/2BodlfsKh3KnlTIBUG2xryAt78Sl0+QNw6xFx3iHk88AL1EHoo
JC1CJC4tWpf0fKBtGctM36g2PoRygtSlSH5gTzxsybKs1Oo7pyHU+SBZtfxYmWoylI+I+pwwY/nf
s9v6TyhBrmpmRj+KuK5EvAW/QNCQPKEk4T7BUqJUh0hiHNUu89R4KDOh5zrz+cGH0sIsDh1viLW5
WHZeCqOU7iT9LJNp1P+ujGJPj+L6g1x1ZTUoZ3xFbjY2ks+CZTcT2oyPnBngbgxFDSls0hv7f2z0
zO7zf1PL5gWOam6mHK9p7QoLRyoMfsDzjMQh98GOyCA15/q5ibKdfqdIFOUZsmSXL5FsL9B0ir/0
IoSz2hAtJ/OlRC60JZFE84NqccCyyy3CsanQjqFybH/6lmCzSEwZa/rhuLAdSenZxgYMwvr+dEDB
8fuXM9hFcMcAiY/nHy0jZ3Tm4+qblgYXvosFUOY1Fk3ARwxLt6a7fLLNfAtrdw/cU1x+6yu9LYV2
sNOUynRsTsdXkuNuU9SWSp06H/Kks9bHAvh9yDdP8xt3FFMOgQsHVOUEuo8gzShanG1QdBT1qzlv
u5W/qQZQWrSETkSCnIuzMag1ih6crlWGEL/fBDc8z1B4Ort2yNZ+Am/pYHoE2yoGbRqmk4A8gynE
m4rLm/k7AxuSKrqaHkFQ/ZPx0hq8no0OXt38AZxgtOPwLELkA8HOPYnjBJkVsNLVwImHOdzH4Yxp
hbrAEyltuwUY3LAuFoEMP2wMSFtL6K25smp+CaMlCwOIQJKZ9LfG5h+pGhp+29bLm4HcaK/mOOpy
weBa5nEoACn+qk/2/DlNxuxPvIGZ6XqjLqM2CfrReAO17XwbU6nDzU+omZgscSvo/ZxUYOUUv8vM
KZeExk7zjI/h6sGvHe0+bRctZ2i0TJoYhFP9RnILUhJZR2XNb53Cr7nQ3jiPS8XcxP1SCb7jAFy9
zWCKqFBUEsQ0Z/pFwqcbatXgQfqehZpnc5J4OHe6/V7k7RU4moxHtAQSmMYtDeplSQyDuL7lUgon
JGwfK2OK0qVEL9p9xgODCD+VOxL5IdfdZv/UOSsm7tHhZE3IJGvuD+dKVhX9qc0pnhkzDSS/sctV
mzfsypZCb/Uicp4qvmIjOHtzSJHQcy60mlOK3azHX1Xb80MBKH9PiQb/SMwTysL9fndo9eVYQFVW
E3Tiim7tmkGQqbApuSwG+8PJvLjg7GTrEepcbE+6CIu1V/FS/HxAzTcSjsHLyQp3Sv6xdbhcP3Wy
+/Rk9KLuRlkxdOFM50WUd9WODB4XekHN+1f69oBlqKuD3jrgEht7pXTxFzqm9iaRq2BS1hCooI2D
V8ruQy0ziKwbkJUkPViLAhWAJtGel4yKoyiDQBJX0Wt2jStqimfU67OIqup2mheeMcga15oNC/FB
7kCmPsRoneBmaP3tNtuTgdu/0VwvYUfwPsEVIZxpDjNwv/80i8DkfGjZmIlf4FNZTf/owNm9VS0D
LWFfl1GbkFDIiUi9QgGIWMqSSulKMYP4G4lV0S3EjUfRDmHEFQlbRQCuPm4FIayh9rg3ff2DpH4E
WnnWJALjhY3FCeJbi9P64XRyVEAKIroCwVLirOv4bEaq/iq2JwvTSrNN0+VMlguAMxZNDVc22/yz
6o6I4Jsk0M+rrIMjDBfPEjW44Tzyg0i9W+0TqGpCIoYPpKamULPPzC3v7u760uLJWK5t2aezVfru
l/84+hmw6RDZ1i0PgzghsCp9OKDg4OffANj/vX0MHZvsyx4kc4HdlnALlFgIKFyHh51pt3SfXAyK
eYjPCocbfqED3ajSkeqjogHRz6JrLqnHd04JFgbPs7rAvDxLszctNksvQp7IKJ+XEQja9rMsXk/D
A4YVOiMnVpd2EoSZFeEpspdz75lh64pP7q4wmeOtS3UOL86YMY6+jlQ54+t+nev+Y0d4rEkuT1vs
YNJh0SzUW+A8ygO4fbCv3xpZYkg9ufuCXBrozavMMcu+/AUEz8uYiedg6/5v1BK3V6mSoqsbx3fM
nxF8nRrQZPWqwbqD4bnN9eEA9OdmCJQYuEuuSWxbJb625xTVkxZqGPKPfnSKoXNHwnN+XI42uzRf
k93I1b0/VyqXtHE0iEAEXSLMr7EJbEYGp3GfOuy1z5ECo9fUpdWqTwzOLSnN8g0/ZLsYWHiwkw/e
5BTrpAl/4HIFjLl5miinODlgboWhXmB9CozHFc8oBSTQQgevI/lUFGHTHjUXS83DEkZKS1MX4k+d
PhJbS6TaKcH7H+0x7fgxg/4kaCh92FzYqO67yl0g7eDDQOF6EHMQrll4TM0IrmO0UkNK7o+FbF1L
wArE52rj0w4Eyf8VLLOLhWZx1Ym9KSWq+rmGPQnbVpB2bui11Qq0V3nzSdzapfvDghawGgVlt/O5
o2EJ7SdM/x3BUXKcuWQKE1choYw8h+nYYqfI+gjQP81SQ05P5QxYJQnyYF2+HPpRkAY4HAHEKRaI
R4QmWfLWYWASJUNP2pk/w1/QirBWLhiKlluZjL/joC4wjGHvXCX+UYlSCvJ86hhcRIHNIA7HLZA9
BQIF1XLXvuemus/gaqTRlNpXVbvpzs1s6dhOW2fCv4Uahcm+2b4BL2cfJeooNYaz29UZVsZuwOCm
cpqYcm+g3Uix/qsGkAxQh0UVFlcc7daJSkRbade6KmMzWyI40OIaOr5WoHa9IBnvnZHTfOGVLEtW
RmgxKa/sxQBYq9MpSrxeWS2XIm1s7NMlB/h+xGksuqi1DZ1/4Qei6LJnlI8JxGF6VAF6Vn6ZWPSl
UtC+FJ0AdOvTuwQaw1+rzgD9iKyL5RVXVfg7aKKiSbWeHqgGOFNns5/RXikowjrUXwI+maCeymEr
soGsyXuC7V/WW9BaO+1Ux6rGw+3bmiVfoXxbL9u4tVQR7rshO+mzRWKbu4r2vvmDf9i7k4z3PGme
6WtsBEBVtBox8lM1St6G2V+bCEbtm63Nh99GMnp2CGvoV139MDqRThknv07zB2PBhIkVrqq2qVXW
MXpJx+jsEZo36KJAX42c6i7aHmllMEB+y7dDPn0EvtCkEWQ9ElA03ailhypQwadWIz5xt/qfiuPB
ODwI4jIQgh4P0NDzSaF1crUVOuJMoTZ/b7hRGi0Y60K5fJHWUN4mDd1W76zWVjuBp5NMghanY4Wc
Ao7a5fGus1FI0PwwR8BljoO/YWCabA1tdpd/1mEFR0f1xrfp02nNp6MuBM2xB+FgGdSwLAJAvOoG
PlI76GhY7Do/hSn9wkIpEt2mLwU619LWfO3m3FUgOdfGLUpOH1ZORsoKSjE6NYXK6gfCkK870D99
Xc99NH6pM5w9Fh+EJjnyyt8SXB6ooG5knUHZ9wwjU9+7sgvCN3OvGp8DXaTYLZKh62GqEB57SDKM
qPoPKVbqjcG6akWE3Z628WZcfp79bncS3/JEd/LDpfNqKgOicZBgGucgVGSNq3az9HkB4DtZiRtn
1eJfdJiaJGGmUesE5sW29Ztyoz0rYKBwTT24yCG1TkA0OnlBtrUTQZ+cY3XzhF3Pqzq2OGYLTCS5
7MwFjQC4MazEsE1SsvFwZMOvcxhyUSA0BRUIJznf8bXHdxyroa6+7ghBe2/YCJWZGMn0hmpV94G5
sgdiTqEXCwYWy6nf/H1Sq/HfbEf3kyyUGeFindugfymw0c7PQev3ReHRGURqshXWpSf+j/UgvqcF
22t5pOGdBAzCZJwEBlPOcqyfSh265vlVE37JYOOamtjREH44SfPuF6shVM3sAbT/ftMpeMj5GNMA
/kB2CS/4M1dGixrUiQcn6ScK3YEVKTkMIQ41SSHAr7QZh+9Q0+dK+5JGBYZU8QvdOn85/tyu8+dd
AIrv4FWxVTIyT5xAIwWOfFVa4/Q5gYpoSNHYSxgrkl/NhC9qbmDAInRALtQBJBN9dznusHyT0csm
k7DGkxJCiZQXjG6lhmQB6GlcTlMbJatvIgp3wrsLpXlzXjqGf89z4/jZL9aZFPmh6In3Zh9QtaWT
6OiqfPSFoqU2ZkYjl4FUZbb8HvH6JegC92zx9ygQmwTfJ0qAU6mooP1FwpsHxyqwQUOFSVDno450
DJtM91Spdkfgt2UQu+x93hOqTU6iinRDkmL62Cv3gwYZs3xR8IDPCblA3blJ7Pn3JgJ8RO//uJxd
O0ykkn1ygBhxPUF9WOjvevFZcinWXGA/OlyNa/UhKQ+Od3GgKI2z0A7XnLlupLyiGqp69cHQTjeX
evBy5L7F4/KDNiWBMpS3F/TCjAZbumFwVMxWS1+KgVNnXYO01vFecdZ5FYvqyIjDVwdagrNHxwj6
eKssRyvDKxG7R1pTKJA1b39N2mc0D3aKSCqth9ItmtlekM7V4UK620II9aFOAnWaJ1vs3wXbY3Q5
Jih4AaVT728caxquj2wBXziCjNHkduGKnn2velWrmulZoR3wn2KhI1FezGsLrV4jBxY6uoWNX0zS
9/XTBeKzB9RVp3Ya9fGjcuuYQYdgH6Sr9AEGgA/Kys96a4+177iU2fik17JaOdiULYCbLgTfaK1y
0RtQHMt1X/xVN6x1Ho00T7V3KUrhQNHsI5pX9QX5bHMwbAsN1UhOvf3IDOUJJv75/2yYY4s6d1f/
519rI0no2EYW5Zd5vD6PXsnM3eUK4pQkjsTnUlh1a6N32wcWZDPdb7icdWYXgvK5IUBhLE5oZgB8
2eVY0Ej1q98GgIkZ2+FXnq5aH39OnseDNI3g8U2pWwTECb6WvX2k3b2Trg9cV9jVYtXTJVv2GVgC
evAy7LK22ypPCQ7GC7qqWmttL1K64lHFI6nJzr1klb/JOkajNXHMeacKjW7U//UDohpluVkSQOK0
Rc/znq8PsJjRSu2j56DLNFNqP6XxagwU4EPDT314EokhtnBMjiCFOCCyxgfIgfhlQKu8Qhv4QFwD
IRjDeOdHmT+mwP1SXLMeqz8KLVmNpSk+xOfYhZNWQyCrx/olneL9Ix0XxSnNMH0+Iu5dpvhvN5cW
j7y1/Dac3+ljGyi9kDCmXCcndX0aC1AUsAyq8lN8NQrWdbK1xE2vV8jRxqOExtMhYRUt1hN/HASR
EBecujVYU3MUOQpU1N6fy17NsbgEJX+j7lFORcDJk0P6cTSJUZde5aYB0E2CkTeoHrFhRfKtOVUr
9JRwdBTdR1ha5/kfX32+zrGpj6cwRDhi0pb+KgSRPHIfoMfbD6Pt0bCCVF3eZQqZStW9p44/gY2Y
+40UiqOHgPFzKfwm8oNc0DGn/Cm0vOAKUQOTsJnGY8T8QrcxwufEFRMpgka/s5arFCV+Uqhm4dzW
4uOKMjSZwp7XcpaTXI1I2DefgijtRK3pZAsYL3+qz8QsO5Xs1UQx672Mpsq6Xb39pY60ltAg5vOB
jZ257uHmpetsfqQpHJU6MD6shIMkKajjnSaWEFPVBI1OEb2N16VpcTOumW82cqyo1DXvSXY1DBFX
1JBa1PSyqDeEw90ikU8PwZ09y5god9tiywHX3bntwbRRnj+x0XfWF9Ym0FYpHsOoKtKqPXM7YPB6
WLVGG7e2PV+svYDWddEX7dprns0RzNU597N84eJuNFW4HL3TdZOfw4n0l35EjeyLkpcR+E1boXhy
DKdgt1PcJtCVFpdLP7CJE+pVwFqacIv/WOOWAD3wcWXnZNW3ncK76ku/041P48F4IeA6Miz34f9y
tk02+9knkXAGZl4Sd16iZ0u2/4HFII24/t+DS6ZzxUrLPDkWlkKLWOEVf2uU+H3ObBgVKm1pxOVU
bFHz2mlv2n9pjfVEGDwvckmNGuH/lx9LSR3V5bJx5E0cNL8hT3EmF/vy27ODLIL4UUwv3uzSyoq3
zrs/DAen/BNaTlcSHKBD5wQUMe6zPOMV7gYDrRwbylwPCqIt7jdgh4TR7mC98RUjBhCn474necov
OalfDziEes0mgQE0KipWNGITHF5ejCAIbEXLHe82FNpQaFGHr/nimaxV9oWGT3uU6Qinhi/0nfVk
gL32+OmP0bjE5ll5PHVrNsdqu7cYqWQzAtZIfx6QXFVbi3m8Y/6qmZ7OXzMUJ4IGx7JOFg+rqwo3
u8w98JlJ4Z5vMedewu9OcJST3qcdVt9CTbMg3pWQGHkkUT2wFp8avfRahEkRdc1C2lEoyHNd2iok
7DOkUQr3APp63QmpRU2dqAQet+d/CiW7plP2jarvw/697P5rkw1cYg4v2HCfmmXSHw4+6M7G16hV
HST7KOUDpjYC2V/LIKV9z3wf7Zg1rkZRo+oIVaSL4azS4gWN1cWjc7vdWhq5uhkykQksBzomiW/P
ersQjxuISMyuY8P5DJqi+to0UBWRobHD4JbYEFOkX/J7ihyTTL1w46IewDoykR6HTFO1nrzy0SYZ
bkA3XcuR7Lfc9AqhwYUbSPEVlQAciZb8Vuc+xq45e4159roGNy6nfv/TvRHupNXZEA3Jb6ZESaBI
tsZyMWPlUBjT2kw1n19PFN55wkxuu0i97EciwRT6YJ8etG+6X5mz+Oh8SQ02CCggEpAptH+x6e0W
0+0LQ7nX8qkX7e1tVslxgm6ikFjDhjYEEAVl8kwaHUf/MAB0QPD7RwsTf5et6Qcwsoj3vSPRiZjL
iekDMqcdymlPeAWX7wVwcGX2cFo0heLuQBimkV7PC9GAn/QN8TgnFS01Uf/z0IFle4I5+V1JaRww
dprDbH0Dgr+ozK1Pw0grq5c8WRtHpQjRKocFE5E0g+bIxp0UMvsUB4NzYILnVqwOJ5mSiHf6KRYH
KAucKEmagCOELuQcXXB82uf1s+lL5m2EdJVPE6m+FU07gl90HkFzAj+roMFcHe5RzJssL9XwF/My
zs8Bcph4vreaj32/VjHXilGtdHM6f6oIPaaPeBipYVA8Vzr39mbDfAsYPITgDq/Zve3xWgSSwmtA
DiKr/yOmHMwQav5jN9BO7nblaZXBqt+DKxMrtuJisDCug4O+bLUYcjAqF+MIGn1Ac12I5NJFnq/F
HH08dRR193Gim8qkpc179Agq8XXzDzxcyh/rIGVhAPaRn+ehMW40UuJ98od++yCjnClkwQZUAynd
mCL5ELPEMgu1odpywAWLqdKGFcFyCRYvhGBfCxOjgcwSDZDSnywbSEfqrrnTxKFP/egRrOQXludT
S474LBejJzJdAeC2xnN/Q7GXjR0L7sHJGn+eXwc2kbIvzgEvGyWAuWoZ5Xn5r2mbXKaBipIEE8Yf
JxrHWmWbBZQrQF2kNEosdzNTEaA5rWlUTMsbCnevTDMv1NwJX27teqAEtQ9bQb5Kro49VU9WIstZ
07VI6+71vEkOV/rg/WUVijZfv00xEawHrrRk8Kx7w/qVqukAICoN20P5Iix/wUNp2XFL4uH+7fAn
USqek6cJVTGZxv7gxXz7UWFT1JneGs9kncWbbewFzlEfd5INGMLlsA6oCA7oN53NFd2gMc0Xr8wJ
0RS1dWrLRlrppRj4V8VGF+nrJohl4nxtcpk77PU7uLOsLYfDN8/4vS1zorTyREjl54uuEl/Unaa6
83IqcTIrQXQPTr0lwJpmZyM2EJ/uZf655a+/4jxmyfb2xtdLY+CZ30wgtgG1BSCgApAEVQ/K9SNj
1wLfPRhPq9ttHMl9goBk7pdfyrtf39CChxH1kKS3aFf3VX1NhTz+Jy+jSH5fwYzpYtuUNZ2zo+ML
cfXx5oqXtRaA2ix5qAGURPQWXgjD1ADQQ/FeL5RwHrlVjfvs2GPY6iRJxXAATKPjeR6dDAqnnOM7
NomyYOVtXAGsot5CFTXhi2qnh0PhaAtPwXIFjlPpku/H6dvF7urIMvNBBduTMG9iu96r9UQStKDw
1o3bKi/6m9ghXOWg8eMt3uIHattOyFFwj04f8V68NcgDdJwC3sbadidiUWcl3vd/5tRt/rJHLxoS
JQqQFRm7EWBV+G5sEsT3jIMLeySUtWjpbuwsOCa0ekYstt+ej5aioL4LtyTFt9FWDs+D8QJleE5P
LpZ5Cc8ZLCe+Ugif7T58i1/d6l1lSqBGtOxbIx9rYcQvDJMy1cX9OsmgvjoSlb+4XKrt6IhUB4ru
A0IirwKoeYsUFBF53D/VqOXi4VJ5P9ItxLe9DmyDIW1s0CO+T/5Cnpki42E4HqSFyZZ3vGDyVjWH
2UAf1WPZ0IJF/Xti421Yg3ETF/G54mC57SqkjI7DBM4tlCS7M7LaWlp7BKmlCKqRzGaZChY6gXqL
U/i8siwRDdGiAZT5Y6ZomrktmP0tE2AdAJ7cdHjmSpdK2+XPTekHOYqQJLGbJ+QGn76dHhqWhh0v
aH64bt+bT/4BKQKVPgxN8gleZlM3CLC0MpeHJ5jlrko2o0hDXtG0qYOjTV3FSS1ODHiCNe1Ko/qG
wECYn+w9aXb1+DUOmgOqS5vmnJu8QfmYu+77vtZ8ImjLFa5ijAPN1+CBcKq1PUPWK/jYlIpaMOJv
bwqdrXWQQCdqx97We3xumQMriZrtxNKW7dPZN4nNI82+NUyKDhSd+wVvalUTzobJtCghE6CRNGD0
/jHAs6+OyyICofadxjesCBFsAK3PZIzi9s3BuE+alYUSHYbRHLtwJt1wJPJbh2ETsDoL70L72tzz
iN/NzJZh2w7HtHiG3OmYmGER2jgBzenXmI9bN4spacYDYkC1ghrS9GqxtT7v5u/AWKoJr5sqPY1d
EvDvdexdHAb+8s+feqQPvhryYUKtqXD6oeRGNlVaAgNn18pl+WAKxlfAfDFZ7DBtSvdl+P4Bd3bd
/RBiK2hg9YezUgzi8LtPms0PFy+Z7JMISbmJFDpc6n4JtKVzbDczyi4ecMbF+q9m9Ag8sHWUVmAR
IUsvxuQ83ytVNs2IZCiWqvCzTx3Bt7OfNvytfVCCeRP47bdUIF4X+XcMKKDstAARrb7kYiEfgXz1
dCCH5VnzbMv9F8GTwCdPWSza+3HKgHMU6PO+MNwoM75785acdjbSB98lo9upkDoq3vdGsp3VaNj/
1y28OVELKy5uPyXg4gpoNpZD4lMYuTGxYOoV6AGc4QcDQMtKtDbNn0nD1ynFco/3fzbk5YTxZ5Fu
Ne5cT77/z2lMdTrx2dgSNJKm40Olo+WmFCXdTvr+19Xj+u9H25pRvuoxinQYNKEiNyIiX6OxctvZ
ajAF5hbraM8SVjTzT0CeC581CXsvLserVb4CYKBxpyZB8PnawLde1OG5Cp3usRGJj4qPKJrTxWSc
OHhanW3Vj+fBBKVM0M0w0YACexZJEKEzBeMgqluguyd+5/6bZbc/Eog47+y5sUqY9fsiOS3VtOTS
8/Pu2ay/2UXqgcSSGzF8757HFbfDInklCu4ej7q1fQ3u8BOEKMaCMNH+9MKmaE483Ft51GFfCLKX
08Uf7dqNR/UvEXNY7xjBMby6XGYlYK5HLj77kuJo71+T+SOZ3ZbphR18j7JwXpEmvfkAG+g64Dj+
9GidsiyAur+vG2XHSsIGD9fLGe3ZiZaQmAV5jmN7rNZxTwlua31IM8nsuwVWAAQsqi/Q5pMYncK7
0oLUzizb4LrvQynii/OynCZVscZU7/Anxn0z4KthFdUwKESg3pJJfYiweHmvVDiJgXW9Yc1ZRjoL
bn39A23cRjLQwm90k3vfDkb9vu/XTuLt9e0rnu/5xrgKLvySB/JxfU6e1gfkbU3AST1cXN9JHgS2
wFxT5jozhk0ZAmM1sA9pa7xOPdDggsE6aAhvqEcC53sfMkiDUMT9HIK5BZ0u1rrVWiJVJBLsl/HQ
kuIDoRfjFOPX6/c7PQDQhvMwAsKQYQfE8hVFFy+Fvq9ffHH22k4fPtsmIdoQXVay0NLdZumw8RYE
HxzHt1btnCwvfCo38Ivzib+6Z101kyyuaTvSNd2/Q8UXkOc+lDPyeZsQdqnlY8eU2Q4hGmsqiMUt
zq9q+9HEx00SBIiNNfFhgRbkm7xN5mmANrx6dSuKEZGzqQNKJzG80SmY7eyP78D9ffJFpkeHIBbx
zjdDyar5yhP+xuDkVH9iNE8FPHBnzfhxSmcqgZIRAF93PJ8CKBc3vreRtRKb2qRrIaszXOWoHTQF
KKEhYKT0XW50C/EPmt5fOQOOEnQy+WqCDMVr0zEabF5aVJAjgC151ouOdpQ+fEjAaG6+2JkEogSx
jQuIo8OG1zD7eO2zQKA0EpJRhfEFA6M2tshAiWm/bGDpud2HyM1UBfeuFeF5d8AlN2nEz5yNnvik
qNdBvM1lLkkq8Xo+Qxe/wkugqjvUE5ODAbx3ZNQ0uHegf+Ke0h0OJfU9kWAGkhLGOpOyvG0yEeYn
kf+AzGONpXa2TwwRuxwhzfvwPV4FUm07jHdqLOYqxfhjy9sKR0M1PX7mJmqQUIF152zgJr3bZkQw
yfXlFLz94gOfRr9dO0Tl10lOCG/ZWeBoZdpQOsuOFy/jTHRYKWekLe8vz50JgGQYLq/Ozs2WVv8P
WHro+E1oQrEytXgGvNOpvt4jBZMO9nHnPbxTxPBls0x9c+ggYsH7n/TdoUFQF5nRmzNVHfLDbtt5
weoUpZijNdigSL+Yxe8jyEeQKNIl0btUb1U+whE8pX6QpHk20FAIhzNrslJWdaSWFjI6E3ttfZ6r
vfzRfkjvHEdIgeFOzymR10fs6tnB0oBPk/EXbS6R1tJ4H59upiq91Yww/S/esFE1LSPiofiJQF1/
AYTBx2UemHNv037euQxFVJICBO+jN2X4sBsgJyG6ErBd/bOhhMBbvqhpJh0DPM4BSLV2LWZUWW8s
FHyU3TVGafvzVbTKXr3F85gGAP4oQuARzFVCq3ZqOzndPEPX8AYr6CVa/4VK6Z81kNQ+KK9iXRSP
ECKKpWD6Gw8/9m4uIGjDm6JT7U5dAmzOP6UMQXVNUS0CF+ALSwvwsl0wBHBoPQbkpjbFr2XNuRjf
IWK8jjN0WgqVv+rfCqr/dz4Hzx+aSR8rE3YEVEfb0lbK7SRDHfqSBMpS6o4o6+/dbLlljT5KRdJ+
ovXzTgVxKAueWTAMMGWPF9e6weNf1DLoDoO3iJTt8AdGo+4E/BRVD73SlNNmnJT4LivIstjMFK3L
bnSSGtFy3ptp0TSpfJ1qkIOGXKGh0qNHgfN37neYCt6AIaExFsQSlvmxaO8yufcdoKZqCmUFGu7l
SeNQNKuHlk8uR8FVaL4Y/Xs5SZDGRBfriBhsjFkQYcvxYYB+FoM7yCSdR/HOQ3rSIfGzK6uz2RH/
JOX35xk+MdVkoKr+7xh/7EqhRFP+3MO76d21GpBUDbbY7+K45lwQfPSS+Dj9fjavSreR4Dxk9OpZ
mP1lCkFFkXDERp30WCJssFvq/iOV+a3aaiuLtSqSkZ/MprZsAQXNdENOhJw4vOvTv6pV5PyTpxs9
qiMN1fyOu2LHWcFTW3uMtwAjZ+Rvv4j20btkXjr+6JLJLVOVpJD1x8DYc9fPRYw0dgXwbvVl9Lu8
g1pwOvfHYpLgRm+qHFbDSqbedT0OppfF1io8YcJQnDp4g0MdWWvXWH98wowa4KQpdlgtpGQRnhh+
Za/oPxYGrnCRcMRs4LwBXpvKzeuHykQ71N1546EvKVD++sD/X3xTcBSWWHpdO1KQCswCHVSq8NcH
5GjHEUaeHxzZLwnkNNoFsqSIms757d36Tx0A9Nl99erhxWplgOaGkWAtTcyZbItn2HRzuhKn4EpD
kQe1SQDYdU6EhX9PrnKpsWmVtEXAvTrBSivyNHVYUJcy5OSb5Nxz0u4FuZ6sJATdiDDdG0tVkwNP
QTAroHMNz18Q2TLp1UBl75Lx/rmQqtqGiWe/ld5HbwdoqcJKiGvUpRpu40YwlOduOYvnuQ5CJiYR
d4Mh7YZheh5tQ32oVLCV79F7g2uA/90LQ/1VIqHlHZtOYsrsO1Xvpr155VZY41/sisMbDmJ/PwVr
jShoiMAImOMsd4yOZ28sMsgx0DeWzdNiJ6n+lZheyFbA5JamdhqwFLXIu2Inw2Tb78e6a+K2twps
VgsQV6i5oAUzd/3KSHvx+tcfbcyyqEHRX2crc5twBQJV378oanRhV2CUnO8Fgnef8dH7djZQxCtG
hHKBBNGr9jRlfWbNEsOV36vqBVKLyo6OS2DXSFEAIigMeiOt2f59UlrgWGQt7n6DEBOoTZhfolXR
nj3glrdK8a9b9/zgCJXVElCdvvlueXilJGdnaAzw59GbYE4ONT8RH9oD69Ho/NOtRueYVanIawG3
XF5J72n2o7i/2Hu+HFM2X7D3pCWoeJW7fns3DHJwwFHFwAuiJRJgwde53Tv3k35KGl1Q7oV/nphm
/kwmi+wXo95BX2AUKvQYG3z1ISNEnF3RizA/8soEazAojZHeXzrSjqJAGWHMorh7gwxDnImPHj9J
osGeBEJ+NkcsmRGKd75FbqucSVzNeEIR4j3FkOgHMo98cQJEJfA+PvABhkr6ah/jn074KRGXky/i
vNa+OZSD8m9fMNSDaX6telIqHdVW62uNNO52hGOQgvxI9N6gV922bswg7gsjpbzZFUkG1pcflLVV
43C1wooEgzHSgHg8YItyrGtd+4GehMwKlrnrGJ4SQuqXLSEpv/rHkpW9/jCrkG0Pu5+WHrZqNaSe
pfl/xPGfAd7BZC+MpTeL3uF0kCgosZnq1tA5qQksZuEuXlDgftbZ3caL9/u0QHGq2fwtWbZGDuoR
NEY1TrglyNTS9bBm/LWysFpil573qEHUKMCFEe/uFqQiq6kgmW4CRWstHE3B+aO02MPEJvKbWr8m
CoxPYbPAso1ThxtKLijaT7q/morT/1p5EMzniI++5mlGzLBrUs4yubZSb4PXSW2fuXnmW6FeQKN9
nba0BFGvYYRIktFVpEjIWgQKiM/vJ6LBdvFqqwifnUXRp1/kR65IgrKncHhA6OPoxVAfopxtqWpD
TI6AI7SkLEXO1YpjdiJK7pJjqWoIGWe8soEi46P5P3YUB0N5Ge0w6F+Jl+Skpp1BGX9//Gtd3HRl
21AADkJkfHX1fP1rmscpKFQ8bZEvS1MDplEOauWSVr9hfLicCjH50ixvAaiXn9wc7lPupzVQ+fLV
3hFp54ywpo6KpgXzMi8snDD9oAC0SE/34yt+Ry1hebxpKCh7tkdvxSKHANn8oEGsEkP/jKwcFEpF
r3pGjv+hGCdWmboBcFkBH8sK54uVQIsAmwYT0iDJYlzsqMQOP8RjgkD61enR3kCPkOLIMAzhrujK
TZEg/fwJvaitf1oc56K+I+J176O0+7C9TFlfej5qrdYnBMED1z7sRH5R6YPDhxjD40lDTFX6wem+
gXDDWnz0VqgUSlp4TE3amcDtbA0m3iP8kDjFu/GDOkv2eNhvxVF4LkiW/+4dT/8q6Lnl/c74s7dC
WTnKftxcanFmCUUy+rIki+diMxLzXoH8nV7bCyKocNQe1JPWkdHixyCnaQAAcinHrPr9piy4oVFZ
YwqYEltVBSsLQ4RXMt/Cu4JJ/FaAM9ypIfd9qh7lkePamnmwhob6sVafHE8hEPQguRckviwG+PUU
iVPKynhlCQ2kBLHTV51Hd4n0FBFIUUpNhrCRcTYsTbahvG2J5X7Y1L1/9qwwpwyZBdk47R7EhGaW
dGpbonkhTf8jsX1vk/uKioOvEmqag36zlPOGlYtqpfhBj7WzbONNbd+usEz6zm0kX43vboFjelnR
VEuzyHWPpmVcHIsIn/VqtDRUBMB2Q3xu1EyithG32dK7x3SkZKppyyElbm4GJUt11vc5yjOgP3Fw
AdGEMzW7wwkDwr6deqz6d8RdeRvCUxl3aWw32oGqq9zWsCLUU9LbT2d0h+F/Dq+ZxByi13FPT5Dg
qrdSSxoRKtDWvHyQ27dD9zveXmK7bGPo39oVt3aBCZgAPXyj0iqjqVC3M1/bj9K1nTHGlhGRaTFt
uVFxAqyvY3mbBGmM/DUlqnvMNkuWh2zv2W/pumXZzxLz+A3KMX3Qx/r+0efCMtvIstmlp0Gr2cSZ
VGgDnDybrejwa8yZ1NwHSEHpFoC0m96TDxmfb9MNh38TyJxOI2iuAe7vpD+d5dEm7Pdr6NPFUdHM
gEMQFEJNavUoZEdkMTcBoZBoRUxKN3NJhemzwZPFWvSxx8zgE+R6mfBWSYONGEgN/6jTBpLJP2SW
50+QUSz7avb0bcB76wc70DSKVVC7JhfWuvSOnM5xaJHDbn1kNjpGRkuCxnMEGJLdbuUZ8uB69QQH
CJF1HpF2uuPty8SdeVLpxOmEejT8TEL354DeTtlulN8XROd3NRe+hWdWZuPKs1yKFk8a+ns5rO6s
Ntw4C0QPyqAGtp0ZmOFftpAiy5pAuNLUanNNgNa8ZZXmOfQy2U7IzY+8VseJExCxLAdloUlMXa59
We8mpBmFGhTgrRTCa9/aeTSPFc9L2nd2OZzBgya1lZx9eq2Yq0raJ6InZgQB+JhiYkaYgYZ+gPUJ
HY6jyzEDSUnK2PbVGmSAqlWSPa/W758aWRPkc2RWWk23mCO8relbInsVl1BgaVIVaMYmVu9F9ewY
Z+fKtTzOJLwpP//jjifEltRjPVM016402euufEG6OLCNTn3xeWviYisukWf9srucKB2mIyfaTYlj
TTjEz4DaxyqH33DHVGd0QGgN+s7g0N0guXQ+3WeZ0JgUlAxm6NbItxHWPMDcqlek+tA0otAwXFGQ
02bjgYN4nxIn9QkR1P3T2QpKRV7HOFQldi6yW2gYYUESMjWzQZlzqDdNjh3zuHs7blu82pLMZULe
Z+NI1mFXfjnqA7uurn7axttzmHpWgps/cjt1DrQzlCjfakL5+RmYv9xGKFgpA/sB3+cKcSQN4ktI
q+oG9l/FnyAUXkEQA6e7MhrB9vadZ6WYJ8Xcw1gE8uOLZxQC0uv75hqwkNwJR+RKHCynByRWiYsr
sM8dX+byZITT8G60vdwhBzoFeJuUNJavrHParV26lEXi61U+L+6nSw73gmt8We/fz3PpOYQ6y1Uh
gf/bq6Zgzk2mowwFKM+T3SlQd4TvLsjazpXmYLLjipg7+MDWb2IcnI0DnH5j/nffXtdoMajveViD
89uEwsI3AGjte9OyijLn0cH5EovVI3hvKfv2aSmrQuqfwmBkOKQiDmXEQRvGFeGIghPtmPYlxVpQ
F/MjZG3owAkhEabgN7LvZx9UI1KA4rB8a0E7slwHmtidrL21EfqFOtlMpu4SxdizH8UYdAmK8bjm
/4+quLTxYxZP7sCQfnQFh4vyKPivhm621NazpVabVMCMJqNgwdjZjWlxeUI21ajFajCiAYvR5uwf
ZkzbaLrd/8LIS0hyMysccNTm5uBrzabowiUkYdR9bzr7tp94hi8b37bDnO5wykUv2OqShRsJkc31
KVD6SExAFJAzaC7L/ie59NPJwVHx9XFwyH7313zKZclry5E/JtyGi/mux6w2wFdBgHNzFIdheB7w
VVwYdDtfZd9+FVc/CZIEB2IlEQ6QxwzCyakXgkspH+ZqCUvyOyvtMz4VE/ICXPBFykas6Y3YduVh
Xur8z/vJdYhn1v/B2/MuhwI9FWeL0WWS9cyn6hdkOKQteew88Sgozpx3NcArFS+Zdmv6udnGeK6c
2mCLrRxh1TZBMPfDvCiQYsOH9s384LE0vFlGVbXvmiS0xlJ6wpvKnRQadecTNU7+Y3LxPj+6OFYj
+sY0iWy5kzKRzAAWACvcs1Vi70x6BUPHV6HYuSX2p7/IHQXlAqTV8RzHtBgyEbvrTNmwh9CgIgGE
nHKRh2oJyC3lBsW+0RiRHT2m5Y537/MiJta/aXhYV9kOAysXRBT9DO7qA4xKCU5zEUiPuBxRdfjb
WT8tvyfMY7GfiWHeNZQHLatf4sy1j+EXEvvnTG7YbDEhK8eOWF/7T9dRDax7Ffkel3lbPV6vbK8V
uuV+gH7mTTzn9biwyqTSDJnn/XEiv7cQbolw0CVFg/hAS5vbcUurTT1FOcYOIX2potZ2hF0ncRM7
icF0e5l65bQQ0vh6keyhshIdtAOGdjauh0ov8UaBEoVkyGBTuD89/ejJGDJASXqLBJgBkOxQ82oL
Oto8QdSLHT1Ux3uvG7aETvNCcdgxHzgTok04/2KfNbX0IL4dC/aRqnqvf46cP4wWTqU0KV6JYEQM
vLoy7Uq7W5utEVQSJSyh2BbN9O7qP5mF89cGeVZqNlJVYMVoHjvPRPBdXYh6IADnUk0j3cN0kMsn
4/ZnNNl9D1n5R6EMGacPUTxpmF3y5eEvlZu3iJRwrkFqJRsvSCNt0LWpEEQrj1exg31demXjWaiy
lDS6zxdSnwHgAfYq8Cchyo1BXKcxuh5C1/qZ8S2jfCULtuSrneXa14Ej0zKnyE87AAPtBztZFK69
0m8U8OR2guoyEb4q7LttUHWD/gIFuT08z6B89u8iILyyCgjKyfvPMD84C9KS19uApbVW0lKRQi/l
VG29FiCs/fQPUbfpMG3eIhzSiqIcTaDpZMEbvrPssJXv2osOHMOl4H60TViHqpdPn6pvOS86ZJGN
Ctmkg8QX2XCg3AqBpy4IbDppxkElBNTulw2uu4D2kYyCY9pa89hWmXjmZs1zbq2GXhQzg83yg55L
W5gF5l7ZXvD6bf4Z+tuHIy1NyF2QheZs5XSKrfmUa7SMKQ5+xKABoPcmuOGAkJ10h0f9OcXCsNgz
4O/IwOqtiuaYHTWCR4uptDkxW+HJFsKFc+YGsTaoPMc2tVJqLmbZBAXdlrvXYiriBNBqt15TFO1j
BArfk2FP2N89DEvdxpAduw4M8BrSU0bimtXu+bU6BLACdq0UDyAC6Z4sz3td7PShBnSyb93bkiW7
CdCeUMPy8Y9dD65lMoz2xEP0l2dh0eVQUgFqB10Um1qcxTXQC1uqwURlNPu0oA9JEw2znKwv4Dao
0XYihUvcNX8ZqJT1fDZunq+zwy7YyFgAYHvjjA7MPpOULq75IODevn3Djab+MSsC5p+CZTpAx7Bo
q5Hys5RDpRNgJPMAJl/mDRRPeD9+BDId/XLt6Z28gvwK8856yxbqvp8ePU7gPRFUEBB6eAst6urQ
EQ6tUbGvSG1YRBkAtCN+HI9kwALJ3Yj0RtDBLAHtGwf4NC5oVkp/lHwKjWD2ynSkfi30CPuHQXuK
12BE4eiuIVswiOJStembz538w8XQ4CVILqhyC+vEDCO8iX/WfjMewt41wkJhIVdLOoc8MiDbnMuk
5/5snSjtPFD5E2D0GZvLUVvVV+1PYiG+9iB29Wr6Pq6zneVle4PNeB8cQS+/AT+Aj5xynxYuqB0x
7ul0bYB7jsTu67NAJjTFM44pUVDnGFCxXQmKfyQYLoas6NeLrEkLtm0aQesAWPPXkHsorhDT6Pcq
Wxw0H04iA1AFJ3H/CklZVZU4wveRrBTgeWOxzX459ZjTt13lSh0PLhytMDk0JDs5r/TLN6qvfJBw
uNNfKe5aHcAOE6VrN5V8C+UjYeyFA6u/uut5u37TJoyJ7pDGTCadLtKkUzhx57RxM39YRr/2jSJo
wl3LecqXLQ10RRHRbuQHFbS/jE5ThTAlX5DKcszbw+dcVAV4MTFKqLmYnHQ3flQ2NAPMaHyFDjeI
XHYgJJWA5h1Xmeki5hUhLC4VtNCdJw2WBn+JNqNofkw+ifNW1wKmGU4W/jbFHaUa9nu4NkyoQUec
NCVNBYnXuexdR8fXL1lCWz/Gn+Oh7Fwpyr1Q0l7JdRDFKGX3JtoRRIkvMovLnI/DWgnBP3KU4sPc
zOkqpVfma3hEnpMpwoQe2+ZkaNWG5/3oH3c9HL4GvxLnyj/w87WVE+7puWc2lgwQ6h8Zo6BnqCcf
Qe+00dwmJRJPYHxUqRyo7eN+T0FijC/7iNNnOXMld+R9OksECtD8o2n/4eEcjOY0XIsewcCE8PW8
xHuKktI3pLSZ0X1KIHJunjgcOyhzz6cWDokWlkUq70kT08wFIWW/fJFX3Hds8rtZy+bvk6kA/bjF
ekKOfSmaiSpGD+Jgg89S6Nnkgf15vlmbxg2f/xlkfBYSR1AbxKN8Wb1ZMq7R07x/a1D1t7NW2/o4
U6ZFlhDV9v0Ehmg6knRtkMgHXfhBdeRSZqzBss0WvKQ2ULRc8EFYIo8uTzkvSsVBqpSgY05kiY/V
EZ73/qkBQGv3NesBhVi0vCcAByp3/Nqbr9QxgDh1Dis/mG+U9jOHXb+FRqvGylUitg7zasoNJS9A
QmL6iynS5fVP+7VSYmsag/s7dA6Dj5XEj3tW1S1N/yeHcfguWmpY0xxRteuZr4JVXz4xjazdDsVg
+dDlRroG4x1WAbZosWLX9aZB/StvPO7F4SgUf7YMGeUDw7W+DFt3np+y9LKar0JLBn467LyOU+4a
uYh+4Ib2Jb568qzsVrOV3HyOv0gFOfqC7453nDuRoBGAwq6xFuU7+MO0WWsuORg+D0qTf8s/vtHQ
2lI6KMvDOeq9rucW8WIit/pTk4olwbmNmgYTH2xbVmJGyJnURUsY/gvpqVqGFvzFFpAyNrkT2TPV
nWkDqwR0C9C8HaxygIQuDTAuWOoTNYl8ueHqyo0hpYT/4I6zhf2NgbF36Rdgb6l9X8rcFQQM8Bxr
HLCK+bmQhllGMoSJDWUjwz31VHinGaz00Zyj0n4VxJafMckzUonTv7p7SMppxDaAYEJUvz8LviDN
IMqiliTodvuMs2mFmlUub+UGW5LmZGPdU4+g5hfnGkfXK6zGT+FJcg6v7+Hqjhh7FnQ1Y+ke3R8o
BkiTzBIQ/t6wVa0qOVAtOB2TMZrBnCpgdVv0RG3RTW0RPJwXXUaAUcUqxzC5tPUfRA+U893aPDGE
0fq+E22RIxHBZPFgi6JyXkUgUlaj8sH1qOFCLXjK0etBrtIB94JRYcnriJxgpnTlYEML8RX8sZY4
vSxAxMhLNDJrq1ho02m52xjpgJl5KTda0xc55S1CLOusKx+6T+uX4VlAgyt9fGQ0whd0EpReh85K
N6kdIf2Fd9lJewtLaT2m8/bl8mJnD08/dhwM/645iXF3f8gduQ4oTG+zHQKzlfsbMjzKTh9lPpat
+PRh/GSHxLF21oZIK4q4ibzZOnmPgQZ3PuEUzuBBGGkB34IyH24pi8bMlPNeyxT76pnNaVFEJ0oZ
NLE6OaBe+JAvqlTHirvJREIBvj9HMVZF50xGoIv3OCWCW4iEPQGUjJR9GFzrJ1ET3llqwUpw3poq
pm157Bj9jia9Q0Qm7qe3yJEHdKLzjEmoB/msjSx4UakUcmPWerJYYj3wSObd0mg1HnHgUhQCsaUo
FWfcQmXsNySv9DpSD7soJAJXdlyuM8+/sO4NFRJXExWqBqRLHZB6hero2nL5MM2qDG7lz7vtVyRP
pJO3n4PnNWPABwJUCcJf1M2W400lc5xhPNdrkjNvQ+9apYEmmv/RfFqnwigOnk9lRqzw7NxHiMV5
/BPhj5JUVjX4rVon5SKMXbZSPONHSuaWlztVHxeTD4mNbLcVJAoGpEcJwlziwcvKRggzxNV6/nvn
CPY5h4W9yL9gJBLG1IPkjjJ7NsTTKpQ35fzlKq0KpA6wJGESo7Q550AMjHCsGBlD7nsRy4abwDxp
Mb17Ck4gsRFo3eQs/RUDKOIadNCygbu/sC8k01chBNL6kHUD+17ALa97r24t9EX3VpT7YvQYX1G3
Svs9Si1lJiEwtphSUj4OHP2VKMPnhTZa+e/yNHy1a6F0a/giRhVMrAoyqke8LhiNMXAd3vXKOXwn
6Rn8ebaNQrOrqcrl/opAFQ2r/b5rH7/gl9k9VdoJ3+7/9YzQCHiuh2Wg27PSTdQzFtyNZmTGL6cg
eQbbasAvBien1TQAFcjfoM8ynTG5x04Y8aKDUl/rXMJOEAHMZU3Bz+Y9qSUtMw+KiPgpmVM+Z1mz
hmaEk6BWmXyqYklBDhj5a/C2KiHsGCRp/zRqFpBNbjC0aQQ+owly05LLgCzerzQ2d4EBDXaRhHMU
vJwvQxEe8Z7OXBTban0w81w7fuJ1wvK4sZP6X+Pu2FAjlBZn2jYi/OBe0YsNaVQ8Xiw4OQZpo4K6
qkREQWUWrhpvaZg6dXtWf1oSlu/PppX4Ujj4HmRThCs2APWqeO3N65I8+fisq3VHo4xuYyijMvRa
uyHNwnR3CBdPiAeTVV9rp3fmjDOnEGbe4P8WCwS1OTKY9SqMppDu1ltGG5WNcRWBij7I57rqu7UT
dp67MVbDRRY/gHldaOnqh66zLlVp4AvpoAyy1yiVXUDefZRYoeq5K4d3hP2ucGqGOBUckjyvr84v
asBRgk+obPERXfT6lJGIV4Q/MvXcuCLmTK4bnzzfXEQCYm90UxETeAlkCSUY1MvXs/mZz978kvpq
WSThYQ3zgqqzwKI8h/puZLdjyNTV9BT5kE3GkNjt4/Ee9NOCpgvJ4MDSli0QQfYgMNBt6jVawQxj
B2fP2yLkQp7SxlJl2zA7oaa1j1FWjhqOIwaCyyRJT7Xk3yyi9LfBlPal7Ycf8cTNbyJnNp5yYcBa
sTAb3cEVkrM6AIDMzGKyNR5V846b58gEXEbtAx3dKyYYHqSq/TjvBMAeByUgz6QXXNxO0l2/NR6b
ZGhxo3MgQQgbeG2txltKVI7ASzJRPsJRH1jbmZFBd3Jr1a7w2IboR3HLb76oORPdDqWAJsiba8Xt
26BLhT80/bZmh/ROcWCiNKcFt9G0Dg5JkQG9/Z2cT/zbSCvTON3ZyTgz2ImC+BihuRiuEZDhWZxm
ZxLKiiy+FeZF0N+x9JKDBphFQ5VG4bYOSzNibORboPeU2FLXOe9gKAwKbWCQAIbggDDdpbtJzUu9
E8tjC8PGpVTOL33w3bpfKOgOe+zndJtBJdH0+MVNbv2aIRKV72vzsqZyTcTIl9tcH+pwKt1EY+gB
RpNjXw2pH+ssuDo8NIzuzbuP6eIns+mgw9gfvOKzrYi04JakHJwk6Bx1hBYHH8RNs5azlcXtxMat
K7TXrlnKESI3TU94KavEbmkUeNk+OGkbVmUvp95QHaNvssWTgudz7l/OBUdSZIo0Wm2Uq9eEJX/w
MoDFCQd9R2skV8dqWGPez546h4uo630gUF88NFpiEM1r5+jKarLAAiKPrhMf5fMU5xNPon27doMs
OVtubxEb1ReDRxYefl/auPTeugbBBYpkrQ4H/a+eLRDEECntb6NpXHgleb6v4phNRzWSODXntcBP
9NUIPpINk0WbdxZcW941+zcVcSAVNVhPmBHMc2NMD/y5hL7as8Qe7eEYPffA7Of9ZlSP36nuN2yQ
KkZtgOnpwo+PrKzO5HY0WuGlCBSr2X4dIfRn4KCFV937tCLqst8Lbowc4eE79cKVlAyQEecF74+L
VTOBc/XTl7GwKotyA2A/ofhZm6WBR8KUaEOpNq8AkqcgtePAr7IVQ4TnpZk4jovlvG4uMcyMte89
7ksM7+BvAwTX8r7ST49oaCaYT3xG5Q3KI6nqftRTzIF3h38i3ZpUfv4glN/dLYeLKLKpU5uGdLcS
Cwi/dqTqFm4eJ4qhriWyDGhCrhn8FBLU+EztuMfqVQaW2ECDMK9QSbDHgOp5WLmqWu0BBVIxfJYa
X2FUlCWlFuQ0UHE5KrSz8CYvyEb3aiyOSVXPkce6EMd2dF2s+9+dJJzyJ/x3F539Msjq1jNAqIlZ
VxbsS6PYYj2R1SjSaAi3YHJDapb3G/9QNX2HKmuT/Cck1t5GejLMeiDIG9JTw27yjPvDpkVNwEWd
HKT2chmvxLkMWHbpCxJKM6/o2yOXf5Xx1Yh7Qy1CdEk8B+WyoJDzjBtsfOpNrXd7XMtJcaqra2wL
dQkhnMycIDIuL/2w2vZKTFDD+p3NitS8HlqUSfktwZTGgvi3GTeUqd9j38FHtZJnV4e/gucDilry
9EIlRq1/Tq94IDTPtwpA65iqj2Ia7UCgqFgBeA0aiM8PGBU/TOOYXvS74izXUcF45UytG/2SWU+1
OE9TXfibnfR+loZMmS+RilCv95zOK7Q0UlBpiu96cxiI2PlpQkooi/QlN9Oco1u4FBh7DQqtYv27
3aMSr/YmEF9RDed4hD+CvYt028Et55XVehy048fxSYVEzu/bWpSCNIIBJdHyVcG9OGWGjV9qZlMH
F9eXOBleWd6lgXICq52el4Ruv5kwaKTmD/GXX74YzOiHr9LCVLCjW2d9CBLxc/PnosY4N3QRyp1L
208RIDu6gtZ9+C5cMENh4/Dnqu6HEDuSuRKU8FB+zrsen7ylXUBNBjYHdSH1wqalZySQPsQP8aqz
Fg971D/Xz3/JhzAleg8wpc7piKLdWxtzeQ7O5qGe+PFl11ruSc2CKwgITQjUNpud0dXC6RfYUIAK
n8dib43NJ+NQIlS58mg1FbAyAsysi8mgc4G4nxXHC+7gOyjo96A7wuf02cY/PH61VkhptZdJjtYu
yerbjK1iUUWksUWABmjRLJri9BhrLZDdecxlmw63Nc3L6zueWdjYmBgQCq18qvmYZ3MW1R5jknQF
NuOH+7XdBShkSn1foJXKHr305fl+UFe3a4OVuC2lnGpYu/WEq8lxIA9EJQAdkeNAhYbz/ODrdBlE
grActCNcLbwS6zx8y0iuoZtpoH/0KF0CfkMW2jaW5zLyWFwIZoiE3YvMaUFsYH1+fo74BNmdf9sg
1iMSBOmGq46OjKisSyakEFysvjpfqvqlFNBhotKLj2gLG4LssGrOC004pvWPQO8KGNrEIglRLeGC
tg6ytgBHyGkvn7rY8+U7VzWrX2ZQDl6Q4kQK+k8eLMBrZaNBO20hO1DjL7zLoZhVds1JT5J1GQEb
ssmkiJon1U7YWxZ72YuDrLtfJJryBaX7f1WlCRCffVG/gwX288K7ns+iPmUG/pYSiX0mbyEdTP1S
THbbVGd51BZYT1PhIL5TJzvQ/76iVM4P75ZKSGqtBAEo3kYi1bd4DS1IyMtmxCOana68dz7vlGcq
ZOTrj78yerVoNLxOvqEoxrlfzUuE47HUM2+hTSVKUQC0SUq1fwwmgG/jva5FuGwaOvPRQiDYBU2w
7Xdw2SpWP4ej8prSs6Iw3k3cBFIPjE74lZgB+qK/XOZQ79IFKfCn0BLhmvm0VGVAfb2M4Fzg7idC
NmYDTly/3ERv0gUsJw81oMpYKCkzFQ0qKXrpoJ0E+jwMhurg4tTE8gH+Sh419dWGsSBBcndVMfNK
i9QQkcfgPXpiLrkkNXQSnz8nfKe3VsW+hAq0D5Ahs2FQd+Mkcb5uIMdGsPubc2Dfk4ugJD9V1sZj
q8dA5VvY8FpZF9Mu/F+j8mJqkEf9Dj/vooQZE4Dydxgv4COG6x7lYE+oIsd2l8kCdm+NPzB33Go2
T4G2R0ak6KshbVX66EsEycq6zBd2Q3ZtYRgHDfopbtstzeqs87Op7HZZ//xWtnmibQKxJpZBXfwE
af6/aiCKuu8mKpt6scgNJibsgNmRmP7LwNmfyjUlaKtVpXfbgu5nFJ4i8OlSn+Ola1EiR/y7kMUZ
krGmACJDxFh2fmbnn7TPhrXTUen7yniGfgK9GETMP0nOLimnlku3h7ob2OnbgZXhbuyDtJJ1b748
on32e/kg2r1u1lq1UecHVIxi3anqkYKvgr7B/DWjouNyLE/ugebyniDEVXpJ6ZEAUh/iq1f8CXfT
qTIXIvQGMmHLAjcMXJL2dfaGHSUKxq5vfrOfviYzpbe6qafof+TTFI4O1TI4WS3l/4KGNmNK5fuB
W6bqQ0aYK4CGsgOn6eJFiu4EcCqNz7fLteQmbtbXbB6odJiy1b45N7Nzk05JsC7sSx9Hl+4Z7HK2
yVngwGw9j9hHOSEayTm/ciRcRv5Z0sdVPuhwHsWrOnSNVgSfKBuNj6YW21ChZ5iH/yCjA3t7k3Je
E9bksWzyDUg4XCEku0/GXHM5cz7bTEhzO3WNzEMFU7y3gAufInEkpaBva64sWPYLGQvnx/VjpxnN
RC7OfEwht/5qxVw7PT2Ppf2N7uUlRP52xX1uIDjoHvhqNiHFI8WpL1RBVEOmvRqPcP9QiNaZlRCY
uMEXaOm18bpPI2B3K8zCyhvWdKpodqG8aHhn4QRYe7upNMP2GsCw/XE69/Y0T6VCQVdO/8WPJ3Dt
3zja/C7WChxPh4Ph4mU38WM8EW7bM/ZnBQlkra5l7ND3r5hNt1RSNprRLMeWu9cLgXyST2Pywi/0
nuirEnLPMVZhjcm+zLHjlwFvP1df8TtOa4guZs+oi3qVO+EGEhQFjdHY6kw2dIz3NUhujMJEultc
irzTlTpJX0oIz5gN22RdQsqsOgHgAb9EAQ1L6keNZegMmu6Wjb/frAAnc3VymemtloJGkRjhNg1F
nNBaqrPJj399mIlrO8yEuWe/tWzSmGU7lKyEWxFf16blRHFejgxw6lZPjzRJyCnLnDDKGaVQqAQs
MlmzHr87oD8X2MSF+N/FqsO5tpaVB7pPYZqKwJcuIbUUo1m8UM4DmIN6MUVBYFAbynBPbTYUoT2Z
eggssTT/YIhZMkMMOXVb3VtMc6oPjlz1y/dRpEEI7EkQ47N8zsEPFFIGm4Yi6bTzii7M6gjRBIuQ
iiIhxhF3L8kj8eNfCanjp7mwpJvaiW/4qsAtWyaF3E2Hu8gtFeQqlTnV3nzf67c3uDa9u0GQ5jB3
KRlcK6HwGRDBY+MTJ2KHgEHVxCIOlyrBymfqc7XWoE5VXmXB92MmCtvM9gF6G1OGT7cVsUnyt+4H
wr+MCUXRcg0JhUUhiOR86pVwRYQDxQs9N3c3bNbxbHPcAJX8ZKRTiVy4ayTuM5ujAYPXrsfeuAG3
k/8Na/dqr0PvD8fvwENGKRxs81BoUQvQ5lV8i3QotHXVLQqfChdiXDSFNv7GWbYdvKhKzLOiVjF0
HyMOrzNK7RWZYswmN8A1cbv1Xw7oDvhaGrpUrq9cE3/WoLJUs/dVnI5L8SZe8Bfh6IFZgiuHzfKH
9bV5W0hTt7swXPh0ABL/bE4VMVrZwG3+0N7qGrTCf5tZoGjpdBM/YfB4avAn4/5qmaAlUztx2X0a
qZeqNwXUXd8sz9UVc6sPIH0vnJmneHgtLq4XAmd4sAaPxDViS+QF+DizzVO0gdX9guByQR3xa21b
VQt5lvufN1opiKl7e3MDAHqzPR1eJS1YmNa1dB/NORZRSi746hSIWY9ZY6gD0fUAT2xEpU6yhYdA
WSALBHVdRU1eBp7JNV3XnbUrspix33zKaWfxUDURohMIAYcwXQyEQOWbZB2flZo+5uQOcuHiYM1c
lwHzpQkrbhZG/XPm859FJpMbJEgkpO0G/rK1xW/UxkADgwdw6vFjwMhQEx439tZ4pm6OOF4pEEKk
HgUDmmrTBky6kOMonP6lbzUXj/tlRTFBcYNmAJMBQJme0T5WSemMvjcnzytUzo8JjMoBBsKHSwlZ
5bMy6dzR1uLxbb3u2XfYMAUpHYZQaShZL/P17ngLJRhBfKtVt4eev1IBYMCbzmnGOLDPhWVvmw5z
hRQUwF8SMbxfWEpLbyTdbPhWYkC5J8rhmtjWLawaKvxo5GiIQV3dBuExZtSpuqRe09A+fso41k+0
K/XBaM6v+mr795jpgdgxdZnBNE1ztxy69Nsvj77YtaooYedP48Y1ahElq6xmB2JOidvuDgK+Qoae
9J0+JHZPtUCy5MKdNHm5BckQQCgFB3OVCi2Kj50Ogeyc8X4EFHQEFYJZ/BZWGbvT4qb+F7p3tkVg
wNwH/p7CTMz0pH9j/XHcJCeiRWBb4m6KmcRRWfMp6hMlSmwMOrfr5w+8dRhU5xnMuWhgyUG5ejLL
Lg3Go7ZHmKri+ANc+YJc27DZCwxTdspJqcMHg4/z4TXSPd7zK/FvDOJkwPqAKkCxA5wjy0JAtI4g
fYbyX82RQXVv0u6Q7KEiPGol8qD3tT2OYoRoi0iHFEfOyYX51yx8L8aYrG4dxl46oHBjCTM0VLNX
fvGVBFdUpzaTeJomdylbA8v7fFrOSkzf9YVUwhcA4IghCWiyS+dU5dAtP3TBJGWVKop1UHSu/fkd
q8pIHgZmBpA0Cgdtm4fF+MIPvHoxSZREWyjTr7OC6R7bWoBOTANdAUHNnFQDrt/2vrIymVQSGfXb
3JUBT8NaG9PNfdswaeIgIVmd/zlM+XRsyBMjm0I5LSp/Nsc6es1zHMPdZnsxQ1/DyVzvbSjb69WK
RbJsU2rgKf2mgMhzYX/MYxKYcwsFvehsC88lXhNsi1Dq2EYMzdqY+NUifc6GQLoFmyWSv20Ku2X1
nlXY8TbjHd65mq9oIXuCMdtNmVTQgRocFKrVbNHmD/Xkj3o/mXb0abSH8AeawElSWU87fne4JHKh
4SMeplmTcdR2hQsOD4JyChoHjO/kj66ZhfCc1L8BhleE7euN/Uq3gXspRY5ltRVUzOGwQ6AEQz2W
EW3c+zKZDJI6YTP0JuPMoBBMVdBWOI0vz6lS4HN++BwkgPL5le8rrv55vNnl+ibREpwgHbnD6D5N
GMo0iYc9prUWcFh5psjQuNxGtsUWJWjdW0fNlK78R3W5dPiEa7/ztS3Ie/kNqp37jh8COUyoGLHH
FUhhqdpofRO8O0EpXm1YLYzr/ItH1JVQOmFga3DZDDCIv50SaWKi4DhEEWqBbT9X5ttOCmqTb7x/
qaY3rX8e5V+l9tiJsh5I4rvLBchPIIGnzrjVOypao8esVrEThjCZMlXJplnGCtgIbAKg/nlWi/He
5g/DmGDycGgmRtYMXoToYw9Du3Vkno3ZojCPdSZ+lW/zhV3ak5sh8+MdEFbfPU6TJpp31ngZuygS
2FratMHJH1XtCBInmcfoCCFwEhwhO8IzjngcKi7h5M65DFI6OibjRW8HCnPZyhfN8qNcpkQh3PDg
WFq6DoeFQIQqAew/hjJ+JGBOMrW5BbXfE2Vv9CoQ0HJB/Jwt9sSPcDm/uvPenxzdKmTb2wA70CWa
r4SlIilHhAhj0mVPfm88ZYWiD/sKnw8W9wggcX/G7Bki3YYAJdlEtXbnBZFBx7yMStT20z1R5auZ
kQv5lMN5MiD7XDjw5R8TB2QVFCXBuUgDoNsHA6QFkpYvIlvbSLR2nkxuOCJalXT575D1vRI1CahG
5MoS32yu5sZi1CoI4nsoh+t2yYMsO+4oXPqJt3vydHXkcZuM98hPSzQ3hhjus4FCUz5rk3E6wpDC
WF/mkGAM5UPLUTOLVFZKrKqRWGe+SELiP4KE8ItGhrVXqky3LIo20sD+4QQG3HI9CAk7A8fctsms
7/+F72cVU/1mOKHlkqs/NS3vgkki5P1KvB0RMnTij4d9R7hmOMRBJJVR2cxopmDal0fC0mv5PI5y
1BnYm7JOI3v0SFTbF0GCg9m2epQJkpK/vSbaSqX6/RX8d2myn1SPr9n6/CV5umSje3ww3evWZCAL
b1Dtrrl7XR0UqSEVsCMbg//wYazPrOUow8I/loQlDfW1eaOcf+ju7LNuB7GODi7z3IwS04CorRze
TpmNwJCAh5mFcKFEeLU7kw/H8TPLo3gMipLIN1MiRm/FNNW9AHKoON0eMn0SduPNf8XmMj+YGOPr
Bf6rL8qikbQ32koLqoIHRmNQCC4s7GzR8FE4xYqxFU3ns9Pp5fdFaGlWqE2dsg9vvY2VdmoPuhgy
nZWfk8P97j/Ul5UCOyxRnRVMlel4cQFA8l2qvgbtIfvgm8Ek2lRDUVYW88njugEeBXkgt8K0y/pk
upWZj+g7xvNhnnDSs2zTfEnXOzKHyW8aAW+23bNkUlDrHyXVYUOBHJNF4FLWM9/ER/fLSP6tBX5n
pGohGI+rOx1nR7iD2G0GPl1tCKD7nRQ/32Ftl/LuqOWOwBbFOhipO57tsaSbz90dS9S0+Bpa4nzB
zii6ATHfCF8Hu1G0Ym7O5bGO9tGDP703Wbt0cEiamvrBC1zKk4mQdZfByiOlP8VJBTDKLbLf5C/c
/TkSxdKfgx+X6MZljm5JWorJqWsbRi/NBlLdi4C+nLUjIOdcqpP3NhiZd63f468dQoPlKNp0bpJe
S32ifs+YA5NRddDeTpiUZkjyKxwJcD9sxLCfU2G6zm/vKevN8unPYFwXDksJJLTtt7tPCu8u6mj0
LVoRQHd/XEmqjFXvJpwHENKcc0PoWBDlaI0fcsGmp2zl8WT/iceNaPjnx/zf/webE0weBrvYQEDQ
O3mEoKlUuEoGSjeJYV699rxwq1xzaWaIJdRPwzpxIYY2D9qmyDKrE0s+Cp2EdSiRbOB8qfE7U7NJ
9w/bVnNbqcED3H8Zrgq6dABNma2MFqaclSNCd5uYCmAU0YiJnzUfq56aVgvP9vkjYC5NRmHQCQVi
VDaZtsv4NnVXCs26xOR8PucHONmllsiHFCerF8JBRW8kWPZFUSevh+pIX3bGjFWA1/OQRHPt0dFK
auYHfY8VjVnK1EjAeK/IX1waQMwHQpGv8lGEyqST/FlvoQ2YfPXZ44n5/4HjB7QAOjZSn6FvYqzM
C3Pefjsa1jdIgr1LQpGH7tY41XRNwLc6FTvTBhXcW/Ecq2JQXlOjHIjTNSU56DDcrfVoh6DCqKUo
1RHdjhJ5lZIMg2j7vf130ruEj0c6fW5waMnwCgs6tLgStkbyX55ElPmRIkAtvFLmU8N77EikO/Z5
giil1F60DUi8RAdBEtHV8lbj+A1zV6sbQSL+FFwbsY0Wb1kCGp6SkuUNfv7tGhWseVBvtfjL5kdb
ucPHUrBwoS+vJb7XrzOQata9nCNvAza+3wiF9gulZWC0Z6xc8hrx2VA+7YBD8Y5VvlspOkrdZ+ir
aKlq8PmJEWy4koNJFakNlTktY+VBrB2f6h3tNPZW2qhRK6uBO+/vA3KAM8KQPtJB0pQokcLfUpvZ
oNTU1IXjCBnGRQ3JW48tMYsCsKbhHQJxU3Pq0u06qp0V4u1JL+rj3rv0e6BeY/9lvlnOnhHGDQbb
3LEnh1BOxZ7cldA/yqYTgWGpVIwThbtkHvbNnPGGHKkUOLJ2ybHakPxSceSL5PpbYHlY6DNG61si
Fq/W9LKYkRrm6tPq2hm4bbLYwcCCdiMvP2TyO80HFvxjvdw/tcRz7nVsn7wmd1E+Of55j9g+dQ7U
om7901Ce3Ki5OpYtFDW2b+YX4bl9BUhH8LfpwpHauvT2RqLBi433P/zJA3wQHDIxNvLv2suYXrYH
PWrxMze+CWcKOBUtIea6F7BrkL9MWhK9YACvxHz2G6mhroR4I2ocC17y5n2ZQHuo+MnLc6lapUIJ
WCkIqdX2uRjphqtPItKDHxloJTGvZ6hKVSn6IWugqoIuMdIoJXA2HfaU/X2LE+vUKA91n+Ps0TrL
qHm/UxwejBQrCNw3a2OynrdlsgvzyT8RqoNBRGHPgdewwgOnqxCJvdc3DMCl9XyGl56CfCoENNOQ
nOoaaYsqPKNEvjmR4Mffrc1UjBs2pE231m1cEdJGGcunj6ODyDRgEtywh6fI9uEIg0sruZ+WTCRh
q4cYEXg75o5ldP9UhOWz9UH9NeXZ0DOkRnkVo5Ct6XmI6koOwTfpYp6b43XmzCWxzvLbsN3g98i7
BCrLyD1GXmYjij/vrxYKN6FgHcdwh5vYQvpdfctGxzGF07BQsL27UcXi0QIGdbUz9NrwanSUTbG+
gynnbjj2uQxb7y8JzP428jx+EJ5KBxRYvZczoLzANraasYCArpijk/RbeWYHQZrq+GeGh+AB4Q38
7c1pR3lJhP/mgVHYAXzFxigMkgmuAZsJB9bkpPkh4ibJTrYek8r1kr07VDSMLL682NSnmxwjlPsE
z08seyismhNxGoBCct7kqtywh4v2zXrUCzHGLkOrwH9vqmlJWRLIVRnwQwA9y3vBsldcu8FS8IqC
ORDGlEeZgLxyAyssYPYFp1RPuikyVUPuuXW9UuHy8o4mU9ojkP/RtlVmRtU4CxqQ7YlkLVcauer4
uTR5T/PgOF6Y9Z0A5ANsi0FXrclfwWiRpTysupV5egwzeXAyeIS6VdWaPiLQETPZUflbVBlUeDw1
t4042M82bOXa+PFgyEAnRl1TxKVawJ6cMdF0T04DkoBmYyUdOvKYDuDmN1IVBh/VfQtjn6NowVAX
ePyHZ05oX7Havyz3X3qCd1RWhJsPVP+nFvrNWX3U1bY7JK80M+MZeuPjbxnmHmS9SUoacvhpRAN/
r28K91VneGSMeO2T/RQaVVvm+kCKncIkD7JjPKDSX+c1A+LcN1poIvghfgk76e52myVa8yyaLup9
yYP2X7kFNg/xmpds1mCTq6mP4Xc8y0V+0G09ff6GtOdM3Jho98q04lPfRhzdaS5YpZ4rJdQcqQMy
DjkgrAFftAyzmUusfAYlmD2VFHlPpyCAFcHAyApXk4kbUiep/Kt1VG5+k8c8k2XgisS81c0okslB
lwK0j1THferpWmDNRCx1XA292XFknE9WVS79fuJXdjUDg8e5MOKeqyyMc2kDvMIJtQ2Xa2MAQRwi
SgkNhhEV0WGhQXvL31GCm4y/Kw0W+KMo2TRH+4cNj17QqwQhvpTgfPEi9IhHCEwOhgrSfvggGOKB
1LiqfLTj7js4IYZGp4MHRZYzkFKMHwkQjTkkqf6xiGuez8+KJPTre+3yKXDTDCaWt1wLZtHghLKG
BBXxQNnizLYjJ+m+oGhFFtSL/JRxFBkZu9pazgXyyYuN/vxXM7YIYmEHNkfjHu36bUjtW90NsCFe
klNs/HLNHTq1DpuSOnKC6C8zvxe2h1VxlAn04ND/gOx7ft/pVQaf6B8D83taWMBYJbY6odScxXUq
sVzMRthisowjHnZVr9ZkffrNmKki4df6Yj8u+lhiNwl9HESDmUvmFY4WQLrbNIvJ5c6Ic6SBY6M+
dQ4NmZSsosaaxiaytYIJFKUlfD8NrSBzR3L5TeAINFjf7o4vhMVu7W/uWNRDWnKECJQ+LHYZ+hBh
LHsMLtthDmgar+jX6A82BbVsNTttOK8YJTjGP9jeyWpe3vjc+M2h7x+KJZ9iWtl6qpl+u7byr2JI
rBgOdYR5ARaED0gr/9rejzijPypRD85B8V7CEHS4kpTlQGyc0JQDlM8imTTvKjrcuJ9rohbP191B
/tqtRqBF/MIZUOM0h45nBkeIdzOnTANiiGrkG7VucDgi6MFf/ilBIYwERigZKmg4C3eOwn6vNGJm
H7kp7uNnBsnXVI3Ig/prct5CHpXblYS0ivLttx/tT8vEuifqi+ih6ujx0H6NUo3FAcUluaEJXL74
bvy0xbpD5Sz+VBOg1//x4KCJ3KRD/6jhxxFwDZi2g0JoYAlNhMAyv1aeuID4u6n5+TRT4tyalJA/
1Fg6zZqUgzPL2vNL+C6+capY2Gr7Kaz6KRqzeDsjFmAZgwRVnJz6YUS1V52DQd8f5jEk0bSM9d56
m8l1JjQGmWaC1OJ7knb59QQ/3RxV0k+92Rt5JlQBHIxFaCstkOZYYW1iJKdJ5u2URuVSG9hnb+4N
FoesfO9mPAenI7/pVBoDhbdlXIyPTbWybKDrp+07uXEOknCSdNpYX8R+Zsd2yJnjht1GcieTUGlc
lVD7s5gNwu/2RpKmj2F5H3BOe5xsT7Xarxqve0ZtRKmHAAx8udrL1G6TTRy60thhmA5Hs2uI77oj
YJckiBlm0LqYKwYQD0t3yDIaF7JbMlLSe7fMUwT3lL1k1WorMLupUuPv6mtnxLereGSIL3z/VCwn
5WqMH6FJji0veKcz9yGVoGTE3grhyBMz8glQ1zztILkkE9vscbLS4Mj+XPNALDN8a6YuI34Gk+vF
XuteZhOJcsvaDHlgZhFT7Zl1hTvW773+JTO1kG+Ymk4ughurG2R84T2RuRJV4BRzJdZFFtKBcAhX
VPah/+PhcBkN2wDc45paEOt97qxUgWHFSVEQZmBTbvmXtgOs8nEbegrgCWygWD1O4O24zyTcIvf5
Ja3nC4TomCcaXkIAnNfXioBB2tgx6XFSvIqDo637j4KwQHYHTJBeTvqsWc8T80r3Loq7S0uwCLDW
5NBjkdg0xYHOXzhTD0Poi8OeS8P0F9YSTCweTzsIT72oMZ/Q0PzBY9MTlQ1X6GAABNev/m8GPAjv
q9E6L3N3j78Y8a8dS5du5dIjfPgT9QOUm3OSZqILYjZr44f50Ohx6aL2OgUt3n/zERHVpEobiJPw
HJG9cWRbRcNNrCzjbNr/Yf2UimJ6hErwU8vMvsTQj4wDo5FS5FnFJwULbwQ8Pzx/nM0lnj5nQ0/C
m9kqJEv2vBWFtrS1h8jj4A1VIvlC5TS3s1ozrAKorIVcCyKRtnVS6rXU69nAHrlfIK1G7Vg2Yfyq
dmEvlOHP9i6HtYppV77UoW2GR2uvaKkHtYE7PyIlVz1yu90jmi48QAX76cH13Jncagz5L31GF12w
dYdbtg/VsRb88gTCyZ3OA4q2SkXr89G8Nh+cChrzwYGK2Pmzp8vnBlAOGDLK/OdXbHrrGnHCht2y
rG59Fq4KPyYPKCmld1p8xDlZNU6uWoD315v0CBreR9Sy5Pbt3Ufk7VYFIqV9dxBwscNH02KBas6R
iXEpz3Fe520IPGnKdI7omU9fb+lY45H+W/kneHq4wYk9gx8UdvCXapBMEUPnIxdJvAJ0F42XBtTL
eaiJ4Yo2pdxhSQpNHgC3pu6OpogijO3Y2coYeNpnwd8XKoEDgf/8of2VVKHc/irgk9fL4jY8tMot
JXHiRVuLhE/vsOOYpXsNsNZ+xpJdIs7pGS9c9+KeFAOtdMKThtHIUYvxQi6K+dfLlOCdnDpM+SJ7
PgQQBtAHYbb7HQV61wRLnJVSaalHy/XMSbw2zxd4kITlYWHL4D+tlrQFjGtQIUf3m09EHOPxgPl1
qjvTKmeWZtj9dopp8Rna3LMW3zGGEu8lZeeYEI5ubiKQP2xEVbJChahuFK4221ZAvezcpzRjsfJe
+CBsvVzU9e8jsfIuW7c2YAm009MaoPsIZWSqRE4cxzYAa9tUyvtyEot1MHix/v3E4Gt+8ZGyoYyX
aAppJ3alPp4GVaoOQBXLJ5CyRMTV2Fu9Ht/rPkHnTkMD6dx89k9y0gmY4FBbBsdf3xgzXo6ZGRwA
v4C2x5g2e7sDm8BfToJPh2hmK/atB5nvHdi61tC+OHed1ecuu2pkk9innUA1St7DWn4R2AsdgkJe
VXCg5shstYSV9ld0k9B2Xd9hZc0TXGzVQ7IW2iYNBWwo5FbKkQEx/CrCSfzoPvWQVbyd4+SvspLg
8xtD04682BjO5HUEwI6EnjR/fi/6CsOS8yYt7fYngj/qHS/Qf0I21+sEJtT08FguxsDGCxYablNl
I0Irxjpj+x8OvI42hMPBYos0s8giJH5NxAcKHCldCHmxpON/mPwpmNMKCnmTg/wJCn1bt28mB4vW
4gYq8Bzw3xBK/3HRf7mhguHJxN7gxsPWk27/E/t1bfiWPtwrv7CQNq3MXnXSuetghMOz0D4RaX3+
nNfEGVu/0MmcFTIeSic+90lFbR3Q7gw0tjVGX45FqgehwZJGdLdZsJ4U7XCtfSymXsI9CxIv9UC+
g5z/MVm1/SV4FwRprSfDhtbehBMdUQZLxgsrqWNugNx/HunUUvD3jiWgbPz865jIgExd413mosOz
GXjxyqw2mDpRuVohVUTueF3UW4KKR/yCNwhMJcrXqZgOiFEEK7pTNM+QitCnB7TtGSxisXi+yKSO
XdoEHrqLI74TuBS3GoyKd9C1qdA86latuLfFrP1+T9sdHEdQX2HAanEtLiABbW8gyNHpGMB6zwAg
BtVaULqeNO5NRwk0Fnh+5mdzUewhYnTJvLKFiYQlhGGm8GD9vhjnQ3uZcV54JYw371xWtZj8A8Ud
oloyKWcqHmOpYn+ervo9cBCMsbMvfV/tQ0QVI0uiDWyryF8/pEB6lY88hOPctLcKLNkdSLs0UVKx
2byYObxJdHRH5DMpp+bspp/V85xI1NPBf0reVjtMIDGw8duH328cJPccr4uyB+SHwPS4o2vbZ9Bd
RbNVZVf57aZrTvYy8YpieCLh3mPEZcT9aSyNzlSsstPX4166oUaAWQwinSXrNR6eBv48xyInX4SG
5mpU9hrqIWpgdS/kNe1asYUh7WkQutnBQCCqI7b2WpSi8y6EAg7QQiFSW7GbWbfHlER4wgzFcGTM
heMVrtUEv/Y3oOFS0h8kZlxiE2ZP0jGkr7Dpci2F1Vg0IP/OR7nJYT6dJ2bAAJML0o+Zi+5xZpdV
i5aYV9kICqyLfyRA5Y58JM2lTA182r5zMdm4Retn138It7+NdaMNKnF4EVIEdYIYD6CoSHxe5Q9X
aeTSg4KooTnz2v+AFe7oMdw3xJSu+2Muoa2zBfOBU3ySPU+QQkviojZJg41n6G5YKKezUNJDjJl9
GkOKX6pmwC+vUIs076MHawgO2w26OcSIbKr4tXxayqRuu3vZoVKfj3B7xfV504knMGWHOaUIa7GG
2hHSUiATekCBHtRF5iv3+cNydHKx9r3Nl7dDEWQrhf+b24lYkGpd8nvGM4+SilBez3nN0EhNr6ke
uq0PJjXuQ+htPmUSSdQC8OnhXaouazhto69q+aPGxVzn2AzHoqRCfkad5aCGlRgS7KOz94m6RaUs
fXvWuMeRQu8HtYURuSHF1ayulQ3i2GNZTtMXVpuRERWxIcx8r1Q/K0PpyYZK9B75UcBtmsdMFIrm
7pU8evJlshuZKPo0FzWsjGXnR2I1sWEKT+OQcsK473Z7Y538ZBZEc3wCSre2XZWdi48lTYf0sAxU
UuW/CG341hoOu0Ev7Sz85AqQK89soBURsEPJ2drB+u7VfyTCVSF61nscqKaiZ7lovSF/AXYQ9DKz
t8r8O6kbuJRJqHXgaXQp8Ke9Z3imzi8aMvoJ/3eC1MR3XvunTzCHNnU3foiApMf74lW6TAJad8Xy
tKOqYsdWuTfBeHJoL5oT1DXR6lOfR7HsvwjAyTapiutb22suky91Pkc0T+87hNHYQ+O+OKW+gjJV
0vkBe1Z39TaLO7C35zowoQ2S/m7TcQdvv/hPaU+Yi8n9XYNpk8MeCTtJHyNDHtTdPtnu5AB4YtI7
vhudGLYV7qbJGpXU/xjGwOEKVCJWZW7W9rh5y3r8kOuiaXh2l9BRgJWEY7tETWWkIgsUjT9isBP9
x2j2SYmSgCnRUrsjQ/e5roLqZ/zOaGLPuhSDUXxm4CdwoRoA+pssVwrWWJEJAQkaDoGjEulEYTrC
UeNnL2gjcrGwEvwwrlQ4Bck0rNKVO2hOPcr9tKQflwbqUzSwGlHWeDzqONwG1ba0g7qBpbSoKIvv
pC6KlxJp3KeD1g1xab8CM7tMUNLn6I59AwfsTZeFMhq+2p7ncysA+LunYkjHvup2+l2xfNEhTWlt
gM+nTnl/Wndkz01Ik+0XcbdA0VKn3l8QV9bhFy+iW2ly4N+WQcKCQuPBIcLZYdmdRMrZ9SYu5o+/
/o+ngWvRt+/96EHSxKgwHILmgNGHYzs4LW7Pkz4xr/IVkmQbajws4ZcelrThlxDOBVb4/ZZY4cct
qaw8OlX14nge4M0gqKpI2VETxFDO1ehDxBFD+bBzhkmtKLUembmWxvIp0Re51/unwcBnlRh4UmAQ
rQ0jrUjpM2Ug3NIDgXTDmySdZHyRJ31x4ys2hDKcAL3tSj/ekU5YnsobKcEbX+8amxJ9xAlkzK2Z
ofQlTTh0pzPhF+b2yZDmTbbma0wGuzbb0VN5Gz6xEBr6oXBMdHetMZTtf9onB0wAT+H7oy1o5xZC
i8yWW73mXJ+kSAEuqaPuAiookKuEEqd3QzrUrmrJ/xl9WsAQVgFUH6C+0aeWHPNgk9o/pugzKxxB
tZoh3d4tz7JQTxTy8OvFNz/fNP4oSQfW+yhAlk52hNz4+7eA7/4nfF1GlM6RF5Qk4vSdrif6jaeK
1KGN0smBSc8N3wqcm4Fuw46m91ZonTLLvVccvK/r8gtXZj+Q48kxuJdPk8Z+ZM/AJlSgveYXC4W3
bIbKwAfl8OPFp98AWD5z4ZyWY6ouIS94EDgqcKcaBvHghxWs8atsvhx7mB88qCn5En3onwiBAR+Z
fn5r6vA7LeF7DFYLlizjKDI3W2APAyAPX15PoS4uRLm0tEiFwoPGPngn2F3QXe0GSU8SJesjLMsY
oOlLIHqcG/lgLN5ZY52/BUssCNUZYjdFibs5aWwz06KlYknDfGyuOuOpeXn0+uXc2UQbl0fZS/wC
wF7RbzIMwwUd9WPWuPIeMS5eZyC3JARE1uCFCF9leepojhKJZqT47oNBTcR/I6onh7DdoFxAeWCB
IPZtNnoZZY7uRQlqoWXo7hwB8gP9kT1BPDR+rwpra2Qed9XlsPirttPTdI0oQapCasN80m23TRWw
/AU6zl5Q9JWeKHE+vNoCyxihMYI7VVGQTp/ny0uflviL/R9IzC257V7a7ZKb3SYypzH2R1AfaaLm
JToMPrTWR+8W7K7sg/viAIQVMi4OCgZ8Tl9FljM74VY3E3dfLQxafRT9MdjHpYZlhw4pZR3PZ33n
Xl4okR/dQUrfdTCY6A/VGmo4FIQn5iSAZDIjIV763VJwD5qtKouvI6RVR6bv5Zk4J7+9w/X+B7rg
AQ20RHUt7CAwaEpwMBtMTvydYuLSdOYm6X/3FZnnocw7ahEK63skmuVmsPob/lc4ONu2i/994JGW
lfPG+c5ETSCpXJ8G8zpcZkEPYMa9xotw2lXxyHrEODaWc0Q9c6NVGepRNQkuLC5DuCeiKf85o894
a+vRXr3w67OoEonrhot1ahkcs0ZE6Kldq6nhglHgi30/LOj9EFI15bKLs/Yl3FMFfQ47Lg5KMuis
N+pWIZkWCDEAPKObd2xy06mNoCDE37vpWRl3HYsh0l5saI6DskogTtBTjZHXwLuvAJhGsQc80Vzp
n/l6fUd3AeHircaze/jwreh2cGRrJCc85zPQOckw0VPLQKIbqkKRxr20KCkFYIkDtPhx+sHM6mYx
qRsev9FXhi9CurT2yTbNYn139QM7iupW7C9exh+FYXyS/2iWeCzfeGvWjgPXRSaXkCbl2MLUvW7a
1CAGSGyoEJhI3sweQQ/DJPhP33h7EihCki96jDTZp65N7a83zsxQJkgCIxO6cUOdZzi3KgdMBKxM
8HTqRMHGRA470VBrtmj23GWQeFYcK4aG5Xnr9P6l82COyT1BIIGZenpSR3T+Q26IDfKfgMlvWVfI
y2bijBzi91I2StIDonf+Bvtran33V7yIPaC1b8QOoeaU8jXUt4nLVz5FI6BdsFqM3iffk0oP4S2t
fdgVtGyQfL2uZ0t0qaVIjRysOQmest6Z/VCy7qXB+X1vq9cat+7dUzvy3h99KCMRMOtXAn5p+bw7
M9H/ofasdvWUVfJ3WAzjNuk5BTXtf47tw78pFHtXSQCz9Tk6XsLUm8Vacm8COPKQDl2uPCagUngD
chhFERoGD6ZYXyEGO/B/GG3GBYgsTeX8Byc1rJgVvBGoYe61SdwYkj5N0NEx2ggzTEYakm7HeBDA
CbgvWchq6xrUorWPXFQEXaTE5ZQgOpRo3uEEUBFM/7mB9p+Cir087GEl1OTsKEA4IAXoZEJZwjIG
9LtCW41U2UK4g7HiHVi1FQ2306TcSqKnCzeSG3YWCUdX9T14BwwOz2IGK7KIEWZLIPTGeEIb7MgW
DDzC4vIWHCa3cOTOlWpvPGsQ7wT8fO3ZA9isN+3+J1ySLzfjWWUMIHy3Twm+vTzRhLN9CgdCo95b
X2FMrkqW9FINHt3jilrvcgSTUtNk7rsChRn108jhhVNBwlnZC6r0rxq/mv5JI/tYTNVRYsgojSY3
45B2Vslgqvzr1ot/7c78baPr1HD0ZeedFeKvH5zeJn/CVnSopPcZWGR9hrZvHyBfB1VTGOUSw+Fv
tt3pAcsLROoKDhUeeIunF1ro6jQ+8kc9lYAGDirUZRX6fNvDmE5lg+wc+OohF6hZcpjLs0zW0hdq
xu5dCl8Vo281WT1+QpxIRcPQrD4ZAkFD3UtTRrMvBgZWDhUBVJGPNRv1AYiastMt5UQvnt6+Oz/g
T9Ty+mSnKESFUzxf5DMZC2VAR0FJZFxz0IUqSjPJ4GvCQi/xD/G4VvJkJtfJsAvJNc2nOibTxBwV
fvwpwX43GKH5ZY+6dDh6FAicc4/fTPfYY+BY9IjfN6gZDFlIobqUEpkeyR9mXlSDHU5a30SmyUTe
wVLElDpYjDBSPGUR6+ZP0Ecsm3yvp6vD7y+mYaYKTtEp8Y5k+z3o4BtgrpQiOo2Q9O3zHxvQQKhQ
V3sIHpnu4fw9yVqzNiAlYO0hzuLzIxdC1ZW96FStaD0UA5v7udiHjDmKINt7kfsHbHog3mxrwYng
xY3xB5CT7aPTvZAEJWtrf/X2mHtjNZ57hX9lIKUsCwGksY2/0ObBbBfEpG1W5ecGYmasyIZ4UHR5
ncV8REHFAfQzq2lXxkxpWuHJFoG7m/oQCo7IqtEwB1BR6ZRlpwiI1YewQPKsugFrGoo0iA+H6Ci3
UROcpiqOZhabdV95FEH0v6+6+nHWtraYlHdKtUctqpuE3uxuoGBfq6lTNER+xnJdKklbZiDZ6vVH
EY33PX8jxgWPqYJXCX08VRXw/YLU1QRvvz21DDQXZZmgKUuXa9ExrAYyz8VPi49lGlif0jvdRtfR
i622zwVN9BVq7SsmEgfGMV2ve4ZeMc0oIlvxr2C3IjEFLG9SyvFM+UjY3kzszBev1Cs/9Z1tyUk4
mwPRkTEKjUKvMK3dml9D8xEJmt0d+4q4pgrGGsHLa8VTtiKdWmF8KExmOM0Shk4OBTrYLCKo4Rsc
W+oeoDNQxLrgWxYEXMNAH2BHT21gn1XvVK9rfqtS+GpyNFC27psjcHgLpd/1JvdNuFb6jfOu3aAu
1uiFl8OfoC8Aatwi8/ip0EgUTCdk4EHB0WWHWVRLXMlYtB49+9mnPHXTzqXWsMVciPNGlcql3m28
LwFXdf40J5/SzhB5TvqQ9n0XbbNMwj004od95vvRYFnhQpA8NAZeTjSuAS7hgJXklwfmZ0k+6YK6
Ruz/XwC2G4YaMLf4YNcXP551A2EZ9F4skNt+OFHtg+9eqE2ifMJRmt2/AqJ3QOUOmL3R0KETrbOR
dfOCEcUMClq2UUohEBvRCAQvVWS33pwWenxbRtaIflwtZZnWyGlLqtuzySsf/MMtThSNpFNlVu3O
pApCK/IzJjJgDsUCZHRppluWwY/Ghasf477MX7QpwdIzhftZM88gsF8OxNmE/128rWkKOyFH0JLZ
JBGpbG1krqRwTeO5FmjCnhSqEAdR1rV5jOnzZ8uwME/pBZsxI6A4NXaPjvj09LMm9YpW1MIceE1X
uJ9M7010/I7t2V3dflRmExnv/yfN6n5lFL6JmwXJ41+9fInDxC+vfw3sUL4EQHaDju9ntc0qIbgC
pswXGK+xPqfNn+Pt4CdJ3pcXQcsuJJDU42u15Lmxv2cDN9xJ+1GIzawmL4zti/DA1eNWtQHtQRsb
c/d5++vfBP2JVEYqS1zzXQUYUvPVZXeuiUuyiF3j/DvrShnOT+3/rA5ugeRuwjU/4peYSowNEIpD
IP4dmTn7p1PZZr6BBrqz5M/AxmUQxBfT1Gui8DUZRjHBl65wKo0svRlZkqn32yCYd/Nccp24Pv9Y
lHTIJLTy544YC+3OckWxYf50UzgEUosNArkWEf7ybo/3Fq7/ruYYylDaD64Xkt1tmqn3gHwj7we0
swn4pks6E4RkLp3QUiVyZW6lno6WTQnii12aE+sQrpBHdrth9LmmC9bDqmgRH0uaJO8c+kVKFzPc
u9wD70CgZ4JuWDTOJXfSW0uKOKgRK4miTc30rnR+duT6LGaSBlV4Gi4IwDalzIJj0bdC4L3hHgYu
I/ifIDy60Usld7gNEXdvAqArYeYhswPzrydLlOSDZqtfbtMiaOeqZR9FwLB2Yz9rZpAaun2clrU6
N6CEZngXwtKZxrsvIG5qpPYNDesfGg47ZKUe04ltsFLbXvSAI+l9P3vTlJUWcpTOlTFTTIH6yT3s
lhl5fI7uAflhlyAL6G243S5CHYCj83Z8VCc8DhPrh/Z3lRjjLEsrLu5RpLFW1Sgj47aXqZA4eaLa
WxuJIEB88KOOBPDzeLJ3yy2B4ilPs6OBuy86hExB672NJQ/A7Qvlh4XoRg+NvtPRXmnYCUm2Bw+k
uvPYk2ztiV85/3KVgtVtXfa1vRhQmHptZaobYp5YuLqSO6wB3xPJL/05QDJKOkCk0rl9CjhuCrau
xJePxQS3WDvXMK3tRClSwjDafk4COKX60rKnYcEXaTPG+ZQ9VYJ1d6aHtHoVLMYonkD0zK9cDsiY
7fiFCDjMrn1LswT70jNZx/ylf+35C2YYUIXOwEppfP2UaSPQd+pyU/AerSowUEMIsPM7ezxBvbtr
qQ9QzX23CR8r4nAt6AGM+/psjmN/+rhIFBxM9+Z8zp9HvfcQ5B1hDK4jy7NAkFUmirH9GXEA0Fq6
L9cb2KH3+1p134+cdf2EIBVOLOuKcdIMGC+M6bQz/FBiDBevjg4l8++6sH3l1v8ok97tmJOXCETJ
8K5u+L2ZUgCeHIv3kUWuL6o7rIMN/psTrkmITIh7utzwiFEavozg++eZUr/F6R+5uMf4ZzT+AMg6
Lfe+ruXEgH8zrDwhpH1J6gXM+n8gL4K1S7RrKG8roaTif+5eyiU6Nfu8B2gfAZ2bMRY3MoJu3wYM
hpb+6Ij/FhtUDlVCY0HVF1glG8FJS17y8PhaflE7rE/bjAJJklzCljwpW0oQE5kEMYbqL2oaqEAd
5z8EZX3O5vA/dTVMhKshjYbKtTkg+PbGKmKCEZRLaI25vmweF65UJes7w1KjeRNXDqBqSJqSprLu
IXdBIQuize2oj0A2ogBIcinYWn5JlmlOrMBY/EuzOS0yGpx4SLAM9BYK+r0ibISXwh9ewf4ujKAg
BktEX3e7x84bou8e65+zVUqiqSd3+CTGdsmpgos/mIlVqDUiCj3PnLOO1vhmGa4t62sP1en7CHkU
A36JpTlVIEl+6y/wyJWn25bi+tn5rcTkN5h4iuGBsKSKIZeky34E6hXT4zXWJoxnyRI1ad3YJBug
kK3HcPBFYzejym1cykDiau+b+KvyQvfUK3Pw18rBy2xX1e+wyoTLI6VLHweCrFx+fU9vD9qOv/UQ
JXUcwdQOU3aGHFN8N5azGCh5FE67FKPoYtd8Ay4l5HdD5RZk01g/EKnEtukhemUtTxTPQ2eGAYK6
nIywhHkoMnqTgth59M3psIzbwq57OdUfN21sgP1lT6btGQ9XvWUWQJPAxaWG/KbVUcW0CeTlomk2
VAmVU5J6cOMvV488J7+A/zYchIw/eoFcsnrSaiJssyMvQkW6CuaUO3yKPZFG9PnOz0kzWfdi/SUu
e7shd/D8PLxAoGYSoswBeLARvOssqeqkNtd/vBXDdzTLZmJzXJsDdRDip4cU+mQL2rALTIy6cPeV
zKYV4a6F++9WaaAtcmT2lyF3FAW8Fk8tuFoBFFd/CXMDqQtlwO5qwWGmbX3oAQvmP00UbqVsHqks
IL2JLWZVf1mxFsyatW1QMAI+0z9+hCRHy2ob4R6vHcjIDv1CL03NuoquINgvgn+iHE7yt2DWH5yB
tKsFx6Xf1uU0r4MfKxAjpkoGUgkX2b48FWFTbcdVnHEs4xMk1c7sQPc5i7ZMMEHwi6IoUa+VVgxQ
06ChI0Q/9DuUVByiUs9tlYfDD9gpeZQwQvrh9w57DCZikWkjl7acSAlewhNQRhun3xLPcSqigua3
7TGdrfe8XQHTduLqikstj1WXVm7jtOogVNtyfs1gJ835Fv3wiAp5Rk/Op2rfynBxJeKmMXJC35fM
8huLGcEbI1kkGUlEfeHHYF8BIu/4lXKayWvWP00RzaBqWxarzWr/tD8u1dqWmTz3XmZqpeP8hOCz
oW5vowueN+QW1NHPfO1tjwGcGZl59omMdy3VItGe9r3ALfJzr8U75DWXql+1Tfh6eNe9ZN4kRcXR
PmY6K4drTtDzKEeB6ucM2NBPAXuoqJQ2cyVQRKWTTle7qbFNxQRs2ZmQuN72/zYFnuH0d+xNd3Dd
XtH6dd6xpwZHdiKYR7kOcTTQRoxqfj1ZzbBcwJwkT/yHP22z6kE4QCgyeoKA4HCjk4tFjmb057xX
zWultMqSc9FLHKV8lA2OB4jtz3LDG0rPTrRFo/wlgKpAHh5uuvMl1owgQKKq0AXmzrJ2unFojbXP
uICowyKBGNAvTm6oC5etWVM1GXmB6E6xNjxNKPFTvfMEJJd5WfupmCz+comfkSZMU5vBZy46DYM0
sE0+NFJkrZxwO0EmobqoUFFJicwhmIsgNuwoJa4+0jPynahPt8AxvfrFHLPHWfQiA4Nj5/2BSYuW
yYcUtA50vJL8O5SZWao+Z89lxWJvl4Cy1CNhgCIzs0BosD9F9cQI1OPyHtBd6rcsVZ5ZkViH+Q9j
+1/y9zn99kdP9EEfcNc7l69QD63jV+FOYRMzLwNcqi7eFzvDbVSRjs3utnyZ4ClbwZNh4rzs0wVY
ZMDQxiHMyTFdjyW+/uPWqtNhKk2Uj55CFXaPNJxmXLJaJ0i3vnBzXomaaJHHebqj1yfKg1SMgrSM
ddjMpe06Q5dguv2jxWm9BQVJ736sNPaPKh/DfES1Bhvx2ZJEliPxhSQkuKLxRsJgQONcvqxdCMjY
wW/poh2Fyt15AGBCgxpJ7GP5Og041PM8N2KyT3YeYADUsJsg8j1j3IP2Z5/oNGDBiiMLA5F6wFKu
99EXo3EeTcyDEyI+pIxmCw5et1l7WtGCyPuI/POFbzgrAej41MCK1OLy0y/Ed+13svjduAgkYFMj
RVPzaCZtyqYrsRyEJRL9+NdhoSQQzx6olDxl82hNdHtakh2b/+gIgEPKg4/GzOC0mavK7voVq5Mu
AV0Km5fXa6ZYFP5iKDyE7TLWSo7/L1Zvp1+Q2zyxyWtN7EnEF/zYEBRZ3o8DVxiKptxte/KbtR3t
xfuKN4zt3uNEWYQar4noGFgb8v+k9+j5JzLh1mm7S8NVR9iwy9v+cvs0seAEq8kzOzLvC7+uGRC+
NLwwDdxuGmSG7pK2u6keT7SgBJLiNtn9RQBJ6Dv+lv73BT70nMPK9plQUwyyqbBAHHANQS/vpt3E
xKdmwNHODXIfhYXmudr6NfhBvWEVFE+m2eEvpeW9eUixNeuVATvZy4uOJMAUQOwKNqnT8YxcJXxt
h2ywCi4cnJAGDa9iu5cF/PkwwYc2O1HOB+5SQjfuEnQ5AAQfFlhaQjSEMx0UMTwccXK6qQTQ6x3N
TqEr9r8yuj88kJnDVuiozFRkdL6MhJUDpQ2HhHYJeZiJg/03usLlRyCuMW7YGA/kALVoJYCgWMK9
a6Izt255MQ6H0FoSfNDkrXDdN2ep89CbBm0tEJphWwXJ5nkIWfZZbErB6dW3rrZt8t+6J5tkSMKa
YCGsqJwfOh44xhdwt3JbfVu2XI0u5cEOthkOetRSnJv2GAihVywtX5KwxanCoVFiyBXQatptKd89
IpwtIMVCFYZUXtMY5saaSkmMbtq3TMZGkeKJ9EFA6XJH78oH3RnIgEqqp7KUJGeJIjBw5c3/jkDZ
tfmlM2al7XB4F+Sb2E/c326Z1PUYrLevbODo+S9BiG8UQAE21pB2nlRChW4OvdoWeW//vBPFi0LX
S6QYnBr99ldaVsZVR7uaGoGweeso23d1Xo1MwP/vXU2p4olCi8N5FWnSdu6LZJ0FrlHXSjShLLRP
0AsoALwiCqnlOKtHs/Gz6oymdYlVuNiT/WnibeVzDsVgUklxhyUpc8VfvadoxuonuyWJ5RJ/zVon
r9QNPOMyusbhe/smDhFGDMqHIMycjWUC+9N25rURgIYs3HiQi53V/v98QYXNmqSWH2i+5ZKs53lz
wVQW0aTz0+As5zHOtjZzqGPhlgo+3oaWKhAwgmxyQAcdPGjbtTKr2rae6jtwusm70zuXlu9giFdY
mMLu5Ycwtxfcu+7+DiGZ3ws4pdX18tMc9XtIzCKbIUYkCVMx6Ep6vsvjLqDIEvADMh+JtMfofiWk
i0lnxec8H8H6sZbznAlrL/nBWZR//PzDp5B8FzPI5Znq6wA/TyefhkMScUt5ZcT1ZpXA2+PSP/QU
s/buhc+qBMH5sZUIvCQvlEeZqPMRrYtn/JceLo4nwY0uXlWGIbr1JINTpw7UNZf8htpqdNJhM7Tk
RhVB8oSd2hhO7nT6yblc6fNCG4pjiwiNVwvXLN/xJYZhJKBX4MWQeKmG5tjaQG93eTW4OjZrupgM
ODTKGa/KFcyrCpaXSUXJIwTVpx8uTUByxN0MYp7Cd+s+bsyNCg4PyWxW7ynacF3GlLgBw/aV1xUt
l68D0yoNskOBfAXfb98t6Z6d4+ZYQvrHFzx6nPcqn5nIjTgggRKrn1m/iV/lC6QnGmtuX6ptBuqu
g0Sofq9BpfZGtyLjJ5n35CUiK+ZWD35dp5gYn1BCoDo6+I/uJJ5VIFVp/kLVowyxbtHm0JLPIbF3
12B5WMZruvdO6AQ2oz8ALXKNtr/DWpdCKpyRjrpkav6oK2tuxkFXPUgoljrY0YA6XNNVMO9bRoZU
iEaHLNwmmM/iv9/WgLz3kvRXQHxuq0TWgPoDn4nGru0OpiQCpdys9deEm7fGB036MGNZeqZ3a9OT
ndMb7jaqvWfkyfishC9y+MpIs9P10/vubuKur7Uun+j+2Lh2s7bb8z3OQ9ep92i9gF4F5Ypufad/
p1rAoxshwEWjJRQ613PLUPGfm0Hc82pTxxjKJt1AzWgEnjTCi/HQ7XP7i3SJTmT62FeR6XRpXUVt
2AUfFZfUanK6JNa6NO4aFKw3KFQh6HLnT7e6FzC+ng9RP14YCvqbSpgEBLR979KNbeQ2s53GDl+c
ivA6mK5CDOQEmQrqPT47rnJF0OHHJhRS7BDwUYLeYSwOGybjfxi9pwK9inxGsy/du/8uvZh202Co
WvCdji5qxysydV57QCfRbkzRxN8vWZ9kfQEfKd0a7BrNAo+1+i+NUviZua6l1qiZhh/GIbO70r9U
XkNfbkrs5qD+LpA3ZOlS7NCoWu5eGiyWpEQtB6QyOmphrRaWm3cZyS4trts3h9lNHKvXUa72PJXr
10ShH8n1rXmCRy47ZWe19ut+nCFEr1dZnzPNMX19q+NUwlwMMNpGlZ15AHwz9DDBL9RAtT4jMH17
nE6Gc8DJOd8HfgiBshF+k+6QpJdldz8pliTL+0vzE12IKoJ92t0BYcysEsWNZOMmuLvaomz5vt4Z
whnzSaTydiO4jpLTRGb72wibO5Ewuk99Vrm5hGRPjjIWTyEdmd3yT8ApkIqZNr4auNIic6dSXRCj
uBSHaZWzxx+msHxQRRxXxPXsgw2XGYedPNaB7DQHZ2nMaWzT0Z0BWk9AiJGxnrgb6HBafCIAqOva
CIERt5hEVsxOAOUpLG3AdpBZ8z8V/f5dsczHtRPJgiR+/TNSx3ui0k6zxiXnnGUxfOABtOzSDj8w
Ocn87fxtSK4SRrn1WAiSq26uDtJ7hPrO1zylSGt90gjHnfVYWLS+eFW3s9WFPljkzdXlg13cEmW/
hfXFV24unEErDlYaxKr9ovgyU4S5fhNNnd3ZWJrzKraS4oomNv0DKmWRXiB70swOiaDrxM42Fvt7
icONDQHFz90rVMvkExftzhTDfQcicSM01RENZVsGn5hyvJkzN4VjHoCB5S2r6/ccFn015541mKOA
ScZ33b0w2a4BNv1yVI++3ykdmfVCNxI48f117UiafHvCRETFiixEtYrkKiwECa65qLnI0jROgOot
pvgJfulb1NW/Cj9o949NjORWqxBVezXX9JfJ8GTVw+910WZyMXN2wmqPSVkkaJiJs3SR/YA1BAml
mPTKe/P7j55Ulw6jlk+vHvx3sBbf7eZZkvI4kdpklINwD1bfy5chnU1I2qAM8vYOxTXsrBS3iR74
Ec5uAiskNbFn0V6XPH8DPLGwtYbfwHmn8oKWaDs4VztAqWAIiGz+4sX//JgT+OUvCPneZysSGvrI
cuFx8CVgD6j+kgpGYZRAuWvWxZlU+VJh857/mOD5ktbCi8NlWk7OlCT/bDb2yT7BZHCZDZw1Po+T
EBKrWgkFHVi99R7Q7pPyMZG3e+dVGU96vBoi0jdn8BH2UaU0xqbnO2cHkKEgKFAfRLbrXQDIWsxd
z++WRLP87PBnZUbZTsc0QzyjoE2DKE566MuJTkK649hXR3REqOWWHLcHYppk1KJGhgOTBYG4sgGa
+lQkD4oErJcNvSCtzIHAQlfmKaUguDBg8RIiWJfSynRmk8tHaXPPCWOuuyYwxIMIeZ9wNYbCn/cI
4qaPHEk5JwKLDG6pK78WssIr+BwMxBKKv5xJQ+s40UghcLQlyyKecOggLrhS9pyhfuLBAdLnf+Um
0gkTggR3KzMRX3hLA1JVo9+iquy1cTs8auagPkuKwteIfzn6l4DnuKLg57bdiAB8CaGOu1ysBu8v
rrkbW+Rkcomsmdoq/nDVCHhQ0BHX7ut0/bds1Xpo7EOtBISvTlMtPzBvyRHDHChbcRyHOkWoQlsz
4YvuZX9Rtz1unYyrBb58qEIK68v1taFe/5Cd3oXMlmCRJvo5RiK6GW+5UoT3G8pKX/9MTnrbokwZ
qqp+y31RgLw8g2VlpdUjzDDdP8jEPEhWqFkbBnSzGP0PGic+RDKkRDP+3mrNWsbGzUYyt7frmvyH
x74SR2Rqlu8i4zRiYBCPNSENXI2ZNva5RF1rEMV1Kqz5Rd0N7qSuE2AjBgjSPUEfDKhFS3Ng1e5o
3m6zlsF6PaNvh4Wob57tOVsJmppqL03dulst0EZGv155WaeiStJ9jIavEctqK3b3Dtf1/yrkHhtQ
bkRiJL95OEs0uxbZasfjK0sbhjWEIsCGkxFA10CR8eKHxyOHOXevLgmrZxjgY4/eg6fUOtYuHhRU
NDIojh5nUo6sQ6lzE01R2Ee+qWV+vngy51640e/zxL81kCXrkxyJfudOaRB1O9r4s6gdDGlJMvWe
mWJ6asKJJTZgGzSjPdP2i7y5FNZq17PbCNMEH9hoUBpfOgjDSZQwwOtNuM3sd9spbMLwp8NPwU3c
Uv0q2qiasnqW15dGLEuHJQXkTe7Pi5r/7fatpLcqOtxNdXeASWZeSwyqNIYLqfghcg0wf+TZCpfD
ZzBBEX+sAFrgzclLyyRskSlQ3beSkBlQqJ62uGrfVBcNnmpeXB7HnXxBb9YYBM2jfKakeUEt09JZ
skWUgBgkM7E9uQsB0H7GsljBKZ7ULmXNNrrjyg+Dl7K5z6N9qzQGWRMj1AZ3i8fI/1yvyhDHG1X6
69wHOLI6hT4LMxP+5Ajy8ww47j6bv8gON5+JJ9ROliITbPClsD+yEZd+slwXUkDzReuxAI+5YFOC
L4hsbfNiDLwwStUY3nXyrGu7jrJtPwHC4xM9YIMjcHm3+gHHQUwHOnhsjCWNHm7kO2BT2l0Hn4ju
khSb1pwwgmHERNrKNUmZyb5vwRDbubgdt+n92m7gfI6vqHEs7E0DteIAcvSTHQlDFEMPuqLSieUN
ODGUzjdyyf75Ok+xvNQ7Zc07QGiALcBviBcC9hOIYvpJyaYn4rPCRrDU7B9W8aRqFydKTxeQj41K
LOFToRCWltrGNOkKq4feAv+3Wpr0ZDEzTWm/uCpyosYItnnM0bwaCMtl6DKmZBxcIPU3g56ztCA6
JJPGHE/hgU9Kr5rZ+TDB7yVO1/roMfq0DA9p6aOes/WBF2lAD9LNhJiXqbMfyvPUevcCNRnAp9GA
JuPMuhRLMQ3/YT/S/TS+UCcGfnd0RCicb7xD5bGZ2BH1EIwT8Qj9iFo0JLOtrdjzAjKAred3/rRu
6ygJqK5YkArKP/ImpBhn2EpB3+Z/5Vz/LiDM7zW1f9MEIBNPXxNSwaooy2ZqKgXMri6YtWEXXvU2
4+g7xW3SWpjZ4+LG1ViroY4FKDXcyaANtzc3mUuTV5MRsIlPU6mnU6Anzj7npDdFkpI1amngp3N/
o6FWkoMcRqWezS3B3nQ1b+N1Fte0OVdiMvmZ+H0a3t/Hy2uNl1h7ABG1YUTyjL2WQLlAgVJPGcLL
BX/oOBKVl5vGlTRQi/4wE2vph6V3zCGhsAYJLRlNOiCSXc6BWXNBM7nTN9+UJw9ofcZVZ0zCgrmz
qtJTMkDGlTPp8tEqpZQMVQNK3yGdpnPTClALT7pc6OTwU656jCgbfZEuWoyKDzXWaF94mYssLrgU
sV2SbNRHNIsojw9QH+avuGWs44luNMKwudXB4+6YXIycOhiOPiqs8LWGUc/UUhdr4J+HMJjc0roL
CK1sPrgU8TorYcjBj6zQ3q547b2qsXhmTLu+e5IYnNpuH3rllDqruQv6vtCMiziwPzRKKITBwXbJ
tACttL+aGo5ZAKJe5i4472cjWu3AY2XBwySWkrBLLK3pPR2tPxPlL+T67FvCPiPxYiRqP199tdPR
bKyqtFpoRvRs2LnRCoU6JKuwBdZoVVyH4tU/bhe1rRJvNG/z8hNhv5DRWyapeBZVdFZvpSvVxIeh
s3nA3kdo6dbaz/aZAeDH3iETNda0z50+vsjQKsGvOt27nYUJT7rQhNzbU53Y04rc+omv3bkJdJcg
pqlh7O4qYKgFRJrFzW705280KT3PPYDgIOxINgh2B7tc9KMb25VUGKf5Ew4O4LbS3LEZvSR1lpUO
Pi641HvQPfKJt5dAbDr37mdT66DiVrRibH4w0YbFFSATONTBjy9WNqarwbshV5Q8nxThierQNspe
rY79qf8LhjaN64EYO8xP6LicUyf61r2VYYj+mbZS8iqYx92oaK9D+b2/ltO8cELT9UdjjSElg/VS
j4aR1jmISXRmjTMwI1sjCgmZTDJS8Se4I6Wqgqx4MSkDl+S3aKBwvztGvUuRcLcgP8L5Qg63sbMm
YR0i9/Y9gpk6kGGvPwxURgxf5ug+X44dwSoRAdN08CKbVdgmb2b3XauzKaIeuod4pe5oXEJ6tEMn
Cx88kLIOXWbN94+7+8+c4QelTw4kPKfk7RnyjnMzqxp4DNuz1N5PaZd0TvpbShdca5U60nf4vtMG
uBkbkec0/TWnA/enClbi+trZg+QDGcvWLfKqVdpVdUbkgBgLDkBwmtZrCUtbiZ1tvEbUyVHKyYXx
w1VYyAs9R7JI+QY+uFqMD7znF0uomO1caogdmsLm9Djkilj8FTrRNcrdwlo4eiWSoD+5KKYXlmU+
4nyTraacSuvmlQ4oU8lXddtJhKrxZngqsgEveOd5mVvFue26uUSwULjq9WsC651BR1ydL4yhQ7Zz
TXt6MaGl24Z7Tvnh0vBTqIZVKeMbAS9wGBj7BLiYBcrXfE8NxueuQ3UPcwvMFOv9lODeB56p0uoa
361j/e6+cz9Ym05QveRlIEHTEIQpyagjkdFQqytAv/IOoSO71y8tqtQjT0fy+w2quTbnJ2v8UPHz
hP2HdtkLI4j8MobyJvg0xKIMA5puXTCjxuVg9q1peYW40MbIfMkb1E+/fV19faJhWQbMKEmfeMKy
7xxB0ziPhm03ogc2N8b72yHXbg6x5L626Xf5KSGdU8n28g3p9myfufQ+OGA8Ohn8jlHntL7sDKT1
16/bydKA8LH4gPCqQtEMgiVZ0PaPWllb/4RCoUOjoyVaqrEPjARLDNuYk4NnTfAoBol/VnFYhzBP
OgQuenfq6Fcp9vDkNDHD8hFV7eNzQIdBrYltRPioED4/E+27wASDXqWHKfsCj6phxSngZYTnPdfO
t4UlAhBUnf/ToEIQxjDr3JyfIIWzjOplVDmolz/zvkHGc5fxqxNjJswnVycHl2EoStR9nLNyM4jp
rGY6tbn+Jp+7dQzxyeeHKctjN0ouNFo5AWG5MmUzpksbob0ByQ+kOCT36Vv4NTrijIXTzKxWeS4q
HMYazpqxTpGtwDG8qxqe5q1Pt6ztUc919CSo9yGI5/ykRyabqEBphv0KEYZbUjOvPZdh0wmB7HgR
TxDvpH/DhWXvmrIEp2LIXg+KHrz830JoSI0WRSS+rn7LzKd2L54ecM14HW6MJuMII8wcvC52pXtP
I/IrC3LSowwUfXYjlIqr7CLm3gbNgvyfFUDjKbUhav66UgJS3WFWhGCeiCfiM7rLFk1qYm9N/SHb
/FbHxTKQHHYh5iQxdAAmkhQmXrPvzv9oKTKIHU95J/oO9jjCYJpyz3eCt/FLOnNY4Lv/rijZmRIX
8hFX16HnJux6UtEZtvc9Z/URAJPTizJsmyJO5ccDxwznMZhdAU5YwJ+8g/ZSHSadp/BxoWLDpzne
QueVwr4P3otv+P+0xNYd6zDqjq+1xquQKjaxDSqhFgaJj8PGvNIFEV+mFf2PAyRC5XmSyZbV3zyg
HEeuKLNVpcJHyPf+oO20mA9D6oBlU+kbOFr2zPCC5Tr930hzsxpHDsjb9+Mdkdwjsvknarockzjo
tyafyaVewoi3B+TUvSMxtaiCt50GK+CPZzM0YCB0puFVT2MsFI0AvSvhWykDnqv0QFx+u1tHdt/6
COqh21vlMXi+QibcFSmbQxGACPLc/5am84gEMVwtwd05FzSKdOstkv4kPVlmIai8NYPVS2j9SB29
kRZGYKvyYW97XlQhaLMiUD0Vwn5FHqj2EGMtXw0mU6bXX99GHEZbL0VHIDovaMp3M1077frWp2Fm
gSs3PyOxka4XLY7koCFTleu4yk51OEyr5DLffO3F5ZSVKcfv4H/1U4OabQrW5U0d5daiI+Ijp1f6
hlONDeMl+g2/HToyqUuVTcM0IwP6E7xGy7z6JEq62A0k2pYFkcbVDUXE/wHdXgelj3U3ZrhBc7Z8
XGVB+es4FxFOBJlLcxu1tlm/T+y8JKN56+nRhRFvTo6zg9bqEmMMmyMcez5Fv3xop4t0tAkbQQ3C
1WoeEkO9Dyri6HspY+Y6ovrqoQyprp2L2oDOAGA+p95P6NX+FPPoa7vDMJCDBOnj6tCz4+1Qzi0u
2U8gsSEFu3pmbzGgltZOrXI96YS91Ra2L/WrsAX8PAPrJ9GHy81p4dU25BirNL+Apd/YDDWVetSt
Y0bJUQkaq/gKC7yW3N6xNpXhi27TWRdUTOc+MxgMQ6ByK8lVCMtsGnc6imAOoZWFkSuXu/ezJnC6
Kz9Y1bkLuO4uZHSCkSdevMTeo7rEY9/eiuK4+eAdiU2DnmUPZYCf/0fmHu5tiVFNyhDpyLFF0wor
yariqyXz8T9EDEFwz5W/Ie+lCbjNR+P3CE+9zX4tSmJnBmZ1yobZZ5/AXCsmMQ2u4nuHlLDDFwCy
Yvlq4ENtppxffHi7h2bGyYdxgq92bZ0DPy4Hj9VyLswM8r7FsjH+M2Hxd+9imJqOEMcrBgotlLt4
5cX1AoB9hzTv4N8/onR/+4jqmhFLe/OBr3Gc34nLQdlvk3g33GPy1vZkh0YFp2jXbp4QypnPe/CT
5H2yq4P0yPbm+yKktm5OwjePDrmIPEdJaVCk54D5eLmF1yYt0yHgQHbnwmjuFrxLQfknGlGo4XTg
KhkdLyA6pvNEAmQC3VSFnRY5x5+pwh2RXm15fUAS1mynVjLQ6h3Xs7LoLsJLjQg0hzQQkAWH9Yy9
ehMvl47ryM4xqTIHNGmn+5dpDgw3g0K8k9r1rNADNfMk+KVZhXYtxgxytmAo30Q+76ppQ9jbhHbN
ea5RZcP6jqRey4pleN30y5MffgaWMjUfGSZN6EZ73rzcEftNfOUNunL/FSAKf0UUKTa1z3XjVqdA
m/EA44gKIYM29TjOJMoL8QGPQ3sed9SP19Hqktwx+ZK+YXQ33eDMsPAK+BvGvb2OWv7Fc0bRHlUE
mlJ0SAjzGPAC4qs4HiXKSLlVIbnxDkD8Viz/McD5UiY8LF84mpTa+LMuoJ/7O2h8Ti+jJVcjcsK9
JyyUQguxW93FmVxHjkdnUKROVvyEpkBl25CFIYFxublidgc67lwN2KD9+Ep35d0C3rdexkbkU7ty
8X5TVxXSg+6xzbY7aJH8hUYCtL8j3HmPYIgNqICH3uWpgg9bFrs1/Uq0M56eZR9+JbrehrTFNgZv
RKZPRRvGUt4rpVV74DZvb1bCpA66MjhIcEtut2uaf2EG6aGR/0KQPOWYIDCIshAOIXkljk3QDz8p
8mcsukRnLHDhXPMayaAIRDpgLstLVovRJNUEi4yMy6j3gJi+PoErhva1j2uM5UPEfVP1VT9SR07d
6/TdKhF9LeR6JS02TjgZapQHEnXULCFF5ZZ67OiDzTyqVoTfAMDHOTrVGeN5Pis3UD4KxMb3kvVW
GA5QsCNeGFzh7IHd8dB7V8MgL7Bt+RDVj/3CCBeT7ObK7ibuRowX1TdT4GlTR6xvSCbaisET19tF
wSRTM6v5pb8MxkledXq5XhnzuzyaV6ykgd/2STuRpMdFYz+sIYLY17S1eyJt3iwG0MhcVUhm8hoj
RohWfyLis3u5yR+mvtfNuTbVN6AGn9cpry5w83uIjPBshEowkm87ao12I8G4cVt/GOeVa+hXMZsB
TFKI0vAEo3U3/foKIXlhTOOIzFQAGXCE3dYHILgUJBc4ulLwOqm5oKQBw3T6T/cyv8S877MlfA2V
zr6/dB+Ri3f6+GIe46VtDL8ZyguPLCr2LT/5Pj37gNf4OtdtM6FgjXRXUcnaNBB+C5VXWJYeI4jO
BudiF0XoverXwVAkYQ4J7iMKpSUldSGQaRCrgWg2MFXIUVnS2v3xbp7jXUjKIyGHhjjv+p8zn5vX
aGGwY7fvINInCDShEghs3YfdhsGKno4YBmbP3MmacLnocl8HKaAhOfrixJejnJ0SM7LInaeCbGa3
FVfBEZxYwLcvE/EBJIV5BvGHZoXHLCxA5avhVun5Z2CGP8Oa+RevgadjSB9YoUZ/3g7h3CvaDZ0Q
PjBCA+wCTeTNUqsslKsYn8v9fK9wCK73sBV1boWGX94tjEIB/r/v51zzSPq6uNwpbnG2ss+Lw/4Q
E4xnUR2KXSDzFPRPNFF8lDkPVkCZLTXJ4A2qXJ04a8c8Zk8wr7m4+LD+i61G3voY9NrYGYn4G9VD
xvQuFheRB+9QcXI+0I0pz4eELJSnCoIbzt1+4x9UTe/J01kU8WR3+m7NU5nh5uieT4BF3m6ZIcoR
ryBtOMk2OGpiSjaIcDAX8OVuYWAB74JVd7Hs0etBOtz/hXLUXAq1eWX38L11tJHBcV9UVed0wCm3
zcmn22z2pAFHAaS61r+AdwFKUMxbUCpJI0z4sE/BFC+9N8B9KEISu/UMQ/mjTF+8OqW0CUpCNrND
HtZ8tQnW+WqGqH44BMU4yKm5JeSYqTVEBZUdZjqvqEVHpUyo+KCeFWuoVegANeUrfufmIe88SCH6
7vV99YyzKy5JqPm9W8e7pg/1/jTLJy+pkDc+TUOln99MA9eDpyMT1BPqE8Et3WWecgr8FbAICGwG
1CuZ7q52b1ti7Kj9tc1hf2J2CbRdoiTIgGFh1huuqHX8eXUNTXyIIB5WXiskqAgCMJ4K2hdWd426
VLZwc+xDG8uZi40jBPiPswUITYt5QkT5z4DkxoA2bxY2y+UDaRGdy4PUkOykFY09i+WRg+j2IYUb
RtMYXi33LDHPQZUnmqrIi7r0+MKFBSC9AI4W4sWYVjORoeFOksH1ACfTZ4Xih5eD4lJm0/nSNKco
H/SdRULcNOvZ955UT1yjg7OYMdufiDDxQkjfgony/BcvUnBYTvTH/pFcy/sr/8x6zlVTGJrTGPed
5g80pCmnzmXEN8DUmjE9mM4gH1vfF+a6sqSA38yUErxgWFfg5bsUaaxQViO5t5VeXz5hrmuqswpi
NuoE7Mpb/BuvoLkR4XFRI+I82NYKo916ltb3+ycy2WSh+iuTJECQ4YCkYwHma9DuVPBjPCl1vT/V
VMkwF82eM0aNA3yp2EiJ36TjJfo6K+FJ7673q/eMu1CHen7cLs263dPor2f5Mqp2B3p9lbOtX57R
YhZk1ytSVHm4GYYewoKL+txTSrLkJ+fSbPMhIO33NrxpprheTGvHu0AQv9LLmjBsEAM7JLg2WloA
xEJ79/Eg4cpdnYxKC+lT5EftdMIvLUOy95/RT5UMwmBau8BdN4gxq09feLxvTEL6VRkefFkSKOCs
Wtpy64hI9RKR1jsDoKV/petuEb1k7kv/+HbGfxCb39HUl35/yT8UusqK+WBmUFQ3h2klGFO3Hslp
27M6Q4I6RBNFF3jXfhwgJBQvEQw/1Tx6G8Zg2gV9iEIgJej8x26K3MFnm5ObvLaF5mu8yJSnLYrt
1wvje8ckxTRa3o8sjbz4u8cno18GS/0FLNU73np8C3CKFaC246GRR6bjorAhBIESt0SG1lY3yInV
KzFT7wyrk0mbHQveeu1vz3FUJ61/NkJTyi3nv6DmaWHKyhLNBnSmtFCub+OOwJTQ9TaxRrRQb8XE
aWkMrVFN6y1TrljaOH9pUdDwqonrVRpWlCF+TdFFVlI2egWyMCfU+Z6RwHDWiiZGJRut6wdjV5XC
fh++dq2FtVBDJOIKQ6g4fOu07RTMxoaYKe/RAvGwVMvuxIjZl0oFEkE6jvZvPIVz2DNBbqB6rEtV
k90QY04vZfb9BeOjZnbCYBjXPnEl2ySzSbFS69ujm+nHwUbsXn8DG4/FxRmumkLWMH2DqUsUSn08
g10w4jskCnSrn8LMFr60MaaQgaqhnHDk2mc3AQ2vX19gZDC/hr3X0dWmAn4coetYRdtTgeb5M1zf
+FWj5tQjRA5eFpzmAWf5xOgY1PsAJKIqVnDX9DW+rPWmDiJfIUo6wlpNrwfYfE+5Uas6AX/cbEpc
xkQTpiqAz9NOhWtzG50zi5chxyEp9w4dXdk6/07oWS5a3S0uIwgIRprJJzfITHl1m9XgtDqqgcOn
noLQuTR06HXzCi6wpVgnbdxKDIHCDo36IKUCNkpgYvByu5MN66Afk8XDtnOxTL+89aHpiq8ppH55
L5Fgt3/Hmsh2WbIzJksuA5yho7waz267Fi1QA/qR9Lh5EqkZwkUdkb3mly8afrEt3IBdw/L3tWyL
0UoMOxreTmFDc2YikntptYAAruDqWHYyyKVaZlGWUZjd2OMXOQKvGhigkf8p0lRlKtXwZwX/b7lO
0DPBqG/cNIE3GkIDB3WTeklCanwpyDPbHTZtc3Nt1TIJRyMORlPQKi7mRNAIP8cVabHLIYeCf3oc
gNJvbV4x9Zrj8cZS3k+c0s8XgU4/twYV5dCkiscaP4+7UBlOIWF5q/yWNuwxN66Ki4Etz+xVAHRy
MuEEYy/rCpmnHIzrf/ju27xMdjkwIP48zAnIKVYFg+BEaEEy3ow55/fyXzM85vYlMK+Iy3/yvrrN
X0yGPsrIt4a1DWT5hjlWENi/aavb1wRVO+oz6dzPlKHn3KB+Aw5O8mc3ctmJ097KaTWL8d9XvsOM
wfImoEofpvM0dewkZAQWPn0cdVX7rtNbPQF23e1DwDLbya3WuQF+Mtghm9MFMDp2Suw+CNeGzHOG
mE5ogslQ0J292JMHB+OYBGgU6+2ucafyKzAyxfXHx3ZJfLjSk6MPBLvduegbx24/INmZZkJJf+UD
KE8ykQJ6RJC7Cuh85yADLZxFlTSt9K3r8zmHK+yHf+o4xl/NvPNvRUGxEmVII9chdR4dPSHb4sKv
X/NbNhE0BIv1tuR3ogV7IFS93GMKXb5DChjciChkXX5N9lm+Ru6x+ajGnim4KlOoJW3Hd6BDiDmo
OKf2DXAL2QR+hQtSJBQIoQKmoxe3imYkazXIsR9anKcN/HEMEDzHFEdENTFT6KnrtfrMY9vHRvjC
2V0yJOvJG0Lk1Vnb8Rw70c4zS8m+CcEdeH4lGRXS3jzC7kXqx+LzhdWXdMyjzYbmyWOyC3tHIMSJ
DiPHMb6RYRdV8OaxfdGMT2R6U6lyu08Q9zh9u6jmIzlpXuKWjoUSeqKqdvKq+gv3RpIsFGUCv8nd
ly2YOcpoJaf93II3887Cb5ToGi/a7R+WJcuSEnLP4Ub5dqFIMEsj9tzldPi37bRTI1gA1ABp1ECM
vlfCSchz0l2K4Oxw8gt7KgSjls+9VwJW1q8+W+qo4aytRvrO0KEYGJ4Oin7QnsrBkRQcqYN4RUjv
b6RHbUlbdrlfOLibhGGWebHUHDYS7Vrbn4DehM0KA7gBmKDT4nYAYOS8j6qMKS2No9YsXrQfgoRG
/wqnx9OVHCiiHVM2KA7fp/BE0Zb3F43xeeevk6Da863nwVWI4tmUStd1rUqOH5YuOOt7+UEwCJZa
WNrr5w1da9h1krLgiF7R2cx3qdcdeYQPcBmbKGeOb2Kk/3sQLRzHUtsSu4/2XEokL1GgJ+l0Gv6K
nbTVtOOIekcXUv4nl+W27xtFWyk76iSFBkkkTXbPa5VDC1wI2tg6gyDpqwosRIVzhBKtliLUNr8Z
R2mea97XOKNsN5GOo83HsU+KHoevBgpVWnxjvXyj/7WToHPJ3+JxN7tqMT4B2dw0do6FBvzfayGU
tCojPewuxlMpfTindFUGnASDsaz+rZdF1pqeLA6Ot9e6bOf5QWFUtIxRqdVjjptTwp9hxk21mWhd
z3Hy+7h5XefB8HL+nvjZ3LJcap55mi+vDBYQ3jpO57fSTglycSEhbRxCtsLYgBiEo+G6uexWin+S
f2ZasCudFvxK530uv+nP1hKiC5dQkBdg6Pb8BDnJA65/SO3gK91Wk6XDx/zQ330RYZfeeuuGovIC
cNIKq89v+8OMg1gACr8ufhmhk+2lpdG4jFyEW9STJuG97LoOswPIDwhskgJOE2L8iMR0e9pc9KLy
SYohYiHYH5As2IdMOQyZM1csdz4oNAVypyMvtIV/kreSkt4YCy+ejjumTHvNBFSH0rR8orAW4J/2
LEb3883L4xPv+OagcYBqY9oSEJhdQjJRiNMsjOwsSMDzwmkg/iZOPbvVteZCtV37IbzkXECKS5RI
mcG84kPd92UO9NJbUh5qxEp8Ys9GOd9TJxot+go4FArm9qTs2Mk8DkDSyTLfEAfpzghkVDK4EMzk
biwci+O8xj6SuiMFuUJBrDe8HaJWzRcCpGd97RKHnhugumVr1X9ZjA6gI/3zWl4thMiuo1CeUYWt
9dBOAqwzNXquRrAvVSP4wxM4L2ErsUJOtmSaxj4fWwep4SFMGevACLgW5qwqJbIqHRxmOvI6xG+M
BfuQW2bPMYzLz+hXf/sbuAxVrjc8Kgej1PtmwPDFeUfp/xk2e9eHRvYYlgaWu6nbz4s0WQpoKJ3r
nNGZ8qoEQvzSTArVboJquHwyhroPmSpFD6mrOtrkb8UW24xrQUNUDeBluG9NBNSKuPBDJcA37TGU
1rf5az1HR6GSzbYuxcfZAPjSAocH3TLQho1jmV5dvQ2tGZ1HQs76trJWN3Y1pcriXSPQGVL1Zp0h
Zh7RX7vSVNqwXblmBWE/OEKVFb3jhe2nGlwe+0HMOssAfkznxtfX20kNH+ZY6aS5LtAsoAMks2ui
bKxcT/196rzcQs5CsDcwALftaHsuZWVM58h/3NLdgzDC07j23a+koqIgnxUpKGFykvwE08dKNOrm
CxsrXUlig/ReEEY6WKKMWzbiglkzk18WO1ihGo6X23tZEW9QpkFhx6iDnlI9Cf1WDdcmBzyYy39P
d+oR1QuveLGPl2dAa13FB/yOaUTbCu/B9bgz7ilZqT9C8k4MoLTZC94TCsSssie9OGt+TIGZwHgI
SXDsh+94bNgT3lPvhGDy27pBMx9DXVttUEZw7lQiOnvPHWK/sJgb+aZPzbINDyDhlV3OnPKd263O
Axz2ct1x3awNpv1BCN7UjsxAQKd0x6wVqTjNz6H2YXgfSAeOqyu+rHCCA38v5PXfCXqSTlIaibc3
MC8MeHGxUDRBOYrXlakCDQPQWQwOZsw8a8OCvl1EShwZKyREbasMwvFz5Qr6/Zr4Tm26FUetHQVc
T+O2Eg2/Fs2/duArhzMMTF/2dcjm2LXTBUHf+JluR3Qmi2ivmyAxUnVY0QzCVXEzbXMrRxUP9YFu
MblQ0V5AvzS9D4hXsYXUdst1vJH47rUmilS9aXYgKXn1IKlJGpGh9Ja/XD2oALjVzwju8im6RNcm
X3uMA0qR1HckSl30dSXt+RZuEgsk15hrx3+hg7H6+8Y+47ZlxZ29giWnUPvQi5r8yTZxtEJM97wI
ZyIF6/d+ZGK9IlAPvDoZ3/KjMP6sQqKgIiBgAm7MG9JBDOre/60SaxCsaB0YYeIfp+25JA3bL8MF
YKbIpiiFMmCdCqucsDzI2hSuDAUkCycKmKybLoxYn496t6xGZL7JnwYzOH7eneI5lKsOY+VvQkuf
sictf9wHzZS+I/taD6l7TN/sGUQqEO6xpYWeu8BkX/TBcefPtx+GATSKqnMAFXSrnjJ67rpa9fqG
wBnCJgzLtxHpLMFjMEcyAT7V6qsUHVzwkCKQ0BSuzWB47hjj2mJ1tGX2yUBj1JVuUqWRHF575+R3
Dq00Cuun1KIH8RHwCv6sLlpLX1qOV8JVliAfPpMDZ9aIMvWVmgPf8q8lieG/eDxAle2LDjqhxaxI
8hKwSXLij9Za2joU7VAn+sGGvAcIElviY+vuuj1JjphxgXo5G3Ysl8tJuTshbKNBnAVCqOItlfkU
+qmKIsUHb5vwmJnNTUg2tbG2nss7tvejM9oZM4iTEWRzGs5zcxVGABnOKznn44yu/HuH+scE1sz9
e1iN5TtlNIqied6khXnLatDR8VwTKWixcws8McoSl5FOErylgvUCe7WPRJRh9S5ocoacCXLccOUN
XixA1m0ge3P15TzqrAZqOGUJMaR4dE9nu0AdRn60TDgoLSC2zyogOVi9Eg8QgQgyUO2OOEiTCfng
cuBB2mq64mFWoY5N71KoQCsG4wlWpu8mfGa4ogeiOvRacjMsjAT/dNOqCnLbVraKio8wuZ1uW7u+
R1kCSIiS5LA/B4MqPPpVuOhNMBSdxtQc3IhIDA5xhqaqlz6N1PVuc1GqPNg4u37FrYn6vSnxySGe
Fcwr0l8pEB5W0tkhlG+bwT4FjLDuNl2pgKupTu4Cl8Hb5at1SjyW4PGmw22ckAiuvq899MbVolYx
muU7h3ro/LgpOlLLrYq/w6+cwNIyaOseAYEPdx58EUBAqfrPg6JfQAXsCDXwfgWO5aDtpdBbZytP
/an8EnlnMBE3PW57q9WcObh1i9Mqu3J+2a6niN1mf4BiR/QN4wOj8lQYcc3fHH2Si7GZnJ/oN54/
KijXxArnUyK4wByOhDC3bvEs0uM7D0sJ+fK+Xa10ZiBmsRF4/uLbeHPRDTYjx3zEkcTIPqJW7d7O
LZ7KF/Qz1Y/LXbVYC/5wYSTvPzsHqH39giPnihOhy1ndznZS5PrUlZSgq4DZGvxSvAC4DePzxiiy
1ZO4/XQBULlPT5c/5C4ZKr1S7RwHIBwBbihxRnqJ6DuQ8fzIYjjjEoqXwrd+Th26AO9pLgP71c9s
Ajf3FiNL1om6fm4v30Xhm/bJyeXgN2OoFTUXvIBnfiwVZOPCOUm6CcspENAKlUJ/MZhgyizNToWX
4zQ+4k5ZcAnACEaheh3KCOlNf8Q5nnRLhmffFcikuOGs1Hq+nPixJnwJN59+O1c6ggeUif3UzEpa
Uq+s6X5oBd20EhkuzEKlrsPi3D2UbeeLdPTT1qJU9YayaSxgIoPmhzzrLEK7IXC39iGfbFZJ2Nuc
BIi58+PTPrGMjdIQQjjq8GZhbAHg8hhpcMWGUTPi/VbTZ1ZeVKeUyNq2A+MgssuDY9QSHyW/qnqP
SgShmfeejtioBd4xGZ+1EwkkcBZljQaNLQqMA+0QKqF8hWxtp73xX+AlrG9A5XIDR9U91sc8Jffm
BYT2gt/sfxs2oR1vqyfoSQ/i8fo2NQj0GrEjfSts+PyKDp/1PBHxwUP+0efGjRQW8oIJTuxCnk4y
XCL0fB82ztUyIysPIEZOUN/FBX6nxxu+i3N5RiXMbmECJYzcE+RGX0m2Mmvxv+b73a2HvX3MQvUi
BKBJq3rwY05Q1Y65kgh8wu3OX1+7VXIebUejMKiWmbZJ7zBmDZ6sP/j+fOUwlJX5ahbcHZA0n53x
nyHEv6BigAjcFbC8CgerLadYvvOlyPjeKyRtO6g6rIGpWOj1xkUZae3fimHBWk0m+DRxBBGgP76r
cK55XBQGcT6HNkiaFVY2cFGt8rwZIA8CwJTc393ke4XT7RqT3NF61zVJTPKi1VlWsUWlFZv0Ksuz
+SwdCQnKFi5+7dyWyicbUCRI1vvL1bTkg1ic2t9YaEEl9VqE7VpnCXKxlL4cnWSgHcxBXrpYCxyc
wOJZcO+aIDdMKSA1CCwIXKAayfrS3fPn8GL5Dl/B4E6tuQ7/yEUFzHLsu2BNy6j30VwYnTH5+Zuh
vHDFcWeF2EWvRd0/npKz2h2w+kSEX4Y8t1fNv2bH5RDGisdNvUrDQf3GX4VZtVE4H3RwYuhYkf8N
uWlsV8YyaOFtX2Zqf374mMvhniT6/JELn98ahvDZE27KdukkQr0hleyUK4k1UiR3Q5f7XPaA/2bJ
c10l5IRDfkc5DS/A1oFQ45fbveNOcU9DHZ1BWonmMBJeZHUqg+gptzKq+zUfFmXOmh84h0Nkq+zG
XawUJhB+1Bd7U1JKpstJUM+3SljDa8Xo4t/cqJBVN0uDKuZvv+lBrhFdh2dJBHtt9gtVqVVA78MP
e3dN2M702w4jjI1o3iskgJCtzX1Kj+AVe6UyE4HdQ4ugJSS6++3AAn09x0ybsB9XXi9jNKcMURr0
RnXGKR0PKPGPO5Wxc7LVqlYDjUggsx9whepleQQ5nptLSxvW7aCKRBXTrAHL2WA4jmTqgqWiVjHF
sENhdFXxFfqZGTjb/uwFxZ+knlIUagkCQ1kWh0+l14qh7e2zgMLW+EjjhmAu/H4CeCUz7D7CQNN8
c3PTwrslkGFpnJAohQUBa2VTVbo44Paj0M9T6P2NoyjyGxCPYxcDTEo5+SCUr4kBKBsxxIUWQmwV
8nTdvtoh8i8IyLDyuJt4MfdD1J3YuL35bocdzZxFhxNrxOaQOR6FhX0pq+uiA+LJ03np0BDxR/os
vBJX0Eh5gKe3N8fje1SyPZ6jooJLvAkgiMpN1jONzANActauSk6+pxXvR2830LBok22ILP8epy8z
heopaTFbf7aVJ0f+jUIZ4yTi4FFF3G7J/9vMiZr+Tl4P3f0ptk0RYHEELx+1gEzVMslcHutbZ6pL
Ls0QW3LXL+EpFv19Yf3BkOE8dxyQ1fjqzG95JGuc5EmQ1yrjGRlCQc9jI4Yt5fFK5aaoopWJj7Ig
KyB7YmqjYOfuRtFm1hgtXkq6vSylm98Z2fT+ctdPFTuH1jw1F8DVPvaH8h60BjNLxSKa/W+BZwBc
c7TIi3e5g3LJW/uRFsRvh6zLGU52N8xVcUHMMwJjMBuTQinB3w5lkbAJgW6XZfru/RUpPBgq16iK
1xQ4dhCO391pPA1jBe6CKiSsKcwx6hympveqlPhbb9ZzHCnpGIFecOUP9iEup4ySkUHEsngfpXR3
Fer+c881qwZoc7pRIZki0i1XzgSTL0ViuHtKOio71BWJNmhda1g3I5nUps8MLF2Z/zGtL7tgtvmF
DKU5ypumbh82cRXNdZ/QdpjyyaQddZFQM7WcH5OISLzwwgRSievdnhbcqcwgxUc1vDXJzEMZXLxo
Z050MqduH+Fqy8nkgmkFS9OKrbwgchudbGXCrTsbZ2+ucDesXc+2WefoTTtibBBoLYy9eaO+lHPF
S1MeNaJJeZK8QSCQWYKZEVDS3ZoErzKx7IZoKeXh5AqwthW4X+RJ1i0tn9eXC3b/rc0eOO26Md45
7AMgrwOU+ja3kRmXeChabzZjhfJiTiE8lJ5e6vFXJvw9i8WQ/658ncZBIl4wBouHJeSbNR0OB6Zn
8vyfZp+I+u9YhnnQFyVbV9TcmDaRdxl4Hv1vlGMynK23uRYETpTKlgGa9wXNuAQepQtanmteXu+t
iCVmNzl2a9ZR8tSMTZCEXwFboWkkulJqii8qmXFYE8rdV8fXHTCxgByzJwWTkkn2oWdr70+vhxxs
72AvYWKCJMzih2UIj/qlNRVPATD9Q/gpB0d8/fqkYb5nfqCYYltP/1r4w4YhQtNBcWkiR57JdTuY
G5w14WI4am3cKFZkODuaAS3DKXrGJ1VYf337R8yeyIqb1BxFmbA+6pZCEKlPCOi2/788oIh/qWO6
Z14MGmds6GhG2s2BvCEE+fYfgREMf27PyPcJp5UdjHGhGZu9tW8r8MPWfdYJ1QMpLMMyQJxoUhWK
yJogBLPUj+0cxCvgVZuOBdOpFz/bT7pbDNUUVMtViy61YOEjeSSYPbjB/lOADyaQ3PUtOGhE/vYW
1ZXUv3gqdNHaKN+3AuBG7XiTj04ThFrEGFgRi9AXWzRg51GtiVZX3gvvSnQLdQF2IIFdUhajBtLW
V9BwKr/VExGnEISvjX08usSmb4dvtqWZlIi0Afe3FXvAnd493lc3MgQvVOC+DTq+zdy1qOF4TlEO
LxCa8qKnKusOW2V7Bg9obOkjuqat8PUGJWctiuXJ5ggivKn26siRRI4BMVk0AkZlULKoQHvaJIha
cFpZQ61Upc91QAF7jCtqxjjo+DeZ5oE4cUFuIDfOSRRRdfkBRGl9NyhL9Tw4uME/3WDAUtCMCPLW
A9NjMU2/o3Ldx7Z4m12EJ4wIMHoEMiVDlzs5DBvGwNtSmFUz3p/1JmBehxhXC8yRG2OwgY4J5K8G
64apRWPOyQWzo1PmA+2Hrxr4jWZwcYS4u5Vo/qCTaa1K+JvZ2lOhIvy5ODDCFvcphdABNI2tllsb
UdVFbevjFYwhFGwRo6F8JWKJRdeaSLryCPQR/ksnUCw8lbjSEsfAuARCX9DVXYY3hU2Dep8bZuX2
bJBZwTv/cLlu4bJXsywqltOkbw2azA15VFx0IN1k4Ju+gZzPk5hmuY9kpJiDJmSZctU9YC5Tk7dW
6NULtZQXdcD5rgbPf7g0G31+JqCLdXAPKkOxYTrGJNd4JKvkCC2ga4pa1i+/CabfwF9kzlnPfcwH
QitUm7+Ao0LnBTwR+ReT41/7GJn9asTuCFuN9IS4C+TaOIZn54BT1tLIfwb2mIoZjrABFW3NEZf9
VL++MaUfEyTMytPPrbizHuKw6i8vIao0yKQUkXzu1h7PdpsBLy67Ii2LwJRKHY0d0w0uv+ZJEvlf
EEDPPcP0rOVkxG2FqjQRfAj4DuXG+pFE3f1XCXmlhGbndO/0M/mXhi/llY4ZrsRZlzWLcGHyQiYq
utqTWbp2Fw+kzcTspxRucGhJiyhDRMDQhNLzqdoCqPbDenxqDMA64bcI0hFQEn2FPFGB2sUfiJjO
XHP/lXo/dHdpxwM7PkjbtqH1wrFHip+rmU0c77gR5Z2PtJyb+cy0OH+sbiA8FDOqc2NT3ewdbrBJ
gWJyDnGBEcsDq3GVwDpBUjc83d8sSfJ2h+jnaI+8OSyBR5qsL0F3wKNS9N2cm1nh1cUUD/jZT3p9
KiK40Wtm9Yiu/i4gPB3S9RKTXJ77+vCoIJg10GFP6vj4nWmXzP7xpjgl4DDQrhh5k1fRz40t4PQK
bMvhniI+MubxXVjYlkF89AON8Vdfv1nSq0au676vC4HDAsTNDqB2wGA8KkNvAFMGtATpQdcA6jdA
VbRSltanM+cLMzbOo8a8dBTUDImgAC4dg6FLMgVsd4AMtHsRkdh55fp2YctvtpHPl6JsGyUeKiGV
wrySiRv5ou1gxRwxJkjaBv38jAkctF1i4uxm3zKloQNvtQs2F6QZb8Kth8yCMAiUvAi8U1tYfwT4
y92iH7D3kDNkZXEe6Jyi8fsZtjRTOZtfqBhMHVkYfoHKPq5WR6ZmEdgm8Iu+560UmRE1s8Jalam8
1p+u7jkqsInTLbm221pQiHTJajP4IVVv452Ta+NhAkmvHTI4E3VtFbM/vkDglotVREuEUsuyzzNu
NNKBAyGVapJGL6yiOr9JKGHQGkNhQJSEBKvHHvgZNoUS7oKVYXV4yZxYFgqcNDC7TIZ6v8fbuc08
IYKAySRjbkci88tq38ZON9UvyrF5WNOaveMnLvWmszL2Cr7bpHZRSMGXkrJNMIW9O9VV4WgZiW6G
uQof2HJMxl4IFvvl7jKU914PhkWdktH52ktkSdAHNfv23dp/wwaGcM0xLBnJ5dHNtKbzY/N9C0Nj
cgl2lC6gyKNTWh+43os2T6Ke6YeOkLFjF8hX6AlIR/gZlFjR8LFU1hlDyglGkIAu2yqFauouOlnV
bbfmGwuvWh/lbVckzprWuYRmQPtvmvJQOgXEOCLoh1cHQvR0weT5Uo5PzJ2kdX+SgE0aZ084Obzc
AAQgf/E/6ZClmcq2+yPq1AUCdatlnkbYmnkAMLGT0++SQbw4ehqUjBN6BlexNTbbwr9fetfTh9n8
YAXdwj3pKctCrxe6EVq11c26m3oq3FXSH8UYaGpY4kiENCOpnLogClS+M0W7vCZT5Fzx7yqrlsuR
l4s0/2r3mIWs+EDU91Tk67oCRvFpqjf8qdyGropuNKbuEV2grYBID65VUSFwUZpJnZtikZPsCkqS
P72RcdnR5bXjoMQwsTydnxAclH1HUHxqnpenIHU5y0eNjUgkWWUDXb3BagFI+ndEpKBMDmSEwtzm
W/F69nK2rO5UGuoLHVafAa1T+6ESPYr3g5pn0eU4ZrxkCVoGgpctFRwa46pdNgpKFQD0OmtKQEaR
5QssLlzAKkS5vv4ZtlL1wmRJ1+s/JZxKIDcPH4J+oXkuQGCc70WY/EDZWfvblEvVbBa9g0wyTaca
nqTnZjGtKM2O1ZP0gGyB2fsFk5isKW3+riP65trGLkosppDI3ilyIWSaCE3u4CuzTimpEq50sTzg
6W77jMZrvi2cYv3YzJoVDdjQUK7ditKxgSaqOjiQv/z5VDzntpAXd5H2PipCdXAqqjsWyMYOhsxz
oFeaE6sK+GfQdUkJOiSIbkfwUF71nFjdj1ITzy1gGqgiToQ5/zFI4mGWV/x7WuJSo4phIs0+ktRJ
cx+ml5h2eyOL6IWMhhgM/p8Ew2QjxlwoQu0R4c06J3quphbZo74FkEFC6ByyvX0hFaZTG+H8yFTp
zCMcgcfwWS7zpImacy9LugWJ61QD8F5CsWyHs6V7RCVHeOc5OnH3CVacmtGIHfLjR+6YASxkT1rK
6tMfC5I7pwN9ep1YK6PLfESx/dVc0aZs3+o1NppfXkmmGF2AKySp0XASF2dkNWVYxZ0krFDcyEcf
d8dGRUzAP7WJml06bKEH3wuj1flwkDzz9fkiZx8ScRw3CcspFtpI7eIt0UVK8ZJYZhW4GSEHl3lA
WOHZa2lE+HMnAHsovq26MLL6Y4GeeId27ldCOBTYm2clhHMwS85ty/3MHy4bKTtkv1lMj5xeCtaH
oFbPVHuOIGRP3R6QzVbU+eKZ+62qlxQ04R0UFzpxhJFsoshADQukOj4epIVzp1bFj5FSCjw9lh3D
L77am7mSzwvKcJT0574En/Ipy67+HhUQiJZNTqB10lbIDQxCTD0Jxdk9euWfAgmUnP1tqjKErFL5
zQrqOT/57T5OLsREPztuhDmj7wXip6qq6lJ+Dve5YGOawqe1bfZRnsQZ4O8mQbNLs0LiE5sRmzwJ
p6tpOfSdYCUY0sSojrRrAaiwejgdrWJfVj1/lAkCK/qGO8eRt7pZo5xk2iC9pUAoglIQE0Ue/4OW
xTIYyk7BSGdNe2sPlskeinzHRriIt1tc905XGSYVSTLoxHhUfzdrRLDXKluNimNFrwbhUaDRusJJ
1maaEV3ZH97zpGyJcnAX38+84THE2Ht3EinhXI1YpeVZphxjvEmSvxkRYj9zOHqYqVG1vY3Gdmi/
QI715OBGOwJJ7V4s1Csy2ylJ9EWkw5YwUuvKkxQJCVCPRwIJEXJKtHtn8bHXbOlx49Hw+a1pSDSK
+iRylXJ2qKXCUa11EK+8wRuQdn68w/4p9FPTEdN8pcykpB49y9et+lRwqfo/fAzDsH5SVW1KUUkh
EKRfF9d9+JUXfTXGi+bE+QPlTX385M8LpOml3QOI2K5t65wSJpoP5Jcqbz+fbqw/ZWUnjr8pEw7b
XDp58zcF07dqGC6+pmlBvbAzgcKrX/MKeMXKOpkv+Co8Jrv0N+AHVR7PwbzCZck4MMo1kzVEio3D
fWwaJ20ZLpcSyPARjgwdcvavVwnpcksNDsK08twcFyBsIa9V+iWdZqL5+0G+RdvQlJc8h31BvqtR
CJKyaEI3PM62sxyWOe/8t7pZuZHTv9TzKxQ/9CAv9sFp8qN6PDNLqx22zpT34YKjGI+Ese4y+C5e
4EJbGl6nMtPom8eYHTrzGKN1LWV2pUnnq4tqs47xXIjV8bHyOsr/FKSWUwydIIdETBgzBZeOcllS
VT906I/dX6otlkJtvfLZ9RxaEkAHvKDxMAFXDFtTfbHb/BhGcUaChs7Pm9MWySy5Hf7NrZFmJ84U
/GclJptekHa1mBoHb9GFh85Fvdw0SLur7LoCsQSBzG2Lph9Nuv8gdynNVr9y/KTmkM8toVj1CvR7
0Y9XGpzzELZHV/7VbEPc7KjyH68Su68+q3XACL7tZcrzFCbGdtfvsOQBcudUUGpGtPhEp5sEQOWG
4yuLRZNx8jhLosWTHzu3w6WD/pPHt1e4ghZUVaqWJi/GoyOOa3ykhC6fWz+JMGSoQ2vEr3xwrO4q
RODz63MqUEr615Ie/91vOZAlQ7XJV+893OK4KZOFvmd5KUarD8S9toDc2wrmji28iJmTXO1QyKqx
5+pMswhDJTVo4B94AMYA6o+Q5RuXN5itdNOgHybTNyTzF02BZMaNckkZr4YoLMtdd/Z6iA/8D/Pp
C5SmbjvyGkZSwICZWqiJk9OQPBdZkqMYuwC3eVsHuUAWhiRu5gBlIq7JEgTarKyWtHKJUBdvjLEr
qIdtKRek7xt76hK5rns3bh5UyG93FrthTNy5+gmLmuc4KIBLKD0WQ+H36BM0dsAMjgeOz1gcyZTp
4KeruPdPzYuiGiEFv58UZnAPFC6oY91IpkCk/fFZg7lrtE7uPg3vWYj5OVuf/Q67KoudkjB5GKbJ
1MUj5kGiwpeTPpFzgGZ0LUFTvcLZiodTmuIj9MnxiNbOeohHuS40TuR8IjuygFGAasNUVHjiXzVS
FuSPsiiPewba7a7PAFY/xVvI0TJy9S3U4HHSQfU8UbTSb1VW//6ZwZP8Ad130YIMgZFYp37Vq4Pq
f8eB9ZtBQqNeOMxuYUQeGoGVuNYbHSuqKQrTjPpeQ8NstEqKePUtjz/iHJayffjBl65yviE2b/0P
5gxlaPqcRsC8lhWY3zDXrsdkn2k2kIgV27GqcZ6b7eb+yLFBo6+PNF12cLZQPsv7uaCLSWQlFp27
mb3mjtnkl0hBEU8Jlm6cafzIFmxSh85t6g2CsgwNkXnE4AUWgA3IQDAR/ZtdSf2MaoN2H3/IYpJD
pmkgxfIvCbycgAnnKTLaeDcZpkDTwuRJ7+svdGS9MvdL1mF7VliAfrCMO8ybyKOpc/i/a+yzggOy
pM+iosZEwXZNkB/fKxOk0G2LD3//r4JRiPOyV8tUHqGopAaA6w8Y+bkuExIVEHJl7rWHTTkyFvvJ
mCdiUavpxvSkEYCFaNlgOtsM/zEm6Kj/TtgbjC2jnVI4LFymmLOLe5sPIK32KCdY7h7KHBnM2GWT
MuxkBFQSGcUcqfwNuNgLtmQN75VaR0ZP6KWpBzo8taBJEwP0upqF3kEnxoOGqcBB7Ve8nv4rVq2C
EAgsZES+rCo85FZ8RrCpMHZ3rRAESuWCZ303hAtnYyWQAYQOIkF//USe4j4QdUT8MPB2tvCGRx6B
+A1f0Jmz4XY3vVqEnNA4aujzqFqmSyz7eNtLCQaKQutUvDk8ESTJtfZeWHmhcBZuw/JtmUm8f24H
5syGrRyRnrcYkY4POYXxmL2sk/fS+iKox7yNQh1CxF+R9Dtwu9W4gpxJo+ujzj1/czeXKVtiGQbk
hSUH1LaAX27w5mSarNDZGiffA6zTxQvj5zXR+F7v6Q920S7TbInFGKEFtKH2NaIYYBH625rsyIsi
aOr/oVtcavblEaU3PWKxY5Avp8e2/QJbMbcPDw0JTX9V5zPPhlLukt4dn12HyfDqYdV/UQs8HVyX
OMnc9hwcVsK+a/pMx5oM1oggqUBzhKMy3b29OlhDSHVu5JrdIm8cgWqa/QbB7nLAQ8+tGkc30sAI
mdNx2e44djQFSGZ6NxEzUECKRhE65vXlT9CElIDI8PC11346lMzvp5aLx9Vff6PtC3ZQBlvKMrtS
+tmguI6wqBDhL94hPD3q6DY+xpKQzSh0kAHyAp8ckeye23wdMdfNPVlPyHLSzr9gLWWzqStZukAu
W0A1Rt+a07egbNAN12o9CNELotAIkdyZ//IEngnyrIyHNJVQMBF7OYIA5Sa3bUyMSRrrYuw3NKDj
zIcMcvs2XKu9WqQXfniNi8tg4iUwMLoAo7ieEn+QaezrTScaUxU67ULHJCzHQXv2FffzmeceaQTk
Tr4e2wGfqFw8YAZ3mVAG0rXI67jqjhg91zh7X7PYOLsrprUl7g30uSmOI8XkYXejWJ8JpWjAAA54
fhiu4wx9yJYWVpcZ4Kte+G+e0BCX0cBraFGlk3v7mzSUsnWX5KfVFsDm7qsyovQuWjEg/lMYuTVF
MAYENLu2pHWkSIeo9Z5rfikmHDuynjGOku1EPyqEvEpkSz1JmP2Zi6js25Llzxl2g05mdOkoecCu
ndy6yAm3O8qAFcXhP0Zk8iuxmp752ses2eaEJ0BvqW04Bg/gAg9T8xsgxhenqAkbDWoAvWIWbxcg
91qIIb8D/9CV4E5odBWYRfFdZi3cHVjLHgGjPXEXLP6vRQ45gPZuHDje8S6mTfdxVaBlEVYyqcJU
20434A3455xzrtcx756JRXZzkxkG/BBK3axmoZ7wvpTQXViu86yofnm+Rop5xwp+GtjB1XOCGUi4
m5I08JOmepyP4a0QLpRnyxt5gK8x9sURQvfMp39aq/uAANFIVtO4dFxskni9d21wXQfHP5Y+c32d
NXsK3vsq9az6YLNrj1Wc92EB118xVBFAQnMUUqM39M/YglBX5xwP5PJqe1JTM2DI13JYiu+zYh8t
2Jv/4T/QVAL0rEpaNNSQQTJSAlVQtN8AMzAgjNOju7n5ETK4nPC0cm3AT3MDMCuu22rxUGPr+iZM
OzCNRVOhU/CmTfTum6LecLe0+AybwDl+5wmg2hPPohJGAXWHFf6+Ubqgt2DJHRwO2XckuL7icTxi
y9BYrBDeI4+MeGM3ecNaikzRkcRyi0V3amrAbS9GICwZ3IbdjZhz7dvjibd2W6S6tCBi4TjQsmHD
OTY64ysh6CxPNAVjjyuV1iVrnV+9fGBMHRWeonN3ipk4YWBuum5vFjeKNWeiJDAz/4rri6D2NvD1
0LwegJhDemnkMvUe1su7K06QqQIoUl+nMam4dv0bRMyL3UpeZbOZio3dp9nYOqdzMKdlstNwO/au
i05kPIm3zLhu4lXiQ+YRFgRnNorYyovXnvJ9Jq2iVZIOzSjHPZ8L6GcfDbmc1F7TTaU7vR2E0Q3P
qiXF65QHeFvYIws2xryPWZUdBRxawSFiOVTjxK7jtAZ+TFTdb786A4c0UJiC/2QN9Jgj9LxnK0OD
GRzlJJmRXG38VdCscqpUQ3LRq6Cg11n6trtzsgbHv1NldxfDFlaFnz7RfqYwTOY/tM8Zr4YWg01Q
5gQa3ksh08DwbPk2E1C+XIDPgGnjEzXw9FjO5K8/R84h2CySAsHFwXsHW6Yk6yVmX+7GdNy/0Cvj
wdOXptCeTefR9Fh0jG+hF43m/fLihS66NKSjhiQ8Q2MvNneTpvocU1ne0fPuPqOXmghWw7gRyaSx
0exEXHjkLf0MdG8mlcgsg5HyL2HtRuoCAWZf1eJ6CP8S3QwhiN17YwaX/mT6izaB3lra8Ikbkedu
v8igxJ44GIdjqlo5JB1nRuvYqAMPu5N565STVsXz5mZRXbEd/I+5pssEjQeJdb7x7FJ287TUOo3j
c777cALRI3hWiVCOMd8EkF6gYsc5wz8m2Gqghwne0zb8gB6vr5Vno2JRT0hSl0ohD6MrWzkmeN4/
Q/dMFu8HgtGJX+BamDTwYTBYGBrNIgc4x2iCjGeksHsD7BVY3pThdOQXBYuYUxHwzSH1zrZhQuAp
+7933p6BQlIuI41V6onTIk2vp2EveXB3g3QbjbFn0NFmtnosSDFH9iw+QdNt9LM/kUPWaHd6s7dm
K8lLHBzMT72Pj0T5W0KF0KLXVvJlV94SytVavybvEsIDRWz5/Z5eRmcciZ8SlMwa/BIVqKFozKf1
gvvszfUITQEEW+8VVRP79ovWpFsVw8h7Q96sYFPuRRrtIIZ3kK/OtvYthH3+8S6jh+HnmOrZqUeS
toX2N3I8evRNpGoQhEwQSV2XSETlj5F3CCiySuBjV4CCawO+NzVYKOsD8UGk22SfUBqqrhePF9lt
K4K1skr88Gt4tyQZZoXEbncrCWZ4ZMO/MCArOImFGrf9Cq6Z1ryL/BHeoZ6Fx3DKdSxcIYObXxYZ
J64TCTBbzLcBVUxXQZdtgCh++0+RXRkv/nL7DaynBhRIVfNkMYAr3bTXGeoFsqu49mayhU7SiATa
30vpVlJTF4yPkVMdbNKhkfSgvv2sm4+5AZUXrVwhI6djGHX59r+smV4zYmAzXXdu7YuORk2DBlJi
J+86Pe5SggeFTcVijSLE28Q0V+aAFgNN8Fmv0xN3ryRG7WQjSDlx3liwR0cFL+MdOZ6lV9pRiGK1
QL1F0UtqeZvvPO4r28SJRJiG3/gcZ0HdgzrrxD8P85xzP7v/gTzH1n1q7sBWyS8Z5rtSOxQaRn5H
PpW+Es0CWg9uu93bM2buq2G6Ha9iSMj5arLtHn3obgDtPdzF2i5309ZTMfvVej/5Hj2E7w4/ng5M
VslcJHG5oq3BwQlQ26FdkY3aUS2T1mLOJvOnY8OhopLieCv+Al7v5e6ZrPzLU7LDL14h9RSolj7c
pvWOq0OVKS12LIDC+50PLERYfteeBX4Xx37lMIs4pZmgAZP0zjYaF8MTTzdCTcwjuy4rABQ3+D2u
n/dQagvRzbQian8L45MT3Z3ujiVE+MIRRX37Zzwysu4voZzMGHZbSSxAKTZ91pHIQYUkXuioRvps
v0NJcRjUw4PEYVA6ZCKZnIT1jo+ScnO6t99wMY2BZhqiTX+Wtj5yl3Lb0EA9aWJQmRLVuaMq1E54
oxdmsGHYr8LcQntFie7p9p2gryUNjZepJoJ0EuHQ6RpT0eAqJxOEpHnVLHYsn57SS6njLUqneA8j
lxk99B8UHe47kKRuZrwXhrki0AawPAM7Q4EGfz6XR0/dIVPio2vdzhir3TXGM8GqbqsEGLkFiNOW
F1NAE2ok6EhrsHMCS1440fwdHA7V0OUvTZJiMgtSm7rYa+ehBRQaaOoDw1rsYiW5+h/Pt9ECRIMM
5GfiprxAH3/l7UihVPum62F3pyE2dVO59RZi5FMRgd+rHaP3SA7ngGXUQRTmItlFjd4iMjG9+3AI
ZEafUZpV7SWpf2rJKn0HCSiEAdyV9NRjcYfZYaoUg+Yo2Bj34e+KT3srgoHYr+TQC8aCFiNDytcC
JJyPRLY1vhgnaUybm359gedOdCa7YjaEuHZ3MBFwE32Hq6NGB9p/8JerBaZllgzwyIYmpecw/cy5
yNqWpDq9LHtrYpm39z0QBkAF1Lzi5J9beYlHxMpp6A6DdFwQIoC1tihbS6pj60PCGw73Cieepp50
H6ovg+xXbXl+upt9Kfq/3qJ/occdkzbxhWFMl4pu5rRV2mMh+o659FYSSpYKBzP12khhCtmkC6lJ
6O58hUAKCGUo9KeGaHMt+89dxY80Xa9OBHrGbFASqoDgl0ZN62cZ9Q/G5zkY+fKEGnHvkAVk4Q9Y
npSRrDm8BlVAP4g3U5e+43BpY2cpJNb4R4wuRgzTgVxDERFRzJ/vaE3sNLJ57CCIopEz+94opt8F
tB6f4ofuUPdGP5vlEM5qQR2yRK3D1MflAmgBNk7Od4qweudKw831rI/9JzVvRoLZedk/nCc61AxX
CszwcEpXVk7ZIFnG5gGEHL1y7eu0ckXRVcnuJXqfiv3rxF2kuUTn6pUGOVsS3GgXo9U1mrfCRWBP
3x8Q//d/5/Nsf/0kKNo/DVYr54TlCZFp96RXtVtezzdKdRxl6v32VP7OZVY+I4Yrf2tYtPVOjuNM
KRtSZg4ZgS2RHhG7jbUzZMtGUhTM+Pd4MlCYsKNpXVH8V65x61bYR4+2TDpLWDvdlx34eOq1GcdI
q++cFPmt7+ZxO0bufvaUolVPMu3uoBgtAtMVkVhbGbX/w8xRZZThEclaAk7w9mD1ogvi5klx/Gaq
DAPo2AzNx6HRKQAUMRTgsSDGkdZp4p4lWloI5yasg3X7IfKTdy7/1OuOgXpC8/JOGiwMS/yMywgV
sy9S1URwGXo9Jnx9Ucj8PaJhnxICIxAejG9fsSjifoAWQ2UOwQlNrhlV3Lu4/kn6Q5VWZPzc8kyJ
14AKagZzpvv14Iu6HxPKwAeVABG2/otWyxl+GMSxQ8LELO5w11IgHR2MSKtXGG9CiVf2CBdx5LV2
5yhNlCVl+g3Nd+jShhGf0KdXy9zqSRp5CMfI9ClOU4BiUmAMNaF3p3F+agWl2T6R5qRKF+0iFkZg
qJNri06DH4mh0a40IxbaTHncD5tB1KrHmgn+MPG3lYjGMalF93qyGtTn9BGY78PmebA08YF/kIHr
XUj8/+In8M00wtQWRgxrsWomC7TDhdW70mZbaRgNTZ6GIBCN+dl183HRQOpENM8CQcTo16LS35WN
Uiwp9LwyQWKbsXViO7Oxb/AlaGpJZ7prl9ESTL30n4HlddHceZszMoUzsGZ9Z6zR74dVAQ7Kiex1
OdKD6c1HzzxtvfMw/3SAoivk6mrYTXjeqSYGLlMDlMtS7XmTSUhk0xfXZWTDRCaCvtcWZiNaEIM/
3BAB3Jn0J2yhPxs7v9fPWtxGO5WG4e152Y3PhBpOe/PeUfkg6Q7wLHbIWUpKtVpz0cvQdj1BFiSJ
iJJ6TZuZadFNnqlcbwHTjCA6jEQ78iHdAiY99xvcg2CloKNYCE2pQGt1sE/Pz8kq2b3DspldHIUw
cogjalLZqrQJ2CgWK/CO4uP8ZOhQXSqEwbG5HkpOlvl6YuXD85RE+539GalH+Yn3qKj6S6hfgHx9
DMwzj1AfpqzyqdQ5xANcqboUv/B+E4ou4DKTprQzIzQftHpTQj5d69z/6e6VfJ2XfupCGkDrG8jW
0d/6IlQ5YJrwgtp5/QQMnLh5YgHxIa19/pOhkSPhU2AwAKgMEvN6izg7FKiGX3hoStvSTkzTdf+8
3jweTJBKI7s0gj6LyBa94o3+4MLr8dqNVeCGznjgs/rb0dyG75vbcbtXy1v0oIaIgxCf1dWxsgRN
IwYtc3VSPHLhl6sTGCvzCnzDeQ/khtl/0ml3G3mmhbZT0titDjkqP++XrP7j41NSgBG3ywePr7ES
m/5pRM78LO0ZHog9/D/zO5AHhxaMcEk9XqsJutoVTb8kpibjI8qnXsznyNdG6ni+kRT/kdI2QPma
MAy4Fvz2+X5ZyqtaTT34L0XSzTnOBASdjy2eNkQNljSW95b7KX6mxfd8x1pTKz+8z8TtvAfLrNUr
p6w6JtmJ9haXKi1aTOgyoNqKP9j0jyCI1ny2m9vbcnqIDGpcudwlxrBHMkO2Hk7bvAaVettIPyRF
c0QJEQmvhJ9M0cSMlN+9O66k9LXiKb/hRoVOFSGSfuQz87j9GQyJOIwMnNWC/8IPSJ0Pau3QZcLH
/el7xAGE2uHCcSPxPhBNLhnOi1ZGmPfnCPTPrrG118xEZ2cWqznA9+hu+SDyzJ5Rjvg0PMAs/NQB
xsKCDz5GrO62WKZ1wWmBLWkorVxLB0Wbv0oTanJ629GCe2jg5Ure4zo4KsALOE1UsJbXWbtXviph
fOwAk3576eR8svvHkZfdJ/VgCRn7b+eILVFtTchfVoitkfvOqqpjySbXcJFFGLXpIiJ/kJKbzGM5
vF6x2APPeUa9O8LppG8tmvrbnDfRFLQvtO8uS0BqbXwiUmOQMe8pixkNk40lWY4dfIkU9LZq77zt
Oc7cPvm3C7gG5Xy3wxRV5oXUnhTfZkpmoeFBFXAVsSBsQ+M4mBGpvFT4B7KmanKm3FslDnbX00m/
L2Z46H/PjXyqE44tlRcu6YD61sC6tuksPznYws9EcvAVOxeiss5ZbPayLp1rTO96rQmxkoLhTir2
D+WcE4xbDI+QHcV1lXV5Gto5+bsxw/jP+n2nUcdJ45SKzBw5aZ3TIX7l0wV2+BaNua4Ys+RySKIt
nBjewQ6gUySpm+xFlcJ6zlCJw1jBlOvzX6axqb7q5dfiLD4sikoctPaf6ruFj0fBMXr1GtiVqmcQ
dkrZYlTerk7maB1v4LVNITMrk+rPFxqXMIZuUhX1HE64FOa7NcpTp1TwgLOz/HguxVFZCwf2QT+p
nBEdWmrw3uwua6CIVX4z9fbteM3HYqVPcYLWWa4bs6vDruKtH5lv2C6js63VMLK82hKcc3UiPVaU
0/cF/J4e6q8vwRh5j4BB3MdH8lWrw9v29DOUCJOj7uV9xVnw+Mipo7LQf4/z1zURHXZKCJIRDe2P
W0pI0QtStJ4+A5Ucoblinsa9KUXR+TIIJnhPpp7LUEMuqQQXDjPI6fHHxyqetk4zxgbU4emuahj8
EtMI/WsCAgnH+4mdYm4Pht6HPVthKWDFvlaL1PLW8R0EbsD6ojkxlgMMIuck8ibexyFlGsdHcJvT
YGMfjRtwYh8S2Xrz3YUJ1uaIdhmyZbjWrMc8hWwpZQL5KKwgepSmAysEG1yoofIpw3aDoPetHBPf
dbPSe+OXZMugZ2fAZGmF1QpiVlmiDtKytrLBsebm8iF51Gk1cz45fIar87689vIHKyzxOfde/QIx
ypioTNq+G1JCLvR8kKP+cUunVDqjWMyEy04pV/PdAyYV3zie7yq1Mo4jUf217DB8BJCH2yeDYezM
GJqR/fdpXRhq9tLpFJf8y+Ego3JtRhuyoGR0cNh9gFrPVoMyhSRezcY4mB7M3vXpfQHZZ+TLG/aU
sZU/C9I83LTlA5xCsAqzdAkzXonVvzaB36YCbolizJNLEQLA5AY9B/1C4yY07npIuUp2IAldQnkD
PTM9+NahGOwPpN6s4KLSDzkWogXZtlD5X51RgbRJpLZ8VDaRbzP+y/ijrdBSzFMiiDR9aJ7Vhhyo
wg1zsgv/558qiAcZ3hi4mHP27IDM8IRorAEKgnaQmrwz2b3tqlE/nD6e3DoH4MKqdqXqMIN63EyH
5cQ9uQJc+XIzf71jhRzX6RGfbrOjiIDfRpIBNtSlc8ueR1ZgzUiZ7Ewsf9h9R8wikLdHQi6lvuzw
kTGSs5e2lSO7Sjzw8VKP++Hy5ZKfGf1Cy3h8npqtky53Sl3A/qkasn/Wrpk9HrIdT+qYItOpamAl
qfR4wuIURbBXZDTPtrZZkpE05IUcysRWba01dpxxJlBn3uQ0an2VtVW4FAbfoBOYh15oGymHCREe
fPEHt+X6TAbV65ZwNOjK3KmB8uHF289UgAl5rHkvXKqjvy1lEHoNtEeZFrDXY+q7QSzBz5doVld8
7/LygzC0NaLTa+UZMAO5Rf4ywnGoVp5OwjFT4JiISk5IKZbf7JTESf/cmiAgtaBg9haF8utDA96M
i0lytHl/YMbLjkNyLlNs/JPzrVaiOyh8fu8vyWRh+rBmqsgKXhmvngYfE38Qi6OMG8Jpox2vx18M
VKaZPflv6/uqR+X7FnburK1ExHlhoLJwQxjA8Wi/W5t4TyjPb5HjevHP4rXzmxv9iXKEI+DejfPb
I2gEX78t8xiyWE6+6MbQFEDf+arwTCTpt2jpnnnmkA/sJD+VcyRn1Y52FUE8K9jHGlvKlxaigLEL
HjeYAzmTXALcXmca9fuotyCoZeXkIY8vFWgRHqSrbw0WGDBaiemOlRS7Ftv229k5pdQloq99QWLf
eAUezaeLapW5F6ZzfoHFwyvNfAvrQFMK3lyamGan8liGKVwHR5kEhaDLTLihL7N6O3N8y//gRMqg
G/1B5HdJJzfb1JVMV4QkWjmYeebwfPyW4NcOaHwE60ovFayJTRLavfJL9yJrCYETS4Q17zVgBLWW
GPSDLC745SyWErFtiBLWBqn2PzsOxtTMKmjbGlZpGBTWh/3Nyr1QVD1Zs7Yy+2NiUSHBZcYn2BJp
U9+OTjBeekaM0w+7C8YzUOV+Nr6BoanC/gJwI+9ukJaes2lUrCC5T7qWtzb9jAs49XBzZ+h4M1EW
C2UkCekyY4U1r+mazABb7GoEbw74bEH/U+QfOD6gilt93Z0oMQgqhsLz2SoWnRX6ZO5YlAWYsK+S
6MBEqDl2r/4adBAKZl6eTTG4cpVKcBwb7Eq+CmHTjT7Inj8/2HsUQxR51iGJ8DzX7kJLnSu0UmH1
4Wr3dyV5OgmdQDJS+Np6lv1Ekw/ufgxOOqemAQkVmUjKpt8tEH/lOJozhAn2DkZ+5whpXQyOledc
moreoVy2I+sRNVWbPoEkkcEY+BsDe7e3jo6DcVbMuOMtoxC7+cAF4UkNlrxkcsSOEufGj9Ymjb97
rWdzgoA/wevjd020xcH5679PDcDMi1hVtLiOzQ/DI851UhmZqy10Xvtbk/vsPDGMQ05xJ0uiUNTM
Zrtvg1LjtO72jErgoDTcSn2vi4abN27rAl3o1bc/OXq8pJ7UIpmq12dCLXJrUKoPCT30GnhFJ/sQ
Ll2isHp8l0PE34M2+Y1QwEG0WiixeAE8zJBvxavhuJ/oCCye9Bqf780PMtZjaXZip65UXTfF7Ngd
mb64TobfvYauOkqpsk3tMkdI3+asEKZcaWcA0I5h3UUz9HO8QrnhcnRJTqCQvI/RppdZDHN4D6+2
iWMUUX+jZak7nLKWsFoa+h/8UV8rkB/mOkz3xTwCo7M34QIDEEonyCaakQsN5WJZS7wZqsjbZ/cE
QXM++56KPlXXr2LPCYW7FsrOEp1vWCnZLXkGFzA4JHpgukfNG2QcZS58owx0oLw+GTSk1LRHdQ7A
NpoGralBVvEV455vl59t6O9ZAiJl4TWXqJcpOoGF2YYh/lCsNQjoOvNPq+ipp1nZDjVFEBXkfcq8
j583anx5zy2ghpFynJMuEg/qLtzUIyxou/ern6q3ot+QjWw+iSxAKUDMCFII6NmE0BDYPaRFuuzH
bx2/HieMGrJiESA5T8K4MhV7ZX2pTIXe3h61XYeUnuhTfHmKqqedC2/rf3igtfWDnIoF3yED5Y5Z
1A9gmq9dsO6Gqq316UbaNzOrqmUa5zkBj1/jWt9GvENA7ot4AGx77qruSOQnU/VF/Q7De4oKcDIT
8h+47oMqFJu2SWPyM/3GpQpM/atsLzORfE15H7XTfUmFCqReSVi0mdCZP2+TkxtB2/WDpSXOV90L
4Mbj/b3ViDDpVI4Q5wnRrTJjPob0PF4A5Gc8mPlcPx6dyuWHS4lztvGKTOP7WMU6g2SFzm6ZrV2q
8GHcMqV3xD+xGJA1kiADXT8M5TB1FMhRU/1vBF0COznmbybWPR+gb8PM8jmcvVzrjAo/AD2DphDU
OlFnFEjEjwT/KaIG9Pjyc2grZZnfEhkjEKJOylcBwpy6hSlyGTVQwT0ujVwhujAbLm4lT0E29cS2
ItGOtBbsYqJr1iNDWQd3zfEJA/rddJD4vH9Qovktx3fA0TXnOPoZUQ2tV/rRLJ3HLF+Ngjo14O3C
ZduGeoUvzAcji90EUAB2WFMWILR/4oeIRif2bMZ1z2AGSb1d1PCFxWDslwzI1LQXOIJyUTQjIlZN
N548t6AJ3dVIe0jhCJV0TsDRewdiZLe3NqX1PItvhO+2Dt2SWFvwAhGA62HW/fPTqir7O82/uFSc
Cf8qrxv5re+9WHj89QcupCNY+kxu18uJFoX+dIGP9bwTt76HOrDk8sik/uURQ9h4/Yh3lJLc2QBe
lZCG+7Djd6v79BM22zixmDJWk2177Z1Ef0XvmWjiXdEkxplvlizG4waiKGKxwRWyxS9M7gbhrYKQ
RHJLw8sJidJHPSGl9VUsgaIIc8r1myKTGVI1uJi+6CaruRJNHWLnRXGtQb6YoW3+VP6KIYGxr/50
/npNrra/s95Y8OXD6eGxf+rkInf+0Gg19lkCRYjcIhl1I/uXd9im8aY8Pr4/l8yUCc9a0GoErE3h
DMHGd9sU7JYCySEwZQbVco/O89MQMvqTdWA3GVQOPFTlq+uLDkBZBdh1V5vOClihlByLbCTL/zc8
KaarXDXfjyaA3J6QH9UTnItnHcXruI/Yzc7k2+jXfT/NXG8AvlsAISQMxLTwLgRvvG+vMR7KDUce
G2iLrhXfMQ0ezXx+IWKs9h7Mq0ZP8r+f36KKV98lahM/yGAvG97na9xTI4ByBLFyZOsPb8tRIHgo
Z8rwNQ0Yz8299vLgwnrIQkvbgG0lpMisV41Bpbu6+56vIyKjFy7hrOQIGniG9BU8qYsGEJ382jVu
mpEEdZNpHpnLzFRH9EZWY1g9pX56enf9mMngygJvexd148i/xuxLLUxirGCHFGxLbTVzkr8pKJ1J
iKYFHbkRXGG5+0wjU+WZR0b5TIRNZMEFxx3Vg7nmXDVMCopYYIb4YNfPJxicB0LziCt5ATh8zPdL
e6bdSVveaLAsD9NTY2WQjoS2n1JIVnIjmssNq8vcIQVppuesCzpr6Ocgz3FJT6Cn55WL5HO91OwX
hjTEZhEYCKxP4KMcycCFybNczlgUIhLH56m35hF5O7Vn2ZCuTGFF04ezkljZU3eepHnzKdAsiY3w
F1EYuNDDfgV1BUGA99mkuUHSHUKCyQT9+bMVszFUhXoUiCcAes/kjdnaDn3RnfnvDrZ1WBzrSxFr
dncTrodiEXkVSV/p4suM+PxR2j0jLOaggAgA7xJvSsHj/rUoKT1DV5nQCKpjWhHaEOT80liVMo+T
UoylEuKh5/osRJ+npu6O7sEwjfLtVDlJJ+HXnKRfAbKeRYjkEJkqkaVqAVfkCMQAB+Wdq5oLUAhv
nnqBaZFPOUkJ2KBgZgEvkAnTvK2euox+gDqNIKLplaMB18aYWxD6sR64Ijeo8+8vOXxhkpri2qCk
izJZ5TOnuFcU2j21IK7QqTGxn2CqmCDZMAAI8h/DqfaZ4I+zaC16A7qazSC9OnvuxWzszM7P7jb0
/HIv628Sg3zelHsyI9P+/Eh++zXNYZYDqRjgMx340V8tJnYT4YfxXcgHJroUjltiDbDpazO1ixQ0
C6npvilKF3FLn3ifm7aobKpbBhhvxEhvj/DRWqbLyLtXxSX1rKO2H6mZrgZa5dejOCWiVoclXqXn
o6aIejYzqhu9d2njc8zyvilMzBXF4Kaz7+pu0rXQ9fJT3yMm1SmcDu+BuYJTmOv7g5MhgD5KkSkK
CihbK+zk/bmt7LlwZ9b6GYYGfwe/aTmtQoqVXbVTysAK6YFRV2MHqaBMlEkP6o2BdssjXr4OeT9W
RZpR7TMnFTGYVo0dxHSYoZ3dGI+FEO+mJWhb18zuyao60tSRgFW6euRCSS5U3e4GiakT9W+rrTxU
UYFA86sYY3EhSTKFbOvBw4bFe+prv1cqeVhzznQvfsHXTsi119Z6H5vgGccSLgbYHHyviikAu7NG
s/C5U/6uVwtT7EBC4l5fQdD9B6qZKK/b5um2jaFdUURhaptMza+eXorhlFMukH+4kU1gGc2IU2gf
r2faIndeH9G8zU6DjePfhA4vjkbOEO0dZepfZxTvzQZ7+XWYBEIg8/I+yd42HWGCsPA2h37UGCFe
b/kf6xfHAxy+rwAYXSyfLzqegvy9x8ph6RP+Hi5IhIBkVLthXwyZLXEsDvHG5m++JhB1G75f8MZv
zy6eQqQZAZfgYvrSOHYOgLxP3PEbv5dmPIFLkZQsdcdRSy6Su7SgvJntymEU0Y8kTy1/sy7nckhG
VYmUVjPtc8FOoyZ4mnxlDD5ZMk4vGVE2XW8Jss5wif0rGMcyfHK2EHAg+YmSjJQyFhVb07QKukc9
8E+KqyKEm39eYUWsTJPYqXN7rTiMpjT4ugG6i0PMWMwCO+KEeD0MB+gS1lSftihdLGEpxRIb6kR2
V+PKIzKvJMYJKvNZpa3VzO3wgJ3V5YddRrraAX9GfoRFu92wpFviMV3wkJsAF5fcZ1GQFTrOgksl
Wn2/McO+pIVRifDyekNawxUeIsvHgrJKb/ZNY0CdgmAd16y/+GathvNHaql57mxTZy0RmKNjLtid
6Og9S1Z9xg4cVcxcTiw+dVq4Lpv6EspY2a3KGXMuvrFDD16FxIshU3nceOCC06NKDXk2x2eJHMKn
XmMtP3CAU1/NVRDQQ/6U39sHD/Eb/LYDkjwpkp1nM6zLXJm1C5ex15fB/5PkDP6nVndOi3ERTGoW
Q2QVzXUePn5aWV3NbmULYSVeTYEDP0XoHxK573oFMQp74WUABb44Nmm1NocG7WfSKkFlLBcEqNAX
O0po6CnUhHiBwpUCJ8a9DRDd3HTShnG1kxdAQU53NAXss5qGe/YtS+kBQtmFZ7DlU1nZR4ljedk9
ZR6kb+RLkyZ/qz1CQNTYiosU+8wjIL9kUfuXiuseoiQSf26yVS2y+xOd04MzC3+YW8TQWcd/k8zh
0DBA7VvMdEYEyiBej5QKOEMtu5RpB1Av5hAk3AyW6a47VtQPYr7UN9nGk5f35LV5zqzFUAInf1iL
Y35yL1PsCyZrwSVgh0mIxr6NMWMhLJpFgia8Yan2qYEn7uiGnRtERxrGh0wEp5IqPE5Uf3FJPNYB
93EU3YU7sP5yTaChmSvAbV6GlVW386KIotjUZQzpoJ94oRqdrraOIpSwv9v+FHsMXJAhOnQlQm/J
sM8n/Wd0sCdHW/4dt6v4siwyVJlDSx+oVNAKdQPxVPC0EJjGd6sBZ2HCW58ubq7UEaax5Ylejl6V
wkswcBzKJiaomnk8wrchZQWUlGwWeQvES1Wo9kYA8GoK8gznZ3tCJbvC16LJeN7A7U5YGtrhB1Mp
T48GTTa6ralgbYFkdFRaHpEJ93OorXV57qzllSw4VvWjdnDwkcSyow9Yj6Zuc+dycrYLNkk6siZB
/fsW6cPl0kp1P8+jE7X5pwAYdnC2+vS5h7TZQznhX8bnk6sHHwm33jzCdH3PsAYgzohQm+HjaSBT
Hg+vZckIxwIiyiWuXQ4UxWNOjpQ4B0msSsyk2pg/ciA3pmVuNloQ2kkDOzkvJyw3PEiLiK+iVG/m
KxUU3mQW89rxeO+JKVuPgKDlrgKoDXlaLxe4ufB0TdR7l/9tiiasn2A0yoQBNwtZQ4U3iZ3dUAly
FMlolNwAzNA3HvtbZHcCjnGZ60OJXKEDY3DFzZ5Sj2Y0YnZNfn41jirLU6whdXWMPgNKVqxGLIh0
Wu7SrdYEyYInh/5VmV7yZuOFUcfu47RUq++Erg9MWefsW1faa7jEvSCHsZXlGMrzrR/WxaJwquxq
fcrrrkOxYTHWoSGkNyXw8AlavaoRhzS8fNdyeJIH8m/BNKL67FcjNghFQdiCF05n81+70O8cdz84
wiCkn0l25ZTXhhVmbDgKXRCA7qUJyRdrJgb4/+oZW48CLSVal97d6mPp63eNYN8TDkvveXTMSR03
tkk/uEIae0clSJJUe927LOmH5hJV45Y/JF3cgsGL2Pb0iqr7FRjzIE+9olWUD/5cpknZeNAsoOSP
sQDaX9YjZvOCvHCfyhhwtzJFgPJZv/Tc5RSUNi9tLvO+YUpc/Y1Iumiik86jw74JSDcOIZWHGVGP
Aeng7kkBoEAiQQ+WJ7+ey+v2xOvA2idOFWd+/5GyalRAAYsylPNenPoSD/4S/KgByPUxh8xZ/6Eb
5bKRQF2zyRFlRRRKe/aEqmNAydSjsX0VI2Al2J3Ke+lwUhLgfKaWASIN8JSTXzHqgdzJ6zqJhwsU
OlQxiE3omYf90OVL4T+cLQoeWv95ZXOHRZZY4uMmz3AMKeNALCtEc8OJeNRkAZqq+XSlgSObVnT3
qR+HKhfGJVttmoUQXoWgpZltgK+2bmWbfzqEmw9SnVlSLT0LaFSDavnkdpEs6yXWNi1+6hKo+6Ps
x4bMUCLeZGLf57Vd9wdoDHxwuwejZgriLTe9/9StvtQprWuJW/7xeFntcscf+rriIXYaP4OjdVts
JyW1suqANYgUka3/2vuaJGbq9pUGIhuU0UUO1GepsWv9/xUYAo97Nf0dsJKzP/9tZtW+xZvA+Pro
fh2mKBhC10KkPuW5CTboX5KKHt4CKGF7YMd3CoXjaT7fBvdgqyXhcW3agPlDjI+P45yfMSXaHhaX
Qo844mFQYzX/bmZNFttdvWb72EqqrP9cHMIf+Dzlggz8Idf9djN7K8doZgt6HhTljeLwukvagoV6
Mw2TvnCS/wb8afZGJV3Ek9CYaKjja3+iJDwJm8fAEFFkqzNUJK9ZTGCbPOCRZDNw4v24JgXVGQdI
82SswDbRLoshBRJltG5j0v6jIg+5j+QyfFqdLluOBVEgZvF4eWX4dKt7SJcqebu/bouLTBHi1I3c
GI56Ylvfuo6vQnDZ8CFSH9kjRHbrrISaTOAAfbujdKTEP5rLKDAfQZ9HE3ysPq+GbfwuNBqip33d
YxekEmjIa7S4U8x1FE2FtTtxToDrxUfM3OnoUrtTysBvfqUDoHLjoYYWOXB8aRQqfl6kG3SJjSNj
T/uL6Tbwy7MPGoveTdxESake5UqQL3Z+1lcWPYOi5LJQA7JWj92Lh7fysQ8g+OtWAswpFYjOjRxx
FuCMjAEZsoQhw/cRvP3ZXNRO6+wrGLxQLYHiSCRoGOQRMs9Y8hYD/0d4S7LL28g6cnRv2p0BMByE
kCWlUFgRfTW1kZlwAORepW5FiwWS9mWnxBjOBqIFjw9oG7viwhxE0y1Vc/DcVXEp0EEetn3Q34qB
e6wcaBkEDEcW8/aoEfAU/wVRDrnfbqp9BEWM6w7XVPopQqv/stLPRJ7zzfsJfh7w8bR408bVRC4T
4py8F+hqKDDP0rFdzkJ3Sqg0FFy2abXTphC9v0lyrS5B/HWyqw5YTRzNvf7CccSa3O/8tEbvqPAB
+wJd8LoFCot9GdKO2wxODlxIo7Npz2QiQ5jOp4IqiJWCBPDjn6Oul4Ia5mED2dmVJ8dONsJNKgdf
TdqsMjBXfOsiAodgbEteFVkPrHrnUrVNZ4yqtdZ2fyZ7EfewZb8pYpSTOTDTjdpvRr2mLUDKREEG
cOg2JWPszqOuieQIryOKbiIm+AmUakV7NvkaoiiQgpkCMQ4Wn6tTOSBGFdgGbCDvh0U6c+6JkI/l
WI4siAcfyTAo/NnKI7aMGcf/E0sfFij89DIcyPjeigW9lAxyHatx2JQo9JEyzbOGJzaU6/Zy1Jg9
2fo6iq1eNIwbdGIiMjMKFzq4lc3w6ciyzxtp6A8inGwOWc085LS8WMV6ccrusPocFMqFC1S8+9na
s9qgUMZXQY2tI5k+i1Xv1LJ44RuLv8ZQMf/jDJp9ysrj+D0v5bJqq5dWdzxlSMSS+XH+86xJnJWc
LNu8AdveVcUMFHPY6byoZd2/QL06oVsfFKxMWQiRUgdon3Jdy1MBiMxe5GrNmEDXH/BfCXUR0eww
F2ctDcisPRiMtoc8f0CQF3QYbw1lTE8F3UzMZ6mLVOddikCjcjxxTTiNrTh9wtej1y2W4UM/yTab
CJ+PbL0mPHNjkxrPC4PZbTPnafEji/vJV3gl2XHL1Uo/L2J2wq3GRmSHQ6Pf3Dx8s/sNZ0FZS/tv
IWtJFfmmev5nNAuZrNlYuSgzmcs+b4OWlyWt1n/nqarVwjxhi14bUG/G86C5HoQKC3Po2sexD+zx
GguleJWDl8rYUFQxYR7WGPbGyFO4YhZLfPhDYevlwWvlu22JmATu006hVwB/ucIpxIuyUxZi9Mnw
pMNId0N2V1WPY6erEH4qmopRm7Fv1znISQBNtCj/dtSESilF7iKUBf0wxPXOjqUC85ydJJjddhCx
txvkms3brPjNODwp6In/aPTpyvoxkgel5O6SDtCSb/3KboB1RgLC2ZMhqdpyARDcgmTebjDzseBr
rBIwUWOjwW4AW85YcdWLi5bQpT1L9O7OfXiC9cDxQEhoXEvy0ceiNprrvrjoUVC2jG4Mb9N8swVw
aCUz7u/nHA29z+c3FdFnlO/wXvX8Y13LMe/JkkNuZRFKiGVGOef4dUuZnIfl0jqmEzBgM9ATZhaS
u2KdqZsaz9Dcd/FWy5VBP7E0afrkTq3aR63//8t2VN6ezOpNmrFREUsnlZndEH6I55Qb+8maE0YT
Cs/IwnMZxMnPf1F05kTUlPg9JNLtyidV64wUQLCd4tZbLYBgqQSlDt7tvTCnNLaR+SCkGBsxBnhw
B9r9iUI3gylbAKhKcqfK1qZDPhkrDCuyIYnQ7V45EZxPPD5B8erjyJNR8sZu4V4XaHz7WAZuj8lC
oamn6tPnOcVAmOmUdf40L/g5SsA0QgSV6+v51UP7lz64j3/+28U/7KFlPDXYmZifYSOf/xrN21pm
Z3A3qYdsBxNYpSIwdfpmw+5jgZMrO1Q3oTBXGY2JmIQz1cU04h5ZsMk4PEHjLWI02F+g87hhfczS
Kjc9gg22NHytTxNKfAZOElTKnC+5Sz57IktEzeo1YB1O/e5avCJxWuecwyxa3z/nMlKXdKBmXhof
/uNPEPPR4OU893WOxklQ8KBn8+pMiRDZShVotuSR3kqQRytGbHczgYOoVgn6ECgrJiazB+Hj+QLE
/5ZIgkJlhdcYQzyEOi3EIx7VmndNZEfbYU1yE0qy/xfZ3xxN1R1Bc15AisotW8LzW7swwsrCSKIE
34dR8WNTHow5clDOopj/S2EcUulEJf9f9tE7zs5lmf65pS5K4apQecH7MV/bfHVGh1V8QFVcbuMW
hpv1HYmz/uRdeotsPqdADpp9opAuU2YHh3vcKaJuXhmaVb9j60inVKyRkXE2aNYhW6osgbJU6PQ5
IOnL3sh22nEf/FktEhxOMAdvooE1WI0nfJQCyPQm5HohsbkRcEmKCUyJ6Rx/jsgCH3+q39Yf3X5b
p/hgzzEQ52LirdiDDAu06lMqog9BrZGID7TjgKBqkPhLan1bT5aOptTxiOCLfGi5nAKaV00mLkck
Pz4g7wSg3dgXlvk0E7Tajkp+BDYaZzckGFXu7Tkrs6cBUZ7GjqxJ+r9b32nhSwWnUiAIsh+O6GFo
18U02610dYfCr73Z56CW15xdGYYnK25FjI75epG6nq7sQ0dmZ+4HVGGXA0FnfTo1dZj7Bk/pyjld
Hu5Pct2heYmyM0/iAA9H/TBPmZ6FVIw/2o40YdlxvslZPbaSlaYULB216k4Km2NtGo1DhoFZ4rjx
oiHTqUcBEKiqQAuA+2H7avAmFxBsgtF/K4jU8yDyMF/YlmZoNHYqbxn8mpykfeuYj2ksfwdTNxIJ
R8u05xDk9do2mpvrm2xp3VT7RpQG5t9QPEZK3GSPlUb6xb0DN0U3/vvy5vo3DvOzYYqhz+YflFOD
kuNmnEau94D0ZwhivULzbdPlvlVIYS9seliJ3C5i+adMVqTdjREltrG+z+6hVOocynLQcZvElTe1
mV9DIdxkTp9KyA/htddRIaxv40JmjRsMI19lniad7XjvdU8h55N0TBWo0OFBk8lxdnt6c6mUjPKg
F31eY4TqdCoT0a+ap15ehAT6PG/hZ3F8hBp2/qdzvKr7lDXzsau8C/OxKwhYpc38aMFNHaF17UJa
joJ2wdEUBJk4KP1MM31of9eDENOiqmaGkoNZ5JZXVVutOtzN5mmTYigh7oPMfbFtukJ2QI5s++OB
xZIoZW27+3JLzJsoDHn7rPSfi3oka7hdyUe2PI5rLB9OoGRspJ+DgN2xbrkLEdIMB86rN8lD8YXK
s/S+X7yWcnFol8VvNMfzzc14TNVGQRstDh6X5Z4/8nrx6ERXa1287Frlz9z3B28RkhnVfjnGkxUP
k/iHqPvTfp7pd2BD6VjzYOdL27YdwxUtwPc/5ydoBRwu5zFeE/Zyijxx1SpeW8wyPfnWOXRxQRAQ
joLDMYjPv/0Zq7awSVwxFo4M3SwhgoPMLXFx4aVjxJ+foigXstIXA9d98uc1Pb+Ked8oYUVJXNc/
VAlD8kRplIixX5kBPKfitmHeeoOteTFsn02wfg/ebLEpxhqFPoHxZQbn1EtgI6nr8N5oDdpwMV6t
WuB56gSirSL9xfAWCwvstg02yelLELpMtAMmk6ooMyJnrLJ1HTNOqqxJl6OzhKPAtV4Vq4E3rafq
GkpRI1fFqFv/7iW/PNhvM9dYOtg36f2UJnn+tUFvMdEsWUEvpO1rurS9wV4NXfnwchPCVzsKsQmo
Llq0ASVSnT0gru/VP3G8LjUMdo4ox0hen6lyLaWLDkYc0+XEbu6GLdtKlJsRSwlmZDSKPjNgC8Dy
WEZPHsvMPA5bkAODdzXnMKGn6vn0mdcbuSRxbwgxPimHQ/w1bcww6WtI4pJlQMsndy1n0sZ811cK
MPaXaMV6m3/4VEqYObwOZaiWnnOBVGXViYjbELLSdCIIgANtjxkRjbZcJfWaHaWjDP+L8+JuS53M
s0fxwUFZQ+5g4tONHRtnHe9YwZcdvAHCssHTiGWI7VHsVvuOZQqfRNo0NKf/APNTz5FK+KxcJHO7
PE+wT+DsKHpW69Iyr0q+fvhQhEAJ+Q27iGEoazli7vdNm3sIVAilZX5v/2X/zd8TfF+bahHR/t9N
HxJR1u4GmRprL8KeLfbFs9er+V6gK6qLIPee0dfGftF5QmSQ0yw3YjdGlDoHW2GK2CYaqk4tmqM5
zJNXK8fAGc/V4bw56qYJwFyC/FH+IrK5Ep+sA0i/HxI=
`protect end_protected
