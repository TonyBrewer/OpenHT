`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AnQx+YisHvu8+qMZMBolFBnZkK/4WYIvco6pWtoNekKbreiRAxVXNyHJfpA0/mNml1xliXfkbARh
1+iBmBAGxw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MRj5AQpaBF32mUBwzcRBZUH8XTwoxy0gve1JDC/TOV3cG0jaTjXIMCJ7FOxKW6ALUDRJQZvQp1S8
6er2te/OsPSlUZtwzXrAE9zHUSYpDEG5uLTYQoj0iH/N6SLBsSLhN/74el0vZhLHLXywIWWHqdgF
eKCPdHOQUJL/PPNarE8=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e3PJZn4x7/INNKY4DbBJcaeZw9sSYfPF4DPYUb9XBIy8eTg0jUTwqy2FVWw72N+Lt7UGbu2bMfoS
fNBY8oqwe12Rdu+a+3997S2De396I3Ql6GDcCReR3P+KQs5L/IRnb975G/56OG4MpzZEVohk/xF4
ft4kUR1oC3Sv+B7ZRf7qo+fgYDyA9jxThnwzDuiorvPKsRiQcQIbqnsv3FlRVdquL3rp1fDL9nkD
6sAXwacF4Dpx6oQ5q3IjRRgVS7XSebq+5FMuOfqKRd5H/yimRVEoFOS7a6MaGpxt/jwVfvJYTxhx
Gk3nK8HQ5nba+Njx1JeI5xKazy+GmjmI5Vdt6Q==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jBN92a4iTsybRj8182b8J8h3EY43JExkAOZXods+TNlchqrzEqta7VoqFyFAacFLmDttuI42xmgR
48h/XyOcPuWNz7X9fkF5rf3fhj7UWSIIVx/tWYV1f0sIFhGqjbzNDegSFJpnUtJN1ON6XGF7tWm6
PUeBLkkUJ3DBiwNIJdRx4bQ8Fnt8DHm9Ssyl1L2tc6tKvxWRGtWv/4l7QUE4LfmbOEZv+QsAe9fo
x3zHemiJoQVz+AMzevKjM+pC36kXoCdKzVusZS0j/c85is6YKInm2JEE1dLY2fGqfSrURm3uJWWH
PS9XZpH+cQT3KO/0mbSfYBNPnTZqANEvMSUatw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tqpCEM9506wOlSckZf+cvJXwZSri1iiVkQ8wMzFRN6A+Oq9RPagZbP0GVieSOFIHh0EIVLCn7yhi
3sM9LhypgGMLe+XTUUvkW4azzWxywQZ1GvjMSwf0/4UoHvKkMkn2DCvbAGLgady4Sxw3xoIezaNI
ZKYyWfdm4QabKlNblcmjUhBR8fLYH5AT38KDy4jbNSo7UnLhGZ8jbGwOwtqKWeudP+WQPzI9utWw
U15VOdQB5eU9Vnnjww2InQYmlg4TZR+blJsoKqke7dZpzgAsgrumBDI0FUObkqKNfVUd1LWq1S8s
I2hEW9mw6+i7fRkM5Hu9nCpU74jGmAboWY+tGA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d1RUy2wwOEnbuF5v9nQkfuj1khqrwFSDbJpWzJuNHrxz5wlDA866HD3jJudmvDTj586ZLZB4+HN5
czqpRKxszhp5fdmQWTmZTe2vZD5d8OWYa484Wy4ibcVSg3u01sidLxPtBHuic0iFb6u1jm/LNp0+
xKz1IfvWcYzJsu1OtYM=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YfIAsJyGbp09vumcNDvZqn38T5Fa47ftpOKAZi1idgKYktQUsuW0jWwd75HvAXmuUMsnPrWM+19Z
4z/dFsgBQA6gjK9CNTOY1ViKcG5TNwitstwV5F2bOApPoW6HFMPI52C+lCJpSFqpbo7JYgLcYkcA
AHrZoqSLfreSrwymnyEwPhkv4CkzMYArC47shKF16DMl6OHk8knYLgF/qQTeCliy6ED4f1GZsmNC
5Y0vn9LiKa6P5rSnEZAC4YJIitvJ5Q0qCQE+Saf/rhnqqTK8EbrAZ0ndA+nCeppKmiL4El+ig+5e
S84PlvE4YJdyzdKbiMPQiAmRnhIg9gBODiJDew==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1065200)
`protect data_block
Xj8sLUNI9GWwitq8r9zhduewLjAuzzXixS56UjXoL8iqWXJp+3A3cpZI9mDrSIGbvs/C72fJQqbX
KtrCUSrF6rGVUkEWuhZJoSMObwkTUxc2TwRe2zupo2KTXfNnOaEHq4X0zeZ9wgLKmJQGgq3QP9DY
IUgeriiNZiVUTktJAbJnHOqn2pxz2GdXSlk/5uL37u8oqXWzy4WyBrfIKyCVAXdtJZ1b6tMtRx52
id2YQzz5pZrjdCLyD9rbRxmvFw2NFaKLu9lZ9cZ4e/Rud0pB0QV9wF7hEuC6oCVOeRTfUKYuQY27
whpQOYilfw5KfYaPTPe2E+uiwYLU+YieTerbiU214u700k3gS3nPza4kPfpMydpAW7aGjVUVurzU
F0G3yugzS7C6f1YyTuJjNQhvUtFUJ3af8VesNAjCwMvjf6ZkBbUQ8Nxw7XaUkQmGOcSGC0B9AEbU
UJFs71KOHNK95IlpF6oat/GYscTbUaGTkflqbmDuVqXCMJb0SvcyrNxPPfAAyr+a1uyq6GPINrv2
HF5Fy3kdFz11Y+ZERYURRHcYrMIY6HfrkWYUdrNNjIqkkHRXYHK9GAiwGRwPjrMReqJiUfTGX16w
8emsP7V4jV81/8gOPV6XBFU98LG1PpBx+iWL3YCaA82ue2QP2OxLb9cgvl2C/A+YcMt2E450+Ejs
EhfgVrz71WYN3jCQ2PqKfBNF2/yvmtvXuw0lpPRx5Zx/6MDLfwsgRB4bkpk2KROspui2NouWt6Bz
OKk7e6rXDME+l4iJUpTOg1H46ZuaSgDdkw7fohsxfpJNdBgXfxQd3OwNVoRW+SiPe6AQgCldSIr0
y22gwOsqnd88WFLX7wBNi3x5GSLh16o0KrvXHKCYYXCsOR1welE+MVWXMAMWJ/AaiYv98BL5xo49
ciPfa/Mj8Fg1pBJd7HmlY6kpLYmv73Yu4dTnjQj2gX5+KRH1fiYbWDXXbq/5gGUMg0z42hpQmBqb
wUVM3rpoNZuBWPgzg7sfzleCnJ5CTS/7wihQUx7bn6jL9hZTB6ki5/6y4qSmvnRZB8SfuvQQJm+e
mmP9ba6YqnVYT2ibKeFssAM/lcDl1b3k/LMuNKErSQYfK9uhYQcAzXOiXVWQXWphS0x2KuusBs7C
VMNC1J7YwEE3Mrp0unc+IPrrH8geV1HMe4Ovt46tR8Z//oT9HZy4R2JALCLshPHo1NedV+5NPs8z
r44FbsX4jJw7Yo6Lje/xp8oSvRgcuVpw+M4cfnYQMjKWkwIeAkSmqrdvwYS2Oatgm5EqkNCk6MFU
ocP3qlMl9dxWSUta9Lgr+MUePGtHTVGiLT365fIs+FkQ9dPiyKAV6pZd99fgDg0J+kJs5iQgy+rm
c6FQ48ow7EKgv1JUweQ7JVuhtBSoyMJ98jDqz2FtYGBYgtBGmw0TmP6HVXrCLBV6gtNxiVQqlkZn
vq+GMpvU9vjqXP+gR3Oakhfsa86rlBEiSC9a3i2HrkzbSbPGtEc7BCLFLW+ZUhIP/XjbtabgQAPO
nFBO18swFd/zin3KEPFVwj4MSt6MOrNhxssd1XKgGecDDxC5zYxK21Iz5fxdYaGiRtAGLTccnCIu
8UdKJCxZSCNuchnXiZYc6TRIsxW3OOryx+MRwMqy4GrqIxfAeIp71YZeiL7lxu2hI1IVKJ2P44Na
ZKvZAErs8A4/ZX3iupitfkhRrD1hA4e67nE0fgNj94YDAd2RiLVwO3rZy0yMbEhkRUVFAM+kQLE6
vPgM/RfS7ixG+hXcAA33pOfz/MUbRJtevvVZR6CgsU2sfA67+CHSAdD0ZhCenXbwRpIbh4BjKqWv
VNl84ZT3rKadmAbw8Q+G344sAvgxs7fEeHj2EauEsRGNbnwJ7P2VrJxD0cYRn8fzxK5mzDQ22WVz
I+E/cze8kl1QXD4ZJ+RP0V/6ZMGLPdnMDNp8AbsuA11l18QEBT+rwmm1EJ7dBQ0tYgutmlVYk04I
9WGYQUbakk8JX+wSk2n0sSIJ9bpPKoCzHib2NBmvIWyWGzqkZ1Zx1KS9stfLDa4+Ufs1ZzYHtiVQ
N9RKmeieCTcdWRfSdKVpXqArJ2eAlfh/FNDkN3f6L0hvR1Bii5PDvl/o8b12nznWXI3t63eWhjNo
5xTNtPP+Ob42zigaO0OtVe+5P4K+lvyi86xJ3hQFSScpzpN5lixyjBPVTFSdU7pejylqzMIsLHA5
pXc3sR9tKBAgN40DXq/4zfuSm8PTtgpA0v0Xr81L/c7vCDn0SLr4QnQz1d/TBLZktBcZsggdm4Oa
cnLVxjDNHFaFVu9jYAGfOqDGQpsucFL89iH8tbq4zS3RqUvvF423dGgE2zZ2olp2abBANcME9XjN
cHHwZbQ05amhl2oBqjzZUL4+FZ9VzO4AccWU/l3/I8K05+NCQbeiaqE/JDXblKqJG9Zl8fvd6JAj
Cnt7aIwwNxeMNOHt8FU8gKbPEYlTQQp+lGNUSVAAerMKNFUPMmHPmOXRbRwzS4YC05rDjdatVQ7M
/qwp2ZMLps9WmlylHHVNfID0cxLMG0a1YAwAJiSLdU6VGSw5izOOBfBAByZM6rKRJHBIuSTpPy2f
PRTlrUzalky8+MtcPc2oSx5y2oHRK2fooffjQI6fHUwukGgCsW9VXOS+u9rbc8IOLK290pcyH/eO
QV5+x15csBrhjtVMRUSlK0jUUuF+3ym5Lf5kw7qqTAE5bFZa2VqL8qNfncB++SN7BSloC9xjkQy6
+Dw3kWQDk0JMps8k6UYOndcIUWEN3lfwy9P965d8oZaKM8e8xcRV9SIuPVMQqfF77srqVy4kq1uC
VVBIowbLQXtltb1cKQU81SmjoWOuTO0nLF7b6JsbIqL4cQJEJbZTW0jsIxnqw7q4vP6vFtHJj4pm
DZyhK2FEZvIW2/0ZunWE2PXJwuT3/JUn7bbZ10SlTW7rjx5yKeExgTdzePVe/jrma8byplUU+I3/
PAkdUT9ghN7gshElK5CEtAMTkyBVRo8EPwmoaKW9yytKlvvCTczn/uTXsXGXnEzIyUojbxUbzVPO
VOt2qH/QxEaHGS+wckWPPNKBQ1i7Oy8Oo7ceEYyMRoTGaB9A6+E2PwhEMveSuhiZhNrscEaTBqyD
eO0/KeMDHzRX872DLFi2QFW0YZ9/aZKPsbocnzzLEn9xoiCJXtIuEOQ+M+O00Vi6F+ixR/A982bz
6P1fVoxhvrncn8s5lza501WYW5d6lfqIWOb155v5I7LXBZxQs/mnHH7+FoVRSUi+tJfBM5uBDA/O
vQ/OU5cwlb4982Orlj+uCvesruoyosuY8dlFH3i4oJk2zMgCkdqyppfMsgMZcIewy9ulxTb8mQSO
WQxFdAZZAkoMb2E3xKHhbu0t9GLJ1XOn9n9mGuOzH/FlQ+ZT7sEXt9NVq7BsxUaCL+wK47tAOnd8
m82KCIIy18Du0vjusmNwc2d8bmzaPRRuTTZQ4Tacq6OjiSfA/LVy8CtjNpRFrviK/1zM4orAmxQ7
ZHeDYEa/mC+Zt8gs2Cn7Yl0cJcmhLuWnrylJm7ZGXWlXeUoch3FezBjOi+v9x7xBSOjvLvmpLHws
doaw2s7WcH5Jj6zsXwYLZJ6H3czVYXp1AGEupF/DShO8xtFCM/d0eFlHDmbsxvwCLXu61eqS8tCV
wh5xgrf21sHWFZVi4P4H3x6yaYGq48Ljjg0MjJn64cWpw9sjKWp0dbZvT9Tv1x80kKFG6VbLiBhz
3WELIkqd7fxn30pN9hhY/Z0K5l/OGiFJaWVpfWy6FwwLrXx3xNkqxD47gbej39hFyR3S7GFNHvkv
yeLdKAreEiy/gGWJOvnwNvkJDzrHx/UGXnS0xfGUHPmRlnzLjt4zkdTRQxr/mWE5VJmmpYVpRttj
MAEZWtj1tdmmIeRmqQlowTSsyep6WpHld73j9gbc+kOEPxVohjbwqQAeHHW/iQKn6DNtpFJ37TZC
CD7IRo7PzccOOe3pHpoYkdviemzYDvizSCWqTRCEzNCHyF8EH2t2IWLIvWYtGlj4/0ToC/s9yjLq
p9NHcKJYkVu0MmdV+cs9RUOZrJfiU+cbpUKzSvKp5BanDqwkf7Qrdl9hobg9wAn99E7e7pCNiTB7
rhthoYbE82QMZ7w/pwEq5FcLYwtvkPluMA06QZRswAa/n0LME7dtJXAnhoJJwJ9hrSJVGakKm3wo
YT0yGXzJl26u90qlN+aGuRTFe+NYbb076N5ZFKV23rxkiY/4oxmaGIH+oWaJw0fbzZ2suhaqrRQw
qd6Z0MDTzaPQYUiaYtkRCrrBnXLL4iA8ior/pMm6gZ/yADq8kw6Wtdnb+0coz0aJ2Tf/4IUOfDCm
AXRvwCIvL/Rm/xp+EuvddhojjiccTl7Q9CrnC83wMlGtaud5hRYVnLuXMFl3IR/Kxl+s67jHms4Q
1tg5cLtY3qRVeqeaeRyGJmVBVy+hZv0RKbp7zaTDws+kFt+5tyWE2cK7RIbmb7OaJZNh7HxazJEm
nhZgsWl+bAe0YFp2JiRXfywniS3ZBjyY1+06E6p4BhTuzOWfuksycP9YNdsznP3r8joUT3wu92js
fhnS5e9yO0dmJR+e1pH6pr3Qr7BR+sskCMFt8JiiCtGpxe+Co8Nc9vUOYkNyoS2LVq3Wu3xpfI7z
HIFojWqABpiaqyWxkGiGCfFsozjTgfnyghTV2SU4AfhMAiDLgbyaLSCyqcboWw5sTO7MBeBFj6An
eW4htaCJpby//TbiwETYiwtsHziogZgJm7H0EwgjMU5u/t5/BSeEhR0bMW3bHLA+8V9y8kIvmTXD
AWhOyRZ8hRpSAi5VX3lYUK6bbCsumjZUFQfq5u3EDcvBP7zY7WMht4qUQTeK1osiIEZv01Lj3iGt
LkHhCqbLBJHz3krBAU7/v80weYazoQkn6iXjExhY6TDmzH+XvP1FLBTfiELKrxD24boNQ2sfD005
9Dk0gjBEt7Cf+mTSx5LuAnnITQhr5W578EZoVnDyBVtMeO24eE1t3U+1jmYUur19Zw5/yOCUdTTA
opUJXXW5ZgVt55P5l9+U+IAtx0lmChPzdPXTkWGPNtRL6fyEEG7tNKURgsVEWf+YM6wXBgRwjqX5
m8NaIfVDfO2+B+tnlwBUmEejHAjfN34YCTX8uZlSyQGavf42VdSXzmeD+Z59D7E6h/Sx9ygMsO7J
sABTmJBsF0BoJDqRU2LOD++FN8Lls6Ulacp/4wriXqE8I+iFBQmw/+D2yQg+McPYEC/l0jnnlpp/
ozZRUu9tHylBQaJVEEDupGr2lavLFXjTE6Q+aVbJoCCLcgrMSkYZFOLxyaB1N/P2ZZ8AThJFhGgX
ok3P0RXZcAjdqjsd8Sb+tekO81HRiW9hU8IVO6RWEcF1Cg+ZVsD9V4UMFw3BPDph/NuwdC8EFbEA
3RqGqpOaFsY+ostyp/rKgb6kQRMcCb/Ei+mFNOe6wAkuifp7ygBgGkJ8yZYKAShPSW7NAdgAZUVo
7YI6joQrPJJIcKSv1pX2IHo5ur4gW3vVYaK5Zc/OF3GvyLHNRl7I6YuvsSmgyHtt6mB7jROEv98W
DOgS+v7QioTRQZYgP/zj1zINyFzGYAoeuvlI+qBveYH5LGFEuNkC7xi/xeajckG7fMw3i633eShR
vRg/f6gRg69h98iQZB4y817MP4R9UivL7W2keCV47uBk4Fh+vcV/0TEAnTiBBYfVp+nOhHGlhUZP
ga5IjEUGqfmH2mYjSETmMcyRjt1gEwcaU5uVTEV3lhkRdPnJcfd7BO5xaKhY4+vPcDLy2Ex36dEQ
c1JBGrRDY2cYtZIFYQlStRU0pb0f7U83m2b/QSLYBOUrzPcyMp7o6mRc3YcvfbcCJUn4pMp7FdEW
rfOFqwG6xygRPB+5VPKOqsT3qYlaCjr39NQrDai6S1QIsHM83l3TsCot6qbDG698TgI5LjHVWK5M
Mebbia2envMgoPFHKEVECbLx3tpgcjiBD2IknGmby97L05fKTRjFjnBGr0d3H8oqGCW0BVvXkXso
pClGlO+HqDCBXK7pFHII0G+4Yyd9D5SQftrDnBv71nVA2GK1fM29tZ/9pnL+YndD3+2sUVrzt8Jt
iysvJ7u2vm50/E5wXyEv4SAAb+jxrjBscfJfQFpGNivH0KIUSB4MEQ/aM+Sa+QtZcOXH0g95uSNU
IEWdKQSZfhsPvW1a9O9yVYSeSrdqJby04vPC1DVfOQdewlcr8esnr+zRIv/+V8FJegBgJjOeBkFc
CNBUmHnLH8yPfUdY/pRXoup/Os/oAduAZUfRr6LPcV6JpSpBQlq1iuO8s3c0mclgE7uJe9rLdptw
+hQTDGqk3/Jo9eMqOfrx/6GTQefwyBH307Axtjr54yQ3UWxHExfTKtCJ2At4Y/W4XSnKe0PSd/hh
nLzKXmn+IyPBjPddZWINotope/IO/beGCcuYwJsxIfg31zuO3ejY3AzCqQntsQU18So81OklA3XB
lf/gSeKa01SCKpATRO63PGFVGERnWrZ+8Xok3TmKDHgCw+GGbyL6y/VIiTNwmen/9YscME118vrc
xO03OEhWNHrQPF5dj5CYtQ4M4sKDTUwiQEhVjKgdasLCd9LFTTsI1BXK3DYxNmelai8dE0+wTTTT
za+hvrrd4wfiZDLk+Uto4v95oXjtZGs8krz5fPoCwvX0cuw0Mzqq1P8/0ouYBB6R7zPciv6qxyPn
YqT4dAbKLxY7YPzx22JDfdwX3lG3DLRvSzyeq+J8cyYl2tBenOpG2E+n1AOOJ6v4Gjd8HvOvoH61
hsFxfkzMsAEocZ7+PzuambH/ha3haWUbilrquX6ES3GU1omSPLbWbtvPcpGLqmR6HCDB3Z1KQ9z+
9GolSDV5AMUTpD+m10N/PO4D8/WySFuMluVNRW0msFIg5gg+c5YBI01zx5ac7vpeYOuyQcbLt383
NDWN1iV+KmJGJyt7GrK79cl3bDi6DGikPE7wOeKGWjnvCV/clDhMRfrwP3SOybz3r1A7jqQc4pcC
X4KvPtwE6Sl55cXUDPfOnevtxcCTCjKTvN8u19aYqiFRfxH0/Z5H48ouzsm45JfMno0XOIZgljX9
HUHh1zIkMknh3zAWuGR2PPA05u+ckIEOuKCxnsfLj29T4qtbCH0jPONRrEVbdnY/ZG4uLT7762mh
AiBP3YVdwr8oX69wZ8vhqMdHV54LV2/nAo2UYmKmmOBUn2S4x1/j6yZS0Ui8n9J6v5tJXM4d6eZs
4RTujnTSTV1v06RgKkdBGaMiCAWOF86WhcMd2ZQsTb82I2WX/4KZ+LBiTMwBpR7VPre42rmpx7R3
4XmgSDswJ/YkvEo6daJqsKZxvW+ETFb79bG2MGUE9bn4WXJBwgKdw84YZBEeE8oEH9e2v2mgNOsa
fT2dktHC0mNbCeFC3echFNn7rJbzLDOVe7O3QQ7XcTChG5IzRthEevYZAkDb4AugNLtkY36Ow+bt
/gUXGTArzkl1uoOGRD6EFZXDoHwfNKvqTXCgGilB4MKj4J4GVGgSitSeOphZUFFRO/MBfAlma26g
TwgqeZV68P77kTXsgran7S5+e1cuFgKiUIPK5RapH4CNWIz2pHsdyvlmILx/j0aLG/aR1AQY+yWh
5Vg4FqE6O9FArCvhmovx746OEuDKemkPLdo2+yK6MOicYncl5gEdj51oR3yptGfXui7mUbradzR+
sPlzsHkiXRffDlhK8DFki32VMzzwnMNtX9ZQFV0dKbOtlhsq4x0ktu+6z8fAdqQa0KWuCPd6UM1B
8aNSqTEfVgceMXj1DPaMFBnMmu5i7fCL5Yj0XsF78qIcWmn/b810PLBPGtklwDoMrf1nhSf+xUfh
6i5viET7x/115XHKYJr3RN6agLPDMFOjIvZXFiOZLt8iblIq/EQaXT7V+ZF1mDgfnRzZ3VYB297Y
XRCgRUZKZ7MtR2zh+/re8Ielf1r5VYtaenLrK3QaikC4MWA1TpqVPtUObDA3rSiimzFw7qTUfN+l
Ex+qxNea8XID8u4NE6tB1QgwPl+j9ppjPCLcu5Jw2eWvUpKsz/o2wdHl6tEruHwn3aEjAgID+SC4
SiaM4rTbmKhO7LCgojZo0TI/8GTxHPCXTIqi1TwrWl/MrCtifJKkIZNwwUzF52YOguPu9O9+0UFh
bvxYU3tDZQiw+oj1p05ZzQspMlfZVXfo+WoMuNaZoquDH4JgUooKraTjnUiZgPFa5J6EuoGpPMZ1
lVioTJYW2YWEcGUl8CSBZmkM24ixtJyuStQVra0gjfRIf6x/Q7r24NqpLnUY/f3H5Dmud6PFcx90
sTFbw2kY8vB6j8yKF6eIY/AQojhrQecnBkVEOkSl7uIDuDqGVVcw/2o2ykUsFZlANGsgnz1dyKnn
updbzHKEGjSKYuUDIF/OdRQ/c7ZM/dYNMdIooS8Fp+IRbDeZVRyy7xL+pYNG1Pzpewlt4KD75pK7
TGR7a4l/gtlJkZQQctrc17vjj1qXOMqwUDCd7lhsBm1bORSWgI56iEuSukWrLAIRZWaDkSGx1Pty
bUIOD0Hf64xq8r6t++7lxSEv4W9RdgoAbFG5MpIfVOPyGY+Xg8p+qfY97LdxE5Yqyaj/12PdeJ6N
brviur380wyvmhj4iveJ83trnB36lqN6YoHHcijPG3MXxYikeE4fx3qt4Jdwykfc/z3CkXgAuI8z
gvMt0LDve+V2K61I4xuotlb/ko0U4NrTka/RWwMJyTpgCyO55RUnvWRC3hb7n8t5pVL7UliCVBBm
aDjwknHQepKbs229u0QqmsUvtCI0NmSud06i8hNn2fZPjHA2MvH7kVEG0fPJW5kT/QsfFQxMtx6n
8vGS2waX3VChSPLcxWiaR9jc3YPae/3rB5MlGP1gagz3XpBiUYw+WDcVC8GCAaEoK6m4iYY1KKbv
dLN7TAS+4fORX7Rh8RJU0mo0SJdslPMcRLFgLAfoI0Al8uv/DGmv5cJT5eyfxp/U0jSHuokIpNZt
gCqzgKSYqV5oHABHEEsWbbOO0RLJgSBb1RviydphHxcSlVynoemQLwfr+Ns3NukMdISrV7fodgDU
Q1Pfou9vTLPsDtB4rDpGy0G0J1xiCKgIKLyYaupGQQp6lb4tZOhiwkJU56q6Iw5o5tGD8Cg81L5/
ppyQmqEaMsoa6hfo7htTkThmFczp4ZXGLlGFVj9ZOhP6canXWtNm9RJwoYJIBvBw9BymD1U6GcEa
KGPyp0TUPBMgzCxC7QHy12yYXIT6pJQmYsWRETL9vKkxgeqfJEE+ZXH9fhHxNs7vYyVfm+CQfLfV
KpE0kpFh3ZhmcOQRQnuGmqacaeR8iE0jePjcc7O+vA1CwtL57w2fsR98xWHHygDUDMjWJs3o6rfM
Rnvk7xJNtZRrZm5Q9hVkbVIBhCaqt+yzY/Qv5jf8n0gOdbWI02XCWyl3ComEfvrSsuu89sZr+oEu
xuRBNc1pWESxMT6Zk/1Z9RdFDhnSDtH3eNpdrk4Gi3klMgmfrf3VMjoUNRVwpx6CukvwRdSQsOVD
Am1WvOxth/zzF9EBxr7SKWaiPgEvwQzpLP4iQM1fB1LU9DgzjhXG9ZmGoHFGvbl3AM9MwdvL1QSu
NeNCIgu9CBE7jeCUVKMos6+5T8Vxygx+Hqne165VwteLxTe3NempLmjnj5Bn5kLGhX0TznmMbx9G
npoEK2vkoICCmN1T6NMKt9uuh0WcGokKmZwmggG/DEK2ZBcXDg5eHxWpBna1ikLkm1ZJ7YHcGddD
ljkbLsA0ki0lmbeUU2hunDNK6qOd1Bg+7ubElJIrJaoDHigJySVNhflaAzfBAIty4BOEIv3jSfjF
de/RntL4uf9Xk268MVAbgoKNjZWbE9cVoPUvHw+CrLs3OsFoNiRpi9KowwtCT2CEZhYaMGRvhhtT
ZazV8doxYLA7Uazo6C71QvNyUKxcmzxnuTeXu3jjucCNVIB9blLTaSQwzj+56EK20EDB4G+8iuwb
qbZ6Zo3KJI4DNTeffgD7gPLCuqR81AX3regUXqCWP9SWUxSaLZfXvmdjFLkZ14ZJt6lVHqFVLncS
+kfRW9Lp57r67V+LMWhysLdzG8kjlgt5u5oD1UESVd8LFHk1gMG7J4ke8CzUu7J4v/9XfuuA99wv
fLcA/omJ8dg4Ie9T/ZYBALGHkeP1wIWUzv4mfw2mjgwNm8gZBzJfh8mpAXSyHsasjUHVl+NMcy1l
EOSIQ0ndxvTJNlU75e7m49PasDCLxdfhC9+Wn5smKTM9RGtyhyGWFB8+SSnq3UjU/TCMvsPPwsrn
UgEMFxWB+GJE0x0dE5S83gR8ijMujQOaWY1lLGGQHgEIcuxzdkljnxZcIlGuo3/QMtIej5nolmwP
/lmz2O2+hmX6MBuJzkHkKfVbwT+z1Fhi4VFvfnkwAaxLnQVpvTaJzSlf+DKv1QkITHn1z22GHlTn
i2RIR29RXY/eS4p2+nur5vfN6iKYewL2VX+SqnzIh/0S+pRU0ExxH7lHiUjYpNUkHc4eteF1gBYA
J1+ONm03oXoqeWRjsqNg00TEO2YQFvV7GejWXeqw5FCLFXkII5mcY9r98vhR83+KD/lqFYDJ2sq4
9ugf+D7mLw5AJf56cYpLXpd78S/O/6p7lvNpC2JRGUf80cF4X60PUInaegXtfAQQjG9yT7arIgXD
rEmO5udPzHgn8QoDSCx0MprSFJA8+t9u3AJ9Luo+N/JDCKwnzhfO77Qiv1UG6AF31JjacF1RXv1F
Ed8pdMGnxSkoCh4b6Sm1VIDJ05wBwNvJhuxj6wLK1TgNEciSJHSeWrv5Sfx28I3/fLUAdjaUFDow
bq51rsM+Gozf5YNuM6qRA7O6kPMnPd/Go8hqyuVQh/3hWnUOKeIc89JPDdMki34wRtpVFWC4cgJt
hYQr7IGuLgMQPnP5SDghZ8hNJi3TZ+2OzLphvyp4DklVLDN/Vhuhbqwu5WJNeVdFjEt0JZAFVeso
kBjr1vRjdAb2CvCNVmtSglUYGtWkj3IZAxqwiLmHATHaoFSlC4Ljjd+R/cUac1SkaqDehehRAZfz
DnWWjG/e8kFzf+SX3Ui419H6kfn3xa9hBpogTx5B5BmKmdGeuKpEnc8WQBIpzZjvcvW21oQ0PQPk
blvSmMrYyRT6Wpst6gdh0g6bVuaFLRRemoSiwOAvIYmXON4b/uEPMTvZ+RfA7BoooAq6Fm7zVJtO
EBhes0DygPvampCHh45J0YRIAg9PbcIPJzTUm1aZotVLwN2frWJeczn6VaKPbTTHyYkjSSrebhgM
ormvOaASFRQ7BI7G/k8bSWm3a+e+K6BQgDUXKpmo4qAS44i9REq2AZ6K5cdEkj+JtHjkFYFxjamU
TN1GFKlhwUQvfNOHLO7STemv7P+Q6BaNw6CwuJpYi+GlIE9Z+AP8U6hL1zXLLIyUAHh719gwMyvn
x1DU/LL/OocJSFila0CdhLYecgbYkN24kVTUOSQop9ox7JC7HuOr47lUpbo8USHryzfVJzeoexHS
INkz9Wvla1pal6aK7zn1GtizGAIm35E7A25w9nzwtzg3vV/Rlu6JtERbir5SEJbpW90BCmoMe1IO
4NdalaH8qYfvGX14gUWVYjyRks7IrniJfoO8vK988vERi9JbCHkoMyWuUPfo6Cv6ojVSGF7AbtgV
+irEWGoxIXKZSoBD2RKlNWNkg0xNA+48jGoJg2lnwz9CI6vipHSTY5vgOMiS92htp21K4TuyAt4I
wAbzs/zV2oY+vJD8wM0ygkh+563al7lN+SuDwJrtiwskq+zPs6Q7D2LpGx4A27rJ0rMCRN4tDETG
9zSIY1cIWcEoa/SYdI+CKjgaxqztBqwK3Mkc1eF8PNQYBSIafuvbvkCxisdTWBj1yI4wRIBhSwhV
0aAYudVsswSZMW/Dc2G9TZsTqmmiUHAJ2ijK5Asza9y+SIjH2G2e46nY86GPvpOyMFkPkRI+y273
ocBjgZhQ3xDPGgekdrhQ/RJcaFQIqK/q5vg2oEyxlF1Xm/PNepTrQYL+ViBuH6J8gDTAOjSszraE
BuxafwVTR1fe2nwM7+acem9JDq35q30epsEglGy0xll24+HaZ+FfEVfGfM4a5WpAAnO9xuEL0hW+
amp3rwMVUGDC7bbneDEKv2N+Ymw40HKW5CoD9nwMsiEyo/c98vKOIAvX50bbcO+mAlSyOPsmRtnH
2E3OVv3b4iBJ56b186g1rYrRt0MZIyLdQKt1x7gSao+dDxmchUYtJfjqeNVa7FBXcCdmj8j/Bx3o
WXAF1u6uXylID/dRras4OnvAD9tZ/jC4rS4iVi37mvwYhZM7pH9/DBvw334JDe12D5mAG0x5rnnw
hxmfgtgKPyzjvcymVuJqcwG+BMiraLwrWJfFnDRMBuDwbV/4LExz1BJex3yG7vf3y4DfYVAq35Z6
XQIwbJeUlNNj9djsJu0uu4p1Zd9q+YSI3ASPcqoFb/wQOl4Ixy3diNMj6qe8N4A2bczO573l89La
/To+fmtkTkx5YFhL7gJkPfoS8keKXGq/JPYJRaNUmKYfHkS7Cs5lDVComs5xhKIJWrZLW1Q62sMt
PM2R7e9p82pMIwKjNYcqyLYdfsw4mzmh/xVad6cpNLS2bTkTpwc+Xjf19IifAvLgqWW0nQGIt48M
Sxzzd3EEezQMISwkXfP5Kx+L/ELcKc16DwzEXGTxyFvzee3jlIlRIB/hUrfpKZKCXrl8lkKCW3OX
o1dXRX5vNCtiDQjTXoqkv3lFbVskO3lIg4wHdX2YKucSGVWNSg7ZnqVFILeW4MloCE0EUMonP98f
mVuRyam9+IrPWEZ0uIm5VoYdnXzECSPFqA/xWmCvSnBfaNxgKzmZvPQ4GkLSFLk9RQo1S6qss5xV
TZkZvTTh2Mi3nFzawlyP5XzmtobEabde+X41zNgbpC3RbPilWHhKT6aQYi7FQyt8hTMwlDhMrS7U
ApNvmtbTYHIVZvn9fbN/vAfnHB4hpRytOLSx2M+38A1ksOxARbINjrQYBCCaV4El7govHVpOQYDZ
F4Nl6vJgUn4KxxMDVwSVSQFIaX3QbZKb9rtt2akr5+oiVPYIqsyL4lTUePa6rBZRNrjE3mkej6cD
hPc1QWJFIbQ7rvdj75InaFuEjf8YK+HZAoAgROHLXFkYCpq2ythJEEGUHIRQ6StNlNAly0nV1j0y
+R65VZdfYPA9cBPiC4CSiIoc2AqUzPYlCKx+6iHw8/HPwtmJiysJ7EEccQCfu26zR38pKcLN6ZOO
YZOOgGLd5tiJF/uMQb68V7qTQFlw9KOE6zWAZy7YZPsUrrDy8O3Ew01ENzQyT0X+b11YBHZuH1WT
McctfIkjdBT37Lh56PlXFV4VVF1moy9+9cd9m3MYlBYqSsynMSrd3Hio/P9goDTtRzsS4w+Tz8e2
W6Wu/HFPjpsac8aePpM1PqM7RMYur4kyHwOQ7rBH45wdp+IdFGWz7WVQh1Hxz0EISJR1GrP3QZ0e
WxSu72rMHawMM1XsbPwi/AAZMrEn7fNxbuFhd0hiiakPoYGD15Fn6PVQmCSbsZnIdFKXKHXO5Dkd
1uT5kPs2vpalI0QCbzCafFpN6y3GvkZuM0baNwmfK7aGPzuVn3Y4dQyc0zB/smmw8vTeOB4R2++7
gtLK8EAqslM+LDRArO5NyDhYimSSiyMCnu69p+6ej3w3VOCV0mWDLoBN3Ix+ry/5ozrcF1+5erI6
uril1THWp2EA36N5R4aoFQkOU1KUilZJnjIjBto3WtBb+ieu08APcYESHUpIaP+4R+5uhxVza8v9
wnMUh7Fsb6UgGJK+g69Uw/QwQ6aWATla1AqWpIFI9IAo6UQ/Ha0Ns5dp+KO7LgCUfys7EM6elwid
Lnw5RAnwYdXKGM9lE/MSKGv/O6s5kfR53kA12fDXqnLluGW2fvD/4aHM+Y/TArL/PA3Fb8+TaaLt
i4PEdnIQ8Mu+1OYrEDtVhjarRm2JGQJsjcmz+FwAV91bQog+SijrghKMHej7K4IElqqubjS29Iks
QdXnyfwFyHvGGNoMacqQLRz1WfANh5bkxdVJU8RGqW7dZTMkiiXKSJr27GlNdcj27UQOND5VbqkY
lxN6JeOpEFvB9JTyboBvVtfXiZTGES/wdHoS7H58qUqKGrJHzWH0bd9y8LWKuwLnieP8JgfXBa6u
zMw5+pmkxEUEeRZCz4KaE2HYbYnxmWGZphXK5voJk5Qmfud8DdGIdbN8M6TqRVToqgkggAiSEcig
oylW3x9yQyUj50roI4f8joOaWsZ/g4cRwSA0uUhN+TPDoxLUrzVXAk96LPEjzjtbzFaiCRk3Vc0I
e8SeDXIEeGp/0kjLV6eDn2haKMGSuQhdJgoc1pKKah6GwBqlPkQ/c49FOM2eEMSZPnyt4v+Iufon
qdsfcPnXo4drNfBArfyqzl0KgeMN1ITjqstLtBtvoQTuGj0ewk9DZmJWEc3q24ssULpXy9k4oqvT
aEMX8HVX/2mjl4FfYhNZ3vkcdw4/p5Y8LW7yEM08U3i8OM9IDWMJi5rG0n3IWbch5c3MSQdy9dzW
HvpbQH8ZH09s9+q8kY7r/juvyGLUB68kFODUUQlKfxVKZZFbBCYmw/55KWOZYa585X6zugVauAlx
KEV4ETUArgPL5AdHk0zWBLvtrKyDYd7RpUXUsK8mIb0LUhKo6rN2OKGuPZ9BcQJQm7pX+oAaXlsq
/LUSIApkeIfcf5BSVdIgOovw1AFgxanK/c4B5EMaQI+nmlQB2lkofTc7hLbB4Gb3m21GcgsRogn2
PMoCIwihqBhw2w+ZwA6dNb3CrL3SHaFZriSJnvew1qPQR7FC6Z1tK7emymeUwyX4DtP8HepkQ3Pg
CZyIxDuS6B3TuH1rNT3+oQzaGyPh5/ZcpbskjqCR5v+R+CWvNi3s7NpYSUkkIEJ/2ImM6cwogRrz
BoVdS5RHmMn7GJzo39RLSW+iSNLESzExyOmBG0fPVZcSXmNkvXa83EGC1WPMiSk2xfXeml6lLvvU
/HGjhQXqBc7a78f8QXKbMxviEI/33WnIjoKmdmsLQ9UAtyKM412IY2c+MW1oM4iL7BW1Jp+M3Oke
xTv/X++y9kU1VJjU/9B8q/2aY0sJeQashp1fo9bF1A5rsHxC8DKT05QcmYsgPEX4vM8RixIdaBNb
yaTjgrlgz12SMRkQYKOSiKTKNorWudnRVCOVSSspnQDBpA4o1BJBGE+j5t3XFCYa88lNUtg4lgaZ
kJPDh4s+7a206e1j07xZG3wNu0zsd8oPm2Sd3flfS8ZRWSN7oP09+iyIkqq+8a/PdB47rXq/mmw+
i822YHtjcaatslpvWEaTxtAocB1q1PKGH/V/jxx3V/FLYTiRVQuVp56t96q1XrAGhpD9RVgzi/c5
9tbdUAtVBI2YgsxG4PwlSwR2wuoSoOxFBKQb3j7IFIqQGBifgCIEeBXG/19gvggAj6VVnWfCVCMa
8nsftfoCwwkWH4Q+mM0+HS0Z7jy5GTGDTku9+vFkubCbKj54mCJMgjtULESaoKLmFfz8IB7R+qox
r4SDlkfIShhpTI7cTC/k5FWf3nGlZ0zfFgDwmbsegPoJnh2gChptAlFPSCiLIMZLtTDlbQAgYYF8
33lqddIJHa9SBHN67iampmQs3hNYASZiE8w552EfSa2DzuiDbeo+TdE7l/9Fx2X8DKacWs8Ax9Zx
x/c5vuIcS+g8KS7u552mLY81HfkpWCDvqs9f3d2jKiKt0lzmNUJYvobsgP+AZP1CNgTq1XN1o/oX
mde1trSsjgbOqRqW5srAVXng3EXMJtnEvzZNAzDACD0GCUvGZd9mWTioETJGIjOZC5R/WoSL4YYT
VTmSxc553X7na7iQAZ7H3WmINYB2w2JoR84ookRkr0BYFJKa97ZdWEZ3dnVLfehwGcd8BUf+o7qn
V8svwm4WL2BLwVmjSjdVncq2DH3wlGa9aCBpisZO8SUYJIGnoZtiYHKFru2fRACeMqX3SegiYf7b
T7H6adlDb/VYqmyVi1FoT4t1TPA5KwdjW4eKbTcTqPn+gQcYSJL++f3Z9RZOjdH4GkXg7+VauNx3
XpjlXVRzqjWJslhCi7GpXwU/IqZwljxir01H30oImNAuMCpqgaLDRMrtIxVa3hiqQ9d642mmSv62
tlL6Kok2Wk+Q5VolqL/QRTuT+fsC/BPLIHSOfTBj9s6VCb7ESUOmExuc0vDiVfeFD5JuTS8Fk9SQ
pD9cNHeJ+UTzQJnJTLUgoCHpp/rqxFlHnB0hSjSTDngMOg7HhWL1WB7usGvdwYjX1O8tgXVeDwAc
Cr2+YcYldAf/4Ms7qZq6bGhOGIL6VNB19w+SAFavD43zVIRKxLGCkbGIBhL8Z57uqKKWAaiWvNoN
EGJj3dle44IA97nJgcksyVLZwC9JqKgfkwZZQwV3LHwo7HimS1TYIaHvyCz9/D9AFBtbrecHa9tg
XavnwBsz94oNfAGC57SVxA/qad7esrn7KIvcMIxWJuScCloIcSvFw6wVEcbkyhhN72HMnDzYVkQO
pRnz8vj/kFn7mNNlMlQI1Q/IUwYWqvTEmQCS+phArMqup0CmAtuHiVrUj4iF7nqxBk2KWkwngb3Z
SrRQgJZrDlBq2rFhrDNiX2DtwmiZjjFp/EGS/fl5iCBeXe9LOJD7auclI2O9AvSdir0CekSOoBoE
FiHOiJua1K9D/Lm819zASH2tG2dwiFJCEF4dNLZsQsFCwZE/zCJjRw0IZqB/l3LlbGFM/Fj3dLSP
L+vkrLIm/zqMx26oSem3BAXRaCgljhq2NELNuioDqCTyKja7y0nam8qKdqw65H00FK+tK71yp5BG
nzV3TEyg1egCXGLPRpeCKbJxxC+sIGmwsdtHdkWXdKKYyvJ0Y9YNo/EBEUHCBqkKjFjN7KmOjKzS
Z+OyBboy29Nz3bGukTLQ7ks1iqbP6C187MDnl+n7MbN2NTlhiUSU6YK6Ehkp6qQHoBN5YUGMPP+t
GH3tNVzQETHecFdzO4Sdw1SlC4CeUZ37Vx77HK4pDwKI9C3m0DiwD284Ax6nitx+HP/olYF0Mqyn
ysROgJfS8UyBTQdyz+F0VmFWGJH8tBOkXPX1JVEL3+25IhwOjhsOUDFDWdNHM+2J6HFXgb7mmJ2v
FKYyAbysIVSMDTfbljHnCjP6HjSDT5gd3l6hRFWYXbn5rJvKiWkOu4bbQ8FyOrS0SZLTgNFBhSKr
rD7K4DyrS+eBZG2WE1nbidVMvJaXCofqdOd8d/ykTrivDT6eNadqxWnO9K3Vuju65VpqUO3EZZP2
80ufW8HxZNZWWi4sxt54ZcWzAmeaOvkLWXE2psRkdrbSxVc1t4qUeeTwOJtrj/9ZbHGl39GqSPpS
HVmCfIWdGALxJBsqBsozRaUCAIunlpoN40ZcPGRd1DTgHJdjGUH6z/uexVg9oMttml5V33yhhkF9
4HsogU1Aza/8Qgs1J6NxcTZroG+XOQjZou3+TvV60iu3UKHE6SEAFHrXUl9uwjBtvkZ7pGJd6er+
ckE199hSQ7JhNJYugHPdpUTnGXJY9kfuIzaGQQm/HPfkJUL/lF6P8a7AuM7+DPWpM3XZxrRT5ptY
gT+EW9wfUerd/kZpOi50uRS6PDyGNVPE0laXfzWQuj4QLrVpqPCv1sNOkpeJwIDy0KrybVE+47V0
a96vPiSm4lpg7zfnc14Tp1FPKXF7DMUxfTSFetQVDFhHxfQge2t+YdXqYVYSydauqAShrXlTz6rA
fienfVoMr+et7OTgKKnBbAYjVekT0WKr5AJ8t3EnAwovt8vmnIXTlEChD11omga0RSkJT9yQON/a
EkPny3QrgxcKjYtwal3Ek+Q+3edU8ThXA9IRY+lAsig+LLtkmoF0zhAM6DYxL6mqmf2U0SN8qdpW
DQJCLPJIEYuqy8juYRxOxfzRMGeElpPlXprzYA8mDpGEODJRk94mbNrdLj7l4uCqZs0wXoe4YF5H
53XFmkimEkFboOQrnMHIs/+aROJS3ffnmgOsU0AN4kSy5vtY02HZ4Akj3gS/8bIgbVnGYimf1BIo
+nUZhF5TgaPLnkm316kAOSBCczMZO1usDG8MyWDmDe1sGT71JEtKWKK9bf2Ev5P6QcQ/8Weg6128
U8tjBBk7pGo2KYYMuzvWGYzuSdZHGkBLwnP5pL6gmnhYhPPgCzcrKD85S0pUyvhwKwExtOoBRgEH
eMFFLxVWpU5EPV4lT+wTjQQYqHuFi/c7DYV+CiGPC/4ircmah3XqLM5ZiCxAyvgnqb6TfvLJAdYI
Zc+RNDFEVac+EIN4VwDaNqPWHRHzN5KZcR72MHPWCkf509WYHQQcELmLLYiY3r7sN1jf3p2tj8QO
9br5FTVvqELyogpUxzEDNCEZCXfe1NTYUsMaY5k29v5/7Bv6/92b//gXIxNvwJ9C5rMe2Rj7yt+J
3h3xEBQbveuO9NxrytnnhwtzMyNfQCPWA2Ms+1Nop0U7lJgwnXZcPRNKyp8Gdehcflw9+Wbwj6jv
j/vparNTwpNS1sHNWpT9rVJOugM4GeGV5q8+knmqiTExk2Pcc+K7OS1VAHhL3Arn45nS7nl6ytGp
svyaWeZPAs2Fv0xc7CyDWURbif9TRL8u3KiHYgrqfjrbv4/qboNDAd+UX4i3ZchUffb8ZkJv2ejQ
1HZsb15PmQCUimVBtY9aspqC4fYrAFnUYEbd2x95RtxLGP6WC0oCHgJe2b1HpTiB0lNkifJIbOjm
ZNTj8clHh6FQyNFHTO+TPfkr1cyqectFiUuvj4jPf5upwkrEoDbx1xcbmxexyUurlO1yDRBzgcbk
XWUW2aT0IbN9etiwop7DbDZ1LwbDnL+iaOdgDKNxdZSVuXMYdIUPXsCePLgv3Fyz+mU+shieJ9M1
CJPGzgsmMVu/A5AqCdnRpSJRscaVm0XDYHYaRwTCZljJMCb+cud1QBuKhPX7Q9jtYg/UYxdDED/C
qDkVYeFkuVWfLctEEfLH0Z6v+tOm5qdOp4xOvCxuABnapYfIk3tak7oYAgVbZT1F3jMF8rAPayY5
k8iuS94EN0nNBxpleEhpVef0+Fj9FK6Nj4u9vE3gHEi/ZjiPV3mNZ8b5U/3K0u3fNECqWf1Ov6Kv
QKbtwa8CtDVXyWAkZR2X1iJDzadzCzE9IEQ4Id3wJ+m/50Uye2++Lx4OafRwXtyeTmiGgMOzmy4s
IUJCOYbJi+km+QGkSH5P5QffXLPd2twuJX0UpxSHiYlVWzAt5WaZqwIFo4cNql+Mc8hvucO5mMAT
JtZ+YbeC345BanPabS7MnWAQ6vYryEqOrhRKHIt8+Gehpa+qQuvTdsZapCSAl3Yb31GG/jUFSjuR
r6bgr5CyZPR1/1pK23Zp5LjOMsiOKj/azYLwMeVj0fMOOiJMtZxDHFxfq0YPoeW8F98SYz47mIMc
6w2COkkvz5QxY5OV6h4n4ZnXM5+WA3nsaJjZedX612Xa/IBSo8RX5Zb9+ucPjkAB98C9aZFEpt48
iVhH8VEZYaL2t1Yoipw0tie7xGBvsaF0Li+hdIlG4CxRZEXPzs5yAhrVpHrgXFdFHwAoGIHMZZNY
+dzq44ZZOQzc5FYwynij8sFbOcFSsO4qadenZuSYu51AAkHETOHtGQN99CR881iPRilWzh4oNYdh
kDpfTd+zm75Iw2082zWPXdBWz8HDpO1Bds/2UxGm536Ff0BKICTOqm8SjDVMQGlF28HLc7LHxFAc
nF7tP637ulr9HpeCuXQZjFn4F7cq4XYVEOrfQ4svAX3h0uKrYwIMLCrohmsMd0xRSKjZORUqb7sJ
q00lvtaKplwILPUinluLvwgU1HS7B9zk18Hp8f5QDYDlgbYrfFXGzmFPURq7FoFZhs1USrirCYuI
srxLaLEjbFhzUnGkbEeEqfdeJ/YcSDv9If/YOZadS+yq8OugkijSRvFsVCNCFdDK0G3kGZ0i+FZE
lhAOclIqT1e1yVRWVZIh/+jLRyHhJ1Kfn/lTd7YWUwSMPjtOlEksBiy11Q1zn0bqoopWl4CjFvxO
RThDOQ8y1yvePCdMZVi/ZeLs61BVOKmEPiPrdSZpQQtOHg3kwfMJ2s58NN5SdK1BdUlfnxP7akQi
QRFqQQAmdAhKtyBiM0KYuAhNI+3VNP3swvt5zViKmjGRFg4uBCSA3iLYSG78y+g4F7qui81XYpRM
GQA92ipSR7MmuavPKusX2DfGmU8kWf4KgFyj6xQ0VpJAZH4+8XLQZP3bOjh5sbSKslXZybVu2jwC
zfCbwHyQYjDy8yb/o8dUdU2wd4JjG0dX/a56+iDMRt32+CG+lmHo1WtHe763KBHjEfFXGWiYbhrK
EdEsQkYMwy5nImUJWKBSFD7kpgHe+Cq4gPS8yF590XiWVXi1nWczTXL/e5YcnOE6UZMJrbrOe6gt
CLbWKvKs0F0w8Y1ZPIxNLih4Dw0FDH97/wNR8XQG3FZM69o8+P3pPTuNAENYxVjxQrJAAs2Dq4J4
e8pmzRfap+SZxJel+K9ZcK73g6Sv5JGZDnmaXQSOBXXxMrJA6lWYAkXvwNQ3w1mu/4BLON7+UZ/A
AkaMwjBuSHofUSx2on8hEhYk/f+AmnGMcjsht3e9pr3hSWGJMzDxjkhEut7613pd//+NacW0JSx+
vA4IfAAbwHex2FF6m8YKDUWLO7/mTYiniTeEr6EgaIRycSXejJSF6KwrJ8EbLfQWK3tIkNG6mwcI
OKkzBK+z5agx18t9PN/M5CqJYLxyCKk8X6FrMOiVkM3wLkCvtpSMzC4Y+tW+pesNgakqC/MKu3rq
IgZWLO+wk0Ezrjg46HdMgHbzXIO1ZcQ1mAUEZStrfgyK4Me+l1JTesbN1uerZhrcy8LGkE3NYWtb
wPpBkI/bWDhnkfsIcTJsED8we4asBV2JfB3ychky8udAOSQbginQve+WJEujiSjTPsABfDBL49wq
sYn+qxdLnYQtnq+d5FnKLGzA8I09uiLfyVQ0/lm4fn0qgJLbJF1cvrG8KIEfGGMIQX/lwQHa1yZa
XNI9BN/pxwMGLJWjmol99KHDV+gPXE+88IAQxKzX+pod3hzLvKT8eVBBV7kfMJno/UyyTpeSuhWM
brA8YLYDS6vpNUPyAghB6aXCv222wWqZ5N4mYCE9kKUB0Omt4PSKXXwTYImU+FGbdrt7H7xDK9MQ
fyusqaLTN5NSi6w35jyOhcSQp37sqEnXd9dLmwn7w/SRtDMl49mRwYkBtU2vO3RFyxy1emJ7iLln
XKJw/dC+Us8dCYIfcnd4Xi1xFJZ4lM7AVzYh0tXEqqRDrWe0Ib+gx9CIUw2rB76vy7Bk+lOTwI8r
Bj2DWkboWidWWsVDoNdBCp5H3BbxSeRKcfAD9dZmW/59qAi37Adpl8YJ2DIOWNodNlKHOHTlwUWc
Tzjj8KPy/8ch59wRRfomNEK8CYMBgo0F2SRlYcnW+Xlgoca69xW7x+WEu/3n+iT9MpGUwgSNEcIZ
nCdVBZwP5R63azf3/GWtiG1gUz2jJ6nnFkyGUGYrL0n39mhYFd6/qrWkdf84FCa4bXlGz4RNL+F1
FmKQAAt/XcZm0eOENjIUWBmNEDkq4A7OgfOaZO64ARLBCiVi6wppu1vgd8j7JpdaCZiKfJxskHIl
kQHl2tGHwmu97Q3DkbnvQH06QycB+kNht0JNnMoSdgsKMAuQ5zxuuf86E0xTQrrflB0uMAwy6/t6
O2w0BQRtYRvcEMj/J9bU/8U1YRPBXo+sBetTHrD7gGIR4gaHQ6xQuYRXcx2Xk7mFSIMOhlQAMOC7
NJLmIZ+gT11Wzs3CRfqyvZIWiFOpUdCvzN5cCA3J1e5dEXIiURmdwbVO+gHl6QQ2sZi698USThAk
iC640gAhw4tc0LZMUlY8ZV3kw+CDtACxWWOKnFbwVVCzmrADvgn6uXljBsiPxd8L2Ijk94j1JD8b
rggu82HUOAgvdoXQ7BkiktBl2XF/bT/ZEAX+V5w0FS0hJBORXd+K2dl7Jf5a/ISn0qgNLQlWx4Oi
FRhQ+oZD0q6j51c26Tcdtjzngaav2zUYZe32BiWIgFTBY2+UNyrW7nHUsnYSw1YDHjIi9u6NJ97u
jpbk30Fe0MIaWBKZDv+lqRT/WY8n9iAUnH8sD9pfmTw+ixUV0yWppOz12Vc2de/Flow6i/eZemmd
hiW+lBGyGbSZeqqVEWRPn8u8pXVVhsDcTp1t+zY5jWmEzacMEpZlFe6kz2LWfV8FnLjKkjrHJPzy
u/tIQGHebQERlbQX8TJLVziF0rjSK8i+e5QwwvLCNt0ryIClSnnQGNWv+IKcnxbIrTzbM4uX/GnX
5qmLOPY0+InaouI5IA51Pqva8S2GzU2LozmJ0x0UGRfu63SBlZv03F3BoBqh63Ly40jWAPIhEpMX
vGTJ43IL362M0l4+bdL7YPnQMTktykzL+/wdAR+Yrtlyp2XzvRHgZuZv0jFme4rY9SMoT+koYAoK
0VJphtnY2RzO4yD/mJuIzQHnAqsn0zoJ/1MgTlpsakfBdwbcRD/p6vs1Jc0dmfcKx023sMfkWLAb
A4DU67WeQd2+FAzJyuImycxuxr5cXGAr1ngK00PdSlxWNrERl+ikN3FANwiUIIZtbhk1QdhLZYog
6ebeR2zYHyU8JXWySF2+4YAXf9nUO0pxW//TUCh4OghUSOwdGHwws2weCcy9vmpLsbLcwuz70gvV
ayFmAtbhAVpDFwaiZkQc/oi/Jmb46pgbSRLybQl8zDIrgak98nAO1RJG5aZ6LolCn5RBqLx8gv5g
fMc6EcxmLkknnCNwG5k4S1PAq43qjcxIJ5/RTWa6KcoQnm36Xo1FsTSxzS35f4ulzAPXi1Ona+Uq
Z7bME7oXti3w/8HDroSWGyuSTqZqHINvLNOxc7w4m/DF5rVNxXrzRKgi/DtU/V62uRi8IDJQUImQ
kKu/6PEw3rRTuNKpW0fPupuY+Js1lMyIYdRyxJcm5V0xJeV5Ep+qdHnvQQC8FoMtoPiwlJDD2M0Q
ujkXTysq+0vGY2p0+pm0CY0HVFiwagb43mDtUgoWFBanFnJjcK9Jqnx8Kzz6KnLwaPbRl04mVbV/
TRPDSzO4I3k4MseicJ/4sQHTTjdKcRHIJL4VZRHPiiPZ5NyWRi/U1tL/1m8qQ3vkBW8A59m5L54X
4z0XIZOHNSZEgUXNKK8TrqcB1YlaLhPfXuUPfi2ExUZhHwvAx3bTyshbriEAafYDv50y0M+71T7W
ovzO8TfWRMw708PbAMxSNLCeryHg6U5Jv7CWvREVgDCLom0BWNFy2iOO0HkhwNZSzC+ITyUGZVEw
xIuVXpPtjhN8N3aFq0RZD+Ygg4THA5Zb5megVZQoVc3gxOIgKVhrTeZYO6v7/VMOR8VAUAwViqFh
nl7Ph2KWt6tRCoI1s5uz4I+3AgHJnoi+NanxRkyok9S2Cxr+IcmTnL4nqolsGDP8Kuo3FSJdl0gh
rT1Dirf/UPerw6zJ86tA+3OY11u6ySGaCDLJeWIoM++qi7QuXqP5GpN3LhyM2uFG4yBxRgb/pebQ
YnW3kmPYWfeSUj11ian8aNqyZwtV/33SgfFulbbdl+z3H9RhpcOH31fEDV8tr++MozP43sl63kqi
mHDxtNR8YbdsIviVJaBu7E0HZn9TJeWb+wrZLcR3kuLz1S8QtqIvG+eK8WnMT464keiU25rSJmxW
IWvno3/16rTK9v2wJJhJN/NvTFOuRiJh4Vpcq7J6XU7PjgDyxrLbNfVp4AIstHJcqD5mDp22Ed5r
pz15VjRs95Al3YyfStC05iDLfvs2MFn+HzDRTWFTNGzf2Jasb9lpMcxtU1FnSFqrF+eP51m3cMio
kRfOmvWizZ37mGAgP4D4M8Fl5AXnpgQfOXgUgTw0prwsoTSzqcQ2nRdQa3V+Pio/kxYsKe1czRMv
LYuOgWnDgcW69suq9qtHwElWM5kEiUTMM6feUhnmfGhz9L3Y2VKBI/5dcdbvW3VabMAjoxC1iQHH
FgyYAbaOTinoxQmho6Gv1JpoCq+ArEiI2/Hq+5ehMcp4VSW48cpJXwla7yO6G38w3GaxsGNX8LxM
SYg0Mg1dSvIKWJy/Lb6d7JPe25x8n92lqrpKJAe2St2FiCueb955l9bMj6fSILRCdjafl+CUyovs
j0/g7WLBpUWJ1rrIzcYr4EMKPsL2cADS/x0BOnVFoqEKdVByLQCToILUq/vYyiTMCyU2TKzbcvBE
NOISs9CjcX4x/o0t1AperLZG1otVElNpBov2hj3D4t8d+aYwSn953vA5WnbbW7bZ4QWuACuCAxYB
BdAZ2rzqmqB4dahwXeSBTs4NPsqMwIUBEDswotYwEkS7ZnqbnP9Gxybi3iQO8aYGNn6dMUgHzi2n
kuPEbVFvadSdRu1wPYrjHTgdiKHNFer2b2N6boX8GtmkIIqzGQCNXM6rmv/6zVR0T0UmGeMCpp/c
dNuG8chXAN0UtN85ppzzrl/HEfanxZQZ+Eth/eBqf694AS4TCHFcQ++Pg71amVQRjaINj66TrlDL
6cW6/t97QjwAMYTxsNAcBg8ZeEmqQdY0DNOF727JGRicCagjaJU7Gi9otrG2swIjWun1dx+Bdav8
mSmRGM3Z8lbYp6LWhQWuQav7KMcWg9y/MwgpcZSRYzVvZ1ifSE1Q+xAimybghmBj3X3T2nj/Yhl3
Hk6ai4y3Osbg3xrbhEHfFyFlWSWNShrC3IWnX7SD4WQ4+ne4Q+SzSWqQnBcAtukfNKBmry5Cey5d
ScMi1iDE9hS8vboh+wzPl2EU+iOINED6pefjNSVHuYVD0NmwElN0PMdL6VH4DCb226iQvre8bGyq
x73wNZY3bHslTYpyE6huCG9eUZw3+r4Y/oD9WMLATeQTCJx3xtJRi8YvsyOaE7coRwTat/Jr1hxm
K2h6I2GJwXtyjFHT+nk2e16D5FpbR9Y67Bol8Os1kVToas+qb1HdPTWnqirR2ziFT21lE2sq2arq
kys6in+qBA8dkCD6rAebkqCh5TyF3FtZGTOs4NbWvBgxci3usWMhR1HYxE7sWsW5ghAR1Vbwgv3O
BW3HHESoUVTvMtCI/ncbYFdgv/u1y3WoeRicbjPB94RmSu2/ZtC9sz5qfxXN3IZiofS1QJRvyngQ
i3WkY6YAm2I2KG/YG/WxoBDZgF+hU1KJnlDkXqfztL4l+opiKE5jWJ9vjIM4r59Bn60+k6W5nV0z
LPTuZZ5gHDZq6OrhE9+tRS82lYerBBt3u2jV3PkmDJ/OjBd13ggOCcRha9Q2SOWtsX0U6EcKL49V
IxkZNuuQfEEkcj/+K1ggXFtupr1tHeX0BSD+pHPdxpmffkBCCltiPht/+81ZYY61dHiwoZK6doKf
WHb2ZIG4rStRJfgA/KJG/NYp2xHwYDspAKQg0sFyG0c3doFarq+pzhb8hxHm++HoIbffmuR64Wms
o4s3cZKjFF8xPm+VBB0o/Yelyv2RhdwCMU9UHXUnQSPJK9oyvUqqC3X0NTJib7hlqzW0lJ5nKfcg
+jUvJwF61WFZW3ivla/cofiKvX02ooFxgYV11MXMfFMHKGmz+FYGqYGs3prwfF1RLFaxKJuFIOs5
VEdR4WhK12VKZ+BAe0pfcbE/YbkcDsuzFgRFGtTLbYUCxnzOVWiaQ6mxjNVO7JiqpTPrARQKRSx7
L6E+tk7VOKNO81Tp/3zgYsnnKdl0WqGBBmguIE8sSFFSVT+ONFX8AgpSFTCI2ssAB+DNIZm79R0b
v4vuU7VdxiS1Ag6MY+a+vKhqRbl+NpBhDjVBwKpuOnA4B0OtUXOPOfJTworyFAb8b4o87mZXfdHG
9ws71/1nZBU4Sla6s5wCNmUETgoeXzSWhso9sNFKJ1DEY9wirQii6g2cJ4aBlzK2x7C3GR4v1KRA
ztBf/CfAJAX+KTM20d2yZJoYPmz8ZKD6EO7Y21chMbC7E0bsi3Xd5frsZdXJyIEB+xGd/ndOqHsR
mg2IzUrWD3RjTomcrx89/ZPeNMtEeiHmeXkNX0WRvRXoO7EnCImKgsIz018MknAa810xvI4Gk7FG
V+jkfyGaWUYSNfRazNFBwNpMwKf+jMgvXdUu0Dxbeo6pHWvbFlJFSLrpfZAl4MFff2U4bDfABeph
tdgjIyVaJwbQ1FW4cJhVh6rYc2rrI8LZ3ELRbQa2qhb1A1yWml5/xo3/POCVMv2306e730t6bOf4
FZjssJ8Rm9KlrC3K6RaQCg2Ia4Fh6TdCiu8uXgsufkZvJTjGhlwnWsuDZ56hYzvnWJJ4gMrzS0SQ
5q5fSjiDWgrwRyWH58jY5aP8ewE33cVujCbr1zeXyuNm3GRF/QkP1ZAadMzpTzVOLI55Ukz7rQN4
zAJcrPLgDq65LNlq8FqioyHkeUTzDccYPO0vzDA69z0yyRujhsAAHYJ+poJdEmcXvDLbM4jG/7K6
r4UA4m74cn/73CKngogMyDh2I74YIhSmThgMojmtAzg1kw9f1AkcM1uWEXArxrNu0VFjdDN9t23f
SWASJEkYqW1Yo1AvpHlRaKE75tm/sn4ZGGLu7DVAQaKVRWkfSrQksr5FvbVR3CZVB+lQBw7tKM72
f9WePJHgdxIMPV/1L5VwLSysU1lt8qOcqIDkF8r/QUrdML0OEkwsLLZfgolozdrqQUx0u00C9/N1
ahrd1Tj4Mcq+5mDsvwfHTuIokfixMK8L6WP3CX17WTGLHXoykDqHg7DIeTrnFJ6XJp8Njc8vVTVG
1oPoDkn4bgxlO8dpCEPArSZ9Xg7ZYUhd4vALZ9QJQwM9IEzz2oUIS8jdKb/NGM1gZxKcu+UG+WpJ
bJjj1CECDWMFwzWM2qwMVqoNWqDzm/69+Q/PLp0tCAWRQygDbHIdIw6R0iUEmUBnGLHFuuPMDJVH
1Syrj4WyIZyMACFdaPdVn69wXMZoznFLtKsQrb+K4g096bQYQiXwTGRrZmSh/S1Wo9whuscyF9IT
oyI11XMbx6gh4TPADFPhAJmxi66PrQnK5v2Wz/1ZysqVn0tZ3dUKY1H23tV92CiOL42PH+uqFa1k
N37EjuNE4G+Y0HqUonkZF0eoBpkgqsE9XHQyRDb9h7X6Pc9vbi8pUPaMAnhxMtX1fYLJaYnX9log
uFWbLT2gGvL3jZXPdYe1+Ed4v56e1RCbYdSykajrZ1JYd9jbztsTaLqiRJnHzhfwaOQ4DydZBNjU
NMfYAMHuqjFwvChOa3VLdza7hK/wmkCd5iUow+d96/wRsGJv3n1GuBrx6QP44xWa+g5WuxyPWuIK
ik+2jWvwgyf7CbPBjA9b/3ySeXX5890RGIsxzkvmnVQiBuyf1+76MUBNYBdKlZWnLRWPMs0s1dpO
CII0+cs/VbzsF1RMXunyweQzZGgGkWdRBc4+9n8q86N1WMwTx/eJ6zAPer5QcA1CUkqlRXswJuIL
o0GpTuc7WOW1Hx82wReg9SrR7apaPFr7eDYSpXXsOVSxjREqRX1yffU/HiZKyed4GDupFZUOJPZ1
DkxALGae3rpdQokGjjwALE1jsmSi5j1XUSd4Wo6E6W30oVQTxNno1Yp0LOuBFxFBD7p4/8VC8v5G
jvoc883fMbElgApqfSceIPR9inx9ZZ111+dAMMHA0O6ZDn7gQ3TUcgvVxxjtbAST389YQ5AXMaKg
o+5R0p/WPAV9FKCwRBMVPIgC7/jj2LtfHWxTSZx/0lrmoZRRRbg6MOer221MkfhL5to8kHhNIKzQ
lEuSmMh2NvoCA4lrUC4Dhx7GbhenR2UToGw+lwLItHv12vXpux/90lhekkifAWwWfp5Gnsbt41Fx
/t6dHLdRIO2UAYBNuZ2ztx9NXCUoJgou0a3ydFpatDVChyFJEiH8UkBmdyLVU4nZKIPRkRlhESVw
KdD1XaZW5I+8br4i+MJr43JPae/qPePPh8qkdwbIivIwCfXDTnReR/SgCRh6lPWvfdbF+4llmNGb
xCHb9DdncPisQdLBOlJilH5MNt2w9kYYQn7+t1+aitEkVzcQoVa5crGBujOKjZ7trfiMn47tzsx8
mCdW9ngFVfBvZ6FzEIrxj7DFGSff/kRKR1ZS2+Eyi/Ezvd2NsnTBBaKO/gL05dIpKJLFflRe8B2g
RhtmmTWR86iJ6okfTvESzm/vlf6t7ThpuNSKQq2PR/SzSoqVfuJZG9Kr9rFHTI6vd4wwci+ZadhQ
//mryMFpSgUMF4SkA2HwyIz6Ae2lI0wV2M1fTjwQ5WWEk5nkUMx9C2N03V/vqZIohVtqi8JyHrsc
tkXt/c33xIuSsDDG9RXwCZPXo3+3rG98P0v4q4CA2f22GRplU0eviE1JO4r25Xe7tALWCl/dTwVy
SYz8/LJkCZDS9WlEuZQIc4Sezu6AuPmV6eXPdQbfnFkEH8CWapcj/J4m1QfPGg19sCDUyjApL4G2
DhMjdIw9ev93xoO7y/9w553yxuY0z5gNp/873Ip+pzTwRvsC62pLLg0m24hi/ylx36Y/1I+mg4t1
VZB3jIHE912QkYQg9ebtNCOistwIzMavMZZLcyKMYbMluA+ofnLh11FxwE6fKrqmKS6LLaZIq99m
PodzqumRBlcrr8yGzsGagh37NStMjIvJ2uhso8ugzvaPUa+fgOEDUMjwhiOWTjoh1S2AoWI0HqR3
Kh8wgDPHuxU722bxrpHrHoCJFZOJffIwVNUeMq5PSl1G4EnrVC66P7f7x5IPQBnzAwQd535/2uvI
NlBCR/qlJmphzQr5e2Ri5i2isCbObMAxqAM1QbgvIN41qblK1qkyDAmsUwnLke3ZKAuMdsROvZmh
2Eymzq8V6+ZQn/helnhCNjkeyneTgUGgfzYBXELBAVSzLcIv/95BeE8WuBFVQNGo2pa6iWD/X6J7
I9Ae/6YO5szYz8umJEnFAY0kdtdOpe0eH0ESO2DeStpyS9OYPsvokAyKUTDxIDc/Q7km9pRJ/ba8
taa4FtAInMGbjzjWMCrpggEvugSxUIXAtGFxgTrCIkeapremc868YDbwcYCOCQpZiGne9GDH0+X3
7vlVm/kuH1xKMw4kQ6aRlWkTwAiQxeD5aRI3cSHO+sEYUanMfgYVL3vNOXuTeOB6AJXdfQKjbGY/
KWynnMWZTQxuto+ffeSyeJua6yyIrOcP3SdBjxpDs+X2PN/2CNRGIRfgNGGJXxE5supUtheZghCw
Hnyq+9VEXYOqA6luaM8c4xurYC6mGYkV7+BeSJKcJwdb7CRzdwziecUPQru8EAENH5ySE8nOnm18
JXawm99+nY2RYQ8hE9HSI8lbiam2aaNkp5En9mi8k9YIIwk/oxaVhXxZjW/+IuQf62Qt5pyBgOY1
zIUeRgxl8xrf8SM3z5UFUt8eLX8t4rnELWMvYsxjP4xkGxxRH99UPZ1bvw9gREK3xSGLlPvBdCia
qVfyqFWL95qFc1lbhSP4beItfxBpSL/j++QJrpQP/QFQIkj/0RzDUEbt6BWujgY1aoszysQmhpyj
YiYq1fF4ZhTjxk1ZSjQcsYKohkzogPMn8dYGjkPw5j+K4sODuwZkAE2QOdrveeTz3fltUGrd8kIl
0pcO8wKr7xu6GkuGMGEnLeSPiT7ILGU45ZroIEOxPeKEqHf4Pv2wE7+ZofRIBtM2PQ81k43DF/az
yHjGqfo904CXTEosiX/dSaLxjE1tq0h7Fi+a5oGQRzl6fxcsiNTBFa3eNxdadOoaBjUl9+L660YB
WkRveCbhyQBqxSaZ/ncnqEM1gJQrBMhEfUAUSka1lVbYPrIv3kOREiSfS6TYtWUnn8MyNSQ/kYK3
4XzG9PlZ15yvJPbz3FueCCl487mdXJX0FLpq9XQio9a6KPNaV6hOlAuR7JqUMmrWsOgGRNDd5MhR
rYE8PE/EVXH61vx8I5yrzlVK6bHDQLc6buOvJdmBetQEwrOE6u1PMYYF0gKBtm+sdXfT963FtBPK
de8rRrkJbDnotFzUrilAihHFwpzT6FZS7cDU3XvUQjJHL7/NncMgbWx1rrEnrVeSF8OUwoP1BrQV
0EoqfOlkvWCA/A/zFy3MxlPHtmU+IcAD6Lxh8BRw6alh0yXZhRVcy9Uqd2n7eM3/4VceoJFpFant
Q8ijAvL2OdB5AvJMYSt7YzkZ2iNzQe3Y6d+z2kxJTTxS/uREDvSpM1VSQNKmIBUIg8NLAFGHfX+W
0tBaBNLm4g9q0I1MtTrEkLR2fXP9PRIiwV7zG7mrr4j09IddYcy6QZIKPBkjO7dfnihSSffZhUJb
r74e1iNBNLEBf34hm+S+MJHpYBeG0DuCkp1JJXlPvBy86OrWxPJSdYXFWFFQWi3KAv+xHE9+iHpr
88wUMIkarGvfhb3QrZZ3eeYzsU/G552Le3T4Mn+0gBWfs6W42qMMlV6BYC8xB+LfYSAOK4IuVbDN
MHO7lZA0eRENM9x9niyKc+UeUcKeNwfkGazPagE1hcADcLMr6kwZJgEI8dn26ML1wbcWXii+mbff
g/6syRpUQKNdl5O9SbcHX9Ce6zBkyKNY1dDR2UqSqVn4db8foHj0iIVH48nBeB3XIKt2VNhibzzZ
UNGbk9Bnv3uf5xgNDuv+nTM9/s5eXJXp/pkfpTra4YujjTclyRr+uOR/fHHmQBvNrSxKelH584Vq
gRKefm1+c+QSmdoJ3at38ntfK6IXG9MxIVz0oy4UB+KApGC0PYIHk17DJHrnLf1uOHzaiajJAsm4
UvnK65A/fTF4fSUTjyTZBdUbbIsEdMb/i3TTCM/g44jCoM/vEOw/TbRjCAZodcSprvUFe3pMXD6X
7bDwmIfHnZkPsUzgi9SybEsFalamcPPUVQ8dX4iJhdlrrP6d0YJFZWgm72GSX4jJjqvkrlnLSK/2
Vot5yQNpITeF0Quvoqg5tvoRFwA346R726mJAWhMhPV8fCRU3guDt6Wm9C4FcgZwdx3B1y3nU8b5
z6pOIKZkL9N4nfxN2A9etpTQZMx+kuYRg6G/k83kB6mdLnTXox1x3bd1A+UUKHiNUJMw/rgDjlx3
aWinUvZt/8UF1cw3YuoQPcymcus5oA/ByTDj/3Aq8NJ29NsZqWfXmz90beIhxrmZqaRZk3uDbk3M
L7S4EV81h7boBuJkcOrhZJEyreLarLt+8AQD4mrh0L8ErmFUud3WyrOIbgBva9f8tc4gLOj2Ltji
hizrQQPn09qlXyN9LVxQf1i4897ZGNi8bKf8DdtHNuznTY6c4YtIUp2qD+X0q0DnOHsTIH4jmFBe
H2xlU2tyxT8tF1/Na4c7thm+GEZzQEY3c+E4uxuzgRpwPFdCvTZ1Z7bIgInJH8bVFQjnNk1PTtUp
lBCwAabkG/Td2a6TbJVPGSnNB1tStCUNmT/Tk19nrNm9bTju8eR/TXONNEgywfzMl9iWCR1cpjsT
I5HDqGXkcvggv11SejxAyeqgN/aGph+oCWQl5u74vyn4HF5LYkxCjPNwehiBYsm4hZknyz8AQyS/
8oowNQIJvuZiE8QMEMZAdfn8mNJPcAzsIiTxNoaYKnOTbKhC1SnGDjlOEomhxBAikaDrc6ITkHgP
JSGZvPwJRC1yV0ry+9mvG9r2osFHkqe3A+R7C6FE3c5zxks6exBDO9AxaD6pybUVK3Rzzd964MJY
GYuGssdNMwShwpoCmbmDBRHRY0d+H/xewoxcukIckX6Eewag4Db2O6lk7iXXvgmEa4BQmNko7Xhw
D9JeaNipAgoKMobId2C3l0pUNYFvbZT1AO0fV7DSUK6NrWNP4Bu79O1cMRpmw544ZlU/IiDRqigL
zjKPDut2iBSBApZmav+zo4U4kszApHVf1mt/KAmmOzODuT47NqNmeXo0rANkse8vgauFVMbR+IAc
dMIjYR4TUMf1fA3pfh9H16Z5p6pd0SjUekSGUALPqHIaS/yPaWq/AyipB7fRaIibZCNvWR2zm5FV
7IL/yB2Q7UvP88n2deino4ibJ4mUW0xr4aZ1IaHvG2RyHBqH98svyZ3T99gdbFg0rWXqIe1KVV7U
SAv8p9HdfRruYvCieq+zrmAS/+pq1a/0dhnf39DuEPXzPZooqveuiRD2gf1nd4hZdGCgT5s4nSpP
AqjrRp1W+SSUI7yLX0AILOQaoIPlVv8NTWptKouFa6tf3nYwPNPrzNCs73wErBFNNJj+Rg2HN/5n
dlQDqBONZcwLqmrUEenR9JxD/tyIx1NYK9vzboW92F6RhoXGuAQ/Ig58d3mDSnrut8ZYrnlClwk7
1y5Jj0iRf+8DgrCKVN//965GmjqSN7nRhkf0BwjBWdDQ6Z2vlMnh6EE6sk/+HNcSGQT9pMwm73lj
GnQ/u5kxulcfdMpyr1GFCWmjPlETLzb6qNiqn2GBmS2hBxLtuYJ6hrFjPQEnPaaCuQxggNJsoprv
xrIdAzDxOqzh0OWMmRkFtfTBr0oMcxJbMHxLWDb3GFGG1PhqCOvgdFXaqE4ysP7yZDa9xs2ZLCk4
fN7V8GPwMipkgvD+VdmEahhbiL0wNCM1ghFdsxJQBMuwmmhF9Jtp0L2UbojZtmQuzTxcBp+/85N1
RBh6cj0KIumSfvnfm5l/zPP4uLA+TuUqnwbAPRjCB3wPCvutrYsOg3Nr/lP/zeuvGDaw9q6zXwM4
Glg1ZWbVIkHrJRc1tRGdXsjWt/Ezr0A5VsYmO/5t71dfhlAvtSaOLMJkM059hkMP6frGu+iJLRwc
Q2wokgrLw7LX07AxIfs72VQZ6Fd3R5B/LJWFyfp+Dh7eqHF71l4HFsL3ZJ98jOCoRRy89TNdO09X
xomv2/R83IK6mwLuHdo9mtJ8S1GNjlW6IoqWmZxPHliKg4sdeYJ7SP+MyX3+pFIJjRLvVAosJkYR
fQAnxYOzzv7zhKfSOv3KmlRvETpujIaTWFVqNnXACJGG26ZsNmYc7AalE9dNODXRfFp3EaNqwgEm
V+DkAVcb3H74TBTo07P3eUgmCZfHa7ndKizHxsrLN7hp2p6T9WQn4pFOwG1xQA+mVzY0E4uPpQw0
gGpXBkuWBm883If7sIz9t8KneD8phYyAbecX9SJr4xPIcAHMuWyFQ5G8wW1Tiibb4MScXcts968q
OBNkLkbEiBQQUlXAyvbvmmDjEHBz34OOEstmczVXQlDeQsI3J5fSbyU/8V0NXS/pMjJszG190Q4k
Z645bCmSUrolvn0JJW8oWAw4lez3aBo8RaJRvart1/F5jH5z6YQ3Z9lvimxrgk41xFLXjTgI+kIm
uIHn/Z1mPxQpPP396b/iiTBurE/Op/pWbRcdIKiM/ETfHIz8Xayee3GfkWyGD0anv2nkaArKKlVr
E9PFcviVuyEaq6n2Yu8Pf2Jq+x76xAxDj0E8Ezs8TnymyR77ui8UxPKqVTZfVdu3sqPLpTpiKSzZ
fFm/4ABD/ploz/o4pQzBRumK5REK2zPpYqYu+v9RHCJUaAiDnBh4tpv8kc+IoxZqKVSp0m1PQf2F
J3y/3plCSytVZifxe3qk+/PqlkbW75UHwQipWY4BZJ+a2goLiSkXYjIxah/qUzStXY6znLyFxqGA
e50p1G0AocH3Vg861/p8pDiRPguac/wEUn6+JtKUuUpi3TMEtiqQDi130rruKU/Sk2tyYif0qTdA
/c2KBQpg+EADgFzoI+jZdMEWMY5HysuJD8/l1ibBgbCM7w+hGCDBUfHws8OH7fVXPzsLVSiUjrFL
mPvC1r74rxnpR23rQTr0rbMhQluvzzAc8ZLi8eCOWZ3kTFh/Bh48W5f/Uh2UOFQyZ3YpSHteQssf
plwn6WVckjEN1Hgs/18eIYgbqM/LcjZsi0qBxQbRBsYImmIZt10vmB98bnzmxE3T2aBTrvAJJhBt
N6rUGFTcW39dVUld6AmzJ4pjR0OQO1L90dntgJwkPeUMkdWYGwR05lje9jr5wK045QMTeohr1YBa
rC9O/ja6z5dI16pI8HuOnup+gYDWp6Fy54tkQS33s0HnvsaxnYK6k3L6uvNx8C+cV2nKVOxOyPk1
TOZzK4HLrQ6pZErXATSJoWRsLIKW9QtwaNUdNyL9s86pTEbyaRdeyY1EJs+s6eEW/98uDJcuqWvL
Cs8UqyLCyXTet/yhAFtBqaoXHZZWW8COBQd/MDWPuWlnetYJgNJGDI5m5E6GuoZsXjdVjssvlxHi
1WE/7XsKC6vd5c/mIZank9p1WzZmvtIefDa8+uyfDC8YDY3sRxwtzrLOIP1yx+nCCY2GnK+izFF6
ot0XoXEGklZRMjZFKZuw9CMlaCYlTDrxJEtcZQP/yko3EtlWp5yVJVB50+AGEBeD6VTD3u6jAt+5
x7y8aRjqArh7BPJqCCFy0v4G+d85C4gusBWlGXj7BHrP+0zLZ7dVB8K0JTiABYlAHUCmlSsZRuYN
CW7SM2cd1MoN3KKeqC1kMG6xxmjfIxwN2HeNmjbKJ98HhOddTjdZ2m2+lnvVoFxHHOKzpSdcAQFg
HpVkEzpmj1ZI1Iab0vtxExCYbW7CMTYYP+Cy+q704hn7rIcI9DqTsG2tLpIRx1wVvoVteDHHvnf7
5uDEkVUIgjoY/MVEC3vGV2LvgGR++M6w23zvLF8e31d3f4B+nACKdeuKJL+CS6FIB/xcuAnfg+dx
0YfheOQMK/chsa+mG56mfhhhJUbIA+ZnH6xWPltrcQ35nROV36o39FGtKvvcLHs7TAXPhporoILk
+8Um5Tn+MELiWHZmdXs7+MMd3K6yyAwcTsCY07ZUQINSIKttqW9zpHLYfanMGRLJTf/anM+QKR6g
jEBV7OEYyHmri/KjFwBwlKq4B6g9IPOIhD0sSreSwnphTgO1aor2PvcO51o/+cssfLbCuoWAJTBx
pASLwXl+FNFOslqVc2sMnramq1BHy3NhiX7VVKtn/JNPoh+QSik5S4eZOxvik79K4IFxzktPFWjh
Ftb9Ug/WTkzo+HS2YKiuSTik6EduJSUB49Dx5t/D0sHUuHt1nj0sVHQ9ESYktpBxImHGK9Ey4ru/
Gu5u+GsUyJs8sKjw0Ei04egET46ajl/+zWVgRgqaEYjYG3CkC6OpP48hQVpLRDt638ft7tkvD4LV
/7gEfqHTkOcqZCzHgeUalgWvSN8oecGuyPmgJEXZ7V7ou17BsyN4UfZzy2ZbHdPlQQt8DuftSGfx
+pu7xG0j5Ll78fY+obAnRBE6nMzMSMoZICfl+t/EGg+b2JW5Kzlk0FlBY05PWb8CLn6KYgaTgqpi
iTnh/uEixKGKuYWJhDvBbAeG7pOnLCuvpg8oiHLfIVU/l2qT8imzWJutUcpxw9kw2gGxGjghsYbR
Kwp9FaA8XJWp4OR/qvx+QqfBE+kc+yoe23flbjhMseNyOLIpudUIL2HIHlByNNiSsLr6zGwt/g1P
+IPmd7JuPUZ+qURMBDpTjvqKWcAaLCSWDYHKW+hJbYfTuP8WzshOpBQEFMezvAl9Cf0Fc0ORUNvv
5Qx1oic99aKgviaE3sbLYhxC2ptAQSQfGllCE0f/5TTngTh6YNuKInEwJSfLdS96wdN32elccXzo
Lq7aciqvKrpFzgGbOpoYQY+57MwCkFutmc6pAyzaxWgymcURPkQURuBdL0HnlsG2ym+6dEo0tIdq
EjJw/JG0s8KdLZBUhKW2ezZvc/BnN3xpn8MjJjZmqqaKs/COYZanACW7/qV138ip5yJnQHnRa5Hc
2qJ1vEj+SKuOMlbLx5krTKtOgbXs7O17jds+3/O3jdgRlbaSNYFFSajZsFPI1QbRLSkqH9l5dV10
rzLdXshXhoqBhN7jUsOVmW1VL9qEpe00IBWN4aD1+ypNp8Lw/ZxGTh9buKCPth66IoFKWyKD1tJR
gzWICx2bXuuAzMFJTgV9Rip6A+HNHypgSVb6ULF3Rv0apaMW7MOKJc9dg4ryNqchFn5dfMlTk08a
iVsnDwSYKjWlp9mam7lH2n8DlTmnQFw7IFoctWBdlTlR8HOdzIQA2p2YozekoArArfDNENn3BOoG
/3L4F0RyO+XJgv3QAApK/5K5bucQixw2q/I6O5uPjJXKP91UHfmcat6tPLbmSwl1xDdT4V3xGOZ+
jRqRph8DWjXrnXPX5i20Q3SFPIreXLPG/LVftrugcCx6ca72dyke13+A75ESykjV7qtKpC7QvPwQ
6QELR15B6ioJQOdwD96Y6cBTyvvy76iQH8wllcBDZvxxVf4r2jsYrIzI9W9BLKyzZSwo+LVWAFo4
uxmUqolL8nSAt2tFxf7i2GZGNRZq6Yo/hxTlQuJ2MdUD/atY2TX18n4OsDxwTKZ6xH9LLdS7LwAR
l2GJ2qHAv+hO61NmtttbqPCZU3+5oEdyLwzqqOEOgVPR6xZE/fGRYrHa72qFuJSm6vXwfab9pDph
CZVjkTdN8+tcdZa/p0GIcRxGsVqzJBsFN+3GZ6OTCLG5VW5Gf6CMDOywgtrBCZwWJXK50VKUX6yO
HoNB4OLoRGwL+eBD0GbR1i3QMohR2mXrZgIof0nEDtnEAKbcKVR+3kGB0UYl4ZLapEgvma18dkwJ
RvmAqiqWX9ZruLn/bBCeEezCFoUCcqJYB5xbvVYIgLroevmwR+amemPV7rMpsF/Ja8NV7rGDT53s
SY1VBnzz8xTZFR+j1/TgrlbTXd+MNsSfDbGX5cxB3qX+5AKhX4IJDkuQWfHKjhc8b+yesYGnwGhn
orGq5aLYacelAk7jlPblkBPgshqMZLBOXjs4zVtkMWamwYlPT3bKEktcu4/S416Cn7SAoAJDC8gd
ppw2wwwsWqQydrkWY7DRCZ3Mn8rjDbFFUlXQof68WVOYWgWHzQOFwUDTbVAMigRbFQh5X/JT+4mN
/ZUEwuuQr19nL3nIGEOb5qg2CYU4XgJYb4ooxslX+NX3EdpFcCOx1xBu2rEkqfhNcQ3NRhdzKG1l
JpTrHy8ABS5Ozt2IqYbd8U87JGRIeQuuP/1NL1UgQnnvrdkxa+Q0ISMqFsP3M6d2mB5iuemPAdaD
HRfU8x2NNRExzGEbfMyai0vriuUNYIPs4Wr70tP3p/CPXoq3TECZIuv4M6V4BWHG2WA0xqCaemGF
rJ0xSdvKPV5KMZCCNzwW4FCO4nrgL70ybseZuAj4kCCIxsEjlTjVw5yYSehv+cfzHFCq1OAELNcM
TJzL1wZOHzZ80gRjrkU1EROyhx6DDgERTLxkptIsGW8OGfRny3hu87D1lYYHRxDOTAcaG1ouSd/v
AFGYnrViUkcsAzDSrzDQzpfxgq5+G+QpP+WNZgKrYcdWjONMZ6cLe44/wvmCfOuyhKWyReHEzfP5
c4CsVENJDC1nsizKqIlB/Kh2ooRiKkERgDb1t2EKQWornEEYtRj4GK+grV0kaPpuwseGbc7t3sSF
/QvR6rw4QC5rNgdlP/b0VmHTjDl7n2a0SVl4eUZgocPuIKO/mgNHLW1y78WQP7DizI0sCY74qG5O
af60wB2VWKzTblCCxCJW4thQXiEsiSCkZzZd5fimQnboOtmK2CFxi+alehEG4RfL9MTuySlKCGYa
jwhdKRZkPxrkxxyi3rN1HAqS+fckQhWFUzcQADkjkmjg7YOwNZym5nb16PryHPuuH3s64x/YJ7dc
F9r79/XAmt0ww/hQKWS2Cx0xDtUdyZoJ9PnxW03DNfAiGdaHLwyng9HBpH/+K29T9ubj1pLh1TqC
0fe2fTiccPOPK7crALP8Zt6wTi0QraXTtzBMO01Qu8xbv3noX1+ncDSlHAS9ftgKg+Cr1xUfrKbO
u2PPaTak/RNYxWleMoL92gjhBwregyGmJV506kMknZV2QbRrH5q8erwFOrpxZI0DxZ7tXLBikje/
lhPg80Ht06419Kwp3EY4O5gE6jDAkDI4s5KABL8+UVG0K0Yxm9bFzBbMZ9o1XAgV4XGRdJ/0WOkE
DHx2Dv9ogESZhwDs65ve98hV5mY31/csTQ/WLAsjXUeMtHBa0/TNf7bHdQh4+wo6vdhMuTZvSoYF
P3z476reNKlDHkBPSEROu/8kdG1xIOh4ZqL1MyRDAQHym0ZFeH2hxyMsBa7bPq130aApkUjWx5oy
uMvD35vHu3SZKsZGpBSzudNGEk0Ol3qDq3RnMzibsth0PvA+pLG8yw0+Cs6ltjhw4lCS2tueWG/n
n/01yY3I6YlA8mZPJj+n1u2aW5jGI5LRTplMvEvYfkIN7v5LDSoKfQcXbWjQIMxLp/E6tjFyLlwY
T3BNWLBMAEPrYtyMbgts8uwR9MgS848LJTppWsS+dDOUzr0gMjEC5tTyWz4f1WUIv+hWOqT7lC4j
kvMKAqxJeIqWoA3jY+mydoBZX+V1D9nBiEM6834UYRi0ZDncwd58s01WYFXKzMo8vr5vqa0MAfzK
gr+cuREuQdL2tCrbJZD5rz2SrLTHjtlxwME88yaHK0r+MM2y4DOKZ/NN/lBlKVfb2bgIaBj8Ar8V
kw2fDleFB8F/bMllf86IR76dWPkgfFkVN7ObCvZD23J9ovF/munrV/O9olyLaTie/tCId1IHevZp
ibX7S7wpBkNEyam3mgTMA1+jQj0KhjyrdOHtgcxCwZLn4yispvUMhW7kzoOxYGw+ZDFib1NnDUFk
306191ILFtFnJkTxNiU+PPzkuv6HCJrPcd6Mg+FAREj4xeZ466lDF6389AFgBHNNYj3vyFGk8BBK
2lkKXPuUUH0fwvbrjPPUtq3yDoNArq7dQCirQ1cMRzT/Jnd33iLqP7tjnggFy/mqrIZ2fw4CSkNq
ZuZSqI3ZN4PnjDYk36ylUJ8UcrUNbbO5PJJbE4BOFfc4Kds+fmdLjpeK4ymJEEDXDMkblFW368Vd
/UdTaMITwhoUK9DxbdkWvzcIXU4UI3sDm+d9VcPYtocxO5HRcULdDA57Ati88NLFAsRvPoBaOfXL
jE0G7RXIoSNZbbELt98CFYMFVnqWePJA2hYL4fQ3vRrpifOqoPBdKVifdVFks8cxYpYUtlVFf4ub
5+DdLcMLAHaJ2XnkGeqsB9hMWTsOhc8ZW+Aa1D8dRViQn2YO5ehIaBN686iLYxUkf+Sipi6rUf4P
LTywSnPoaff54DQBVEI+OhhyiA34ptSwCZ9TA7vZG9BwKeDBrY/JRfZfK+Y50uDbA+cOyD+AzslI
yl4B2DzTM7EbGCwUWWXKPHg1O4bitgRn+fadqi5lJ+KE/SS3HHvHgheSk6JSSTyFNTglrLa2rlwk
Q9mAQ3U28tG15Wn61AVBQIIsfB0jgvs2Lbi62FsgZ6YzA5LmVAabG+uXE2BhULpni71FCvzujyDP
J/SNsBQqq+l/LyDyOFJkTpa+KIomVXscynKURWE9h2pw0VXsniuaCO8Y7zvXM0gXx5lgUoSLyzAU
q4t212Vs+vyRjTYqRVvqH+sCMDLJw7SKyuwZWzE1fHEN43mgdeJwmgf4IkK9YgGrdloINDSktx4U
xfkxqprsmT5DdEUdczM7Kzi02StUVNK9CPQj4AVBDe+6MaJUU4SGQOvFLUlWNNsihNnM3o8LqSfd
85t4DS4PErcHnmit5J3XvOW350xz+x/FxJQ1I2prnSgYAy0w35/7XM4scYgNUAu27FFucv6uuqO9
cYnUOk6TXQ1/x0KIMPG/WE1d9zNYP3k+XrWwn+TDXI1t951F9pvzEW1p2Cj8+X0f7NQaOeaZuD2A
k8XxI+2LPZsIXKMXfAk8zMA2XBzk5YhpWfT1JBJm94DHDCH0Otxjpv9YrRKd2fK5noLbPivdYP64
/4zNJ6+4VeJbxIJjgK5Sp+yzvF/hRA0YQ4o5wytJdN2+t/jLmeN5q8gi7QmPlA0tPELCzkiHTHV+
uWkcOUnRllduQI06VS5/PqshgAoRn2b8TadPG7g2Qm+Kp5CB8vSVgLB938rNpS64wz5E4CKv09CU
6hV2LHxeXuZFt6bVM3QIcUGCVMM0UjhEpPLSY02IgXTu91U85b150oispPn7DRFsAgNG9CN3Xnts
k+lw50os6mEcVzXc2+DwKNauTapApBKkqCsQMbzdcaZHocLtwRtvIq2ksPNqB67kc7JZfZJ+M8rx
07xQUPynQGWdhY0GhkJCcc/S59/RKJaLyTfXRvG5MHLCkPHBPZ+cz7b4krOTwkrcLu+wOUjpAL5E
uQIg2vwcVnRQxysoRyKIS5THHwA91jgDwLw68s81pOqTRoG0vjtD1LgsUyl88FqX4nPTNh11LgE4
T3wBcOQRz3PBwloz6ID04FNcbPdtF9JSBdyzPPhpBL/ZyAWC/EgTAOQ1WBe4WKBv/0Xcep1BBr0Q
hmpKNF04vXCrxOSCPecPNfedmYnT4R3Nu5ymglczJr7pOnhsk+gsr5dURmyNBSawrjyEh/62WsAg
66pe+6PLVg4S9UPqnSOMLjHPnVBgGRLeOl4b3VE3GhBDENxqkc7c2wDNOf2LeqFr8AHUWWj3cvng
kAksUncVDHtHrpKvn9u4BuGYitkZrzPd6xd7PPDUZT+uTJxxWfarLLBR8Cau04cOZA7aaJfOVMbO
qnks0j8U53P8tMi7qfenzRWhFr0Xng3CmkvFTFEu5rAgICJK4uHAeWDh5NzrRTytc284Txyg4Laf
E3XrzJL/ZJNv49iaie1D9HNRNTT6omwVVqhrTN9bJnWMdEbc8HsmkmLWi2qH1FJzw5ggHwKq0Sw9
IFPOYPyqUVSOK8XoR6/50g7R0vhrr/jyFukNBelXm9LWYAzb83yKQthZL42ODpllQOk2onVeRI11
qYhwVE8sWR+dXJBThyl+UO3FfDz5+/jb16UBERfG/s+pBlnLj7IYX801OvxXTo22hnOcc5qcylUC
kzBSCIlmrC3aicpUQhWM5W6NqfcCUM2lkj6+eXpQM6JqtCA6wicQJnuZZFhkQS2wB08qOuieO0B8
Cv8BWiUJUlN4gTepoo9KLY/Zh5lVq9fiWFH8AvRLFcsnRXgAMVwBbmvhPAUP1qUZNs6Ers4Wt6FR
ElkPs7WRiSH9B9fsUZJksven0OufOWMfx4Aw5SZbNrKEB1MBDmfuENsj+3ZZeXDRWDQs+3ifSpDA
VwASI3k6Z99OpoGuip8GiAwQK0pm612NqJwQTWT08OTnvk4PwFsi9kxa1VsHJuKcE0UV+d2buk16
M5yat18ecSCnJSA5qTkKeKLmtnYnCKV4gEibSlcb0/2QlTEG7KNubRy3Wfv9nSi69+QFc0RlANjQ
hKXY0OkwZ/mn/T+OzcPbFT81N0yRd0HS3Zwu3QCB0LeNsrS2j+XvXodXUOeT9LX01zXh1xEtPEid
nV0Oui6bc6Z+EQ2Dft3lhQ/TwlsBzrHogmAYtKdZJP66q+BmTBD6JNzNzG3DXGCkQcxlf9lBK0vM
Kl39PWG+enqGGxZX7S0ywwmb3EqPunruyNYKbpOesMSUf34jGJxw5wfAzoHLC2H0XIAYyFW3OboP
d7gBqrQFPykCsbnOMOn1mIBKSJhToARgX+TEi4D4puspt4TY4K6UGzdodLk4Hm3bwyK37wYTHtIe
48HP+znuOVXvnRxfyfrhjf2kS3m4gUHW1Z4UxtSHSUUnqqhZmGpyWEsYetzpCB59tgzC/eiN2kwG
ltZuJIEKXtN1PnFavW4GBWSnPIrOlaML4VumK7uXaD/8M/CJF7QcPyuA67302/deDTDJiwJ1LZfW
j9BAM8TW7kkLfOxYg3g4eOw6RtgQLO5WbtSO0sJ1fYcrsKBvMsWMOwtAXnKK7NPX9/3//adKVmW/
HIbKV/Nlfl35MXGcbiZ6ZPtqJWXShOkraGNun0ZFiGRd+qaW+Ci3xDEbksd4DuDzBlNT1S2wa4Xk
9csDEPOhMRRdie7+6EyKGqLBccZ2AP7VOj7DwBsqgKUI8FMKucj7DfM+hJSS/SqiQiKjCdDjf2qZ
UwRU8WU8PctIBPdZ3N1tneoZL6AT9GDkBTfk8RfcajMBq+h6SJmi2bRQ4mADWaP1QdxXAF0zsx/V
RhPueTrQ58A3TX0oCNIHS7SeMpxiMSeZM6JPa1rMxgYpbkPgnoSfQlM55ShcR4Gspht5EPRQHfZZ
56JuCtz2wuZeiD446oxWSHoyIqyZWg7W4hF+9FwL591qYj68zilrnR/asG+xrv8YEuVGPs/gUIzS
pHz7sllj7BnS0/BSuady5/LJ/eMZ01mfVWtqPmC5nRjfPRrHB5ZyJQICEWXC+MX78Fl25dPT3+Rp
9jgyCNxG8bKZoxCyT4/4kLpjzsh8EptavTSqMbstE3/iB/uDatjvf+P2gj2NBoJHIZwYbpVBOD5T
sLwsT2Dwd/RHs+TGDKLgVKb+ImQ6qq/n/Dk9HRWe+gxFpqpk6S27lJ01x1nDYPLCvfHnbP8cX4pp
cKwwfYQGFLQO0Q/wHjMnMJR/9KZfZaRcxEpioUcA17+U5XKlERZDzZKk6avrD0kio5O6Tj3s7B+X
Cm+Ar/b8Ciu1e/m0OLKUKxDzii/oLPUM5l74+xljjwX08YvJkv3RTHqC/1xpYOx5LFW5yAwL+sM3
J5qRUSeuxLu8qnPpfGfK/1IXuFkhxWpB5zqFipBAuDVrEHWk+T6VhJoJaqenWVVwpT0AF8BrECCZ
14/4RTGTmfHiOyIe4qzjGDvIcMy5Q/zOj1tyQZgEjQgWBNZ1s63sLWemvpXrrzQfy3TOHI5YwcQC
qnVnHghcEbM6IKwK6VoqKWI4pTgArNXL8SYgFPEc6TSxX2mmeWvKwRr1rGc15Nw9rtb37uQzSI39
Eid8wa/i+WU2mOBuGtB9qRtojY470tRsDgA4RaGBMIiwcMwOEeJoNUZKBgcRCyA3mPDC2oUUovPn
w7mft0zWdReZGAKWF2VbhMFI47ynNIhyqYRQV4D+t1lFhdZy7gXHrWkhF6IesGq8RlQv1A1djCj9
Hn5wRxSn7O/M/m92mJhaF6xocn2tXoDBBYhFMolLRpy/ddx/aJ83n04BN7Grx+EVa/EKeyXLhv38
U4FugxfUFKX3s7xjznp6k5WNtGZjOz2MPHQmoIWCf64fNP9grsXxNH3ARKBWLYKzhsnWAqbtuGIH
AZ0ed0UptwdCLWHuEncQXjeFuRC9Na1gLmRHL0TYgwf6U58/NHf795GezHrCFgADZ6zcsZq61O0j
eBZfTc0K0yrRegC4TY7OT0adTCFucPIJXb0hstRS+rGEp3piSFE0ijz9rqu9Ob6xy02HTVDQ8GNf
L+4tyPACzfpcPcWWvkQhhfl38LR28rLPRxR81YeBAfbGDb1hwUllb6xEdWx088yyrg3PO1L9wjsQ
5ZkQeejSEZ8U3RuchsZffGgdBqX/FdcGjZ4arGVMFDMHx02JP53b9QvtUQxtTazKrgsO5Zl4WzNl
t4UI3c988yL46eKY1h4D8DHlED8W9CMaVwpuKO5cuzT4RrHPLaCN8Zc0lTWa9+OI40bcrS03c9Kr
DN9CIJiffGGRh9vRyQZpm1bpxP7wzRU9b1HFf07UjFgdkIlOopIHT9aDtBq4P8JpCAcptcZRE+Y2
ABQwzEm5lpceSYbMw7EWR3f5s5WVS7GsbfbNMhyS+NtTSMcbd02ASo4uoi92okXHNtWoW5moBoKf
i9QM+/gUZ6H+ilE47/GfywIHYwA5p5N3UwZ7ingOfCTmy3CIBOrsONddMX/7NgVEs0KjnFpiLdUr
uWfMrS/O+zxZmmP8Pb5SFeLkmEgOsqAkoqB/U+ngIVFP8Hqk1QOWCqyi8+t5AoUIiTvyQOPlRahA
0Uh5NGW7zWwPlUKv+lp2xa4FRoMWHGSOdAzZkCnfxYvt20XgsM2gPnS1IKVNSEaMeq+j3rJQOh1y
BvcGNCn1vLuiGe/+kUBCQ5MALeKhNBG9LIeOV/v+0zCfImh9uJ4uKqFGLcMyGg8kxhYU9v3Q/YoL
Exww2DK0gDi2wfQ4xPdxWDMVG7L3Q+y/fviT/8RrUSCfKKurWaigvqEkMjfMjZjB8/TnJ1RaUzF/
hzcVrSmB5nmapFA9o8xII4gh2k+e4B5bt9Y/JSco6PQN5eu7c0mE83royCAQsLYX6KNDV9cGbAGS
r/V4d/iPnLbq4A61826W0Wb4KieCceFv+0f5eh4NaUnNshvPyHzdiCm+SaQwSVpZuapELQHH7eWk
3P+6UAP8LmrTzD/JrRHRKwdPrMACUySed/ujIwtgDu9MGoE30odssjrakUYoKr/d4JmorQ5cIUTW
RnWKI3F7QQO9VULk8ViQacWTqR3Jdz/Y5BJQnHVNMjkPzYnWQBkQ4ZOQYAPJBUrd00I56lBsRIwF
HYXVAB4Qot6BoFXmBd5Am5RJh/h3BvdE0a17l7qfgECT6bZS5Y0RWAAR6DThS4C8HypETYXue/WK
xBdbJXeF7uqWVtype7Ht2yWO61fVsRycda8IzpAq11QBWdY86jh6ngxlxoQ1SrusWBguFy3wjJGG
JYnVN2jBsvzkYDc8HDX90uoUqMdizw/J1rVCmfZSH8jy4m6OqUeL698SG71SjNKP7sFMvg2LY4sP
vxxcf21p+XGLn/k2L2dm/2hWz5I9jPWlc9/rXLHyG5Lr+poG0p5ERfMlHJ9hjKrsrZgpnKRaYHgf
Gk2ZfRVJwCfQ/klsbQ9jRFtb42IpW9mfJ/tHvuJiqSLU8COD4fCkwAlPrayqV/RnGhfqOLfBV6f+
8F+QvlvIrQJ3HBPIXgjmAiJ7NpsvCM1hUtDb43jXY8dV25Xo3BvUMsLDhNkWfCdfzFq4sxJBtWP4
AWUAiyZkC5+GxmTgqbabgyaFGnlGlSGAm5CqKKeABzqsTXmtl5H2nAWA7Jo+gQ5feQsQyL2IVVIM
CDZJfQWElqoYaSAEzFkxEfsaaHgWKjjfJqwXRLIojGJhj6lcmjQVp4B3cPXWrNdWiFEaP7O2aiHi
FrMsayTuzReBZsnVlxMUdKYMuFpcWgrP7qZ424BY+KxFAqv5Zi7QZ+rGtYs3CZiMV3mSLcWRmQ+p
xBYGTPIMw3mqizpAAQXc7XK3LqXnEhmtBe40+vhv923UpkGfOMhZ5EIyj4Bfv2fEyuiioveMrPIY
1pFt33YUwVFqmW1VuSo9v1CGzVscOYeHGD8qVNh7iLM1ypPEZpSs5PeulUxkM8wIGFXSuar8Wj0q
PKqwb9CTrLcHrixC1zUT0HAZP2r+HZQSlcnHiXeoyJg/3Jp6EZ5i0ukVZbCxx2ueVL/M7Nfp/LL1
Gtp3rST2qiCaOaWW8/0UQbcXBZJXNl85McTHaLaHlSmy3BpQ7omNgZ9L9x6cFnsh5SMG4qRgV5LP
jUrd5JD8QKz0yHKWcL731eqCENG7dwKAMHGDq+mfI5rE9Ahi/IGkyTJUM+SmPl6sV7o/r9s0C+Xy
wFsk6rFZUtZHpQkhSy+uvuAmQJDvFAiGSZ8iGSVXTVRoU+BDiyyEd5GzhxPfAiCe0lTHwhHU6taP
tyxNBqi0uVVDK67V0jxDGqY2Ewk1WuKzAC+pI7GiBNOSIaQ6i4fABlGtBlqE6myVepWJhQCb7rrd
KTg0S7FTStDDA/stsMRRvR9+/OrCF2rN7iWSO+riXlO+qcC78y4LfcwQbwpGODVBe86Y/00GiqQE
0+TWRMoTdvRMXwMoMhE6gd4OhCfbSRGg9miW9usfgmEWu8dQRME8JY7iCdborIR/JKMFgUzceqYl
WB3xofrvSubQn5yMm1HB3oARtmbSo2uNejNB+9qZsbyPYGNGvigR/nRqUfb8TIZqKHcNjVF1fyG4
ejNYT2S+69/qlcjhyln7IWH2pjEAcSTpndHFjySKaY/8ed9871C1VlWmS+E6LS46hUbuQvHsEJk0
LD27tR32q1kX6ObrJZh7mGs3DhcNfu3wOTTJAFOOavKR7HhfWVnM70OZvZSEo6Hs9c45OKRUg/Gq
H+KGMvI5dPApBt7thQw2mNbtPxttFIaT3IGKcTJX1POWuWJbjH8jTuYY7ozoCZ0bgxjPSHYYRi3J
voZ1tGRCI9BXL06Ac1DK7UP3RbMXHAAbLz4RWIIcbqJHVFGQczK7tjurxtqXpfS5MeRMlvNf5EsU
Utki9PNfwJWgD89XyHFbrMaJP3LkSNxsLBEB2+rps2w24HQl1Uj4FuoTqq+XS601phy6sKSSWEl5
5dSW4GMEaqwJIyQD7BIPxvpfbbSXfIepxv0C7qNniHeExfmGmM6wLeuzZX/pxU6TTC0K+BlS5IQi
jklIM+vImPh6s8bx27ivB68NQ2y9+zqRTdAzDSzdNPMBlrf2CNrw4J2Y+2dcCLl2fJQC2SgRrgxs
iqEpBeKMIMFMkUPTKbGoBza/qJ2jbIglj+tIh2VDDxpY6ODmTHxdMt4om0BIx9ZmSe2eri3kPuBG
WTrNrQOlFzPfBVCglJHvLt6AsJ3KyLQwrYnE3LuJEUIiwAh0g7eWvIABFXTyOGJy0Tk+xeEerCpj
wy4KFnlKDpWKFiVKibJXXc4w+U1RSMlzyO9pp5im7z9kyudE2SQ4HQbnFgyqB0sjwq/YSBzY2Evn
rHWl49dwTU54XfGwjMci/m3SZjbmoic8cvC/OU8sDB+aRSJdMEej+qj8cCBc3XZSeZldAUpdWP+A
LaGderLp6nG5OX7ATdHja/K+sg8NdKp0CqIE5MB/iswGQXjQKYvVl+Pw7MDsKqdwVB5oiMocdTlx
hUjLoK1T64xsXSip6JVEpNg0q/YeMsgRt4UtAJDaJ/RGHHMDqvaJyjQaj/MJ9CoTDj+Y1hMhNQDp
2BEDcKRT/5itbnQTiRcoDFSTI3bYsgJU4WeAVicqeBQrjL55zI85niPRTj8IZJT3BLc5S/eFUrSq
SmvEiv9+67ZytUB2RN6uD/ZKQYQIeF+s9J5y8xlp1GEL+7qNsw3r5GPwdeV4tPe6m0q6c/P2FR9R
Mw1tu0DjHXaQ89lAprFORJokrlIYfO4Zoeu1Xtu2zicxYr7JG3t21Bncl1ozRFEhOCJSSgN4Rgjs
BCO9KtkWk2HpHau7OGLaFSJr5GgNZFiLShoBj/V64qbDGPOO+u36UqLXiug03oHVpUCWwJ+DpqpE
8gOfiIjsUhiIwEscmakKIURgpr/F0onYhLHpbl8oef0gDLv/vqbuJVv5r22mWUFlwZipUG+ATC0y
yab7uVfjUcV8uLWRivD/Tb79IriAIR2jzM9YSPDse6SJm8/r5mcpQH46U50hStLrdduslwmTzPu5
4ZhQjFZ8T5zPhOfQRHhJoaM6jvihuH4sAuLLU9wefKVdWpJS8QeIT5CKCJ3YfNZVJHz6mckk/BYu
t5nKHzBTNi26A9wsFP16mafmrLO9s92gbHfOKJB70G25/fZYGV1wt6C3OeO1bp8IpXpMIvOmakw1
IfYzPh/IYy4q2eS+1djKl70Op/Q9iWwrffS33Q640YRuUt7ba2iBMKusTCirzbLidLIEVvbUYzho
WJ9VD6zNWBq/PUVe1Mb31mBxBVyDeRxcoqHRpxV+JbDLop/id9yY3PLG0Q/twb9uCMW3OaF9Mjyc
kmKFBV/mB4yLpSDWRT1RraDaNFobAx22d+73PP1y/Gc/TPGV2npm6YLuYfs6bnKjKS1iNK3lmWZs
P9S+JHOqakTP2KqIInhFV4rX61Ei9hcAPhZVtyegwSNKYKmhfEWZsGbQ/R0fN6SSxohYhPg5dCwz
+8lVmm2ksrPiFmxXnBXbTrafIvrsnkAwqP5lbfLq3+nTdiFebff8jM4Z5WxxtuGC6+cA0rtBObKA
bobHO3vvEMyVgayk5dvbkOHsQVQf8nKvMAASIIJKbqKke0H/ZWB+E1NFj6QwYdP0Z3tLNnRFWLho
WmPFXICLEx1rkwevU81qex30MpH1ZKkejaH9MrpP6Ka9d3RCr1K2jBeTY3UM0B5iAP6XNVNR18j8
cfqk8YHyFI0cjYRVnobVk0Gz2o9P0K0m6FIEuZyY+2MMjngvC4FWLxtYU3YMojYxcV03pMnoXR58
PgpLntF2A9wTikOInnoNHHHjxWvsZxSWE9IMLSSuMkjWbex224Z8Kj28ew+qiekvU7CFt8Aw43nc
b3t8TV9w4dUnVc0YRaOmuZuKoWG8YeVMbKzSC1JJuRQazLbCEek5B0QQ8crOCShkpQEaiLm4cf0n
uSb6sf8xu3+BlX7uLHBuY34AQTMJTRQyi7CMy38PQkSx4JJ4Tp1zvjefi3/wvq/YAn8+FJJ+LEwr
ua2/iIRfh0+mIhxE+9PqjJ7yclY8obsRtuwMCAKKcq4SBkh8YM0vSKNiz5mau6S6RfarVG0dYr08
HKLpa5SQtUjzPeWPagWIc999J8TJDYN74ffgbSAWvMhWXcZI+KHAkLiKeSzTo13l3JTZf8xnQfkq
hm5As1MerJ4zSWfPjkhDYNjtK19xNuaNKWHJV8AoENP2SHCLzH6eeRLouww0eNHxalX7kr+X+Cmw
iTnZlLqkDizMh4XQMByHjTf/bzeRmqIqNF3Y01fyymmH4fNMB6BKH0K+tAoCu4qi5CF5tONLMhNR
Dqvi4dYV3vat98UNOUnTvS59vLNgAEXGUc5b5n6KQe9U2bURvjSNgPyF7BMTy0p5oAXyIq/rJ2ZQ
Q59pE5UPdFJAupF3/27hT47VmOeYBGSl80I1JRG3gHc0F8DtBP0w/guolwyX4P5x2FqQqY52b0VT
O+pbsjRLiRKDR8qPJDDL6jR/M0iON1agLhTEYtbEBgQaZdIYCBMu7lC7a7LnijCvK9mQyIK4HVPJ
hqV6EiMszXmg752X4G1lnxkM1nr/zYvMwpP6yexdRHpx3tcII/AiYzYIwj/leueDB/+D59FKe9Rf
6Q1qr0tjtp7CoJWrRnzo7oNzdoBWK60bjZPwqYR6B8FbWepo/6gC9sIqr68bwmuxdsxZyGJ6kuvt
ft1djTjqt+fABm4nwnineq7jLRjWqMoOsxT1Y1EhgcsKX6AaF9iqSv1cw7Xp5sgtb9dJhOM4a/oL
yRlf0pwP5TFPZmH0z9dQSf4ssHY914wsvKEDCXICk4GWMfkmiTb0DUVFXV5+OjUfjtUyWnn2zBvR
gQslNZU5UnD9r6Cu0qXpZSxu/r1uOZT7y+SAwczCCAWUjnm+vQhmpozvp3M5+cLjEJUJH7NC36go
oiagmX828UA5tB/RYuSMPQZvwprltrrwghwq1OEJMlVZcFRRkht7q3a6WscA7sa/yA0c+n+wjqs/
a6XJK/jMyPxyE4k/Nj6wbbRz5ZG7KGT1qBf979nN7uY48TuXZckR16jcR4LdziRdNOwQ+5scsWt3
b50FdOGfX3wt8rHsurPOsIg9/1HUdUwJg0L2XavHUpNxL4HKAcTfPJoges7swNyIJNnHG0i4UVLS
kWsDwpPhqz24xQ6khg8QXfARRV/wWmWsNHF/sVJlK9KywH8OSYCYaFIw188UgsaFmQB0IKsUkGTY
MEqny7YdsvleDOnZkGJDhz6JHGlYKFg37tHfhYPgPPUG1c55d8QMaC4FPA8HZBpvQeA1qV43uqpo
nA/GaP9PKK7bcMYbyGgYlEjRfTOYQkEBlyu3OX89dRwvvwBxttDo/6YrhUwfk+p/mTONlxiFwPvE
B2rVDGHIeYXHZqSyE1O9hdDbu6uK7UPbRmHNDAVCS8IAD9qR1qtNLccv6QMKWhuGDjzbyXxtdZad
FBqqevQK3ppX31sXeBGi0k5KAKIOoqnV7HLJW94foAjtX2B1V1noUJyFEIaIIDvZnLb7Js1AZrUg
WAsfLVz2alkFZB507/Kex+oKV+miAOG61d4iKthaWBuTa6lmjCUxmFvTlbxVY8Wz0IrAdi+2hQOk
wnoaZq+9hLPeZe966Io9N1CW0KbTyS0/OLoiLvMLataxgHjxFE4ZmVHomVk3YTmO58Inmh4BOak+
eNkcsYGctsT1+evHfCsjzOXCWF0LDWj/MFVtT3uC5XcoVk45QnLyiVzPwDg4JrwDICG4fPzZ5nOW
vwJZ5yGyU9xr9bTfArzB/9MwRsE8kGIkgvtanaZjWQfzq1IeC6I9zkabKpDF7RTd3894JVdX2pKl
UAIe34W4/uQ3G/oLw9O5HrgCE5EmtdJtSgfAWMSiNy19nMhWKZnGJ5sSrtwfnFWRWKUxITEt9Gf8
+0Trfxci7JfInjBoX2YPhyBmpJLxP1B2SOtnSou/24R1/qBe73rZTZ6PuDYXXcBNAvcc0n72YAIY
b0i2rn+aAIA47bsNC44VMsrdjuiCAvrmi7WfpDw/+aGD61Du25IOZyfINgo+nllI9eMlJKfoer3C
c99JGyDCVIzbuB7M6bcrOYTfUGNzaj0oqp16cTIjxvJKAA/ml84WaKr8855NwnzTbPe5F7XeTWR1
+1U43OwCon3+p2F4swrT6pcsazt/ad9GYZAKEBUwWUz0k+ycq6wsG5jujlNcOyMpOmuaJRw8E8em
8T9yHc2HQlgDg/jJUlHPVx9G3pajBz0d6OjY0YRwZX2EL+xtPSD1G+D5QgPqmAvBUwREQ8b26gSq
UMe3eszIv+oenoDmroH8jbl93PYiakFooy8DCSNH8eoK/5cKtShmdPKxJwX+Xu52fNshYKwXfGaW
weqV75UNEGKEIs/G98yKI4amzSnN5XIecnkg1AaDwGC5E9xJX/bP1WLsOJjPRP16jDUubnzZwBHM
PL/Svf2BpwGWxH5hPDOX1xsUlVsJSt9oub2RjM//niAjLmVsPeTpCdrMOQNJPVaLeYmQvYBp4Dwh
6QsfBRH1XgkxKx+Tq0sPbzrst49RTMACez0s0VtDmZANcaidCdL3yEfmi+xUwsyU3NbiRMStJfBS
BuE4ys3bgxoIQs33IxCG4AHKk6HrgkI6S0Z1kBM8gPCU3aUInk3lqgXTizdG5CWtp0W7FHiNd+Pr
gEN37BRQJOKxRrd8oWHKRVecwrymr89KwMmW8niwO+3S0J6cIGmVUOypetJR+uvs705hKOgH6rUL
P0zhzVkHeaRMeU5Q29GZIzaTYMtr8Xh8/JOFykpeOSBM6UGf/JdjChzqbWP49rzjDpT0QzwAbf1/
1iBTC6AS9b0XdhvukDyndC3HZiPUyVbCcGHNxrFEwUvMkN0sjmAPrYHfKpfwrnQhzVHvekfOzbc3
FSy+DaT+CWuyeK+WEMYNuwNJqAtQ7bQxK17FvKYdBPHQbfZpXNDkE/NkWcuoaMBz8TIPLAZO32ZF
HHHV5JSByA83s6oc+mICJh+V6Xu7VkXkmYjwzOk7Aqf39LTjz/Dq5DYzksrhUAHfIRjUqjdLSO2T
46DXTUKHJOPne2hWrThg5mCIRguWCIauVRpgW46ON0MtTYkDBLhBr0SsJIFeMtEro1yTGV5Vutww
HEz4YypbweJ9eWv6uXlJg74EILElV/RZhV5Je6aeADZXGj58Xtu5bhCRkKrR2mo1Z+CMARKdhBrd
IPTrZ4lNbg9aVB+5GPaloKbNjZA7H4nllVERTUU/SSNPl9XXBJxIpoefDjhNhMMcRn7gvqaSJjZk
/cKdTSsU8zkldTcpLKGovjds+3TKZ2tT4xtOW9SMgOu4/DWzo2SHk1ZkrFuIjnBTNpeHx7YS/CAX
2sIOUrr+wfbIQEng43aQ5nkmMlQ0G4gJqRvMglCL7qFCqY5eQ5qj/YlqY4fbYxVlJMnOvD6t5khT
O2mzTbzg6baK5I7tLMFN6DMEfS5jU9ZaZZ3Qf7u2qyq3wZYx1zAb2x1o/v47VKsHiC7JJlOOsKJB
V3g5mlMLKdrFO9VQir0/VtAvfdaML13CD4Cbhbr2gdSlPNqPHaAq3LlHpfN9Z9nCqjYGz6GIIMxo
SRTeKnGPNHfDRFKIbZab/F0x8HUbhqpBGGBZegynhPkEJbHmIkTOx/2Xny4mpamqYW5huQzADS5s
7r4BHfMIvHbJZYQLMqHA604P1nymbQ5YLfUBnqrXUpoYVbeCCDOIBbH7LS0k5WdF4WYPHqA9LY8w
YjJptlxhRbMDqVPTLhiANLGdhK+jvAhTlXVJo2NcK0MIKsuTLOEcEcxuJWSl3PYk7m7+IQroKmjW
Rn0T1xMJbis3HCw3VzbqBENqdl+0/YB2XM2uJKIU80ePIWEXt5AWbsrJ1OPTuU+klTB7wTxgjNUR
2GLs4Jesm/2htyfl0Yyb3ejpAcBaM1ySVha+r2OlTeiWaSZ6MjHIhNQHBO+abMKFTji1F9T/yzEY
0+L1vZVD0YTQkPfXpAhEfiMvnO+PNIjOt0WRR0KNPFAY8U3iQCTHSMMW9EDMKshn+epYJfjm/3iu
iQisN+rEvlylqmASpMCGsXcl8KhM2NjjAG/8mG1CL5Eiu8m/tPnk6M0ldljwSWltObhe9QPwQK4H
BgcxfOjB65L5LQ36jOSmk/d/gKw/xB8f4IigIUBusB9VdbVJVOqJtMmSSaTQqMIN+xSz5wppSSFi
hm3tx5k2uriQAT9Yr0kuyDFL/gi8dhZwruP0rKdPQPYtpi2TBfME4agzper13kt2+Woyj53BBrRN
J41OBMEaUXvbrBo6XBcdulwxaxBqdR/d0BgllF+AKxfwm0O+gAhAr8etLZgM6S/JpuM0IPJ7fwXh
FCmggmSuo2RcxcOfHUYKuV+PK8CgGGKrIwPVC79W/nKA72zmdxCeSPMxG5o/u9Wb46SFOq3Qz5gH
z6a9toD+y40bfHUpkx5RqtRNyDgBdPZRDiJfj3Qd+PaErvBiYdUf59pOyvgE5xPEC0BDIJ0Y6MW8
uG/9lgPYrrauPCaTdoSUMcQk2gECkFPxtR2vk07Tr7T9cbr2Iw9rz7Yj2p8WZfONQyAjFNQOiGLp
MkjQf5e5mck290OI/achN+4tzlPgJw5ge+BFyIiRDa7Xs13/qe1Z7rGagB7bO3Lj88tbYvskg162
thJRk+9+2v0TFc4vstMfMc7jZ2DzPK6xGIqnN1UJEP8abFmz+AQ0IdlG51zB2SUCS3QPDjcjEgZk
ud15t2zNzD16sgeDw2fUmWudhT1qtlgfcsEy48kV+g0vkdrQv5nzHeGuBj63Ovt+yGdrzUnpHhSr
hfBzMuE7M8eU4B3snN3NdaxvYYCUTefaN6rQuuHyRAhOy7Bs6C2HjAwW4ohRrIMy+WdsAjUmjEem
XD/aUvtO42EcdTx2ZbwfVlW/t6glOVL4yatLf0FcasHBUwg4MPBH9s8i7O47a+GcxLRELoopbjem
ZHsn0JyAWm3Fq0HGtX6oyay2D9+HKOu3nctj4dxFK+3Bvr0jQQwtZNuHtEzBCABaPUNTn5dOZPZG
wE9Ih/fuvX8jJwKxkOlUtkb6AnFaHn+ivLMBVJWwlfo+EgCTjeFDw8fvvNNE53GcesfJlKyEMGRg
W7sKV5J7CTAkdzOjNb3JTdgd17r6DDB3nWfEUk3DwMa8QY+uKdBIrClDlMA98SpWkVTGPByfGEEn
L7EY/Xcw/ngLoZ3FhvwF5gZK6RP0R+pCkx08OUbXthKJYH/S0GSYIUv4TMVU2TAi5APbehma+hr9
kC5EJm32v0Vi684Wmht8OdAEZQgAftj/MKvMSqcCydqOysClJQDNrZUnniNeECQEKlS5z4lukhWr
5GnfOi/GOyuqrG/7NWcyumoFOTKTN1uAQaQjDsx0FuYI6+MjVo2jS4qZ7dCYvKuVekk+BkROK5ry
FijQjd8ANMWMSbTpxNrX74gpO2rURSQJTj4z0nQmyEu/mPtgisntYBA6qdynTYd9yR1sHqEw5ovy
xcRveuu2xRSrgZVoUVTjHISekNoAV/kMiDOnMbC40BzyWmCk3k1aD5USSrgJcF0is01Jb/37cCMv
jAt9hVoan7+/hG0Znphx6hl+Uf55f1Vq1hRJ9nGFx/fnsRGn6o66P2baA8NpOg4sLSTect4KULv0
gD0Sy75Urld+xc5ZmRPNtQ9lTQmXt7MNQGrJ1CVJVAfOlqLbgQsVfFJC8TnNgBKyR8rEqokJ6mux
TtrQc0CPBGK69ttfNXmgaSBVhtjsN5YRV/IBON+PjyifzPJamkR3s1j4vCf61Q2xsgJ6fLzMsQeO
nZnNmWs97cjC5PljwXB5WHnyGm4GIkRhnN/Ys9XHiHuhj9TfoFLtuy3qYP3UHsKwczlYFrQDBpT7
d6iiU/fUWKU0EA/IOWZWI/AZ2kFWIHvCfXy1sYxG12fimqduaxrfvA6qrtkyhHvv8KTc6Bbgra15
Yn0e/hgA/W48CwU3uK8bZCEAjycyjRbiXpKmvBttguUsTZ3RHcO6oH/gbX1Bj4cVirOxzxE5dvmv
T+lfMrUT6rs8LzfpdUj23rfyGHgiGOYwaUdoNum1eBdP5x9rDiKpml4B7VvZgZIgWBNiMbt+JmB/
F7S/IPMeTr/PiETwjZ0GvFafn9KqWVP3ZKXeqQ6o0Z2E0flWsue8kp6upWuttQRwexXcVCsCK7DN
mF78oSigkGYxbMIk7XCdwxOzXFr4qd+/vUWDEEnz40GDun2oelRLAarIvSjCwGSQ+GUq2NWdQRUI
2zlxoL6LrxUxhPCa1GkDL+MzX171ODXzDEggX3ekWYVbcuCOVd8nBxeApVr0W+eZLI8bcmqadHOe
nG2oPiF5WAl7bvY+fvUIqdi3aeglxoSRXPw7WybCA2n6mB4fROtcs01TaqA7xZ6gjZyBGVNg1n84
s6RQugx2cFPtZqAiD6rQaXwTMggFonENmf17xvo8Ho0G51Om1IgzxNk6E1SiQv+kvierWcpZHGhu
iAQldOZC29qk/vExhgnnL3hTEJVMMLjo564adZLqa+QagEkjWwt8UOHLWN4truJN9fLTOzz9EWnA
u3+Apdu40O/AnRcKpQUeyKISFGLudVWfiyWNwBHw+ff3nhM9gJgyrU+4DEXL3RoUTS1R9yWyUXgy
gLvoS4jmOL1tWjrJZstohqj3FXwgtII/bOu9J3TwCCc+SO41FFM/K6ZIgBozTohjsXwRHQUexc78
PuY685U2leKpDw4SRL1V89Lell38BiTVQZyNu/NQ696Uao3YeWIZSnhy8pDVhbEE0cqSO/VkoAFn
Ib0FRnl8yNYijsNnyZoYzOd0vP3FXMeewyEUpKV1IA1V0sHAPHpU7j1JdQ+YuGPhaMs4C5aTFX9f
4LdQeu8s8acL7w6IDqbvQqcDvQeCzHzBoCDGvPlolQlLh/+4+REtbDCmybMdFKwrLOAx1WIsKIAq
J+bTc1HtCFZzBTie1ugaYcUvNYOQ2AqfX9l4eQuIhxjJplQ5xG0CxCTsMjiX9mkbl0WoNsSX1+iZ
iw+r05TmlPUH0XbiWCXQ5LlqrfJteVvplIjZ26am6Z1JoyycP+4CZ1zk/lJ3/aL6Ay8DbFGXwTwN
SNI/z0Y7H8MpniF8NE1MwOHmOYkNLh11iP/VbSjgSJGEXKu8nDu0COeTj0zVhVaY4xxDcQSlWIsZ
divb4WqHLZGGvy6lF9VD75tYq5U2M2ebj4bphbZUVRPluugOf/YFPlFf0XGutSV3YmR9c7Lx+ECG
WYF8M5v9Q8xrhVQBQD+ji776mvtGMH8yV6SSEJT4YFLvLwNrGcMX5SW6gEIg/H5YcMF2rYcKT0Jl
jKuT08/jX0l1F8uIIFqH1qxFl/4u8roAP+garTN/4PFabHXrFnq8FDELpNuRoxuNSZsqUBmCG7E1
uUKYDpk5qE0s3MU8Hq+J64wpK9hhlATo/m4+wOKFPrrBmqSvdT1e8V6YHB0o8PkvweOVvqGTSpul
VeBvwu5ynf+jy3y4otrCIYwNCi1oqibg62ng6sQwS+uOLk1xtJICAlfXpRXwVA4uBeT1LgjuCkb/
5SgtAAElQJdaHV1vRwyOPncC5rfcRDaSLkMlnGKn9g6T+5yv/xDmy7sgrWVhScifpit1A161qFLO
/cqdbtnrIUp8tL5btCbuShXzRu5B6mVtk6IP9HQsx2Wbe51yMDLBKiDIgQNrCuFlVP8vDpHtb/DA
sC3VVVqbhTFVW1XGwJr/9ip4M9Irrjv+gxoxqBhtorZVwCKF94q4FPP6vj3IWboPMd3yXD/LbJ76
7ovR6BFtKFWuCrdJ7F+BMiLSJ7zsOF+LyubLY+llHtKQwmkPNZNLg4LwCHPW84XUhT37gToVwydA
davBCD3YuMOK9gA4RKreQxCUC50S45eE95i/o/riu94hOQXwN6HFQA8CXx2IkGfvKcC8E/2ImDgE
1Kz4dhgkPCxO1rZNyrfM9dKOg/UG8gr63Be5dW/WbK0qVbolifRsiiPwo5ymcYOlfhrPOZ7auARh
/TUe8lxcYBsjxNiKYhPCYImbVLZ7VVXlhYeAwkuMTL/i/+Qd3FT80xa0hauqoINAnx1f1beXfdrA
FfNnxoTz6NGsYQqGaoVibDRHpO1CcybK3/9pBxmraViDnQfQQw7SuWoU6C6unV1U1dXpcLuCagKO
4r1r56nKEn7qFCLIPeTr0J0KAbzyd+76h730+b/ippWQWia5fgE/bu/oRkyWoUL6DnXOIT88taqq
uLIX6QaKZVKAuPrtcLaXn04bBGFSeTN3w1AlDZ4YtYv4DuEYPak66PivQM42jgdUH6lyG5mt9Fcx
vAvAD1aSmBpJhGg73rvktUbKdGMtR5tvBVAHSXvx+hoUlp2E6i+2Q1ToRrjI8PyBrCIVidcI/FCr
X0ZPEu1Tm7NlbP0Fy4qk7VWYowdfzv+BCtOUng/oyLqh4obmalAlr9RWArQ//h34a95dwWHq2dT9
UoJi+kxB19Of6IxX4AUPw21fvfd8kiqEEPlJAip9QPqHwcO/wjXBHMbuXUhnIwO0xbuSI92Ve3eO
D02N6P+tBZAFFstxCmI3yXA8vVJceRph3rxBMVHGplSxsT29Fkt6Wj4jHU+S3zGdRrN6eG+HdQwF
3c6E4w9nIMpBZvN7VruGtqBeBt4LXU/DY/Tvvo0tygWZPCOK2Y1llTiEywQN5FpRoxM3Awa2n7mn
B9fvJgx6b8Wo7Tdb4TDPAIXbrgZA+0TLYZFYBzoiM2y9RnC47rTMMsdvZC47MPtsI/+K5q0CpU9F
qMzl3Yk6DlljccxRdrNQ1FC5OIvxjuvVz3BWBCN0LTH4aF7lh19eYlA47qTiqm4g4FF0MOvSrFdr
P317MZXvn7ADD182VGcj7DWBtCKOex1afpiY2GVWSX81OGP1buCMUqHZD4K63Reveu/SqxDsfDZD
biJV0aau0l96DyVau+EnGg7cbRoisAPx6O4F8Nsr1S/eZJKgQBkK5HEBDBJhipkIX/0irzQKfUrf
0IVrG4XROFpYMh8uzfxNIQNUvppHAdb2OlFOh5PtKHWGUj9eqsnI3Ke8h0JldA165pcfZnMtQiW8
/NFR+GoOeFYPjU5as5DTfv8hCMjFDTU/3xQ1n9nar5ODlqkOK11uI/+5HH70/vVgA3jYFYXCtuE8
nVW9nHXoQWVbGB+IKsa5xQh8ttQZuljqr+fRvSwBWYZvGMg9tvrqf+3YiBt79NfP0YVyB5738MzC
3cz2Q1cZ/8egJXanLKFTlhxutAbkUyhRwvL/nrDY6iD7AkS1Kk+VoPLzaWVIpUaym054udoHHZBg
S/hAD/88LwzPGnzYK1UvPQ3oTNYonL6vLHcnFYYXnA2IiWaigHhPfBosa1lBOF7yLE040hjfUU30
obR5G0pH8+njLczMhfpdeuO3ZtTuCK+f6k00cAMQ6y9m5LvDnrJOxlPkCJU+eRRi9JdmzyWPdvVf
KvvJImtR4J6P0IEEa3kp7rYCCgEc5hhOYeKCvvNmXfDnE8UcDP2xCi7tPzSIFOmVQima+Et33QBX
rL2x8rsMYu43ABPzNVlwlIMxIHkSYOP4aDTF1I6Q+mmCY+AQmUz4iqAT+NEmVGbVfDGCa54t6mzY
/BWQRSMh7Oja6aFymJgaSIOeYL1uEuEsAIWLE3tebn3V5ICgv2bh6mWAjP48RtqRKYbnRfmc8rLI
zmGhRmNqKAi5VQECg32KRxFrbC/UlAppKn7CZXiHLglLJw64gGqH2y+LIou575sG85d4IM9BvGll
+pRBLJPSeitkIbCZHO0mfXn1R+vyqzc8ix1YQnrX5EZtx5erIF7JkM55EDn82yQNjDYzP+Y4c3Jc
6+ir9pHVr48btZoBiVuljiNjuEtrukrSfsmNMz4igZ2y0AlxFzXXYgV9aWprxlXetkLUtmHLfUwg
0AkxbNPIfYoDkXNcEikFaQTCdb5OiYWhdC883ZJs1IrBPP19PhTDJJ/aHHzO5puoR9u6YPFKVpd/
vqSd8b7HyyN4rRGhd6g1f1+nbN5m6CkZLij+Sq7hfpAHcgxco5epqX97S86llj1/7QHjGL1ZVt4X
7RraSnUfmCrrOaCVJD8GaxcJDM5zKzvvqGU5NhzNpZDldLEiNttOoof3NpUiAplVOXsDulQA5VFm
JimxM+jGtRKH/KxcEtZtpa1bw8K/h8Fa728hd++ucQT5Szo6dR5pcvAvEfamgxBI4IrvpgCXdNk8
F79lEicZ9l7etCFB0//AoyTdhbHwXIzzMFYxWa5xsyqneS94Rnxlb51kz3l21Y3c90sPuYo+a5dh
txv5dL6AGMlEcArakR65a0q9MvWASMqbeZU3GJQjZ4MQMQXYqL4ezhJaikqS6cNrPamh0uFs02Ui
2hJ7VOc9UzLCLATTbS1s6pLYk31rLeX7GCv0RjzOuDkN4y0racux/q3xUIVyl/fpaNkDeQKuRW36
hbfL7a3+fKYGnjLuY/0pXwkOlfZFXRYYi6VzdGQXlCFkrjC+dqU8cOzUHvTuyWa22zM8qHmA7DgO
0z70faX699gGCEhWOdU1uurNwVU5Noqobk1qhelnXCrRdBTAd7TWmRDtLak0qfRUeIenLtETG2sv
lfLQpaxfAfL05GlS+DGBGdW2fbcELp3Wn7T6zaRzZjXUp5pd+ErzR68Hxycwf+bDP9syo93P/Qiy
2W2zXRmN58yWmWbyNxmgVOns2gvd/sWBRMsjQeN//UqATppq7si9/IjhLOVt7/0I+WCxx970uyrG
7OOl4fTyOzWWvZ5ozUFgX/Ezwx8CH57ZXCn9LB0HbGkqbZGupuEucXAxm8oEpn0By5q0UiJEcku1
6QQl8KGUAJ8h+YDzwfmopL+1cEVIrKgyvbdaUnhuxTCtgFjM7ifg3M8iq1NCB7zwuy1gwqdPiTit
NYez67FwCbBu833p0uxovq0TfreQOXDAR4D9d+0gDgv6YZrd1ddm1+c3kBy670xMCOs6v4XArz7q
pKtPtTqLbHg59TtMVGms6Rx0GjyT//8fZ7WIli3j7DimFWcxSoKKNj6hg8rCShwbXOoxgHue5NXh
wKvOgXUy6PuiXhRGk/HE8Zp7WFJfB98lnbCajEphStYzhXB3MlWqLas2lsQWylPX19/g0diPXaUg
CYeDa/DDwWzYYTFloGPM8L/nlVKmxcgsQVxutBAfn+G2rLq/mlZ6ftEEBwJFeRKjhunL1FumrCGv
yDbDImZExIIX2Q295gliftI8f01PP6uGNCiC/xLZQmjhyH4FDEjpeY9IO/xBx/EXnk+vRby6i7TH
pqlXmtyhT8wC2StAcQjpOqTa1sQf37jrhwQxhS6beISylOdFghZ9s3bbU61G8kIpcsTaLl4qo6AO
auVhIer0a+rSJjCCNM5GfcxXsnB142rSNGnSgZPR1j4pisE6gl+qs2d0F8iXJXA8mCu16vRPxMYp
aE9yLjruVyyRwZTqSp0nsITPp5WAMKN0URB3KH/LQk1/vf7RfV8B34arqXlXFTEit8TRYtHGA8/n
3TFbOOKvRoDjZdkAq/4wAj8hI1pq3rgqDLqwlC5Q5G74W2HvH3gl2GOpk8bqJCj9unPH44YOVapv
DgbsGAWf6uakEm7JRHsa6ekGzCXNNhhjJSwQQ5TXfatwo/WP1/9Jex3/3CaZpVVJEzm/vx07Gizu
Esesh6Co8ZTZy5Rv8poGgK6K8AtUPexFoV4XJ4cNc7/S2mQw7sPOwGjjOoEfmil4yq/bEcNxPQFN
JL0kdnKQrHqQuFieWRSlkHCBbo6zqKMY0KZJvXfGd3qxJVc7k/GyhZCSMna4xYYZf3TEawOR85EL
/2lOjijJUJPt2weWN93A5uHzY1/HT/gJg7eUMcSvgn3NwTX3Q6e3GJbBBIVB0WeDV2DSr6VWTNjE
h9C6tVoOrPCCXcvqq1uvl0WKjjDF6GelSuZX20yuKRUbdvzr3DMQp655vNXaGoZTtv0jXEulD8gn
xDetYkOY8CumtHjvMRGrE/FfPGih3Vc/SZAsC1j8VOJC1mDkcUiYuH+6V24qs76MYf3AJXtMyk5R
r6WUjM/J54afMxfHW8CSDYkbA+AzyvNUSpXdfHsqPe9EFvaWPFKKE/SykTnXHvawT332CkgEpoLh
NoHdIl5GlgrFZeAqJd9gvQDCPXZuWaC1MdWzVCTJ2MZkAYde2J5cN4NwZl5JNHpkw7djya9pXtKz
0UArnsqAAgZQrg2WbatindCYCrBKs9BnVq398gzymYC34ZcHrqCzHugA2ECsGo4EamTqUYXSN3cu
hQ1Y1wE88NsTpn4Y66cLchZqztRMpcjCF2mxddiqkxO0eJHbH3o0dQ3g3OWm3ASwEIB7Xw1xjrBR
3OOHIaweE/4PjoXgNBfJ/ixGXQAqAYz1epmWuUV/GK8fRbBFedBhcEbNph2dUH/EaNI3yXn2onwo
TXi0yFONvioULNo8khxVtNlsz1vxbEYLBsjihp0QA4Q1GHLqIGzOn5pluYUo9jwcYL20zHqeuekt
6q9rzNXFtsyBu5Qm2AHiODfUNvYArOmUV0BlioGJ6K8ds/mVn/ar+U1sFMGzgShyEP7tLNI6oMnB
AtvW8+BOLIEObqy4PH2lxgjragrA3DxAKZ+j3W6gyBzVzhln8EvvEBeoc2ujB6K3vqZdhUwi7LB2
LJb3BtEgQuoabDQW3ULPJv8ZfPzbyNaMuZwHznuNV2hMHo6+HVtbZX8LcW0r0Ai3XWWFeP10N0C2
hp+B8kQcSHHl/xIcmCN/PLCf99aldN1P1pUeL5GLCGZ4BiSRl931Ar2Yl5L+jpLv48BoquZKb+KG
QnFnNDsvGyA53JJUz9YUwIR5aaosFG9WWx9VL3tmko7WiOiqViXZ3AYqdrnaYVilVvB1jW/oRJkW
8B355PTaIntwBcpHp1ngUjeMGX1jbHMt7LbIfR2NdBzVH+VNP6AGQt1gEyajm5z6Cl3IA3cI41uD
RVno5XRM8cS9+33ComTuGfWxE2aTXJ97UM0evW3hmoWaCiOeQHIYmkgjk7jF1AJGjsoyGytwsHEL
R9aCZ72vK+M3UZT2tg+knxZLKPvUoGLKuaNJBJUXyxNxv9okAi9I54v1atodYCsCVL6C7O7DwGVZ
kUlvInU+dce8YQ26GJEPITejhXMoU92+GuhT+3AOam+X8xONoIGB23+2ytj/94VLknleWioLg+3q
RiAwDQrF5b6zOIWMROtTv0zxzVxrhdYzjhWje7QkH1GM/BaPUCjyAKTyCzNntyzLLn+bvaxeS2lt
2GA8IKInjsM+VRsNeBqNxRneeaeto2RuM8LaFbLCTPKBnZdoFYtpHSucJGzJGbBaUL1USC53Qhkz
JWUAVjIQkv7jkGBw7AmH6V/1zmpRYCRhcPQsrARvYwWkd+uC+XVq4Bdpx15rFEzfCpcsrlywklWj
DzdkJEJG4ph8eWIVopyBMDrbqJRO8+m+K3QvoxfOhq3XmCxLXrea2nSBiqVCXYkwWr2wO9VAeaV1
XuLCFBM80tDyW/SR1RusBe/8N+rSNHKtpx5caWj6BNlauz1eAzTrs+RNuhFFuQ5kyiMhT5gkQiws
vSWM6y3jelAtrYmbxFpgp/N4SgiW8JDRRlypb9zZ9IxBHl0evxXNq1IfFoKdUbzo4eE1OAMKD0/a
YOEKju/LR+L/M+41lNR5DO3cO/BlWxr60aePsaIf0oxjGJSzQvgYN6RcbXZEbkHnXY5RVtL+goAD
cFR4gTrZyAeyHtLNGysZgnBBhrwq7Ef21aKswarAeYkDHYJxqXMeLgIHeCMA2C2cXOaYg9uzcS5Q
znlJZk5hjaVICXDtNffdx59eVFFHdCEP+zZbQCAHJZpjHvy+T/vQGm/LfEFuv9uIsQic8HPRsqIg
9V0EyQ0vY79DiGw+R8NgW03jra7QHphGKWjKj6rZI/XAd3FxrZaCvyjn9T8234/lG+0KRyg3xmdR
3fCIonZwXZ92WOUwbWlyBkHsxDl3NzcdB5sk7SuoHdiOzMO/jYLOzmARxrZ61MBIvbnQ36V8rUFn
pg9NKWL7fJ0Ul8Ardq5gvacaiFuTouqegCweSVZKW2S9wYwEYzq90UEQzzacMnQgCkb2G06i6DhB
M7gUdcsJyqCbLuPlQgwAoCXpsXNuIp0EQV4EAbisYW+YjjUKVct0eULVvwENSqchcdnLhePWWc71
XrEAgD8H9Uqs4BDkkBE2CYPiZ/aT45vBMXAJG0B7kBKQuGtKZomeaLz/voQWzmR3HcjRUR7BA8sa
GWPcb9k/06PkUWleMN9Q3uD09wHy9MjVFgadrUfqePQLt4YJ3Hlxuti9fA9PZ5W13WHxjipo+1gS
ShNtImRWSjtQEP/DbZmj/7V+zs/cKlKJOQnQzoNsZ1IA2/cw+tRvBHcwZ+TbU9CLlVB85ESNTmrb
QLqr2U496/EOLAZ9frEdzK/3DeSdiYIKkGWZ8kWrnAhH9QHHHUZCYYZBVblfcSkBQ5KVhTFWVpGH
sF0fp29gt43qe7yCQ49ikw2a8h+q5BRAXzstd02vJqt2Bw+jR5MWlGKPbPscBbQiYxzLqYBf56Zx
WtQDRRCKiRDRVgX4SfzvOnUJegWCdI2dXFhXty00ndQ4pHydCAkA5X1gHZKIMzhRd6rOLNCWeHwK
DEJycVAjrcTRnRPA3pfa1wAWeg8T++aU4X2ZZIo0DkfDlp+nwAfdN1PhhNpV3DZPr9YSnhbuBtCy
Oyn9kiRZJqpO2UcZQJwbYyugcn00jS92JT9g7puR9r1ymnvrhZ21hYT7LjlJdUAgzzwcG2JQ+eLU
RbfVrcrVDpcxuydrOEB9cvStA/JKMDXHN2wZi7GQH/epKnLQdNH44NNk96jEXLr+zNwo9ZmAvKwc
veL4lfjboY3BUj5snYPjjeKHJzDLFYZMQ6koEI4nSdCS+ITQ0TmS1DhH3uwO8/pVHsaY9LYgdw75
UeLBctEiSSn2m+rdDj8A6ESZuB7/2WYUyKKljZkjNnrzrOGNjfNwRqFAYwmXN+sk2UgYKrL2tQzM
INR+AvotZL/Qw1xcS5RZisOpOWj0NFAYfXeMmG+zk/DdurlJ6hpD9ogb1R7EBIdb0ckJ4Moh0BWz
hKROs1QcIFvzhicti2TG8nl+OMNv4Vvfeay84NDJjFw346vdppWGsZu7EBfKIoIa1zhMzE2auGf7
P8x8OJxoX529Jzesfr4xPIJXk+okWkjHipYQQIyq4gm+J5vdazV7NwUHRadglXRB7VX06Nv9efpM
u294R3x8052kO7oXnq7wSylEowaiP3IPPttVLNL1Qhx1dLZOIICJqEAfQ0W1Mmeshj7akf81huho
TiJZiwK0UhaAaD86mw7SyLwzXkjdAZYtNyQqcIWtYusgQaG5CfQetLhIj72xjkgwC723GvEG9vcF
OxonFI+gSpwc9lQdS0h/T7CZvMy6bV63def+6fzY0kBRiSZjqJz/hcLiDMkv8BcTUXgmf9BZjQug
VOTrFLMF/ZCBsaM65GolPaL6Jwu6IVB7HP3W5bZslILJYs9xVWt9lZk6bYeg9M2ADwo72t5noKft
x5OVS3QlWHJBe5Jynmc4IKQ/uRqOKOIFnZGqkN04SWQcTD2lAqJjP/Jk82otrc2FYTB1vdojSJlX
Lr894/Y/+XBC+jqmszLU1mydRlvZVHD8Y0yqlp0WlhVIoIUG3OlCFmDUR/uiJjijzbyjKO7N5Skj
RUaTjUfsWh1cJD5ltCRk04X7WgqdRA0R2u2XWf2H0tO6IqEJowwrVfY67hGaus3xP4hsdbSOxJxB
ryJDryn/vfp5c8oyQWRxRZy0u0V/9nA6/b6q/mR+lhmeUdwZlD0oLQgJdoATD48DDkjPVtCyMe3E
NOzyKd7dIMDGhSk6YYkT7aipaf3ctvvzB4LI07HWsHkoH39S2e9+caeJBtHgRwc2WeXe176yjs/M
xEEVbCJkmwv6RKebX/cj9QuqRYmNqtaCwl6riuhrIxgMlaWh/8UyUfeThQKTV5kW+LBxqREnNrJu
gLaiqWzyJeZIrR6BtiJvCGAYwPTfRk5KyFAZT3e25DJaQ1GoHdSB9MTwJR5vgXrLaqJDj/wTvLc9
En1VH+0Htz2sFQMr5EZS0IOlf5k7rO4Y7g0bAf1mwu5souBUNeEcAURqhq9jAuyat3lZQn9hiopO
SdsChTdwQYzwHORG7nDtFye7vDbtKPQhgb7rY0wF9wW5KfugYUPmBn9z4GEwGTGYy9sjNTfJ/M26
TftVX4c+rEOD2/ljxfBdmodOvUREdvjUnuuayVxwZ5gOFUpCroQOwFOhNAv2rfXrakjKZi4c4sS8
Hk+9MKT8qLLmoM7h8QVdghTfR746NaGHMApqUWa3dgJuXaHbaffT/+WW32btn4Yl0t7bgd/SyeF0
kEz0cwQMJiuZdXF5M+I/TCRAmKvwBxSPITwH8N6Wm/dLVUE2Ay87sDywHXI/Opaqyk8c150rcbjN
dDP4vvOtv77DayHBdVPO/QVy6V9NxDDaosQOHXiDzbqDpr/joQCSmBUjuOTyjQVy3feDLiM7O2CK
5as5p7FM7y1jJKySEZ4Rk3Dv3c6v0+VurwvgnMEAzRog/zLMAlbGI4hWC0FJAC+yoPvrp+NwwD7i
NJNTZzjeOCVZvH8FGA/nTXxeJ8yrkGBflMroyiZZuYVfqTgPG6hZFY4mwxK+m2tJVXz2lJwgFLoj
BpLslA+I8E7CDRCUR990TbDuOH4D2WFQuTk0LrbXK7tKG9yxO3ZQ57+YzxGucX6lForxoQ+5nl5F
n8SuHQDL+9bD1ZRuYN761xu+C7EhWhcnEVazbyn0XUrydQxIK+wcewrhXjt/dG2iRTrdnQ98o2ls
4E/KFRtTxlS02jBHBGs927W2yULeB2wvNWVay1ht2RqkSJv5dIiBfLgf1yZEKXl/500QTGTc/Bab
WYIg/SH14Ax62bHv9fbUO8avsyW/zt2nkKHeOeHUPBFIYL3uWikSKe3T11eIYA0L4DfQAM9p3yC1
8TvIxcAvfvMlj3oAx5A+LppWcoiTqF4rwQD8DOJ3Foa7wXZdWpyiOy4HxI4MvMxn7EfeKbTTkT+c
zmcQ1AkUUj74MZ46rABEbl+x4Bujlhn2OiMPt89xgrqyLmwT+xzx87DIYIJwzkxjmIs6rH1hKW/+
iwAq856yegnDUCvrvb6qARu7ICaZD2qEwrvaJ+ngzcZBLbmIDcYjW73otoTxJN9zK1y5jhLFAcpV
9wxX6NyEDrWqHI0WeKsSghxAgfDfKbldW+tnGlXYZ191x9KLRpAaRuJBrvY5+B6EiceTk/zEXiEw
1lwYJrGH94STUOScA/yaGFmtUK/EftyXrTcY3+oOt9d8V9FUXWsLgfElkxWknN4dO6FmJQwNMoA4
iLNiTiyongud1+AFhirbux037lXxNrFYaHFgkUW3dUn0p5ClODxIv/cbmX5B/dIWtFnwx+inBR1E
W7PMxlL9JlYw0MALtTG1GXU/4wODozdJKvoIretgAc8giJbvOJR17X3CAHjtjLcaTj2vhi9S7qVb
10MlYKzNryKU4s9hvNbnIBP4uQy2koJFOqaPvdzVm0R74r8vsakcaYjc7mIxyHebkdHwCrjzCaSU
l/7DWnG1n0DoXCcaZfRz+p2Aq1L4wsCFGrSb56+s8C1rAXDCcSzdFPLstjUhywVerfYpyaOjCFwy
W5FfXoFsXH9Wso4rLzv0CW7hj5mIBxT0Jowd7nvqBPjUa+zICV1hk2r//cgaE/3hf15fQkOpzJb/
KaqlOlX6r4pA+UK3EMqXXNcT2poNFnfbIh70EyEYs7ivO87qa6XRizwdNon9dn/clIEpuXVvSVKS
q1E9ukhTmwDXL+edOYXkMWyc4dkBikPcjPMItRtQ0vIqPP055cNzAQkMbWnc5lOmqQb3R9kqSq6t
7kZbVRZKuitOMipHxFb+eony/xDvjPMOvNfLrHIl4lEsltnHUlz8ZokxZHcw9c53LQdZ/e0zTJFQ
ATADfulLcj1gFrI2vmXd3Pz0wLga8MwqoJsAwXYsNnE+HmVMuGtwYa4JQryBBuksTvCxvB8/sTdk
4LJypgmWE9k/51Po1ZRgudUUAApztnbByPssUhSSKbh0+gCJHJoW43k7L5cI5JwTdNiKLRyUOS86
bdiDk8lOpEO/mhj0mop5yonEOrpfoZgNfebSkWDh53g/DGGVSYh0ISK2aFkbI536ImOL39vFsobQ
99rSOjUr29TDuENGC+gLoJGd4beCPKsaRIRIbACP4HbeQKaE0y7zwJZnPmD5GACgq3khd1gc7AFh
rczZqPgV1V63WJ10wYWSowrYwl4JORkuXX+9VYzvYBL0f2+L1OtF9SNw/r5dstC0F7rDS/87Q1PO
CF6VzLZWWZYhGu5UhZEWqaE2uVZdahUeh2225QGqEMxiz682BxajuWOVv0yC1EzlpM6MPyaMdntG
o9HygRU0IVprxGNqFtMA9byoVKp7yIfFl6D+PJ5IuFM3AzAwpd3VU567h0gJz8JNGSMADCcTaj+O
DBIGUUEhuVOg98v3kpL2/5Os4wOfW8Te2FPxpAWa5H2/ZOPY0v4XLdUPk3Se4lWsDlOx1OLnKYZ0
YT3EtG14klsAGtrgiFYeOK+gPru+I1TsAyATcs0of+WyyFmDr7YYingsYRP3Mkhk5mz2mhXt/qiZ
+N6z7FD9oAhafMfghjET5uRTurJCFTIPrk0zYdPEjLJb7HfZoJVYwXiuGxzfxLty0qIZBekWhSnj
yufERc5BQ90pOB1CJAaO9HBWML2tzkSWZa2NU2l1DIOHEijYe4yVDN3RlIOX+P3RycsJqakV7uFt
YHQl4gms4mR5J30KEor+ZRgSGr0D+BoYzjtEyiq6qg//sk34vZufvYquIkihbwkjEMmvNHDAf+tr
pZSZnaTZH4xUdyTOCtHr/LDDJk9l1VrcwWy0RMULFzcY4fTto1q+o79X8103+bxjxWlrjIjAPQDt
LF6b4m0YRqVltbIppVyLA/g2gxlnChgH4Tsn4VsHwpLGnUQFrBDkPUJp1hNXRKX7tIvvU++6eebA
9EbDYIhSqBX4dOlPMZZIek9XMPGn2LkhTYGjRowPBZxoiyYDpvW5vL84vWPhvh5H0cKcdEadulct
ZDvRAwI1y4hXWSPayvN+msNxBvOyIuVt+s9vdU0FYTVg+Dh0/aO4k3RJhMnH4T26RczOqeGbN0Mz
cmztj9+exnuqCXwAAwQKXZRhU+atrBaWuR0Gsw8tys4LZM2b20hQ+YKUR4nABWgdKUU0Ao1JXaOl
H4OMR2vsNOBc/5W4sPUKPXmPcmMP1RhnJCkyUQ0Z5Xe97AhCU8AovMBZXkb+icTLnYLcWpseWskT
Ca+mHjFdLg/DCZKwDK0tBhNI22v7D4HeC/qTlI9T1x3WebOaXllynfuBz/1btxNVPq5CM1YBLVov
eLPhCR/AESjCC+eWdqvzlrS0AQiz1NJifT9rfMYuOAyoRGQShziuom9XnaarJ4npgHSlhBJpDbCA
x6L7LJtIsmisJQr1LLAorkS4r/0v93BMlD15VN4OyIDyaiTCTSU/HXERIPDYozVIRUTZeNofpEYs
yLNgGmxLzxReMP8HMPTUyB+Wjd4PPECMuPTZxSCqa1iIkOx5MHjuw4unZ8Fcyma2SrG1h4PmuE49
R1lvLHQjDqyrf4PilHS0qVM4Y+5LaqyxJgrOsagQvG6dAQmsRwpg1FLYQCnvY7djO1Cp7uCmeK95
xzLRdS9RN0fT2jn8jt47WNxOWt4kdlH3S08wadyjy5zJWVbBgrdFhyCVKA73UvMqlwT8Mj6YB4jk
wrYsJcNKwip1Q1aCMWxAK6hIkLS1ia20sdrLSDn7uAQMJ3nOhYhYvGZM6Rhuech2EEdohBmdNvjP
do7y/hzU6/wcfdJKQ84GAmIR76Iylre6tsYJM50A97XR/Kv6aeSrluSU250lhs2zoUCREQzTSn+1
iZ8PEC2UcMQffIJ/lPWMo8Ff1FNtrMg2aL58hWO9OfTO5gOF4l2e8olLmWNx+DCgtQhXwSwTyA5+
TJOLNOtEe/a6q/aZy6iID062BvIv7WxtnSCVnuXuPZm2dFq8ApiZCU1z8cpdh6T+gl/dZwmh56TH
jYlOJbZ9ERxwaiEUOIX7BRcfHNOxQAUtmMnpzv/FiEy1IniWiYOzFsOfHXe92EnmsSPRJwcWRW2W
riKoeOE3bFfbW4JKiss5IzZa3VjBXAjsBj0FPTwvTCQ7T7mAjEBdT9tlyYCrJkBATQ5Dh2bbvNcZ
qUz50NeYJuQEFdwGaMhxHZJLmczWmNs02cNg4HhFPhl5iYThmHqRhXGpAurzr+2/M52MvLpGkDUy
o3kRdoMxroIZFvgGrq/nrRqz2Mb/XOfuAfU8KgLNmPr908agiWZNkEAr759VexaQdv5JZ0zLgRUb
rCuI2FYi2NFChPNI4ub1H/4O2KVneW5Lq3fIVtoLckI3hCaEvXpscwsp6MlIRHvZj8SXBE3Y2BUC
RlESEbcY6qUJbdQlqXPA09iDQVqtKJuHvUAT10NVQVGKL5SEXy7Cr3xjVEteN97AvyLQdC+ivilT
xUCnN0Z1NbFJTmOd9MfkYNq2nP0x49s8h5X7hn34jOESYsYjIg9nrQBU6CFthkLvY5xTnT4yTPgz
+vimJam2FGJS2iPyHPIlfZQ2EAvbjx9ocETcYfSx1kegJ206Yy+5ijwm5WJ0YFU6Hv7VHkVaj2fA
mI1J5FkrM0jyYuOyyn+F9Lu+3u8Jz8qmzxfDrXnMKsOHuHdEdFEBxAVH+GksZj8XbbwI/KOQ1/9C
WQWF3Z6dg/m6VR2O1dstf6jq0WI8VebGPkJ+BWXRPijoXSU8VEVpFzIHtr4bWLB6KaRZ7tGj5NBv
glUTc6JS6IezpAzMuyrmmZMPKPlbhRlpu4HFIOff34EAHDKorUKEIMaZ4YR6Xj2uLIVXN5Yyh2ax
0OJ4P9IlfW8ig+v4ilxhaXgSXibXvUAfccurVS0eoFT+IJKCrzZNYh5Vq4IAYs4ZOz8cHt5gIYdH
Lq+Ea5zQtd3ucY+//K6kAutapX9XKGwO56Skt04zFePDw+GvxPeqa6QFFsGaR1NHhUqZ7iS3Bk/+
t56sCa+U6rjgiqB5htCir8qNduhxhcyw2nArwLKKfWa6z+L9CFqOzwSxAKOWQdRV4u2Q35NboCEb
2sryQgDGmOKLwjJrx4KcLxUUaDwmtEUetYRQPfTK/yGoQbFQny3au2Zpee85+OJgdSpsCRfzjyzG
yTWI8ZUHFRsPJNa8V1sPGYXYH/fCDEIGdI/tnJgYzSHw1QTGrGjPhLsO/UUihX8aHg+HLbbfYjLg
MiT2fbfl3gDxoc33zf+kHyiIygeIo7eW0WfmxsCCCuLpX4Oy6jPuVKdC6AQS6RDfOdH9z3W2ghG6
ricgtkn7y3SjD3pPXSFF7LaCB9hg5wU0y5dGWr4c1JBdQc+458dpYtGqp/D0tJTERt6ujJR22HpI
1PHgKLbgNthv8lCML4rmJlgLxmtX8rwpr5+k+LCdqLc/a/EYz/OnJRCxbo9zd/gDBaKoqINTz0a4
PHZhusi0xRZ6X6evApP7gZ2H0ISNdJZlxAiJpXQCW/R/wy6n71VOIR+aq+reGYSI2IAg1pabmxPy
pdBh/TwWkKsHvcJoGrcARxXh0QYGvAmDkwfitSTsh0BSRXG5o2dbNZKj5fABQoWh9CD+U0zHquH5
SqeMlqtvR+HnBTdQwpc1LgxKDrCCAZNI+oGyWSD45lyVy5PEiZZyIWsYm52aRoF+/rcTNrcHjR6v
0VN3hChu4lQ0yU07S2HMNudDvL/n0iqHpiDZx1M17aO2e6gnmFKMIn+cC0BMIK1McFGVBtgLJCAm
Y2OaY6/+1NK/8BeNwHFSq+/3lUNQlWCs5pIa+QtzNIpmAKKq7kNJ9DQSwOSn9+OH/8gkgal3H92G
xCQXchXl1+vwYTwjnWvkKt/7XkBrxTMPorSyg5z7lFdZbt4ei2AOTO9vYOn3VOy3IL7lJH8jRJJC
naCpNNmRlFj9IRUAnIeqTuQl8ox740Hr1OBnQPHomkkHapSJzhqvvMmzObE4u40JQYi9GH6zZgVP
XF+zH0VtMG7Jz2VeNNyIIrxBPbIEWi+32jwEP24j4GGQNC8hiTD68uC+XgD/YquqhpNHY2WoLsJe
pKN9qWiuuB2gvvv3ee6CkQPQMOEBgnqHWW6zrKtcz0K6G6i9hb7z9LoeGpwN1VULN672TFyo7653
qKxAYk2L4XnYGJ/d2/f0ejQ+wFAMbnxutuj2TBRskXGf/PaK3bp+L5vaEmrEDnRqHJnLD9Jh2FBp
nJ1fdZqHW7NO/AEmHPidvWShHiz6LEXP9WQbHkzbINjB8kI+g0T5X9WjkXfDtunqleVIxrRICrV2
+NTEu/nDV+NnDYuqsSBhzE302sCgoqLF8S7FR1HKfSBGJ24k0hkKVlBPe/FaxNYcUvjd63F8lUy2
qCx2hwqva5TfX0LI1szYWbf/LKDpPTkm7+M5+aLjWGhr+MXTxHrIxXSxLFv9FqpKzCxXBexx7dDP
pEV0zoy68HM0CpvBSjj705ovheIq2Xzfjn3FoQYVTnl5O6eMOmXiUQKBDjE1pzMsnYbLaGGcMtBV
pwbIRH/2uLRs2CAss2jBi6A6fBhyNTOkLZEKK0WB5rx7NfdK5GN50gBWSgZGekAzTO3m0tDaMpoq
Am/++izinLYf17Q//dL7RkFsLEkSodtLresQoppiG8QmnWbq011nn5K0DlNNVDtaMiltfOXlQclE
fewYMZp0NMZcz9xvUl5ASsd2HI6glONRvrtRB3nQ4Vl5o3A60uI6br58Y41orhCiS43BUy2j5pmd
8pg2wCul6ay1w2TtNgfD6gCL51NgOAouixnl3uYS2Gl9aju6LNuEphB4Z5iGZtFneznCfrWGx6pJ
LFamcKK29IWpInSXk19GPSCgBv+GDMEUs795dlRUCj0Ol6XBJUCR0DPlK13CA86mNu6ZlVzO/P9C
cP+0rs+KEya2hV/GBqXqJM056VK1G7CMX+Q4SbeypdtD2OErce2XTwaVXdid8KA7DOKjYmaZ1SXq
Ge3FAdnRjO4cNrZfQWC6QqSk4QVCFmqQMun+t/smYCQn1OROEnii4kJn6psrXoJ29M3KBok18zic
N62+yWHz5yQPQD2kqt9g0ErwpOey9nsc8P6NI28/Qnzo0Pw6ykBZsWZGWQS1RA4Cb4IlrjZjX5PG
iogvHBY1lZfLiLFkXShoGjR0ZM2RaWncWmyiK71AfQ8wPDWR/XwOkE6YAdg/YEVMQRp4lD1AUSZ9
GF7wd7HSIwUXUZ6gXbyIIN+6aIrW/5AV09AEd6D7PkSbp6jlIvWVUZEhryiJ5yZtszj0lZBeNPS4
h0HucgZ6zVbrEiyY8wC0w58jbkeM3iNjmUQkKAyVhUxw/QP1CPJ1lbr8siqRLkmWgcc/BBglEpzz
CICt3Kw7GmS971HT8LAumcyLvLoKWhTl2DFYlMFc74+AwDJXUyYSszsp+jiS18lHHXSE1Ut//OIP
j51TQ9LRv1tgEqNFq9NwTiPqnDJgqKRF/uWsmVSHqtlKYlux0hyl5P2CbD9arRJrrhI7JGEUc349
kqf6FeAKiN6UOzA9Cc9z2nroAT15B83PGgOadRsjpUfOUWK897Se44uwP17+JDl0slgU7rmfKunT
3CvDrkNWE2F88rhttLVEhA2DyHj5zw3TsPJFB/jBnirAUucl13qaJrCzqdVarEuGPX0pu9IMJ3fN
xT0ltOCEkmQkTif9Nqcqzpsi3zCEe99kyuDaeu3tn60uU+Jb4BOgcr0Le93Vn83oPvza3U4i8RTG
g/CutPm0FZmoSuBiQFfesGM+jRALS7lqYZ5tCKTQ+JapGClqehpz49wnRPepOIunHwg4uRG4a9dn
hVebUSYBjaBt/MgfDZoCybZljFWP+N4o41GQ/EQOJnsudiaSZGHo3LB7q1MIZ1l5Sj/ojrxVJAzx
AzVfapYOjtpP63E5J6VBBFXG95r1QBhp14v44T+euHPL98LU0XmbZzti1VX4n9JNippzzTc7LkPq
8an5YnOl+gdJfC+r5g12T4yO7LGxK3g5SCmD7llOjjQj+KVRgQvNC3oNFEFXg02uf0xnD5xSv1NL
dANtj/kvZUy+6fSdFIz3h++iR77uRTrVjGpNYXJYXTem5MgejW1q2rDDdwzg99gLbZacEGwkiVUY
zxmVLPuQhy6IpP0XkrlmmSXcPcGiS97O8oq4RiPvxx2Wu7jV9fxs5zg2a7KtjA0L+SJmFpoTLd7n
Q5qisvppftAF5fMc8fcpnkQ4Yc4gSRnw4HBCoEC6kr28uBYCOgiLDNucg408owKa5BBjrQsMFwnG
rP72JdNN7Ps4WJpqvmivcd+rdSvfaBd0cnlAeTonvxTDRXcKM7UdUd53Q/eoKdIWOofJCgfsigiu
W0qLXi1mTgjE6IPHkqZjbby5+uo9ekLeJHofifUIsVwO569C7tsD70qFRmG46MoJxkj1FaLsyqL9
3gJiINjlWF94ViL1f6tpMk7ipLtpw1+Zm3T6rE9BHkosrBFNTyO5OeV/6ep1ZJoIXUMOSExvWnZW
q6Nex11gcTel5W1HMLWfQf7kENc+K+sHHnfrJKZink1n47+A6XsmvscVdSpG+VIN8XZXRrV3PxAP
8AiV9HK1FocWTvG9dg0NkQAYMiqfhM1sSOdI7SiVsJNAx3+npCv+S66ERH96iWfVf3Q9eYiCbWKr
mukVSI0FhsONQ1VT/btYnmRzR+b4hxnnXs3rt5XAMOtzut0nAq5q72PnMe3Qit7YOP3L84fHB6z/
8syQQOWW4ypepLa+qvhcYD/DdljFfq9rmNGYgrtGeQm2JJpx0+/wI4OUN6KmoY6iSZulZKIWp39A
k+SV0Nq1v/PnrsBn0kUDEtEG5wAqGfBiX3TukUFdTSD5xZJe9XZgBW/jFIh5HynDsZADGkVYNjbO
ACtkMyeCgyOvY6sxlzjjeEyHEpChSGLiXtSwJCbpLWTQRBEPsoFoZlTL7sSq4LYdXl4TxObbDyvE
at5ck/ET5ijhmqcD1W6Hq3y8dMRALqIr4sO3tqfbrJ20cnrcDEe8BJgis1OZh4Eel50sgp9GacJB
LNcN8UpwDS083pKbtLtJ9scvWmFEV7BrmxFlN4JhihdLvt3J7GMNajOUFUKQEqb3qeeJbJRuB1f2
Vahu91MV5Ll+4XU+enCz0n+UFDnVTvf5MfxvoogKCBFF/kp2pSjBaQHnXmeGprZqHIgt2ujaNlJx
OLB2MINWkgcKtyFvBuXvKflhZgJI/BYR8R9KvinR/z8mGWSBHpnpnRJdWLkH35t/TIGNB9alDT4F
JzrJ++HrizwOLbI1RcnSC3vvHRmXjKtrobAPJ9c2jlgvMwHE8WtakSG9fFWz6g7dZanikZAiedGk
vrTQoAeJS9BZNRwF1GzjOv6753saCmQHh3XxMDVCVsAqm2e5NMLZACK0j+JvnRFHib26+OrJ/07B
VrGjkd5Sk/fNV9kFLxD3Hz6fmkBKjqr1hRIhouA2ha//v36fMcT437cqaTpJooWD4k+k2tD8xZz0
/6JGjb0olxzvd+JMwK3idTxcutLCBMlDoqW0N3xQY2/c3LOyl0YhdlrbwAO47z4OU1DWzWy1L7sB
9fgvP94PfrFOzyfZqi0He/6UbTTbd3gPtGUdZ0HpGywfY7XyYJXbrBBlDx4Ae/ckVcTddKMEiQA4
PgmIvoF4c9fmGLgnF0tPLlkoqHQsR93pu7qrkeCxSCmvlBpvOpNgMQaK4uBjdb819s0V194CvIEB
mMIpkdeyvJyTEGsPGrxXW044lzFOD3hSSJ0TCt6g6RmOYWbYBDqJHarpmcXvrp5k1BWA9eoLT5dZ
sAcoF20eKpzDTE4g3+cAXF+/US9DSp52c53jj/IboMIoGydC1wz9qx4xV5NwPnSu6FxmTxxs3XGN
RAHveSwarjkc3UfvxnCvKnhd4I89EApzGN0gVg+3DFxuFisHQa77d15sG5h8vl4DUHxs10k4W3yp
XDuh7isMX66sIvjHfvfRcSIK0Q/M1uoiJaAezlI/B+wPuYEBvfasMrIgkQpY0MydGCYRpnt6BB6V
rWkVCgY7BrkxrfXsm2CIQlvyy2POdyuBEoUXOVXudStvMYfat5EWQrP0VebBypJB10vZU31qYVlW
aXEFjZDe53xUz7f+AGxGN8aPMkOs59Gpq9pLJiK9DOlUztQiNAhbou17oTyZuqVYMvCt5dV/pDix
s1pNtIKCHg+UTwGdWhoAwkgxhh710eL1TmLXJzLsFiKEbH1KQxyfspIuJVujXa+rx0yupgyDvy8s
mZEmhha0Brk465Gwbv+JkfG8dKokrEmYJGhH4L9wavrf3xjLQBvY8EXqDqJZaSeU1F0cAvpe54YF
SUFdvnL80GHSafZ6mdxp4DlQjZNQ4XRRTF3bBY5QaUKQ7Cvcp0FV/vJa+mPLbjaKjyMNQMizNbBo
9OEJ09s47L6YFnixZFew/59SzR/eE/VzeLsBVXhxJGb0NdB/RrFSeYfc/bndooiODiQ1molF9DZt
Yw3wl0HmzgN4w1QjMRDMk0uXMIabHvlihU2ZHXPm5zzlnNw6jW1hEwD2nAQetMAKmu7FK5Cm4lBI
Tv7VnNfgp6WTnVaahiS044y7H4viFEb9/b70y8V/WHa5s9tFYDJ6iSxUJGFtrt8CXH6SubBeQTzl
Z6u8KWcvFKiXulktwWRzqi9q77KCdfcmL4mRFgHiZX3wgPdLikBXm9cRx9nx1fcdM1CJW9Y74uh8
n0h6TUe8Z9v91/VSg7JMjdF56+wv59NNgyhYJgmm2PQcv8/pboxEPBaMRmyhGxGzyeA5ErA9XFTY
TL3lIroBj9RXo36KLPFuiDVCRI2EOEHh3V4PduR3MpFaWCEyXkVznRBzJpyg/0pA/6iXpWRJUijn
Y/I/t88Iki0/wx7REzaooAZ+seOrUv+NuX/PSzHchZOgH/B7204S8Z07b/IUMO2fCbPjw8A0jh7x
F/Bho0JmrQ4iCXG6ozovLq7CJocvirvCZVwtpH7QF0hyFZE8J3pGIbYmAu4m3HDbilLx+Mfgh8nD
tVnypbAB7/pqgMjRVTqP01g7+//ry+spCf38tXaYpT8sVkPbvujCkgqrZQkIbq4deeBxRfj+m0zp
IuhcSGDSz29LEH1WFlrxfupuxXAISxL5iBg20zB0eaiqKBjyn2sdeLD59LpQPeKmP8PZX/X16qoS
/eI/sLP9qmCB4Z0GnNUOJdNISbB2R6BfkMTEIguw/CxWA6vReUAenBimjQBTUJaDwWGORI1ubpNQ
9v7LYgEehEXw0JjCEeNjOSx9VRy/WMLCbGGu1sX5JTutJx9WbB71JlEJz+OvaP7Q7XBeEH8tpAHP
6eO7bVXleAoEUhpAYSfEhrL+ueU2Sh56wQMd95/qPQOAS5So2EPpyT5fx5ywFnj+TRkRlKSnHE9l
AvoTaMf4E+L2uk6rpckbV5uWC9HxZYB1HNb9Qg1PW7wbVgpBunSjogYOmESyguAh+8JzY54vG4kY
d9OEyhwoQ1OQ1le9waJX5UgPsQv8IWZErv85EhH2vlB3DBOnJviuy+aWnmVCiwoHwxSFt7cZfEoD
0/KbTawN2onHd8vRo9ll7L3AFPkA7jpODgmaWNexQz7RLJZ+UzyWGpNw6PdwWPcUGLLjcEit7NVx
gJi5/zA45k09O5hU7vu5qF4lSj7yhon9gMRenqxM+3MhuRhb0t2Pe6mjFDW234Y9pghDYNcgwGOQ
9VpwWM/+WmNfUvdmCatE6KCOSR5gTjkgM7HhRgmn/oRe8B5ymHMiHm3WWSHHOMQ8Xz7X+78xueyK
G8v3J0Hy9WOQYkvvyVV20i1Yyva/i2Hj6D5hrjwO/m6pg7Z1yLpNBHd+T0cBoIqChua7zKXIXD68
+/YBn2MYpKscKtacahkGcd2YvFH3M8q4zQsIcOQGhsC8W09etcBTlSBp1YPtxiFRombT+Db/YpZG
jp45GptcbwSJdUhqBBIVnXxebGKfbf6Sd3ZKLW6WZ9211XxVwHqEUwn0tb/k+i1n8N3atyOFeqOa
wrLCd8ENS/DZe0GFKNm0POILHsRDmwTxXSrqvjr7msu7Y6mTBUelGzK3IGlEXJtKy55CFvPo1V5w
zUYFK+wf8qz/iptaaHylxK57rFsw3RJqVxfEh3yO0zhWSRm+HN/W3nohSE25pF25+dfhjkn4qBqe
7tiWyniSORMZnLxrJt+13mWVge6P6yokv3Ea/hbz8KkJuTywHf4pFgv/wfSF9P64/0drSuT74KPv
45y2COA8wyP6f0M6F8aCLaz7WBk5pdDr0KarN/fbqYnvELfCm+5ZpXv7rsoVojtZhwFN2J6eqydF
55pZ9zCbNBciuV5PWGAx9mrQPMWga5zteBbozpkMf4nXznjgW6HWjBnXPO8RXqS5C21TxMhGU9jn
NE/qsLWHq2FBPiZ1tVHSmnZ8GYQYe7Tx171uU9fVPzbiFih44Pzi/lJngJ0uPFxihvEGlTaNQ6Z5
4XAShqq5t0BVP9bQAwdakyJFuzVdD4ckqSiO8q8iecvUMIb1UUPGbYtP9TkzMiHNDVYGv2nsKErS
mfBtvxnxxaiHN27do9FDvaXbtG8mkUj229lLe1oEmyYk0oSDpowjF0UbkEodL4MZdR9nTW2yavxY
sz6apzkqjSH8spS8UfIJlZ90UdEZu/XB1m1LKtxRGY1Y35sZxqn0gJ6VQkmM/UvJRZkdHGGOQxph
utnUvb67q9ZB3nRmsO9l4buo1w9uPEogqTXiu529tGKXEj/95B45g/ecyWMAWy3r0hYY5AuVQRR/
YpS/7WUny6q39PR20oocFvRF0Y22BZPAmVF9ML5Y9jRfGGd4ke5SyHRGUl9xLUDXCyu1vl+3TZhq
JDdTs4J4AGMYZEO2CQgNklFFn+81BeXdwR+IZ9ep8/8RTU8OmrYrcUm+QfTmFM3RMZNDWh6eVnI8
ljnBM45KadxhbUZV8tdmf66b6dSgdK2QUFe+ovfYQa4esdCG8KOc52XS7VpJKHeVQa2p1FJLjgUv
ps7w5cW61BSM6Ww00aUVWc5acjEp5rdRF8qJbezQgUivOHUlj7wHF+SV4RKwrDS5IE7evSqWZx2Q
IYr6PWFRrbIQ02kDZFl+sylPEUaPzKQLzlMMznroLP4HsmmHL31AbIEdCe8LDhP0JJ1GeQcN/eGd
r1BTwog091b9DIp73GdIR4LCT6Z3f1xCQYpflyqm0Qx/dsWEqsmachVn0eqcnWt58RttrLZu/yUM
w33cGwsy9hIColl+kvS6CCP1/yrT7G/g3tL7WnnhFZaIRHcdYWdgAWKkMaJHOl6bOu1DcFq503qR
cH16xi5fMZAmAQWHsHgRRqPMfD0VfUZ5twHfdd1aDiwremC3WTyZirqlJNzlNu8diXRBivxXJrmZ
8jSw9MQ97SpvSzxwCFc9pxr3pmDITiBQ3AIV64lL6nwTvOPRuAj/h+HzrifHh2hQB8D3paTSgdul
HrgI9zN6HUdpKHl+wkw16yzcacTmMesffg+rgVfX3VEtRPyXl7yFAbWorVh63QxdajHp7VsH7Yad
TKC5EgbFU5nlpk37WcTrvBJORpYnwnJ8lKlAVV5BF/XYJbP/KVcYpqo8PYRNCoNkBvbEaEVTTonh
HDKgrBS7Yix5LL+aIKXiSKg7UcoBRXunl7mJSr31CVZhjq5cAi/GObdGQ3/0ItHABlFfD3OQ+84W
+njQeMCHoBSe8Pc5KUVwITVO1co/x/A+k4PGdVjuweU8nPzskV5pAvhb4+PDA2rgHtFZaYeHSAq5
ZDH/lyf9u1lTIAc15OLvYsHWWVIfmTG5lX2LOnEIi4m4eUs7qAxfnHOybKCjHx0A0CoLw3qEpJNF
H/qB/JarLV7IbCzM06rWLXwmXkjNUJquRRSt+9hsQPXeJD+FQIw25DE0MDJ8eUUZC/U1HhURHYcy
L0V14bDgfZ73hjOnffbqJXq63kp46wGMRCXnsvc6Ro9InE1yqrn5VYevGazKvgxJ4TvludK8mf23
YwNhMIxAKx9E9VnzaigxnYk63m1Kiq7y4e4ZXnLan8bDLarMToPMiCLDXqVMvsZT6B7Lfsl/d/8z
eZif29ZKKdF8RjOu9TNu1upBaAg4c5ReGVKEs+YljjDQTurUdTwTDSQR1szTXpJUhGiYbqupKELf
8QR2C1yd24Zzlr/XU2YMRJlBPKZ4sfDf8m/U0Lq5AU29jY2Vm8nV802KjkZkrkmE36kdJQCWZlxt
KbccA4AiGgCXvbXTyIbC22U5c2n06pWdC1u4XqiBXiOPPKSHvAkneKllZ4fIfiVq+wDGkBTkfrqE
OzjkHfqmwvvlo4iGdE3uU35NdBgNpdOderQa3oA6uEbNGMmwf0RBbVxCXPaafjsSlxxt96/Dt8MG
vnMDlTNksI7kd611mgYC7TL03hdop1ThXaxI3/y4OwRlcglHfbXepKJLw4p8TMbIXCRgGHShwl56
v5Jx3uf4J8hWciY2t5ds/A4mXRzLhuOguTHJxZ5vp9LZ9EUeoXiCeqkFu12RKrLXx/7gjdTf2gqe
ScPEwCVmYMi0L+378TL9RrjEvKWAYGKU8a+FeWSfmpL25DeQuWVg+bB4Pn5aQSRLRU0FlemsNOgp
O6JJiNXKNJAF/4fmNJJefWtOmT0lLEdDJbX72m9DW03lxr4Uh1i/xltXZkq+Y4RsSMx/wUu74ymU
Vgjd+I3G3cuE75Gfo3NAE/2JJTxSgTPtE1Zmc17zatCpdAyLyuggHPtL08z6JZWGypaIHuBo02/b
rtgPbp/yVyQLuwHIj/e/svDYSR+PB2Ch7TN36jl919vWi0DdOg4rrM62YrH0m+Vpqrats/4CnCMe
fvaHl71QR9pyfgtJ7BkCxjpqzixi/jM6LnhVwQirt9r4muxtHfFB7XMsGK9BhBFQrXX9Oh6ES8WF
Y6AzQhCJXO/PvsOs73HsHkpE3MDJthIixhlqK1jQM6SPAkta3XqmIUS8ZZVe+CRkH+GZhyAimbBh
0Lbp8kWZfwN2jos10D1CINCdJbFfADUvVZqwUJmSOg5en87plpXSBw5RT/kpeUkfwdU8LftE1sp0
rqktk/Pu5ZJIw9WcGspTCWqHNVfZ/lj6XrArzB6q37UwXZA8Lr/0BnM5WmLsTjEhXS0HUGXzYGm9
R8jhG8P7BIxfcro1PIX07YHN80aa0qIQu5gGtWf7AabPvgeL4N20djhJ8T2VMs6rRECmT+vsRrmL
eBv+I7eFnFD1T9gg8xfIyKXaMoQNC6S3F5kQ901GjpJeLh8yEVnSyGxLrxa0dRX9nYnBaNw8/OK2
qlVs2uc0KjabwqlIXC5NhCprgOnSsJwxh97RGEKqBzE/fjTTF9axiSAJukqu6j2Mqr3Fk3mUKlmb
m0rP6n7Hkrv1C7psu3o0uijPV/3uHVvjioLvD7pIXk7EeWF+0Ay+Qd/kIuw6iDYP6qcXnFZe7Re0
k8Eq4h2UNwcuDneOFZKUvTqqjaNX01VtG1VKlA35JIjlGsLMBUo89ydL3DQMRnl8y47Ysi4tPj/N
P70df9QB97Vg/ceAyZjiI11md2iZ0RTJeoqZxxmE7IMfrsBKneg6SJv4W6veUY/XvMYRzHWDUAYv
08GCE0G52YsIo9uk3gXj7lZ1DidgtRhBw/sFk1oYH1/eY1sewnmZqnwAB8yFlrcli+bOr9bb+W5h
34vrQmVrynDFZ82rYd6SYKEwro24oWK4/+xLrPM5oknTYWgaKC+3nshx++mM9v14ybRrg1ubbTKb
ss+/dbYQUkcTETvZTZAoLG/uCH8XjxDjvfYanzbo9lHh+xlHxaZVEOCWtDsA6ShHovavz2mDjiPh
iNL7vlzWjLUQWnbWALl1Chvulo9NmusZ8cMcTDemZ7Co0JF3tDSoeWUZSjgq/HTuUn1sb03gpxAp
Prf4sp2HtAWLcUswE/MwyzHmOE3RRZD3nDtePv+9C4lZVMRzz2JEeax5LKQbSY1qQGuPbrMjjDw9
0ejzoeqC5b9N9DU7ZQjZTEcYQ5ihR0ZcJ0rVALeBCWTH0UyoTN6Hc58axxc2/ptMf2bvPikaF3KJ
l/p4xk1EYUEoFLEfY2JH2XIK7S5BZRMUIjseZK1uX8pMdvj4uIVp7VRmQwB/EJXd2Xmutyiy8xdI
Y4vKd4yGQIWa8DObB7GJc4b7syJ6A6mGF46SQLPNeBmotVdpnT1YDJS1EU5cONYi6Caikk+lrHjT
hW1ybVYqO2zCRhA9fhmHm4Sa7QdWwNjXPnz3E1FuqA4JFa1KtExsWRhTb2/ROY9+rjoOBdDRYcMu
M8K+dq+xSUn9ROzQpgx9KMG6eYRkoJDow6/h//2VTSvrRTZhG2OQU/z4WhZsc0Mr5jV2Q401cXjt
9EyVTceAyBJ1gEG3x2M22ZyOXoOnvwXBn9Ua1g1k18bLoD/cRwnA0BG0fKK69cNGtd/TmJkZLoLj
bFCcM07mfq4koN1AW2249qqet/u2INomanlsI8t19LU7TuEH6AFztlUef5Ja4tynnNCr1U9+vqIO
Fbzy4QrtHKCGt+hhYOGtlJlIJKJ3lcwn/SMIHYvMFzXgQPSsLuhSRpXGvbgs8al7cj99aA/sm1F6
/rQIJQBHAclzzcFmQrlE+joaucI6jlXrKV4LvOBA3KO7I02v3jMKQqVyMeGc4B4Cur1DTDwpRhx0
FLhnlosd5VoKwMZHwITu/sxP4OvY1EwdFHAbm/Hui5+iR9L6iPnlCPDAx/LzV43Ezineudlwm6+j
c27UYbrWGKekZi3+GFBJx6hhC1iMH+S1tOlk20tnK30L9y5vSVzZqs/A3a/Gibr9ReFZ5VgNJguk
XvKBF+YXRSaW/beDJUR5nm/4g3Oa7znJrNQOPWPkLS94N7mnj8cRWJ15YPAxodZFktcUpZWN/f7b
y8gEK7yj2J/ryivWS3DKmbwj70ciG9gwtuTYq/LZ2g1E0ak74cBGwcQFSn5VLk1NjA/RhpQgdNWr
4MEeUZNOhqFvv73SFYw/iT9OWGQKhrEb9QlX8kJgfya1qwgXbFh8JjCh7073faDoYZHLxuO2tud1
GEEfws5198FEWS7SbU6AM3Aqh9EkatVD3OLQ/MpAvu9UjGL9iTZf4eYiF2ZCnz3uOW4Sk89TI7zB
wVKOUo8tsRXmtNui0Z5GZY4FL0qwoHRbpksmkeT/UWKH1VEl1kl0//3tp5T5/gwQQPZ8HBRHEO6l
Fe6EzQLukHmlhwalzLRpTDIjl3DrO0t5nv32CvRV4AiK1ko2lKEzDCdKvF+Aof8b9lui3XUm5FzN
LJlvlAyWORhrneIX9EOwEr2R/iAKysHbtJlP8hWsjApnJKYsSRF6atQVKhqRXxjUcMeIUyOBI1M3
kUJMY7XxXLhBecTgWOqB1nwPnBRLPJpkIfj7kUl7XYsF5h1IynEEkdcMbnkWeL+5RHQXCUM0PZO1
QS5NYyp/hnxoOJltqJfV1+50Q0b0nQHUxtsQC1OXjzDdTsUqIH+qb3x9Vd8u//vaOE0kEEbi3NN5
sUls1/QVGqv32dKmheGQXS6lZcAOuijlXgXMDsOK4OGnR5lbsBgfiGjQIgmlsVrsCIhSrO7R6tPa
VxCEA0c8PRxiEN6XI9tBQPGXXL5RR0oSUOid8QgYdpurEoLBx17HbJ+cUjEJOXA44Xi1sdT17nOv
35KjgdBdlaScsoIDece8IYytcUKcR7KnovuqRKz7GEGve26x9G5327STTzdHhin5BrsUyr6YKbMA
DLmnYzx3MsPh2MUcDpc3m59S0QTkIXBovOXyHHbRZnmiK41F82gnNmNyo4XgLW+qymLlOBqpHMzl
aiCIazkjBv/aW/4H4y1wZIspTqE5qCe6IC8LRcNOgYTX32YwjqvJGxAd145ljZpPaNdl3FEdc8Ox
ONfenY5cuPzcfSDEY3eyI1n0t2Tf/oJmMD+eA6AaQe1Jv0B33clxBDQeGeLCFahhe5Q/E5UsX2sb
OLDxdpU+2HeagP+zGDhJUaDacTKk23jXJqqDikMwm5JoeAMH/RMpAQlMxAebKJeudCf8yefRx/Zj
zL0BKB2hZDSEFTcXNf32VL5z8uE0x7WaNI32SO+q8hL4xnXqG64sodeJo4F59HLhYu+3TmICE2Ex
kjvJpHaU/zbIsQybBrSEidCQTr6IxuzNCqndpN1diQQD0yJxB3Vr8r+vn5UVX8T37Ev2B3CZeP7K
B38NtGF/D5dhbE5PdzlU1TdxO16nmPmYjOcqIAjMyTgjh2GVQP2oXy+OH95Z9Pu6sCxpZa4P2jN3
cB/ZZMEQEDS83K8eBtY85Bl/PNUL9pgz4/IJMYeaYmwJMr9M35EJn2869vAgTNmCKeIulauoCxni
V08RHgJLx8mSJGXOztafQtUybOMpNzrMw+g/cuk7vVK06KxbLCtCPrju9dKgKuJYgHDEZyqdzm2Y
oqsv4+vCoO5M29+aQnS3tnyI9OHM5sONhpjCk7Gtk6NCWzsE7PHGvJBM/2gvIb0Y8ySAQLiMKSey
R7UYMANLznY9+jWwvbmnW+iN0ct/LSPdZJuuJUEkbSSF5xOPGYM+ftvhCK7IKsUgcMXFEK3OD0+m
Sozsjq1QIzifvNF9lnPvZCooiDtAhJ14yfvKeJahppQLTlMlo3mCwZBNAcDWAx4/pDnfae0tYccg
naU/czEaqdz5xjsWVmlnuOWTvWPwrGcQC7x5V9LALnlfma4LgNg187aenXka3kKtibuxRuY6+kIN
Zvzdg7rukdOlfuJMXpWTYDFeCkV5cay6+FLglVeOw3ZIFvbcScffmAld7VVbsQCcnZCQjr//O7lY
DuF67vmq/4sMX7GS44EdZXj94rZcvuhf+tD9MBmlyGqRyFqc7hHb7RriYSD4c8Kq8tJ6LVigLdcd
TcpYBKh/pQ0PYtSM6qBGitPzk75k5iZMayJnFTGuLtEuWO+9EIVs7csVmbSXykrDN+aNcRoa1Asv
LqCUkGXWPoe2QnsTwsM8b5WmXJ+hcUMyxdBAuE6Sl3fLsxuqnaC+jk9xpRVNkGY7aVlPo4CUvMRd
LrEwpwfyYyJWkCOZ7Td6QwYarwatCcT+fu9YAS3JR53An+hRnLioTXYE3QXnFIazWL/8XndS0QhO
g6b/pWlsuu38bKwr5KXdCGvf1n5nWj12ZJKcwG4pUT7Bo6Nn7T95gqN7bGX1bwxGvwBzn/TRFNmH
16p4/lSkh28Ybm8BEhanC8xvU6EGf1kLt3llzc/LoFc9wDXs6225N16/tDWP9ey335xmXC9pBVDY
humX2NCOKuDntR/i6QZXQTia07ixJ/3uQeErYIE6pvCgKVt7+2Ov/YsBqvnVsCg/8RrEoVG/7r/y
b8DXUJ62zrMOTxY+Z1fn8LEGy3f5UhzS0aAbtgm0Xh6z/W1FVuFX/FKNlhOCAPA+FSRsmZ4YWNsm
3jnCybh/KUm1avS4XDxnSe4Y+ICoEzBByj+eG5Uy9r3cRbANUVKSN1AvBTUe4A49l1Gb3K3GB5mr
G6dbTWjrGZu0XV2ItomCIFiMckN5wg0xIvNcsmkmvaKMS9wepyrdTLWrhU2vRsyZf3HfHhPpKAbg
B7U0gqQH4V4hLD/yNL+SNGaag8ogfgS5tmVpaDDHsTeArpQ+OLCyVChGpk/rUpBwHl/V0BdFz9xB
h2tJxdEzmFmwmqc9kvdGosDj6dtcFvuegek4r212l9PFTYFlL+WpUHCPAISxaN3MfTOshmvusVup
MNYm/qEmzzy0rUyVR09xvIQCs7+XkpnnioM5IieeXHXR9SQPOeWuWGbI/yu1TZJ25fY8hnNlaqCu
f+f8FkAYBJXmvwYxf90A4TZUCg5kTnxWYvDik9SxFvJr7ukUQD+qLrjrwFKZ1YZLefpgX6WcCO8t
TLX+jQY3M1nH2gID3Iqj0CEZV56a0ZKPRuSGXvTmF5YL0KK1weHMjk1nRMEzuHRa/zTOeNRBXG33
IX2VlZUMTAf4aESCra74LFGDKuDTbH2/thcPc9XQKH+wnHvwIpuj4NVyjnG0gMzK4JUfJHUXqgkF
1s0KimLawKaA8gHYusFQUK4ZhHrEHwq6P0XwUw/TrA7xuocVWu5MeDx5Gqg+xcKcfea2dGfqNYY9
lYO67H0NAV7DMmIpihE7eFbN5aJd5kqkxnIyItsUoZp9rC123L5jolCrTrnKLZl5a1ZwGIZT1JNJ
pmrkJ2mPAfbruSCjkeJqtZe/DqiJ8f655KCH7Q7CU0pLP4xc7DxMchgyBVz+nWSe11mdM4PinbfX
dt4A0b1H1eahTOyHoDlY8BUC4jNjYDitGucJqbI+vxzPqCem/l8D551eKE+ehBHzUVKZ+hS5Ov67
L3fayW2yXeLRexuELn3kBlqSyXUAZMhUtG5sdQSHV8oabiBkWHwa8a3CpMdvKe5o//8kahLLnr4r
84e5om9f5Fnhg/jmTkIzTqTHOPdNPZf/cH6Lkr1fixZqtA+F1s1U3DjWUUPc/bcDau4CmnMLrYWN
NePQFB/yeKejUIbsF4vHc/5bz0stq1cPnUYBpMg6nph7JNpeJ6A6EYY6csT24Qekg2DByidwCpqB
Cc2k0WQ8E9Mh77kSl7mGRqdaYyZKOy3QGsrFVd+0hW0jkeFkOxeIaFvqjk9lq+vxCDhguYVuDldM
hMK4jvOYDIf98nMk+KdKI0LZkaIa+nhCY+CYPkGQesEDlV8TgCcykBb71A0hnlEnnEGJKY93wD9l
ysMhBpIxDlShVMtTwr/iwhsrqmeQTjyVjiGP5O0pBMGx8j1XYIkQLqxX2zDLbitb411TIfb166Bi
DPE/C1XRFYEuKZtg0QcfCvx4HrP2Gq//u5jM3GJ0NCoj5Pe+FEtbFc1GiK0Vtz8i6P5DdUT/tMWc
301MF48DSVSOvsWIjqHw5R6HDuBgwSf2pq5SbwtQK35VrtVw03nDPDtYzhk4GuAubSWlpoMKl8c1
7BcQ5xGcPn94EtsfbFug2ne6ZCUjjK4F2lbH1Ib1sCf5MHVrqid3ArkdLUSwfAZ2mIVjappkTE70
6VV92K1prMXcoL1qtTqTkrKQ50WU6WX92qdIT2/kc/i3PkDfxESKs08nveUo9zEGclPmNzpEQ8LD
OrEJ3z1NRrA4YrsbShp9ToNlJbzCVdVKqOTPKy0vFrgYB1bUZGL+aYmUtYgdh9kK9+dz0ysxKZsX
kU5zIsANmkNfyCVm5uwxInnqbmHZD8XN91TP9/Gmzt8OhmzdB5M4vqjKtLYJJzO+xUIIf45mqLsy
aZkN2Www2TBmgPSgk8wlE6t5OHKYlHI26GKapcSujwJ5zG0daCHIRLzLSILGfb1e5L4jbG7Z4JFR
JEUKObrtA40orHDNkZ7E9UdqxIIJaHwyLfJk4FZ08Kqp1jrVc9wXfEvNFdcNm0rVFMAFEgyespNP
KdW8hj3nqltcxTB9AiW9ql9PAuErlUpISLVmO6sLcbsCf7nQTcKXKaNVeKjihE40tqkfT58Sx9AB
FO6AkpwQG2O23wZOqo1R2rX2SSp4VYSdBLZO5bi3mg+QI12svFyI+PA44vJfUBZq44DUFmiW9ayJ
ZVA22fGiR7qa0S1GdG9LhvPipGtySPpP2YEGzAQlyG3qr/6O6/cDeyE7GZvXK7LNYl9f+GYJX80C
N0LkmY1cNv4PS9l2lEx3xba7FTIipmuuFfXC+ZBKOCreDZKd1AeE5H5zuNLIJZqCGZRpIyUSO7RZ
v/U7sl4xFG0wxheM5CMywbhNDcD59Ddu9807vfx/24ORIDxFfqSLamHMq9X/5N4+Jjo6uxIFLVAq
jtsSaYFrSvn6exZ7BqauCTz6z2pdoTrai/bAPXnSXQm5/fMrhvszv3Z1Te95S5rQRv8oakWEGaYO
xfQIDDXrTAJfdBnnzUk/aBOL7uclmuCHMN4FVDL4BV/1zxf6R3t7KyYHIcURaswlqNQoc4S0iZy6
pG01ICCa7ZANP16mW1GSXhgFIybOCqQx+SPcMqPFbWkL4tlgwbkZMa1NDeBhGChRio4lOEpZYWdV
/FBhsfobRiDQ+wcqRpjZffhSmE6TDYf6WTHJvueMz/jAEvMF+Z0clvFj/UcMDHtIBwI9dTfL+bba
yeddpBl6x2Job/69R6EOnnLe33ywtCi9WQVes+aDW1WqTDHrSK+Me8itUAJ4Q0kk2Katv8QpAZl3
+2ZVzm8XQW9vc+GdXrN+nNqEuSoK4xIOeYKot7d6jokkzwsIIujoNkoP/CQviAUy7Caudd7I+/KF
AuWOBr2cqUA9e4SUxmuCla8CNUDtrulY4W62yihfC5sGF5CyhOgPUVbdMtsDi0fF0xDsa+JvHqp1
MnaoFtyKhrZcDIrhj2cZhMKqzJJogE4rzdwZQmD/At/FSaZkPpyWip1pFDq7YNMZmbz9yI2i+EiV
DUFRKb2Zo7Lpp68orHkgQAdTvzSwjku4gnU0i7Zfpy/ZG/7Ils5J3oNq3FJTP53jFnzqirMr+gLG
tAqeBykKK+6A4+24yu0Kx0MOlcTmnWRgMCWwJP5ZjWPudM1gPhxiEKzWlCYv+cw8Zof+z3MhDMDD
g2yx+Fsio6HhDtjmJ03ngql0u8ch+XM42yPVcqmcK0Kskk9FxwjSP0nU8lghl0OqbtUmOkbz1q3N
mpMaV7gwxI12xuR/N74SnbdmHOokU3/CukfFVg2I+wASrcnge16BjC9sscK72RZMoYbZzpnO8hC9
kLu0lHYaFr2VrqMQAPjVs8iaDK/DGy2H08GtUGkmKHMuLIIlmqLDjxuHbBeu9JbqNTGIxB0JWtkE
tG75NeOgHt5pV5dLWansdgJawLdETXjw4ISquNbcJMYqoaGltN4BSSbYJDFDV55lG1MAumGZyoQl
WCyadJZffFH/n33bjDyyguldrhbsX9C0IRsj6wmNM/ANtpIZjM6L2+XbiFzAWXo76z9yfLSAryF3
Zf12e4LuLkla62/b3pmdEV3VXGmruksDnDQtKc+Yf/MSuXxvhpTvRECMZEn81auQUAfhdwI/xlbA
v5NMjMt96ParB8806vUpQ2ATZ52dN0hLSw9nvX0fpKwdVtuLUzr3K5OduRW8a0WmwQJu0/dm2P+f
MOSYCMhghntxC3aIvJrcjQdI1o5u+HFAak8CPWmD5dxzlheTkRhS+0PudZIg3oQkA4DyuXGzInMI
aJWgW3T8PqMOjMtSV9q0v8/QcFGkecKM3RGollM35lEj6JIu3DPNF+7cFkeceamdeMU57UZRXso9
i/gwlpQXncbqtfvW4mo7ZsH9mBVxUSO+fILYuXLvVtRnZRSi2VyY6oAsc1EA9dNUqDGU4GdS0noQ
kMuH9BTriUn7liD+eYDQ3/DZ8olr9dJKCtYDEO06ZeNmJGLghhvTs15iK+frVlQ3NzscLyFjEN5T
h634c/HUg4btpU191IDx68ZSGVgpc/+1ds7RXFpCm9ezT+ibfdhEv26WK3gbyQ9Fx1VmQeoEGwz4
cjIf0gsm/P+6V+ZXubjMHmR7/oh+3iGCdGTG16afiTFOVqATDymLrw4bpenDPNYx21srhf0jvyFY
OpxHddef9NPo2f+osZMSS9nt++3eadmL9vAXINRKV37BCeseqGy8pQd0K8CpnSsu7y+n8nRfdUqA
1wY6y0efebgcOJacX1aklwGNLPu8J7XVSx2TBbhOhySoIdcEgN9mjjc3MCdpCswk4vL2pB2xc/OT
mdzXKzMyQ5hmaW0ZSDivHcH/HplflMHL3VQNIoEnIALCICVGYGxZJn+0fVjeVGQ5hPKyTkD035mY
wCI2Q0SBjTeMfzj40byk7NHAN8a6ojOV6QBILU7gbP1Q9L5/9VZlyTDrzAHYO55oTvbSOKFSEXb6
sU00i6vMfzfzLlDcB+GFaz2IHCGEiB++P2KV7GqW6IiWnq5PZXbsVG+F7+iZ5itvP/czbwu2p+en
uw3PvCzzHFiJ7KlrH2zAn1QniJYvLErsCd+z9kn8Zo30CrmnSOGByvKqSjkYO2aw/c5Yn1wcrxPG
Xn/eT946wbrbJqU82ndWj2Ay0ALelt0IEDTtyreF9rFX80i/yNcg54kIxsBaIgdsv0jRnCzJ9jC7
XsL+aZJfoIdfCLiR6MqRxjlkmo0GgSq8RESVftk1XroL1EmcBT/4lAdUfKKnG6+kAT/pl+mveo/5
eByfnMYQEwwtDnGwOK1Iu15m4y4gkCD3xZ5ovnozeaQ1vGipLgh3ikuSpG8cH0yZb95ReG2iBkn2
Laz8eXaj6d3wZLXfTsG4zpGly5Y2MeJ24vkwC/tKBWuuO4NYU6gXcNC8S1da5Ql2wMc402q+HOXk
jgiMgRfZly7kf6XYG5sJoiuMsCnFiGh6AnrZUNnfO2I5ktsnqMs7nZCf19PID8a9PfgU6NmVCVT3
D1KbheaY+5DzEWYHMeJ9JXXAshRqmOsDMryvVFKE+Juja4OcfOqaURa1aOXTy+iye3l0iYEm+JNK
WMlT8suKOyKI/ttiC4yGIiD8OBotAwLrCi0fapo6HcnHEInDbp+dI/6b/POTxcARX8ZD20N0GIYA
5XbaCLBwEPUzAqjYsVl97I1l0y3bQQSh8w2pCUfi6mMbOdRsGE+h2cgsKsEl6WV/jBLJJEHFMIDq
b0F1pUe9liaF/hKzwHROF5gkSpA1l89pJ2TqKnIJgU42IAjNVdzoW+6c5T+raKHfYs7LIVhlFikc
3Y1cstv728eAl6zfAfsevZ5jqKB28RZZ3V3+1XetyL13j8pdbPprLid9qZwtatLF6IeN38rbfeJw
56Q1dA9CHwbgUu7RytMX2G2YgUeKUSKgkRibUnjoVqh8/uUYV1ET5F9Mk/b2y89Zv0RuFUK7/QlV
GZI0HQ4jj2PvLUogryZ1l3F6Xjw1bF6ZjslVCGK63mr7/nyVGXATz4GDsQMz0dKBvGVMoLyG+KYP
IbqwO5PWU06A69BKVTyyc57zEk8Nhx5hlkag3mYipEDxaycD1CyAhx0bmNB/b7AX+jGT1umuzN6T
ZgTtJ4PUJOfF6NxmKiymntH58vta1phORJi4jyJJVl1o17tegF8N2MrILr8PPi8zdCG9wXRMmdGT
LQTGYxZuW6o/tcBkF8yvzm+8P5iJbjItQJRgx3YrO79/0j7Z44Bo01PkCvJo9Zyw7AMu5N8y+JFO
FF2rh2bzjq/eGFl+iNHxjW0UdQquOkEANmlR21MZZv542JcBWcDw2re0BEPGIm1kqQ8QFY2pyjTP
nugVdUt0ZpS4eDY4vocTQ6UZwQqw+xxA/AvXWRkqrHbhX8bNrD5AnoYT0AUjQWgMeksego+XGAWh
UZE1opkHKSrCMRR6yBWbUNA1SkO7UKDhnNCpueA1l9AJRU8/FLMle6DTfRM3vHuc8kjbcgoaiUPU
aoZfvGmpT8enNqrkzZMJcFsyfuxzreAwlx88HN0PWp1u0SRvSGaqx0D1WEDEcedm9vHFRWYyspy+
tXCndqOXgsKHY10q0TAJHP3wvyIWxIDiIWkGoHFG6PqhaK6apf+VAfb5VoHLpjYSQ0pIvCnbrcQN
ChlvIgbrEn+4sMFnjRLz16i0iySDT1HHGzi0tjQx1+wwsaD69VlVrfYu/BMVCfqJK1NNF8kYe1PW
L1VGd7B9ljEQvFZzFKmnMefOIycSf9UoDpDRNu5UY51fQm/VmWD/NDFbmVUBKR6XFC33tl0djEz+
0nCNEV+vP+/ZKfsUoKGh808DJalzwkVPsM6a+a1cTVAKBKbmIZqA5Ar8R1ZVzL3NuxI2+C21HEVZ
Bu5mkUgbXDL/aBu7evKZkOScdSFyigvoOs2V5eiEM27mkFZ07LlK0iSv6NWtpoatUl3AMYOM0uRC
msbBV+XFpSdXXbkTgHDc5LoHBms2+tFE7KOVQt2nMZOeyhEuqkRPxGhQtx8zkdwM7HPqxyAln/93
2gqu2c0NpgGV36IAMMvunjnBgQz81dEukj/isOFZ7EC/vfAE8EIVy+D2ct2bpfefYlZ5Yon/w+Pj
ifHpgUOhbLvMMdvgZHkceafbTuhu46el9k3NwcaNOqajoQxNyW/Wp2EXrx/sYRWn4HJ44pT23wqW
JnqgOQUOiATbFzrhxXodidl5c2YbQ5V8jwccrJO8YQRcGTDZy0Glx0PumUNieDpg9BASAIfpW2KC
LY90xqQIdu8FHMbmvYkGPLNhTt1cNk3/JkwNMEQt9yXlr/Ow0Qq6GYQjARb6GJsy4IzlkDM4iqt7
r48M0l92MY2Y7V+y1/eKBKypYeLPthwLdpUUbEzZ9C0G/ljAyz5MOrdauYlVQYePZUaRGvMMSH0O
mv/ESDCLdJlewAkLNqJvyXeljoVceyBebWaMBgopgbJUHL82FsGehBtroTCHxXnmK5hdyMXqkPJ8
Ui2bzPHiSadLnqIt986kuBLYdTj+oShbomsp8art0JTN5rHwxBUk8vYJNiqQ2h6IuxJMVs/Di6rc
XTBeoITOUHjkV854clj5QKxzpLJ0SYGKfbo2IgxJyeHzEcDlnCeO0zrm6b/aBrQ85XZJTdSAHMbX
dEL/DVOXZrFZ7blr0sozqwL5YJLsK3Ouhfaxx2/T6heDPSQ+OHSujZbb2oBeUnhGaj2RrEfFraU2
5rnlGrzsvBKfKUPraM5PmlBb6kbQg6adk7eS0ffwnnSfm1bnuL4hhESThrQbkTeR6v7k578Xd/8d
ijqYbp521+2IDflIGJizKM1SIdzLBopCpUo41l9VlfzdiSP/GgojVItbjd7IxHlIG6Pzy5oVWw8s
fT7u5+e+OhbLYSMGH24u9R2lKTubRwXzVTXi8xox82RVo1wl3QQ/HBuEKIF1eHWiXmuoSCeyOFA9
R+LM4g0gHyeQsf4MR27/eJoYbuMXMJVKRjLqL3vAq1q2cm6eX7/bC0CkJk90Qb/X7KytHSCiyxym
HIVq91QXDETmOuKGmWmrl9S27FgjoKh+04OQOrprH08oIC4iOz9V7X9dRzX60Fk0K2yPpLayEGgu
UsMm/jdQlkWkc6FOkKWH1t/LCDjskDQC9dAkureYh89pFf4+zBmiUUwRKK8xP3TXWCRgeI30wnaP
igVrOoISsLq+rgCdIaAcDIB+ka7UcwJt5oimin4woGRzLKLbMkNULJGHkaXIRnUbk1LVHZ1VpEYf
ZcHfWUyS9CYHRVug7MQf75nnA0ZjkAEOwbB0uPa07hh+OpBZmPTwfoNWkhL2Kn/phM2VCxJUvr9Y
wOVCrcy8hpdzATEDW31ytLTlEiv23WeBlFm9KDtw3/UUyWjoOFxpEnKGV855y+dK81NCGp6OQ4hn
Lwg2uh1H7P4/0nIk0ZrBu/nDZOQTHn76eOqqhHGmfmWiOVm6QBlNfvj59/GessiH5CrSeI1G1t/8
AP+kPtghJ8XEPeR3S3jQavYIztOkJswI40oND/xiZSZ/ELei4dWF1lS/VEhoTqZ7CK1E51S5Y1r3
1NCU4ba5iPNFyXltdt2qcs03/5KocWRDzQwcT9U23EKNQEk7iTC/xuQl2rvfoaK6gWUQBl5a8pSc
SMM92qsaeLMA6gV14tRnpkAiTtw/88WJDeRcZ8lxwEQZYuEFW0pLOdOm+kM4zIKXagcUWI2izm0E
n1MSGufpuIeHd5gzR3hXvCsSePKqD3ozOdf2iepnVsEotBBC00f+usnuxS5dyas03GoYm351iM+9
obUYWa8hTvkGrWKV55EBOi+wKm5qGFdv4kFl/Prt4F8xxkZWD7F2qQqvsVCcmkuCaj4pmJzadbla
mBtMXb4NVNzmYIjKrVqKZRB82StHp4+Xfga6S7ycJE5f0AjNcmOJaj6+hI5qDPLxegnaaZBOTVYt
v6SNgJDZpn59HahvMfyjoOkEPGFG+OH2kIHvBeZ5hgmaxhT1UHmp0Hftyxsp8bTZ6mI8DISpb//z
g7BF8jcyXpTyDR8K4siHvF3J0nQ2TO8JNSIlA9M6BpIA+wSlhk54KHJWekgUZ71LqTqy1FX5jW9q
OVBR5owDXmB/MKa8/aY21yZHwviJfaf2e7h8YOhGEbDEc5BHYJDsAUu1EBN1J6oVSIumoeIgrR/b
+VSUmWUPzgkpvTNFAb5la9MmbtJWlpy1iRTlsaVisGpQy2ztBuDILh+1k1KJX6PAAGHxDGr3BdFj
2X92kq+jLF5A0xFbdsblGGbLTQPOndCrOSBAkVQJcI6NrGEU4rQ6/cma8Q1E5KSoidvC3KR1X29f
HEvjBj7IeeB/cM3aGKBLYyRtzpY9cyc+vAVOS6i+3ecIfpquow9Mzljk6BgC0bKCMmGh071kfTmg
giuaQ/76OsZ2RtqvhNNddPHPy08Lmti1IBKnPm/6lIqkYylpjt/H72YCvzIDscHTrxJS1OPB7hhm
xOwQokXhMhOkuEPtvz4solyDh/zvsyaQOeC+sJH7L1nb2MA1Sc6Cwo228ZTaLeL3R6K1OFaD/iUE
OIMxgdVCZclmBPEQPxf1ja+//vxEUcStTiLAD1RhST/ogNNwzzomd5TcugE1Hi+CrwClEiOWPJNk
5DBwVbx02qQ0nv0LuqnWIBpvnSVGE6rzT6pct46bNYYdOpAm43OkrxDkFdPmRVdgDBxQ3uVrLK8S
eHT04TIxC6OgxpUAF327uEEdSO3aKjKGuOIvxtVwDyzPvjYUHrGLSOAZ9IHxa+rPEuQcOs4Sl7Om
C7JObsYO9tU7n4MIcXbotGjTJ7FkKpp+l/dXr4WYB9gNluQddG/2SsT5fF2WANBbnV6VtYOqvRXj
/yTrwLmFlPFGSaGJPbnJTV5T5Zc3w+xsIvwkHn76TVJAhEPv0k1gJ46oS9lwsHW+dssO510C8+Am
EZajtNUJPfc8HxYl7wvNR++M0eDtIEme//5/boI+harHXqI/1fM5qK/dN5Ld8zZpedLgsGXIj273
YPXzbduQDwEBWaD767OpfDG+/4oeyaS2aX2FLlt/Mdx3OiT/QrBQG6bvjGggS+c4sTuzjOwvKKA5
PIiDO4Sb2KGPj8qsSiY2B47S9k+p6BvAFuxlM0im+sM7c17kIZVObOkHJif2htd5SKGuizWyNxHp
QNEO2aTjLxsWBcwoWEFU+XHYxGTtnQwrwe6Bg/ajk7pXlRsmGhTQbaqXwiQyBOHDtSbaxgtCuPE7
jxesdsvdgl0MGaSH0Bttj1KzC3osCREymvIFGNd95QTCfs6Ft9aS/vq3RzfvO1u9VZokB3qNe4cX
s47PkMuiGhr0O8C3E+Q2Zpwg1eFf+3zdK8MgVkZcrDqV8w3a7/RTMRvmn2o980PaP8OlDGeBLx2K
K/pnCISS0gc1zt4J56XN6LexgDgbg6zn+DrwuStrHSlC2c97yKzwCxxkHj77vje1kl7kbd2zde+r
yvzP2A1Otsx7WNz+Fme/M/NRku9Qgr7B1XF0quwP2v+0La5gv363+ERvzNybnY86ku5s2vE7n72r
UOfBshHPi+UEP6j9QTSgeQbk+kI0CR6M56yCzLilg+oIG0INxmNjjVP4PFcFMnrabORHuYJHnf/0
oaCO0dX3AWSI/QAnDhWbOaHhK45jmVgu1AVAY96uKlV2kPuLVwCeETySnK7hpR1wZ2I75VKK7PFz
8x/eGviSTA7fGKhW8emPPpZyH8xLFY3C6Rk2hYI4jY2Zxieo9IQYyF9qu80hKbrXyDqydXpfNr74
VQa6O4WD+X5M32WC9k9iACnAq2QBCDslHE6eblD0aL5WImicmYRARn+lmjii4eoaEKHXteiUDtyo
K4y8t8RpskvG3/l7ouOjywE0piYVtkwmuOw84OILxXelpD0rIvh+wBIikobvTpLcADA8L0Tsu2AB
Nsvd97Hl1pNkTTEhkC43mXDYx4pNae1SrZom07iC57VHK6GxnMFIuVKHkqN8qvoOe6kEvgA2Bnqs
n3k6FVw3OXBNzN7SfnB3Agto11KxeGrd2XmWKzremBY2h/Tn67Ttlt6Bb7U9clri9aLnpOzDUCdf
nrB+Z0YbyyAijxfvAK/faS5dhXIC+nR94KfHzs6vxx06L4YIauKL3Hh+P9oaicmonfKFe1Z8yTf6
H/qNuEzZ8tBd1egDFwRwrc8YpNOiSmeahljaBb8Ws4ZqveKCWLMlwdwgO7QdfuHLoi1QwXCNxC55
veMDRfm1Qas8OcTIa10wMjCa40tOEranqkn8J7D6p1cW3mW0Pu5ViYYmp3fmyAOzHnGc15uZ2SLV
xQVuF04ztmWpA1DxcHIUlmu0yKUSQawwmb+gGtIJq+EEv1zDt9yc/vaIPpoKfiq+YjFazX4wG3sd
elc5Oco8gTWZJEUir+rAxwyBA9jPdwK5QBbbDMetXRuLnHA1cZ6XI6DYe08xnG3KdFvygxz1dmu3
2xjPuILicBvZSpEq81XhopTMnF2bcExvTAzsFvgkyrqQlBk8gTOxpRuLEnMk3cpWMlerbtY/mY3s
VsPbo/RcpL1Rf4pW1pgroxCmDScgku774mK+6dV0J7fzYjLC8PrrKaihN/3+uYtON4dbpEt+B3lX
MwVc466VUZbVpYgBxdxWzoT1hIxJGz5reQXZQR/jpO/ZMsYPLs9qsJEmwQ3cKOhOfbKfs0PkERDe
AJqCBptm+hBeJp/tYJdYXz2gVIjVgO8WQT4PdlV1+9DiiLDBZPGtT/5lwkg7C0jKLa1e8NNpaMsT
AVaCPzO1sNjoMYLMNhLjaiOw/jgnu5fOrCYJ7Oqs7q8yBqf4hx2PgBSP04lkRXblkxMnVwfj9Oby
5SWYNU99a+/RD+IJfGw+qjNdZ+tO+5P5BKp8KolpBfixtd7gIrf6RqNdZVBLv7NZztwXz2CjVzac
qWuo2dsTihq1zSP7p2hEajHZguMpoLcKber6sNdDhOslsq078XHujd9NIpOaQJLfVi6NFYfU5Wls
nHkUD4NsW9Y8dIORWrpEy5AEarMJsg/W/YjvZT663MmpbuHFv/0LxvTurMbNjqxiYyQ6I90VLBIK
eoBJYbp2dSDbxdHJlD/8nZG6JDI6k5Cqn77GEZ4+fIi7/OlS7SH1p6WlVp0cdCcyIXzULsb12uKJ
6desAnWr/KGyJ7OkYqmULvRaPTY3UdeMY+3xEnPtQkYd/xP3L0rxsKd0quQYWYmA0T7u8ksBmR6G
0M5ssbM/ywGPdmmERE8/HcVGyloLNc8reVA3TLKmOOqTAKaTPc5vgOdG1s1K6OUkyX0YIT8R37nH
pBSKGpdvrjVZKH31ZWFgQVuXyU07vHHYkpo9ppHwXfK1l0zyWhH1WvY42auLhJxhVQLR3x3QyBBB
SdwmNy+nWyQXQhPOoDrb6hRzVOgXQ23zyB7XoGWRiPdld/SVC4BniclanEY0UiM7/bkyHu7rag7D
jqPM1gQgrjAgqECGFASN3/wNzGVM9mNyCRG/og6xBk4ZdDAGl4RXkhH8wf5MiA5jwMMiTtLUa44I
IByRaD9oWG++XnrjO1yA+QDmMCYnIYpTolqWMapmFSt88ExWwD8rMEfoh+yTnW3Grp8d0lE8k864
Eg2jxduz8PDy2iyw/jVtS/QJmYgZ69uQaUKaeh6ur1roJ8VjTQ+yZ3JPhvR0lgckzYo6KMKLHWU3
7bTynVJwA73+jChe4itZujemwo77HRV4JJOp9uTM5aax/YdkQlmDMWmBjV2orMO0o9gL+K/k6PTd
cicqyHh3qn68aYn/ahhFllbJ2T60jHeXMDcYmsECFd9sPcklFWbF/8+e+e4qwc3nngJDRwB4RKXS
5z+UWgeQvhQbATC/XVbx+YjclcQlSBtcIQfhyNwm13/zJ9TnYrGKLb7J+gcNrQp3ZRZ2GbL85NJb
Xe1B3pQ5rfI6cqE5APJJxc1UeWRn54P8jSz7oWLwqweeP9vwwPdf1gMXj6grm/4SGtSwJcM/8JQo
AOLSpirJ5NHgwI9jxCCujPuO99Z3QtUoDyYnMTDDPp5wege7zjKTELrajDHmomFRZVPVQY5IUJEN
xXJlJLzM8kCSf6VnfRUN1nWA0g+RqKsT1kHEMRrk+gTZuc4KRbkrSjuK971m2iJ513N/q+UgDbjH
igKnDd2h2ZXLwGeyWYBRTsjLqr5Sq/FrwaVqEdztUQ3YlQSdUjJ9pNOb6VLmrFrrE4ppO8Xfqd6A
MGESG6oxi3Jph+GucWe5PE3zDdV2EP0Ms9hBQmSTS528Wk63shOM9KUgJ5DvChS1AqSv5/KdSjuy
BVKdlqpl01gQDU/KjE4J5U4UT2JKrdPEnrnr7Py65WEnlFKWpKgeh2qQ2BrYiKCVHkGVo6uMOnXo
0w3ndIYrJM0E99Kpbeeql8Y2iCa1jOOo8DBo8IS9e6IV9kuhyv1Diurqa5mlakjUAoXEPOUPZbxR
P99l1e6hH2KlTs47T319jPOdYL35y01vNDIi03rienAHnLuslXbn0lE4T483885UygPjcfmHXjHi
dsb+0qPuXau5xAEwlgBYP2bUIHTvtPDvfs3e1oedKbsXDhYgtwohS7ms9oIWPbpQutLGkZpei4A3
UgVqWXb7KQtG5zknk+tyunPjo3BA4cXNeUB+Yjnxvsln5adedHQMw8wNKArfsM2ex3B3dAj/rpL1
ROPjcFo5QtjhXQ3ndQ/S0LxfuubDjC04wUrVWH6iI/HWdnOHN9xFY1PZpCEL3hEyJvZGsLaX3HOE
ivTWWjyH9A8oG0znxv1Y0OhrB1rckMk1H0qEVOmMfZSP5RhqUUcZq5BgfPPmbxLHuFOjG8/EZmju
OKm88z3UCnlUEEbAxbVGARgBDlVNVDaL6vaX6XAPpL/fgxoMvIWh9jDd3cpY2gxamcaffZ43gZH0
otHPhpAzMdxv3bU+OYFURv+vPAKN/OQqCrEN6CnLJ5SmFRdDwNcEIfL8dn/Z6WunwxT1AnzUuXFV
ei7ohM8tOs1tLWGaz4NvezQcRuzWW2BWiH78pY5ggJP4jIuID2FPf7MMLWiq13muhSUUoUt2sASS
qSHaeBlZ9AR4TMxMhPYltSs3oPHankcfl1mT5cduJdmwaCVfnrmtqxy5k70G1KzSBsu/T2FaV8NA
wp9O5+kbC4fBkaanKHB9taNaYZtFzW/1fsdaQa0fiVeD6TbwKktrGPolPu1cJ/kOFZybOFy0j2r+
tUe40TzjSXZh0QbTrT/WphslrgJPkDfqUiOm1AcCA+TAS2pcJ4q0w0ItF58DS4jmufeljqaslqcF
i6c12ma++grE472b3nZpqhWP8nUqM9sbsaO2pghzXKAyKxoSt6QYQx9VLs3OmtinyIjvhXYoPAbH
WGQA13+vAvXvzLbkPnOXhrx974kZ1mr6Qxcd02FvmyctuoIkCFjCBMNUx/l7wF53Z2Qpr2Z+ytW/
BmRe0Ym1vgMCvabNcbUC9fVFggMmNM8xbl4M6g7YFQl3lN6t2/lTTYfMORGQSXliIWDAvHxa/6C9
pvbBi3AIF+QjX3O0+1uNYzrJlwv8GFBv/9ccQmmAvyEVgGmvE61lEkbrxK9SSNqJqofivJZZ9hUo
skGX+acP4YAdO0Fd8NSu6XNCI+tns2rMiRFam6ILM53Z5i40irsB6wN0unFMOc7/1nZk6Dj5ZYJp
s73rSSn0Z6TCVa+UIcRvZRBNAD2WSCkY21LyWTgBJ6wT01RRFj/Y5Gz6iSj/14XpjVYdBQTbf4eb
l4Z+EhjF1YBpnTXx6k5xFlTcQzMMMRAlo4fCmkoGWvqFBTrD0wxrZhToyQS9EglWdDvM/SVlPDu2
LEJ55qsraAKnYNQCw664jR4L3KWLfpDk+jGc5KJqb5iGmxDsu7icItwaia4ndio8X9y7v427gpNf
WCmkHaiGgyz2ZxmrS0F5h4miKidhUuLFGE3E7OeHxs5jGht6Ce+iaUVhh8RYcVhonQMMXJCKhr+T
VB0NUX4fLdS9Y3EGd8MR1KAdPWTzBBhDO5WwYoBPo3uyoO48De83ismEjUAVlMzBMTDb1ewIgp23
P0Go022LYScHSCrszofrf0wSKIRupaSFe6f8aCu6RiSp0pz/rY4yoTHSaxBjOMu8XcD0VaNpIwMZ
3L66D9fz24IvpqFyCMTla8/hE0wEiuE3qAKC0OVE+8RI1PxdcvWXKNKjQek4xG5DMGm0gCgJ8sJ8
uei+WkJ+OZ0ESHrrrTytnO/MeDOMCyBeL/Lqw1+lBFpBi4ahmyGWYUqke8MdULAxzOcBz4Vov0zF
F0V+HOFn63DpMoIvS4Wf8z5XKgoB0iuzCUplglUCKUV0i3Zg5PIde8KZOsQ2KFOgqoKhQMwqveH4
hqTXBiSAesdLnA1HumVsnSETbc71e2q0H7/CjqDTK3G1FJCA3zO78E1r+g8/ra8EpgexVrOUQRSb
Bk23znEcl7Eyg4VjArPRwLUE3fSpd8tvX7WN85P/vit0rtW6QmqrvGgPGiOW2r1goIvKn8JtYu31
2XwrmHoKbuIvqLvdVWA8jQjtpZJztxRNh1CJ0raPyDoDwc2SJp1AQ544KHosdZKtUsJaVsIyABUl
3Zk9ckoBVS5lMW/U8bWbP5bH1Md1zETMAnSG7fEYTyRQwrGHQVXhgph2ERT3DCFXR+Po8eBI/z8S
VhWspURunf58w0IMoMnDyGtHWzESP45itmFFkIcaD/vzPyMVHyb3UzIQoRMF6E7yWKu+U+kV7Pwq
rZZyKAB+X5wv6zfbSLCK8oKYvOp9kEYn4teZ9AgA0cxWm7suAMiEeVbhD7oEGJhHewEG/8F4VGjF
dB680sIPXr11V73VKbtGylFs5KPKQo2xqbxekuCJxfxCq8yVxkm3uzhukCTTzfwh1bnlNfWO3090
Df3RkSG9pZmodV5OYqvVnFZM9MvaHDhiplE/tp8ippjOgPW0l7W6d7w445vGj2G0l5hkF0xYgqG1
05hY9jqYdfM16ta7jnxmANvfc/MzU6g1bX5hx9SryfO8cEThbGZyIV3zqEihKFZQJlja7MXdyXFu
sWw2Cr5RFVejUWrkvsZAUmpoASVHleV56vPnzyoNZ57WTz6VE6DAfFmD5kWXym0+u9qUn+oWBL2y
iqDOJ0ci8jPn1aJgdGKwNHkauXHftzbqMkq0+Bxbyj0xBT03/NcPgfEzeay93xEblGpupZCDcKQP
3O+9PkJCHMIKNwRdVRb+xgMHJHqzHPVPZJfTOK3R0RJoXFKhB453f49mtSjgn9Ih9arNPehUz4dm
v+A5ERyzff9WGmXWth1Y4NRPyTu0Or5mBfJnUNrn9dKtwcm546EmL/IT7Cpj2v3UoBs2E1FGUMSi
tqT7IjK+LMShQs98Z3MC+Hry50ilKYVJVVALMCr9fo4nQAqpfKWqftmQH556X5BC22kWrrFDtZxg
zyaBkvNOpuVcq4ezAPuE90FoA1CW2DJneNVbgEH9tn5Y5McUWpa5vTq3671u8jRFbPddWKeOxrTz
fS78acOl58R50QY27EoMHgwe0RKgLNupeVGjO4gt6QqhjcK6T4piz9lMHYV61oFaXp4p/DFN7VrK
2zkUymnFCw1YGo7P051m0KWj1BeEFD+vTwOj+F6o13RDyhA5i3z3wqfpMiiKDhGxB7w3RWFRUD7E
5H+7gTYgtymNLj5aENbkBoAM41Io6phwrE2tJg9Y0lqfzvWjVL0H1cPiaXb3duw2KqJ05c3tKGFx
8Y+cP0oct2DD/6S6RPGe6DhdMmA0kTa9y8T+x1QonpZlyANED4znFaSifwCzw/5VM4UuR/PMvAQl
dL6wQ15ZciW2i0VkxcUNkJHivOFADMBw76hKbomh88FITsZSh4D9x4KmvrlJf22kPdlNnDK9yYu3
MANz4n1b6lM+nGYvmjdiUFi2wNkU8Vvspklno4XUg0LnAvqBiEu5/oN4JgguD8W3L9DKIWp3Y6jJ
v46efR0f0gjz6Yx5y3YC3Eb5KTgGVV6X9pyMVJugbOPOQyuU5oZc+7INDUPLmMw9ja62oSh5CJTk
aZtw5fLsRtpP/ZrHZ6uBrG1wEtKKZdk46jO89pp/CaLdYvwBL/mnf6O7qSqN57o3kqvRHIIjJG83
W+iWX7fmln1LKF4mrNpDarBEKd2kAWlwrObWAL0FlbF1eyXm8DgufveQzlyMZAl3dchWEb3UeGnK
LYX6lSYM18u8oCO8CJ9vQ8gjLfWaiWr7X9jGKWLgLL6ehyUO87Mtc+ECXLMSYXv3kMFtKKqxM+7X
shdYvJ4b2187DEXYPOtvQUpesAi225JWdEd4UhHfw72XzJpv035Giv5lrhDTUjTBWBHKhNxXBnfK
3dw7TrxViULcAi/oDl0wsWri8SPqBUfsY/kKCvAOc1vkQMUdvDS1MFVg73LbF8Xfjw07udnOknKR
A9cYmb6+IyIQg2IVQFMxyIb/GIwH1a07q9txhuK+PHEwpeDXmVikW0u02lNwn1C/NsrT4XAX8wKE
3vf3nc4gQbCT8p+/8GczwfP558OQmhIQ6vJhQqnvZ2bkXscsTEGOqPtD4GRJlS/J6j/sngi8A4I7
QzHdUs4d2qs103vmoo2OsmEGBHtvvWBwQQ1Bavx9BFn+Sqieehpqb7El01IyhRlLEgEMbhi+pZ7Q
iRqZMnW7MsjJciBIiau8yOMQ8xDD+5J/vPkLTG0SzcodSUNCACqyDwihpXfGKbvpJut+4oKz3oMR
alBUt3Cyaed3zQOwTTdeUyd0M12t8/oP0KU/HVfeV2a2nmsYMdisPLtwMtrj7Lm9zuKx2UhmbfF5
sVqyoDE2PpD0PP8y0RiJpqKhGRRIy8FLrhJ/lcVmkbWc1HBu0s45SrP+J7qbPOWINPq0PAx0ibjt
XS088GgvUMJur0yEQx65esUv0oJFuK83byEYDH9kL2BlIe7aS4D5ONOnnZEtM/GnjxY/epX9lUuc
ck/1U32kET4rMeKcBtbCr1PljCkQIbib2c8wjxrOYpHIhAyzIQI4fAZGW7CeabMZb7JffO5gp9TF
hMILq8kIWZQWESGXz60P75+NpuXrEPPKX82qvWujf/zZwAX4W42Kmh4N15sUS3m5XKvxLmcJKbfV
UJmzgaVTeiexSBMZ2Ezc8x7uuWtsJdFwRD+N0m989DSdN3YSw0y/icSzLtWNoFrYkhopWDXhgYjr
hMx84s46EcAiI+jJPtNa4Mk/hAf/dKRL/A64Svp8O8RkshtQa04ZC5Rj6JiW2aO08OLhyapQ6RjH
a7fJdDQDWB4HkGHQ99avtOxeBeBMvlpIZXnddz6Hp28x1Bwbphbr0vOeyZBGB14vxektu+uoYWY3
75cbdETiM/tHn+7z42+RBI8JZO1wHziGnMPnV7AAusA81P4cHPH1/Oi5TcJPcI56V9nTlWvMrT4v
BDi+zUveWDtlDXCfcaBUfxukMcD5Pk+gX0sfOJwxXQhOs0wuqrTSjOE0XIC9LJWLAevcmvcmTaut
ICzbJRB2GwhQCbgWuJs+RV2Id1LuBUrG38luTeTS9qIGTi/aOQ3ngqi/9U7EOyEuAAwcVeTV9lm6
xzt4AEVWKLbRQ35FAzVOCFhIqeA8m1WdqUZRvVWpGvBTQIaRHUyXoap6fubRV5FBeOAYOAef312J
JlOo6ToGJ1T7BDv/ywngVx/SSAJz0ntkxsg5ma2Q0+zlTdRHClfWdCkZ1zJGBYYthAd060JMzea+
c8HENZoKOrtw0akeNbsTF9CT4tYqHYHwycUDcU5KSrCS4gQIaItMUpgMB3mYCViXTCk6hJ9DCOBu
MmVneIELJiUgISGQ/4DtbFZfl3Y6gxqxuOaYoAV2K3aa+HMVdmJTg9TGLuOTZ1PeDZoywVOKRbu7
ibt2On0euBK+uyprNFY/mXwIjKqHvntuJaxnEio0gDop9UubDOLtTdVbBohvb+T/K8v+LPchZcgt
4sff9DPb4xb/yvlvpENg6BHjBM6LXKosqf9FDfaOK9pTFV7qEOU8awmTNZiojI6/SBQjvysBNj5x
ZKMQJbXuzdXRw5nLm8cmUXw4i+5vbqYHpjbJ/Xu/S+7sHugOs+RR63YHkhsfQawIe6PW2jkgorQC
Y4IJZYIlusm93GW1CDnCs3FJa/6kWRLsrNeCsTuS30hf7lA14oWMlcpw5vjjy834zShYl7wnUHqX
+xrD6UOo6zdinCsPzDGXxSNhKbiYG/TUSkNzVBR5ZVZu5R0fikxQnTeMNeyrKbdwlLgxbe688R56
miGdMNLUY+EiIDqVCZRgIeSwQhtMyzOedmeM9TpAUTSSkO/zhZ3fdfAevun2P2vygqI/+ErkIBK5
859k9Ras2xY3gcl466W5DTtpiX3I8XRJ6oFrC2vrDeOMczCKkXbeUc74idCF0kdE6IzkQ1jSkYXe
pjbzh1N+Rs5C3V/dWy83iyBadrx5MOXcog1tkmckzDYxngihrHmUce6WmDRAzvzzgr36xkDfCYwV
PGNZwUXMdGEO8WmMLzK7sN0TySdO7zRW0lJwHFSuo3LA6dKN6RlW74TqbXBvBvk3o13k8JDNfJAV
KkVzrazUtW5GOsojoZI9v8shf/caR4M1egYzI+G5kWC7BK+SIx0vPBttAGIjqbe//CT1jg3Q6oqB
YT7haIecjt6rFYawQvvojqnx0ElEjy26B8ukL5oRkBo3oWyWzxhQPM/xWDk0Htu29WgOK59s/LTC
0o8zs6phM7bRU6NWxDOoTZZimbLyjcOPUKft+NlUN817EPI/JX+SqUQ24Ajhusbx7FtNuVNacBqG
YxwtBoKCWmAAK6xCs3NtvoV4eGS3fjIaM4Y1SHWvXIUJjd8e2s2+cg4MjfXNddMIc5ki3FNxfg2f
QMcGcpyurD1IhLnI2d2wetWZvKg2jq2uvQHKL/015lgu5KeQNpOvj08wIVX1k4UifKUF/gQTHfCY
mQjbLtu31db4yNPbROBAOjiYJwtNGWKFNG1pWStr1Dh4gHn3ebEexh+Cv/luYoNrNrR6w0XijQBb
wUtDTbe7dSryHpae2hXK1S4tfg0ZwhzszvRudzP2OnM0DjLVvKJeBWYmmNiLXyIdIU1os9TVjo9m
uhn1V6A706H5wO3wJgTp0Fdv6JH57YChqYifhmJhe0AXwDa/5mhUnmrWSI6KgJXOZKBpdgZjKYCT
pkJeOL8LoDGphkWwfP5cLtZXz0jMZysnku9IsdwwbIQ5lzlD+CQF6A+kmTS8Y/CM6tfEuTcB9wD3
mCUnWIy4jXY+nP+iGVe09+/yV1VBXDsF5rUEQ4MX7zOwyAyBeeVXTrQgQ8urr35hvlFj7o9Td81d
jNZZp/kR6RT/rUN8pKW9kCstZWq/HWTySwl1x1FVZ7Qk0dRymOFKR6SR3RYMHIWPPt37PNdd3ieC
O+EAb61VdZ7cXpjsg8ljPPKSKBHaL/vuqGVPKK1UybRyVj5iIcW8QLpTMeTuKge2CubNt2TzwdnE
k2GkAaqEPCd5p3pwANvG1NcgxzEw12bGLHxUW+p1YH1lZMBWlAaxV+ZsQ6RxYUUDdYMTH54F0bG8
q/+wNYetDWyD3JLI0hdqJrTFc3uFfaKnTWNONdw6l6INbxk9cqKBS2jo+43q5r9hSz2orkA9dR8S
8ZPIiIfdLv5JWXamxl4jWpCFEJfE8raW8t4j1duInZQzvBcJi6R9ksVh21Ry8DaD1jzjiKuZMYky
3GuYD37oR4YJcFOxa462RY98TU53Yx5iOS6tH23GUfKq3NDrc8mbmoF2zQT6/3MyAX3bnXCscVi/
Mz77nR/IL5s0Jss9y7xHQtoH6aUYMCeGohibM2LSXodd7vW/Gc6Tj4vb7UNsECp5N3LlCojXHU8e
4qMlhQyAgUbtFrQDtdbTYOeY4v0kh+FsfMRGd3ORt6mDbQ0B0tW85mB+bDeX1uocVAVn9B+iuS+r
ZslD/s6X+wTE9uiDVtVtwru7ciUdVal8FN9fkXw8F+gbSXl1pLfgdy05r8kHOr5CLu/t3GvZedvG
yiLMvFSiFVGBQR09egCX5AsWbGvZGwaK6C8vAgZ2/HNkctb+vFzrhjO4qRbXdObSIUOW2d7vW5Bg
qrZrLMKx6T0UoOxLAVP8sdyleRmT2yVFB4gguLGDyEt9foY7squwy2dnTHWS7pKT7gkSqnTZVBFI
tayyTqifsdltKubvE0ZtG+A/7NanrG2NPDqRw46RBQ1LH7RlKpfni+m/7eaINxtQohGVSqpmQ0uz
mZ2iJAvIrrv9n33dsj/l5/7dYFJ4gkRgnYZUuKQzRpVVqUcWatEwuA0jeAwvgF8K32jVkWXISj/5
X1y5/VOg52j1GAKlbcltb4p2mWMpBUjwhYisdgvXgHX294I7QQJg9nXkxRJLwLf+ErOA8XpFznS+
a0nXJgtfWLmAv8ljw3bjQbpAoF6mkn3/OqhT1J9mc73YPZYeXPb29LbmF8RfAdVIxJBuyQNsi7KH
OM7B9slvzVTg1g6XDKFoDoty280ynRyf+wOvQU4Ahy3p2InqywtcD1feVPWq6e8w38hTWxqxa/da
ID3lflzFud9BL/7vIskLyVQEy9kAeg3wirNMUrV2HC5/ZxMq8au3JibdR+MFEI69EvrrQW0okHOL
vYy1qZXGKPG2mhV50+F4pRuKX8N0pVU5G+yW4UpquDVLyeBAJLeyk/OWuM1NllghO0l22ur8uXEv
osJcdVHCvrPmiR1j1wrVUPXEW5pJVMnBCCbb7eB0tAOwPeabxhyMBQf1r/n1XGYLl0ICRQUgoG8l
eoDqSeP/885t6RZGhg6JWv8YbaPbTFTIgLLtpQ/jvBk7w/6t9OZQYEfIGq8ipIBu/zDkU+78UdHv
GaZzbFoQqyE6WRYDDzotx1SMSdsRilM7Ywhrp6kp1o9SaAJzIFH/rO0qV4loYWaa8Fr+ti61txcZ
6Zfu7JPnugz1uFTNoE7lRKfRUh7PIJh69q/sqKiMC2IoeUsq/s6HG4vo9hauBJ9aASvdOrOhr1u1
bPeIROR0ZqObDouSvh5bcm3sDEiiQSkO6p2Y/yzXQAzEWiC7qWqK7RIMeMrJ/b5nOx8XJNKf9NUz
+885jpdkTigvdWdutU2GlZeR4IJofeyjG352VVsXLF7mp+IdNTa3jz2oMlbPbKQFSoYBYUitI1Nm
/ognBNs7YGcFjvFBTllm7L7chnI5GQ35gA/g2HwWonqCQX0pH+fONAjMOgcq8ha6cNQGJAecP/m8
PEjtOexquY9yVzZvq7YZ1X73XSz+LIv5MCjKk3Q0Ot8V97fdMpZwLckj1FlK+rv0pY1A7USGFVda
BjtlK/1q/ks41cvDdN41JoFCvh7CtjJjeAOB73xkWIh1V/D/VMDN7TvZ0ncVFOmu147kBK9EOr2m
y2DINZFAA9EQ/Q2Vx4UC55IuW9yWW8eMuCyVFQaEo5Ss06hX1aUqQS4V+PEn0WZvUqbyaN3J0AuZ
tF+yzR5SDBrhrdowkKuypCQSh+Ys4qbxeU67zy4XFLk8y1RbyZrHwOBAnVXiovMcVa1y/APsn6Zt
y6liquhIez2eOY6d3UvK5axOjdQYOtFuMMFC9bDC1o2MvYIwt1le5DbS6xXkX7WUX5DD+1uhr618
dJzCbbOApM5UCATGHJ2izSMrJNWkxNdqyYXAkLggCWg51/PP2lVKIT0feqoGKBOY/nohLPNS0GYl
Z7CnfBOUVMwzrrKEHGbHygd5yLcn2HpCO2vyk85QUCQMmaCBJE4wnOke4K8ssgh2RGw1Epy8khqM
C6CpNgT23G+3/SWH5Uk3506ihZYBmKLe9SwnQJHwqwFAuqJWiGhYYKs/gB4RJZ2ZrwuFHXX0qIv+
MQ+d9XBk5AutsI2nPvvZX4e4V6WsB0EdSCz3v7rm/FksVk0fjW5xX/UVQeqe3kPaVmbfLdWprf/K
IDSpF7fRTk8srVnc8gs+J5waZwump0t2Fk/ASHgweiVT6mteUEL4VeYH03dkEaY6YU2+JTQHONQE
LnW+myufiODo2CsMTOaLrHvta1Q6hQR2nAIaSFC3TYNIQ+siV/qsbrTbfJIV+2dCH0mtRv3NOYo7
8ahyTu0ptJBuu893q3nlal3K35Bokd0myzoSWPGbjbIk+1SwnXC1KNRrLO4QZ5TF6d1ZLu+PPxiy
16RlR2b+BUEGkpL9Wnn/82HLJ1L8M3DP+Iq7pwgJn4CSehoyQcQKEa7iENDy7kC2OtC+XcD3hhQs
LX2ScI4PZEHo7LsmXiNv1wZU+i8++ROgwaKuytSq267gT44bhPGWF93z77jm98S7XtZIGTIcs9/d
Czt90K6mreolp+FrleLfzHmOpzCNLq9hFyav3Qcz8QYup2yYsQTa5/I2wZsDhXRluO4YR2sz7m5k
bIgJwmYK6iLs6iDuV1QA6z/CkA0GZfQW084K03GOtok6YcbiHxEbEXHWdW2SlKmFV9i0a0DioV4q
wXiqM377dLfELcdTl7ZLMMb7Hkrw8X4csvkgNbv5TswoO/Hi5HUonkE574Gl/pbOAqyTAdJnQGRO
++0NERDB2PZec8bJdR0BDFYDCIeVDKvkuh/+mY+/QngDzvtXBykaZ4W349cAj9quKbTigelb1sh3
8A4itmGPDJO3z1M7YoK0p2d+8SwEwcTadiPEdkysNvbx1clSRw7S6um12QKbDNiQo4UW2WkqDbvl
wKOFFCArQHAZme3l5O7Ny/tFArI3ZLd/TOsifHoyPUmciFzMqb2hDjZRp33hPxGyYdZnM6QVj2yI
dLhvn45tHYtnhLuBIG2uZumrzYFoGm6wbNOy7THb21kBdc+Bdao/ux/VHIUvzJmyg1rhhOs0SGwc
mjQ+/G7mLvCHPpSzndLuzEHg90qtBTgxjsqTw88Ga+/g6gx6wn0AGXWBP/4H3xmrjjOfMa9PJ4D2
P03ejAIbyKqzjEsKjBCZRz+UOzHhTlLQvgXdjUskERS+vH3vN9rTzOd6JAyHcVASTZXUdeFn4XUa
rYcPyZII9BPLGA8ly5+z1dyFHOawFEmnWQWXGfkPWVQG+MNe5Hp3QwptnqS7GJwSR+mcVNNneO3x
RqgXHqe7U7S2hy3ZISwef9WljHQr+zyhLGec+TS4AE2IVtyM+PJC5FMiVRvmy1SwxFuKemT5aq9t
2h8mGUXO0ZzHYtu09apgt/SROD4Ug15duITxqRDfDM1M3aWlFmeYO5pxIAmtkLtg2imrSHaxsVYb
+KvUGf7ux3z8xLk3kW7hjxB3fYCniIfrGvE4JYJ0oc8Am915qEb79DOji5sTi0wkCoRQ6KRll8zj
uK84fDEH0zNXBUEcklzde7goholpSqCpq6GxLHxdEZrB3h2esaZoCdsF0Gmd1qL8g7WcKuclirbl
EApKFyW9lzVASm9oZFCnwJZ2DWt/aVc4ccXmdpX54K4B6fxlBK7FtpUOtvAdHD8V0na+VZqaIXFU
8cMncvJ8AtyM8fcPU6290+VkvAR3bZHjhSDIYcZhK7S5HO9m+AGVK9Uuod0rSJn2EuOvE0IcmVAs
LzYigq/YBU4FOdgC5JWMnuh/9KPmyyWUCI1f/JX/51VpCYq+PuEaGwIkNuibWwtVxrzVHvv8C2tB
otlly30rlcVE0R5nwQLQ5X7drxz6TvkW870QQlyjiK6p6ckILob8MgpkhR6uCgb12F/gZNT2+uXJ
wpQru2SRKrTpqI1oM4kJFhSkES9PsyD/SBtXLR3LbHQXt79DMiiX9D8UXz3m6HXQLe/owAQpdgxW
Ooii9lmBIB7b7hINQOuUQ2Mb73V5UP8Oa7Kvy4C7/fKTwVjlSymIdYzKhqdeXTfHqvcxQUIm2cx2
jiBAQ3KjKnga9jngtEk3hvd4mknq65cXQOJznu5g5CXm6DMVUiR2cCDQ/XGeWtDTmU1Ga1qQrOh7
qIYtrjP8xO4wutu/SW7MvgriaT1bJjnicC1KHYX/ihd+oNab0rs8vcUBB4JzRxR0905xmWXkRc3D
Klyn7aAi20hCHGEUBU+0VJ8Ch8juyRiqaWb0H1vIKTnBplM/51Ta97cdktdP4P1+gomJ7b4Op3WC
XEOhETr/bSzBXuaekWFZ3NC9T9S89rd+MxEwMNebQBpppRzYqcaIxD4EIKaPCnUgxRIa/aIdPVpX
yTsfbWWLaFxL4awiZWZvxVkpRtv7W/SkzDqG42Kr+yNnD2/WQZYExMNcwJg5RpNjALtB17brF05O
CEGSz7hrxAwCTDh6CzCM3vishhel7zejsWHtA8+Z7Y/vf+YPxWFvyXrJnMxX9ceRrGagLpRJO8vv
vxUGF/fEouc42BogytQkUzfGRAHmZGOZsISm4+1bT2ZPPKDvhCJXWkSXX/MUvyarfQWrMgF/mL9W
3QrSmM/MvSlx43K/uat+TXTkLHYOhI+QEhV/9fIrDXstaOHm0zBmEzgKqWJpUZaYYcyKRUePrhDe
VBi7GIb35PgVtFF1AhizLe6T9xuGsKa1eF6fXsLuMebCGrV7ENDWEqfa/f+HVW8mGZ+2RD+j4jeN
VVQElq29bt33V8/9vjnQwk3X3R+jOkZtUDYuhrasJgRFkkYPy/PWVTYeDgZBhHGZKLWjJvvz829q
gLiB9we0X5d7DdvcbPHK2wI6gxLbFeS+/TkGtBOb25G8orflTa02nhxL7huZliVX3GCqXpb8ku7/
t5n2EMEFNp780gRikekQhK07YrmRCS7ZCEJunwhMCS9yhJ2kmtZoVR6GMGQhUZjcSK0Yl7beIrXD
4CVbbXUr6MMFWEmS02BsH93OX3llwnYdE7HpA4CiuKlpQh/YfFZ9LB3qAy83zwBtx9Nxa1RBdovz
6cuPiXG8BZPV10YmMkoTRZuPzFu7TnP5dcBlhiTxCaEcVpShmZj4B8+38tfC+A00FlUnPdjLcFHS
vnHDE83m60aXEyAuUt1q4tuhi6xKtmYgg7n4yEfat7c/vUVe0/ZHa1oZWsee9oleDYwHrIKvHeZJ
qeUVC78I8K2tvR+fi0Q3htzew/3ITtXjKFbj2i9gjaIDT9IprYNpZQGQuvxM1JbviRhr3rqtl8AN
6/lbCtz/PJnXKamn/VxvbMCupmcSHMu7LvNrn+99TXZSCRcDzRLcRgOcNapBqmqjmw2Vqp7dMvYn
XznRq2mBLdpLdx3TD0U7m6H60GJ3yAZaRV2m4Dys3aLb6JTCpeNnfgWW+AUqDc6rBU5TEqhTZzHH
qG/mwfTjwfThqNl7i/t5pOUDhyz9fhCrDckuKxtPv1UrdjSwPEem6qCm+jOyQql8BLaUekBAY7RB
ZIYf8OxKhG8PXyXP8IRuZmOWfer02mzF/mCxBqoy+vlzfTDkcRpASW6VGDiVhSROAKnVjqttVtqj
BsMveeziq3v0rOJNC5FZs/q6pf7AQrHiOxipx49knwUseXCGlxekdCeUg8akfRFEBO3YpX9ItA6O
Ff2byEgQazg8ZhB2Sq0cpylMwNP7EFxeVBpKrPa/A18g6XakWSJWzldgGDe0om/7kC6/UjGPw1tk
ZCKa7cilZW7EW9ND5hOaIu2814TR5WRzOSvpwMSVVlj3L2m/JmnebOSTFm5MOzjyPPLEaZvur8f0
bIyYFQHQVFqfYNy3EKpBQbw8mvQQS9xjU3uhB6TLB88LirMd0NDWSbv8BwnH1hNAaVrK26FH0Li+
AL6/6Wo/MikZezV9lPy/rg5hQgQ7bOYHd9MjOr4ZKg3lLZ92wqrVpID7JuqI0UB0kV1vK1+V1WGa
oV8M08p3X+V+8l/a+ldyROzafrs+JqO6/zc1CfUreZLDFsqaydqiHMooegIrLhhGRuMvvELVFFUb
il4pa1Lwu/R2pAFGt7vfmH3Ob28X/ALuNG4RWO/TeHJkmtHoJbeLvtTLYnNqgI1RglrkS9B10Cuy
d2BgdeaI6ddKZ48rSXnwhG7/utjOcdOko5gAwI1G8K/NAXWkNfjL+nLs15a5FTSjBmEU3Lhsr+D/
ep4QP0H93EeY/lh3ydcP36+hvKNU6lHTMrM3dde6wFVhS4KTdtgB7RPIMth9kHoijBHzMTz12Q3F
sQJ4MEr/5DOA585+zfknCE2B7HWqy4CdcbMUmkzgNVBAIrAnu82cNfmR4GBRRdsnCW5lXvN+9FVD
/v09D5mlKjlkxIQr2T+fVSlLpR/ksqYDmUenVakjZ1c0FOOItjYE4OXJ/rX+3YtVUZZNq3Ply8H+
IB+7Dz084Ldk8frd8cucC0LKU7zqQNThoCr6VWKhIgd7bX8ry2ZSOn1bCRtMEcY+Eve74N8Kl5Ad
oQ1bz5Hg1zrQwYakk7e5HPKJDJFiaTR750Lgjh6lgtYSrkt2NwhdrGV3iLnzifAgNpRVufk2H/GM
tca2LjSNSawt2KvnM1eFTIy9Ldm3q2AAJ/lqrKtH0R34OYcram6t76Fp1KyXxTZsZdfEPORLk0T9
GlOu6EuEoul+/+vRxi8HXP2oh7Avd9nVoqCm8BfOqD1eLBDQ0ZIEK2YDcEmPrkQC0Su+hsqByYw6
FcExynSN5Ps8kwQMcEC0uemNePp500z/5a0Zbc1Y/VatZ9G1LAJ0/Hws5CXkAdX9Q76R3uv91EfG
3qE5BQJ6zgWm4kxSEJGobxCsnh6dG48h6wHKpC9/Mr4L4NMWeKU9nmfdhC8Omv4JLV8yzEqcJWWi
hHgOqOJfjdXYSfSI2oKMMujnfm8FjZ9C/QmSNLBC5rgZ6nyRcBCKnzZ/BlUUVNhNXHRXyLfnPo/Y
WZnw+Haj2DDVFWkdazbc8Sg0bkgoanfRfr3Z0SfQ2BDy9E84jT47o5lauvCXF/t3t5Ic94asPcZL
mRnNJAOfaxR7IlA2CJBUuXdtosip6pMGLiyaTLoYiGC9/dKF8XQSNMsEYOH4opQSaCoU9+ozb0TY
5e1z2DQp1cP4Dys9dTG4dzarxn+K5hm8y0rxqUToCfzek0pUqUgoBN0HwqO45cK/43AOB3lWgbOo
zmR+PWikscrVR12Q5lpSx9ayDe1XZDTsFh+He4Z4rTnp6tIsnwsEv8oVGK2PxXn78e0qZuLKu9Cc
r1YY7jYe/+GR/NCmZLYJ+XWuACSCNuO8+/wuRbrOFb8173LwbIOnDWFhtile5YSr83UdOJVo+d4Q
i+QGv8YFRuWu0GqowfZmhBPDQV1uDVFNkGbuSIx+I9mdoBU1SXVfpk9JEIIRwcQ4k/LO/ch68+OJ
fdXbfy6v4LldYX3BOVEwswFgkHU68rZApxY3OGl1VzhN3hf9lXLrMoCY5CB2l6aE2RN5YgzerJY0
f+dCHwv6OYbpvh/Zh6hfR3Fu07LNMIduuvEzoQaPrA2WYUFuzWQRKPMZWu4/HCJFWetZWcJ84O87
Hb3a8UU0868C/VgtS/YalJD4BRxK1YsC3qC+wpVS75N/L3OPjD8whCxlM5DuhBJuEMzFTdZXh1OK
kpg1ePeenJcq9PLqAxRPmYJv8EO9RmC81T429zyJr6ha7f458yBy7Fd1gkALEz6zXVbe592TROvA
zVmp0JfGWLKMUllMy+5bhnA4f0hJOBP35QKwoCRhqPRqaQgVSHYI0x1Gi7iazrWbJzafs/SQATrX
KRWNgLTpcJ1Ry2AruzbaWE08LLRzZE9oWNLMMq2v0lJ+QDIPxb0O8jLmxx7Lcb6bWGjbb2w50RZe
WPDCOsZL21NKuo9zfZo9TjE57++2w73cN2XKbRvpCOm0LMIJ1Y3CkhKKr9oLVsdVps+usT4vACYA
w7Fng0CAlUsrFJMUojNTo/tCeiQDpKG5j7iDNFPNKe/sRuNRYTDPGS+4qiIwyCtqrSxI1WUbbgWR
bkRzAWnO9GgjUJTeZY1MqLZxKf/cjub4ZEMS9DxQjFtLiMIeZbo6NI217fkE7uudD7xyXKAZRNnS
f23qEiz9K3JV6FLB+v1DiMK121uJUMDAJlLkzu74gIAqnoVmtlB2TxMmnA76jcvtcVhN32vW4E97
zA7BD1zIyNgOzRffBUk2P5IfV4S1FFcseuip/7Q3S+u4At49LQYIunR/14eWnTGGLahCgL+ogAB0
Q1RazFryMgTP29UpMjeblZm2vGLiKDFS8Yr6GEvXRtpqTU2JvCjjq0yR4dRM2pq92cJLk9Etk6JL
/3PPswdmeNlOXJ2x/udiwj125Nz+q9tYF+JQkMz5z3QvSMh10j/5I/S7Gth8ww0LqXmiao4TWsTz
DpYk4/vyybxWalheITZMcqkxUaaQTw5u9PvuFeVl9b/VrOi2UD7a1BzWD/OP26CU6PBx6ODOi+SQ
aW3Xe4CQYmF5cQklV0i+STIukVFQItrWQKfsjaaucVkoXL/OLFwMDGhd2z6uusSsJFo90YEqr9Zb
4s4xFNbE7rClfleMoPDrtzQaRawKKDRlTYcHMuXuroPslMFhQbiVG5XtmaaRY6RQx9+jUD57RGWw
0D4csZKSFVpAQ7d1YJUBT1n+LjzhraMWWKEU7MpDm2kb9QrE7M+6vLvB7BmyrE6931nHfXcGwBpp
VGlBJY3lseATLBXvawsllxaf5f+R6qAVUTd0jNESSPuefGowf1lUPjpgJ56o41Pz3XUHOxGhFcGh
+ebZp9aj2sdksNcS9bqaXjSIIL2QFoBL1i3F4bc9FlI7Q9oI6Edxnt+sF6O8Fclwndw3Nt2o2oQl
1ZpaDHTf+gM0mYTx/Hyx8UG8FACD2r7u40yvmSLl//qIl9bzLs5rRWD4sEZ71uQFl2bZ2qxnOMw6
ApsPRLUjbWXvesvplEDVgePIDdP8FPLIIZZLJvymIvfNJzGKk/sCKfK3cXFr0WTRWAvYno4/LpPc
6hquTu7w2MH07LKYdwuQaE8/iDimVGfzZDDlHqskn+Ts5oFRN1+YwYYJsNoQSuigmR7JNooddtAZ
WVn25OhHQzV7mxgrRnD5Bh/Adi4/BTqXtDYjfj5EpFFC2ukvQnAuLH9fHYx+0Y5COXollAGcC+MG
Xx6x/yj667RiaflLiWl1uzgMAvojrjcqkh4e14z2/CPATdbekhcVFiN0UF68BWUkKgJsdpJlS3zM
AM3e29Wl+K/EoZN3YpuaCWZGsBVFYsvQmAkKncnMexpLILvJPReqgWrNqsKTetzeOuG/h+fL//zt
ZDSRr01pVXLrFaAmxO4k1v1dhsF0H1dYfj7SuUpP3W+Saol9Y7FOyPQOuplFOyGTuEzuhHKT0HrC
fLnJB9D0fR10qi1YSH4YKWFQ3A1G5DxaRAZ+rb/RS+ryBZo8vqIkwYdulbbqvNfG3DNsg5ZXuObT
oNfHRwiXFtGGyXi+ykx99Ccx6Cy7pAF2Ps3jRo8JD2wJXGdLGrTTAdof8stTRWuIXIo9xKT0qBXE
Zt124iGPwz0PuVBB7mbQ9/BK6wb4Bts1kBr0MzQuV7k0YjEDxKD+xa0gIM7KXMZoaH6PYqCM8OQz
1b3UuxulihAXNceOZVyl0ui72s9NhGtj3z6IZOY24eW5y1c1boIrhkJVGwhvQQT9BT0rKkQx5VNt
uQSL2at8P2aQfNKRMVX0LKDWn6zzRlJf/EP83L0o2eJ3UaVAG7bYOXvB2W/PaKC/6GOZQi7suPrw
oNiu6VLEYIs0p7YvTfygqqWS8M6i7bapcaMHTJPM045oADab22M4NOgeMJeoDnXhBhV9HiR8YpeC
6mviXMyYTa1yBiIKpD3ocoxVTsWHPNWh4Ekb2lS2UIPw1So8sBg/cXsBpCN9LtINeWcPxYvrjzlj
26pvTLZByymcVzW0lLDg99AhlzgnrbnKRspOoP7mWFEM1ivBOVfgIX5WeuuoOFWc3Pcj6g5gsZW7
tyF3WhBxT/O+wce1uFinIGCY/A2r7T+rkx3UqakA0x0L8b5wBGR3DAhCC8DcwVYQmmVj9tz6YAg4
p6iJMvmKlGAIyANIyMMHkIJa6uMg1CfH/blQqKCEWJmZ7C8FFgEBxfwb3zz8yIyhPMXrZvjjKjak
KGHphemPs5ad31bnOES6yVBvLKl2kKda4v5JVHx2sqNVxg8RnVTcriZ31tBMHeVfu1BFd2NVSw4y
Xu+w145eJfz227NpkzSRwufbIJr0T3Q450gn2ufkhp0V197sZFVMoX0RPD5I6PYAhtZhNSWAj5h7
mRFblQ9jjlWAHl+4aW1P9b7pe2fQCjIrhBSMX7VIqXO/3YzHpdsDiOjOa0bPrumSXWSroPMUGQR9
SEhTt9gDHHBZ2UfZlKB+wM26fhhs6XoN/g2iyqgXAMDSD/nBvxTQf1zqRfotiGmTk2Qt8NUEUT4W
2Bg/rCPG7170aSUrPEw9GbS8CcbYrd7iAxWLjmQnxfa2bBrEVo5nxXuswR7NE4DNG3KwlV9ZEbwb
IgNJWBy3IBoWtTuLKo3iNHX3xWYXy28MNAM6AwKjmdfxShQZSJN5ZwTPrQn7SUApdIWrkSwKTbMi
k8/WcPGKFrIAMs+nqaPNuApTvt2rYZa6+jXnnG8teGr37vOwFpWSlnNWGoNQbfPqTP+gJmQLMc+y
CjMsQmocwZ+Ue9YkeO95IbkC/c9UUOdIpHIRznyUixZpNU3LhrWjjokdQnxV67QghiqYwWelUuN5
QJd4360V+j9mQpFnOua/ncKQLpxc6B1JgFSGmT0O99xGgdc77ADGeli/7HwO7rD54vhzVqHoaJHi
jxDiflSuPVWc3fcNQ90/NEfzJ/f4XnY05nS7ubfSGCAZlZGuk3wcXzj82Hi38MnupBJGBi8Sn8Mw
4K+RPP4s2u8L8plHCcLkvLUNRpkyguAkwGyde54r2ur+F6V73m34QcA0lQjtZAU/HPNHQHittRMh
FQTRfg+yL3m8M4ZsFYtQwgRAWQpKKwKSnUTLb2uhwIpIcVdwOxM2zmZ+gqxNDlYRA3Ak0vCQQrka
ln+MOhSO4ZU3o2a3Awy3S4Yj2vcoh0WxkkN1suMWYMeyO5sDgvDQ52LL7F9x6REJ9Dbylkaw6oSR
qFQ77oyNi3Nz4Of1/gKGGm+2/+lWq1Ke/BtFmgM/9oVeEBq799shq+iib0VbT0RKLOSrRhVy34Hh
nR0zYqDK/bjSp0zr+pmPJMk61dqU6frboNdVf2L1tW3IuAkC1J74v0q0YfxXJYRMBCwZmEmyxmUr
W5NApbUHfQ9wb1dkVy/V2PUgq9TqFOVAZmLfwo7EYnsHeUATRKsJNacW9J1uMhwHfrzNRjCmTExL
8RA0eJhYm4MNp9PLLV02TAEffN1e4Xj6HwDWSo2tl5GaDdxwXUknd7IXtffvibC587Yw3Gt6q0cB
ClbjmP/hSSxaE8c5T1heEV9307ZbS9fhVZ2GrNAPg/w6ake2JONtT5dmuXD4zhS53F3WPIp7bPRm
I0HT/RpvU8AC6vbX2p4PZLrYAghs104xvE3pFhK0JT3+0PEkfuwn10SO3LxrESjV+Ww7lxkN5BLO
dYkImZ4ZuZtDNq9yGK0bhLSKGsajUWc8jFSHTZHGeeArmmzJ6GOdxxg548KM7eu60AG3rQPXTvwB
JEvVNJylIUbMv7QN5sFjVBb0yvLKlGjqXVXMgNWYl7xztDONgdmE/D3F3otq5hsnHOG5/KwEfikJ
uun32jFdG19ZzVCfpnS8DP5I80XICVn5fCdG2inrtnlQMhtP3e2y97toQCZehCQQ7SOJn56Rv1L5
HzWLGTcL7pcBG8r67Q663SI+Wsr4HE6ZL4E7CduWR74+Ct0xfDoaEr2DEvv30BqykyMaTYK4JiNq
Tk+CQoI3sEKkUAE1Se19lG7XWQ8XisB5EJdd0JTVKFTXWPGDReOPXr4DsIdc9t16H8BcZD47+lLh
8xB+fijB6qIEDUdfOJCEMz7Lvtfs5cqR+INPHWBga47ynOrLF7+0SPMNm5PKNtBCeJdPW2xnL2wz
F4OZNu8ZjgD89Fn/0pdWrJfJlLsb39LkOxUda/HT+jQw/zqPn2hgL6Qr5IFb1De5/OVCAyid7USE
iwovzsG/1ArWNd2Q1EziwDE+/ejJrZVIA63CVRRoPQfRAwfB1e54zccWqDFkyaeTe2/HGMrmFMH9
Xxh97XbWlrW2hX1hs+orELILHPmp7QJk0MUy66nkaojQgUchjjRchyXjsZmDHNkXs/ZvQiu2tnek
/ULzqzr00+AXMQax8ho2KoZA+hI8OcAOw1x2ORH+Cr7sbk6jObIzgOGqqEdbIm3ZoBwMOOEc4wke
RTrXYLY/84CrmLnNp9cy2FquwuY5FYXD61LIUhYhYDmkaijLs94znE/eI/ko6UMQBNfdiZ3U4MBd
SknM02XMI2sA4gavtlJggOpuWvHQ68DMfp6sByjEZrGawhUCFF6ScZmGZfmeBt5Zz0kR4bXZ8REZ
yigbnfSfIIdvouIHjVeiv9e61+W+nLUfoBqdzUNfpJLYc9jAuzF9mYPHDkm7fT7mKMtNZ7VKnF3H
uDxceyW+Xfg3H3bkmZtAb7XOOACFOJJ3JIMdq2gPmRLg9gN/NHSHi1+JaimqhlSGkt2jCFW25oNR
S1Zt77/alyr4FK+sL+POjKqy/r95vVkxhAZLVSo+HPmJdi4rePYhYB3CaLAGolmDI26hPItdVoVL
0wB2cBpx4pxVZj+P40fj7UhRA7PdBIWMG6FZvJTi/uxbQemszVOtXKXoNohd/GIMr8usb2+Z6bsy
4NpDZ53Yphg8QzQWJ2MKqr669NzMhqCK21XSWjFq6C4ldfwnCz0YhmKlyVEVsRXX9RHtVHT+fDnE
NDC10cNxG1ATbHDXPyRjzla6fFm/eNYkMP3dcVqvv9ml3xnivSBrT7gZoIJtUNEuo7g3Tltr6rhB
1DBqstV2ar2Djv1ZmHwJgHrDG6yrmRVhpo2DBIKHjWlDuurhsN3oRJelzVCXNEzpZbJnjNtxVTf+
Tp6BRjtJf1fTN2ay+z0Gh9g88YEOfA7WgZOI0nKjS4aqAbF/Kc+ftaYkrJ3+mVqFIqa+88xWOe45
MMABo1DPhaSzEwRPjSMAv1497oIjKivO88sHU11rUVxPgov6Hzjvssx8XC0r8Do5fqI55NP8I831
8ByLrdUU5O09gFQCv8OfpKH+deZQU9VoC3udc3L1gdkN/EpVpMiJ9JZ/ObzpsByosr2bTmsSa/xg
AUtnnBcyayx3sxmUdTf+Eu/+B12rejXl3ADVQDpou+QzeC1dCKh2IKJFGoVD6CgjfFGbHgLIWU6i
bsDojUXV5t2H2GX3hxKVhfbsewsFbpEwT/e+ZU2Lv0hjSgWriqNhyx0FwqR/nmnVynWv4fpQaW1C
uuB+yhJBUy07ScO4ZDf277Z0EvfMg5do6qHCc0cKsZAkVzISpJt2P9BHEq2Sv2L7PUhJSAud8z2B
KKSMq36oSEqee8DFS1i4uNSs0uKOWIrCdC6uL3hmFqL34aHOSpyDn4hvuImiwChO/x017cRq1gqI
OxKHgG84MgSl7Q9K1O3IZ6N0KaNk37y2/GaMBtmP12KqUILHCpA49rJbc4OuyI1E6mhc9V1LRne7
C4s+6iYSSfqZ6Ow+XT1EPwQzgsH9DUxey1VCBHsn7ScMGaUyfcrIdPzLqnygZPNwxPqAsQ9a99Wg
2snndHzhLkDjQBSAUBbfWlzu1TZdNvIki4AwKnKz4l/R4xQiMNHAerfoLzG238O5uLaxM6cljMKf
oMu86n3LHnQOeSdQOP3M6gsg6SeLHU7QiM49QDJWTZ0vWwFhcB+5NfG0az2HxMPcfJ+xlG88t7Ue
kkLtsg0ZELhwKINRVa3z7cCRB5xYvzm5WxC2bkhqcF/eH6nW694YJwQ7qhwfBdTjbEByuK8HXcYB
ZKmz+vDmBBjEkAsTWetXbPng1Y8VwbwvcxOgqF7enpspJrr50s6wJ+MpaOp3dKThrVhlVA2LjHeE
Kvk93/AMDLayzmFIDWBhDS49xEgKGLW/sfB1D8stQyVENfApGo8wqCqaU3VlexQ4dsp4JvgZSis1
xmiondBJbQxnLeDkhNGl89CYWx7tFt8gvMWt52GdkO74i4pij1Z0dcEkdAJqu4LbR1llgEWygWKY
ebOo4pUGRxDw3ZFPj41n7MqmSyUl2dcEnTI5wYOGtz+RL8YsjDQaQ+16DSm/ro0xIME3wLGVKpJL
ghAMVaDs5sRSXCJDmhBUUcHEEvPSg9JK9Znp1O2o8uh33/JtFrWl+MAbVPVQfcErGD5acus8/CVt
fx/4qFnlrWpsWTjEjnA+qxqbCjuFEZzHq7/a9YqXEty2B9ApsPXIy2F+MLF+d4Ifa4kWMWBOiBnY
lA4bOJTWxPCeyXF9iLg6BuPUjzssZcfq4XmDDiDwTSFk+L1UL1lYXDZJKF9NoFOTpVWnPlLjhEsD
FbjLptfJMrcekB4MzNs00ABFG14XN9CuPYZ99eVzKbiaqpI3JQY0fshFuoFqxdijPpR9gSKLAun+
cOlHp6Bli4+0oihcJLELyqBqEY2lciav2Gb7ztg/Kfmadsap+zucz3BonUyY7qCokoTVYxg3q6l6
RHYbgnF/MqKmGuLABlQoIuvNEo2hKyHnSo4rgeNzqarFOa5fg329ydx2Hh7qmvi3tuK4mlWSqHmJ
Uapczxdon4VIslcsosxG7UjHvSKAnE/Tel38hAnSRZMitPXN5OQovQrHgFYkTMYLS42/kFp5Vzi8
Wg884PGJmRmm0z9FrDgzSg2mKSpgc4mErL67IN1p9sf6toDXBEXQaJOVfpFFBMVOvcgmMn0I38Nv
OOkh9dc/6pSq0VxWcFGeUdUkD71yvnFAhS9O1GD3apFsSFLRqpS2Of/jHL9JmWVRphkOWUQw6Dz+
DbuTU1nBmB0sol1QWc/nXM3amMiltSPulAXG8XRpuFZZ8xb+/99m8tS4b9qmklVPaTkVVBLDPpFX
e7l1P9FKw3zZOYBypUdG68pq9CVa0/uLzMA4FhHZTiVgnYmmQGZZKzyxsV5XpZEZSzdexKDk0vcT
qCtdVuf5/SWtbmtSQfB667RzcvTXSyUm3DkzvYDubIcbnOost9YKJu6t8o8PN3Jj/+LN9szdi7lx
Z1zF83i8BB9fDyj5331C241NtKwaGIz2e5vpcnf3on15tVo8LxLrY+BsslGQZlyXDpc+PDSQVMRJ
ObgJrc1AR+y4XkNb4IiqXqYY/m3kFhw29zhfk97TIjR1z38Cr+aHR0uor6IUC2XUr6eEFFRjXDWK
Es/OyX0n58By/F3drWCWZ5vmKYgLM6xOcmSnxmUeEWRLzksSnBYtDdiEzutOh78KPJlY3mlxLRse
fwoOxBPps6fsO9DewTdvWCFw6KDWpzh1op8RmjdJUoHqptyz0HlaJ+eGh4TTiaMXvcm/moPNstZ/
kWyxsT0pfbwvHd4nMCDnyDi8Uxn2hajwI+dpOTvsVax8pCSMUtcGWHVDRCwJR77NVLiDIUmp5EXG
bu+egDD3GxRxavddWworRjrGqjBJtXIWtkBRx2OQJiQJmHEbq6FjHr5goakFiIVYT2+3A0u0K6pc
hitR8I3AhFJmt/VECo70UR3qTwGRNPqav41UlGwYV3j8QHVl1RFEdK7suCOvEvRmqPM/Y3OD3rPa
0LaZWW/xt5RvU7frYQbgDOqNn0XWbXB98fNMWrqR36q/1wg+nxOBim1iqSkRnRNS5yeRwTd2FjFd
AXgYGiylfBzBUiwqKAtE0acYZmBZ6kSgZMqnKLj8wsU47GgdzzvGBp2RwYEePOLGRKHirB4qg5BT
UZMAo50KBP7lUbqJGuFk7hqSS+Y6UgD5MkacS+0WygDFDgLHPnowXJma+8Xjp12qF6u5YnVgv8gY
DWRPt2H+si5nakhRB3K9zD3zUc7FXHR2V4j+L6InTAgq8wnjWG00o3tkSb4ziZZRPkJzBcUm/BZe
g1H9IGTv9d6mXVuHVho0Qoz5AFGx/VunlveTDZRuG0QAPTFFQ6H1KZRfvC40O46nYsHqaThevdYT
4/HF82xSdFiFOo/bvlIopbDw2ymACxj40g+PXZrDujaW8g1JoL5YQhoV0x+wQ5gevjQSwgRuSteo
SCKe7DC4Wsud9kR/JzAtixwlvUgoE7BmxD3pvp9r9QrqiM7U1ICyls92DsqZk8sDvm0hyA/91gUE
8XD+V9q0x2DacBF7yZ+G8gXM2mF9PXjkRea2SM/ZytgYjxdrMzpljq2oUj91AYF52ZTanSEJ4upI
MNgny/K6v/Aow4MA69kixyL/TszugTSTPss+tk1K0x6d+ZAtyt9v3yEmUIulWGJkjTLJF8kT+B6M
XKrMIUa/BL0UHDC6eRpxFX6A6jBAjTghcQHuEtsZQDL1yZkJpKm2x/UPIP0aSlb2QJ+j02puP8tK
10GVv+QEX5WTKxS08iyGEUC+edVXKiApVE1+pp3pOFJ2jJqyAA8IsZY6BiRGv/BXZ/7MskVPkm22
q1/u1mMnlbnEYI0KDeOkBNq8/XHyYt7cPET5+Srm3mUsJrcr786/jwHHlrVswov8jrPT/5xfTQ4W
Lga/+6gzeaTO+Gp1TeG05qjJJ7sFf1h5RSWiWiE5mgctca5THpA7mnNHUNG8/Lj5oXswpV1w86rR
hSDDMGpKBpglZhunBDyrvFbwdySkKTBT2HbdNmxeM2T5Xmwg9CmAJ9bJfrhZ83Y12i1MqDbK3aMG
IyefclkNIm63ee/IOF/TuxD/tLerxzHYJRGJZIF600y3etst/erpCNaUMtfJc0vUEUNtttJup+Gz
qzFKoZfAdAx2Jz/RWEL6dImO/AZxyV3z+bXsIP4uSI2Kh1uUb6CJ3UCh+19cz8CW8W6fmGqNZcxd
1sqzavmSO7dE4zRcbkrfaFIBaM4KppKIHBsJRJlg8U2KDaQw3yYq3TiGBpD9OkFnnp28e9bhL3u2
ksPOEMuBplgHGEael7Kf8IuLLiMoX8WU2muIuYhNIn8q+KrH+i2BRD5jk7x6xJqI1anh/dhHE6xf
95nnA0w7t7OLchFLzhNrVRy754CZur8SUfdwFmUZ22HixY0HAGkHa3emDG6TeSKcNFSTg+8QikF7
7E5IP4JRLEmU0yjsJIFT4X2AMT3eJXfVnwbsjwSVd+bqjCg8FWyt3/XMvHesOnezURw5MS6pBSi3
yPgwzZwk+/DpQeiUYV9mzp5Qgq250KwQeJ8a8Jgv81IW1aQZV/HNFg9R2V1ovge1KH8sWJclBfEJ
ysptp9VR9lJKSXuGdQBGAOheNvoudpe3tdWp6CvLd28kgm/9uZsAfO3kKk0QSxAJz7gt4d+/HgOC
NMq4stH2U5vRuYoiu4RWUdrMFdU2PN3U0p0Ilqi2Yixdw15vxgAN3uIyxOP1ojFWdANkLb8h5ars
DToT/iUx/VL0hUUH+qozrvTu27bBKbpfSLg6k4Tw1a8s2vOeo6UY4gk6RQlOfLVGbgowr9wa5G3m
3LdToPTvx75UQqa3U8WweNHmBSzQ0ckHJaPPQmxf3phg2celgIc2VM/UaZUTjP1qKwgqxfMIBZCt
TJyO/f+2Vw473Fq5Dz97tGIeIBzhH6km2w8POxGpZ3jYYtgca0cnDxFvVmmxbUFeP6vVl2WWDKy2
jfUeooZkiA3gp5YVS8zR3siAskZ10aVWlFbT/1xcpLwwBhf8ZGdwkMBqdRHBhJsc0n8Tazcjgg5G
fmX9JHjMaSo8YaLZqbDoqbWvevqHpZdPyJj3kls00tQZY86JfP2bpOfiSsp41rUqMaVZr4qZbESU
eHgPv5zH0MUMqd1Yyxp49KaGd83ME2ZxG+iuwbSF0qrxlNGsXyxBvquBAxfRzDAC2vYF+mon8jjp
/vMcpHf3PmtypL2b2Wf9/YGuVT5wdP0ZOG/XPf65a+43Bz1ceRO396AVUFmAfmStBe147oLrzeSg
2cI0k5hnXMxgev08o4Bk9n9j4S1sNXs1BnAsqUeDqR+TWmwsERC/RdbjD30d13Ory4XfuvRqu/0K
NolOmerjOGfoRAY5ilp2KfPqchM31bfuCuGucUr44ZeG047ArB5ZERRkcuu4TvbAjtZGmv2qsaLs
itClxfLd9s1Idc4ApbpYZjZVz6gqZGEv2xQXPDPG7GpMWgmbOpMR3hryEONcHmmSO+k6zyxEPNVT
PNaI3a+Nbn9/H+P7HizVmt3Z63Lm2E4drb/nYDvpkngOnfdBrYOIGecb/o68WY+rvEIekXJ7iFQT
44yVVpN/QOBy56uE6h0Zt7UH5nH82eZzxE+5LFJ78PEbio37BArUm2mnKZtQc4zTq4Sm49udQ07L
VQN/gpz//2NIS5uZZfqrsvM2fJBYDHmSQ1oMd/jsJERphnjUGfFnk9Qfu/exI4pG72XGXSwy6Jz7
UWmH2FG3gTQkg8sQpw+NDqmqDrZTIMebnOZAhUKhZqB4OlU/Y++UabkNFVySvxRtLH1JVJBg1JF/
oJazrDDjTiY3OHNAXgKhgieZFMDCkHq3B3ypaM6qb0A7exiyj92E/jHvJtm+rtYc5i8F29Z3yXMt
iWmYcOeAGEHHkJgo7nWTwA56AcNwxxbAGQnvzi/LVYncxE8j1EXQFM0f8VI/rcKiPlZrfupRhS7I
8VQ3yr4GBlLK0NBZFEnW+pI9W0+s4xAdVVM3hcCkLpzIHIjOvyQPcTzIRom1BxyOQ+Zb5iE3771D
YABF8z3kR8D96PaEmxUXlYITanOfB0NIz8y2OpPRW6zCpu9NbRXDIar4zsRTMqqMysBG/Hodk4uU
A9u/vH9DxNqmbFgS4R/FG2r10IwzuQJFy4u5rGaOi+2FWK4JgsTySk6zSkG+t8erqxfescIp6RAW
njudOK3xU/v3nCkJFyYHj07GBFvv3nEjsoYhBn5HENYhnQilMPcxh4lsic0wSjph7EffR97Isk9l
rkFawMG5JNtAjBDP7Iiulmlc+YlUS2TJrD/4qkzyqVuM7XbvrNt04F4dBhqKezhdXk2FRWYsHY+k
Qj5gEVQrETfaG8yo9GSGaaeYZzmFdMGXb6IAkvB+I9OLr3/0Emzq1cyQJRaUSUGLE/6Jp5ritN8y
VtfxYgM6qPWj1e9BbmaXndL+REPmN6HW2CpZnbBJ87EDTQfr08jTijLsHwOTZpdv6wxCCLKsbWZN
81dvseNaKICbBKHecTA+zFNC3WmWE5LmbzBL8kMeHo5i+Ae07gHClmjc+mVOsg8uA4WV4bSQK3JK
Tg1+GKb5zSpC8uNTgZF4KcCYYoXXT3rkn8xrN3lCTKvDb0rPVPHp8U0iPZdpGGx+gctPuo3YizgF
vEuoKQ/fjHq9svfxZzwxKY8e2OfF9s4CpkNOKuJZV3hujns0xtFWGUkdFfg8Jsd5xYLT6QWayTFL
Beh+dnqqMIWLh5jEPSxUJVNpWU0rmDzgmy8D7m/1q7uUK8dVtINw10gxMMkMQQTFDYMCqIOJ/Npx
50DsToVeVcou9xJ2QCzuKCxq19+p7VfiyWiFQjkLzMApNy78YS1mPTEhtQem8O37wttmz7EN+2dg
uXevs3edUcfD/fsaLxn7YlfYDgCDl78euMh9k1R5YovJ790MrTYybD5MG02QWeG3Clkw7AFZxe4i
F190BFnGfZJSzAs6zjgHC+atxsQN88BxX+s4TldoW7Op2wQqa23pPfYw8YUqH6bHg3JP6joEhWov
4uIrQ9GXbPkocAvBzRQRih9Z8PTbyhrAOCRlLme5JgwnMjju9Pvlx9hmtEiuHXtLnjLwAPGtvXUq
Kh4QRiUuV2Y++pMVE0LoS5uMxNWgRPUDy3UPevRFZ5PO5U1EKgvtcWBb3OwKxY+jvp1Cfh3K3xbB
sMxoGwy0Bk0L/XGXedDJVONVhN10lo/hcuS1u4Lr3NK8gNMyJfLHtbwazK28zagAYydN0h7tYwBG
17tHZ4r23+SlFIWMyqwNea3rFJ8gntI6llAKWJK8NzHnmkQ9mP0HNHaYSUq0ch472RJ1FIW3FqhQ
AaF4IHxpG8qSdUmFPxQNo5FUGm6m4jKJyWo9o6be7E6PXzYxRNIDB+AWyz/ZmGorS/djGdTZaQTa
KBPgeXP2RmJB0XV1+qWEmdXlO5SVivQLECTHqnPa7vIx+dO8m7WREE97lUm1E5w9hmkblFUhe0p6
gDE2uR49n/uxmr1wVrNCItrENxtvhQ8KlCIkY30EyyNOSBk/FdxZtVht9sdky6hXD6FzwaJBvoj5
jcDampXGojoEDgApzjzUMprmE8KHINcHcnBnyJJftOxwGyQ/3EcWTsYb+uLUP/RiQIcKAfE41X2t
zRkWg+7vT8Rd1pN7wkasgNYO6gUcnaVTAij2/ct2TmqamzzXppWdgzqPeCBIc0YGEUf0IOTK7zbi
WyQ4P9nHTVtS1xoF147B5u/pI6U0OqPe18fldpxqXp9JvHNP/WTIgFeqOd6cEB7WzqceamvPT8UT
fg+M3b7rywT81VLV8ziZeOKteXPqrPLdIA2L8wJZCThR0KG6UHwha7NKFZ2CqYCZQJ7DlXFEmnTp
OTXbhhiX/mOeU3rE8ny9w9Y0eJyV8jQZlZjYQRWHuzGEOCs40LaNf/2RhQ+jD4JhtAtSOiqmu5Tx
DBlxQdbSZF8A0cPxzbyed89rQhBavOzVe03aTxEa0LDQ/YCLHYQHD0oYUNYkGYtr4cGPHCxsJiSY
h+F061Hlgu9XzbsdCKJ0Ge76NH8f8pO4oQAvZdk/lHXF+8/gSu6gpcBe5GaechzRccgN1YvyYduT
8/G1wHgYoYP8iwYwU7QeLyD/qA/+cnAW/TvclrRb4nZ0tCIOm76Yj4g2dO35WdVCGvXRMAi+9s0l
waQEJTXN3BKv6OgwUsT9xFzVyqWX7Kyq6OZSS+LFAZwG+Nm2ggCgGgJWWmIqOTk5Tfe1uyTJdW0W
IQt9k8ml2nJu12lYW1PY9fhH4JaO994xAlFyoqs7TMGnUNLl1HOdEtGbsiu7wUmVSeV0hrF0j+bT
YRSGBPvsxxlE++SMna3M2mdvCi2gFuZ/6wdbKvqp1U4vylcbVScDNj5QQA+U4p2Q8CVknEoy2sN2
+xnOtnvkKSjagJXS/bNxoqTrdpCjMeE+O1HOZWB4F4Z9ODwkSPlp80StrstqcdpjoTJGBAQ0Iiyv
n8wDInxj5xbVN1W3qeiN0G8hEGg1gbEIFQ3phGMVofFyW+ujt4gZIkWI7DVP3eqM2hNgdKae/lP7
4r46b+H8fif2Pzl1qlUXZLftPSCDdP34PXJaXMUzty20zLeO3ZQdlZQW/q1KqtUkGcOFNc3Z+5ov
bv1+ya4IF5+YY8MMoEC5W/DLxhq4xkNZFC2cuHj3TdL/BmjPOmOM1sYozi3uac0BoX0uL+bDL4CL
e0pF078EXPk4BKBi+tqf3QoSrQjSiFKH+yxUI2t+7FzqOyMN83cpt92637+kFseKfGgDfnpbKXiQ
Sw25VvE3DfidmSesiJZMoJBAmT2XP/OMKL3d2VYEUR+szS2V9pxH29u2F4hJnzN5SDBe4ka6x9V+
piM9r7Xm7aU/O7W+PL07vujRyefr9Z9JqfBJSuNepbr0CSAeSLUqJ/A0sp2tm/Y6ExPP6lTr3GVX
Gm3el+0Hr4S0XDiBlqSJbQUmvmXDngURPj6yqHgvG6ADmAZxsDdsXvnkI7bH4QcjyPGHDF4CYQ0x
iKZPDHSzdBCKRJKbBpWIn2xiYSsgdxHMjEZN9R2pTOvIowHhsKlLk7zBjFIhsQKI1coYyrrhlkON
Em/B64ENIlJbvUAiEfO909w+AiOkDM+iPOD/+hipIltiwyUCeNobn+NbjIYJQKzISFhCD0H3THOZ
1FYy8DV0SBVT63KcqqosItej1l7L0I4I2MC2/cqDBICqHe0QqnSzg5+2Z1VHslPVYZIfWEzSuSiC
qqEP49hWmZcuPgfQlYi+zI5eBc9CDgv1a1sZb9APHbMOEmR9PHB9O9ZuCDcN1t1EfgQD4zyeOYtY
kohpW2yIQacd3aNqWmZuEw8bT40p2FtG5K/nr+5ddz1cnOJ21qkxFKXdBj8cI0G4X+PVlHhzeRVW
IyUkiUdtnxz9rfujpY1oD3kYmqnsT4Hg4NAR5cQiEKZZ8ENt8ImowDNvSDbT1F4UQE8+xsl7jPQ6
GtpyBltC96xiEK+QsGuVZ4MuKAE7LwwUpiFu9KNNblymSkrP27q/Je//auDsMkJe2pV8E2vP9XAK
4tDgO+Hj03cfdp2hnJFyTczlytG5l5Eo32BcCF/G6QymzfRFfNgExg3LJ6NPUUzB7l91+n/St7r0
/e5RSvCEQWXrpfywmY6DPDi0VRXoCNmI/LbpR3x7OC1sRIPyHdYJc+BxesfZFoGaECHa1TbAh64n
QGlhEKNaGEC1vXntN47Fvb8FBzEPyLWmyuXhtPncG9XJxNKIDoCR5lBCyekP1k4640dIm8o/CTWw
Z0GDeUpD5gufmK8c+bu/9s1h6HIO+ANLxIRgOeGTiI86KytVeBQbgTbudZ768VNoBUtl9V6WqtV5
kqDR2YOyau5JI0Tqmvlnj/55obFV/2/XCxSCO3kIiqpJ2vAT1STcYg0NCEdzQk7163JWXFV0vK1Q
0GhDQhuN3XAe5nnJO530dcRDnfv3FeUAq+7jc0sIPGx0Uyno5gHVc2UZBmVsoMpJLbrKT5Is7/Qz
og35jfj/cc+5jyOdg9DoBfKs11zNWze58J4A5uxkJwxV0FAoBnW7UbkGknNxFLQCFe72ZucwYzJB
UV8Z8zfaiO/wUlh87X5ov77f4bBEGXn+4fJucc/kq3tXbYZIC2ALA5L/RvCHbv2Zt2CQDqtMNia/
485tEuzH9/XRi67VA/0LDJtvPo39pSa/ytr2YMvor317/rc4kyV7Op/1rFv9BT+Wt8JkkSi2N8rj
zVCcY8aHkJuxwgNA2QUY/5mt+vUQVnmEoxvCzNBU5DNulRPqFOxtmEDTVz/oRDT1VvQUvP2kiH+A
eNqy4EBWNmiWS+pNrSKor3NvkxuQ2WLKHFH29YO7ld7EG6JtPIKyU2/TdcaPLTZ0AcQ87TEczo3X
Kpfi6trBohj1IItDIMstdeU0m2HTquAu1VytC1jybWqsyUTJp18QWqXd56p/xyUqm1V9tvcv4kFP
fD6yRpzJbb+cSrPw+ACt2K8I9DrgUR8gt/eDpir6gqY1xWOD995nVKgDYLSmXaSbKItz0jTS6aDc
/T4DGVm3HkG6QG8w+MKoeAGtXmkxR7qNCIImd+5BoLIqXHIBgKQUd/fqCkt7DMq+844cejJNQ3A0
0jM3lNfaK4UiXoV8Ygh51rV5fWTIMn+V7Afm8GP3phVuZMjiYqyqnqIJPyDCdkwPXeT5cT+tbR2G
FMOpvhfu3AO66U3pOh8MDaWOWj2rhW9SN1rHSvJfoA1CVAJXIsSj2Uul36bR2wc8Sy0WOc4afPDU
IWuVwtxfdD77kKJ1YIt+I33PJZPHemUrtp4vETJcJBwLYXwJO6br3UnCBcj/bhFCX2s9tOCZ+Y7l
vCxKlLP4UXjSHOy1mQIaVpgBjUzgXWuAQ4alCj349W1LsM6OoXiIt+caFsKOd8qnLmjcXkSiTt83
4C/32Oip0iL4SQ7yUo+bTdNZ2Z60+k65fnt4umY0Lysl2shtR+cqjWfjiF6kLL8p1ocByxE+hOsC
1QXToXIjND9VdYVO8imD3aNZwL0PYGn0HV9x2jn6EuoIIEDLW0isIs/dboACtC7QCu47pbbDFWYJ
3OhcMkUOKKagRvIYR9Ihx1XjiuWASCNM7/nz2F5yEhUtsVS6sV8p782mLZn0Pmb4S+W4c8jEQFj5
X5YtpSdwUeb1GNwC+A9xea/twEzRd1kAzEAx7del2UjJjxg01SUbDpBkexSh7JODfFoCgDSTKhfG
g/cITIgR/YnXSptT7Wo1i6PeYsCY8CfqgHcAe7QHpr4ekNpDWossb/lGo66epeHl+ckWFhcuxhmW
h0S8HxBhmwubEdez7+edIFFx1Ax93UMlGOyGqQXJBKwacL9YbnbaJkSzghFFkTFyPZ+K9vbZz9l7
k1JO/z1FAlzavR5f35KRHDmNT7tX6AEi6D0gbvPhuifEkxd5Yv+VvCDASY3pGUIYC/gN0XATbky0
b+Vk/kuACV1jrdHasTOQm62fMSZWe4p2ri2Xj0HHTe+djKziYwfYzdHokMZKvQ+Ics23wQOcwbM6
J5JkIxTXm/fKGPl5mg+gWSn8YS+d14oOLu+rf4NP8jHrJYeY2prImLMsmZeOPOxcqCKHVw88pag5
qOB6NvZWZvVJN4kM+bH1qHHRizU3UwV0IjvJ1uu1Uv7Aqkv2lTV/YejC/pso3C32XW0ZPbRcqM3x
HcsY8ypOJ75w8085t9wKPM9thKnqXBXcDNsyqaTnp0n95gaFr63H9pPRJ20k9L+LXfy18D3vwxIo
2AnF5/476BbqqBvs3xXXb9d0h/kU+nGOT7EQrJjbyn/ErjKTJQUTwRhPTZMKqqiOx48XeBZC43i1
ifM47RG200ufUCxn2Gt/xCBpNkA3mZUaE4OlI1o6UtFu8NAOmFt8GV10URxlsw7LJBO7O7dA/uZD
G2h5OKtsTfY+BeHMYsMbPIwQp3o71XzHin0fSN45V1X5zDtM4x2qOAGngWin/7tA+XdpBjg2wyna
QHbOhzDHxOrb9PfwiNT+hcFHVACAxYONTxIlmgDd2B2705SMfsjRw16YIWByghx7uVYSxNmzw8A2
rlxKaKeSkzg+pZRluIM7UTcZ/L5K0EUuocSCtsOSAeE+tlX+gFxfdoYhM0Z8m5POn251xrr5K4r6
svmGZjWe/Kh85e7tOl7BrEqkn++bFYkrBLG7WHd6Sr1/hOClE7VWTmTr5jp43bVSwvnjbBt5ChTz
mWPBtan3jS6IZufP/Zw0f9iFq+XYdbGN1zab3A2ZdLEPTs7IpVP0g0KV0O5tFAunFYvS5+0EN0fW
CoGFi77uh7suPkbXdRsvJRgzDJTXEfG/orAd3Uk5dCMawnO9HBdJ2ky0+isnafE2qb4AQH+KMBjJ
n2M7cWFSXiCs6n60vDS+uzPRBPR/UmCF8KsubqySnEx8qVSMdFy8dCXTsSQi2dElhuq9aB6cIRy9
8HnSv3jlIeblg1jYUQft0zW8iLVubBblmAlI9WtVVYlaaHW1fQ8GQ0fn4jXEaybc9Qkn6MhjZhc0
h1lYMOWLOO/xh4YKVvvB9+YmFfPwyGPYt+tceoWwKH0c2l2Chrro5H9iF4RQ4D6fwUSX3UxYK8k8
c1I/m9TuZTJ5AY6+jYb55e+Lt6qJd9fIwzitXlfgxYtgHmU4Dhk41GK89fSelGz5lvGJCMn/nY9W
XIhBYRkGNaa62iKNDxCNlIru1jx3j8y+hwkotqpL2jvjOOGjmKMsnlx+4otw2a/rgD4Xx5bW+DS7
J+dmTWvSg3UjNZjiHs9q5+QMzjvVbFdBHL99jh/44cYhE1Oh8gXDEL3xM+/64PGnQK81lUY0W+hj
dXnLkQhbaU0KBiU+oE94AzUPnEOZlNEVUfGlowz0hQoNaoV1RDmIB5UvpyKK2c/ISra/RbPLCREO
t9GW9ODR4Wp3PjjlR9Jb/XT1WrWSvM+ueIAXlHR8/7GdBYLm5x69hqsZc88KZWB/iY9eG3YOA6XU
BL3bGSnIk/RN7DqGtKCf/nSduMYTojbLHUn9US5tN7BpG5OkFFXO5xy4ZMBSmdTxeFYvAwyqV+fA
GVYUAaiUpcJ7kfn5CYShSG0WeP5MBWpL3V1CshT+PR9lojmjGxOI8PzrJOzUpQcHilE8L+F9Uakz
oMT8fSE/dlhB5ejoYfQhWH1pmHS0WgBDXVZtiYTdi7zwr8LVCGdyik1iHQ3x/zW7Rn0AINIfYwwW
zRvko9lwL5wc57YhNPapEYtwPcvnHbGjDFJ+9oteBbiTS43I0TYP3WyMDDl00SEqhRip+CWkTrF9
PvVQsy9eiAG/JvEYHTa5mLmsJdWDKKhVrrnB50scIk7ACwMmbXOJ4I325rK5hxKUIrd7ocjh3Lyd
2WRjI2dKsiLNN7sT/6oYX8/DjBQLVK0TJBDPUHaCbP4noyD/dni8c61y6jqsszc/DayQnNjzSuVP
9SBe7sQIc+Tg4EiUN1gcTVmVD3zIIQdc8Y4uD0vPQxEXyy0VdZCjGc/GKN7v/h7ZnqZgVMo5LYzr
GxkNBZ01sdUHTVc4tr9+Vv7RTJ6zKUiw1ULXsy7D63NYuhT4+6FeBUJbbyuMpVFhPJ6hwmjNJHUI
/xOMjRP+ZYL54kGFyCXudGA/FWlE0C3EIdX7Vzse2TkrrnWu+Modtk3XpmEGosG6/neGl1DcE+JL
m/uVg0WnPlpWN024YRNktNJyeh4liEIv3tFX5n5301y+HLeg54oI57cAwROuKBbl7zQ9X0RkaX4z
ZMCWz3u8RUZEHcroM3Dko6RSjgU+2e7Pu7PPDZ0PBwvzU7vrIiwi1E2JR/2v2AOHO9WH9OW/xwf/
u+SI/NUUQ9UoIp4KeKw2sNb9E+DYoNYx1TQjqG9QBxbZnWOkRvEuCXaF3Q038HEhipguzcoTfADn
ZZE2sM2Td5+afQun8lkQNZ4xHiszys0XiQJLj2VAsfL8k1qr8b2B4i0aiCckAQnsXh2/OpmrwsZY
JRE9KYZgfTPgfOE8rr8mCUSjIZBNxDINAlRg5mdMVeUOnwSW85Ao4soksvYj8UeVjjQ/QNae9+aF
PC+g12czAY6XZK8pr6/aEgINiYDvr4+bJR3QRpANPiJGxWwCQZaBm5wMsx5WCTfQZwKq+3EDQNP4
kEtNSaxDOijzsRtLnzeGZbd++pUoUpqrB7gp+o1b8OLh2ZcW4YSSsJf3UzTyYuOya1otxp+6HuT4
4s1FGkp3ote4VdDsP5nSQf6rXgOx3LbK77/kDKJTd1j+wHGM+YvXyYQUqcWCsYPiGOF189dLBQPY
hIjBOdoL4ZlfYXmzrVfU080dUHMqJOH54Zc2uOA/b5/+W1hxNndhx2cGO5nFMegXDcqRjoPvZ8e7
8y3J5bpf0PqwlsicQzU98t0ujpTyuFT0xPbV0pKMqWLmhRpy2sXYCYTdIP8Y1dXAXSFwlacMxy0F
29YMX84629QnFX0BFDPHAyNhwABmdN8nJYe11T3+hphtFOA3flLtXilWrCe+BDBrWiti2HuYKSwT
4ysB8CIL7dPcEZlRqMwqgiBkedixK82xFiLYmvsOdIcNChixdAj1dkTpr1FIZj5XI1tUVC5rCBA6
fGGj04g3HbmQQXAf8voJj0Wlwh/t+hUkHr/d+D1AJ1vBQGnHMHYu9uV9bZPhCSDp1/ALEWReCkqo
hnbFUYCGRpvF/gPBROepHdBQLRhw0IMrDAGlvtVMGJ5eizZamxASSdV3y1LMHTXrUlRZY/hPuz05
ipmrNHoxd+tcWt4rWx6PAz/prODaHTEYE7wrNiccxI8GzYiPj57LHlWJ1jUsn90zddxN8v+dBLWL
SMyVWH8iwVGe40GoqMZ5V/EYbR/HZe0sPNFT6WVxwsK98nIJSt7A58n6TwDBI7bC6yLHzsfqTaNE
C1EHpiYEWdITyNGtJy89dA64via6pkZNLKW2WRVd363Q9eYVVZdj+wXnj0moOpnOhzmH9+fo3J8n
qVv1F0P4948Cp1vbLbTCdYfZBsJ/r11+M6AfT6/opOGrnGpJkmX0fip+JKgHX48QY+Jx+GAh+n0c
vLMWi/uycetYbO304hDWJQZz7CSnuuWFJr7987SRYUuWAhcWa7Y1QtLrXsQRdBr6mkkCynBR1XAX
kah7nmBkBh6aymMVBhhMSlgsoNIBDZ/LOhFQyY4rXpV34BBYoO6nGb5q2UWDiUZ6bFHbyi5jdRqN
2Ctkdnn0Xj1hU0ejR6vLabkx8JpGyJeXjIP4RLc1fjPygUz7cweTNhJzxvtp7NRhEkAIq/+spPuX
RSqjaQp9oOSdJSuS8axe5z+KmT2NnjgmbUkyQU3nMlK+8B36gbvRZo7vZpu6xzdVW4yqFvWycUS1
G0ehOQIPezRHdXDAXQMkkrpQSHze8rzr3k49jq99NWQc1sX+/cTMhPILE8ScWxwBBS87AG9BDKQN
z67pAuJYl7IVYMAfSal12V9wYnwkt/O2sybCsgauwl86Sa/BVIHC7pLJpP1gBXUj3fGN1UkoEaKf
nRmvMxsKP483n4roKJzJRY3XO6LjAmjC1DE5U+qJqv5ak2KKT8stwnG9dA+tVsqIUnkGBHIqmbXT
wI87yWLSQUlj9l3CiTIgnebS54JRIkS9yF2Gpu7LlwdRyajzO1yVbsRsmwz753pW2oiAl8VL89CZ
FXBZJUF0pljHc/WDDnfral9x8QjD9tjVd97Qjyj256gcppUIgLTqVIhBYKeQbShXRKahZyrkxZM7
+1EstBstxelJ0lgMTPIw3EGC5yn0diaZ209pkkcg6Qxdig8V/6QLildgrB+oWKyHygMZiYC17AE8
H4HHUC0U7/yCzfRPuUnHhbZsugiff6PjinMk069WrbxKvaNdLFzcu/DY/7zVgS8QkVpqXFkFbcCa
sUWJ+xf6+Tjshcn90ilaZJOstSOUPAb0G3+9qcZRWUCjellQZPMxEf1PUJv3Nfq7LzrK/bDlKoWE
bdAdeyIvRg89VEcTJpImD9XcnvvyLAoGHUWsCLQAr/QR4xbtGGnks/j0VFWxMwRKYHB9B51qMP54
hBuI507V3pX96bY0Vc+BeWWV//44Ckx2jqKkBUx+I6nRlj4QE0bpTtltKnPnaGJWX+TlE11MwrZp
9m5U2XqT8OYT00EMtJonEgEGqNiIDlnb+5YYJyrwteeM5CoqSjb31gDtlRdvCyT9JDAkbTD5EM1Z
BUc/yL8nLX1WC89SiAQThB+gXmZZv7dL9qMPihn2fFHgud4aJW74+2Gzx+D9yBCE1gls/EBr+CeG
wHUacQLXV2q+WdEZ2ELq/Mw/OrvPGoZRt9xkrtJel3aHPemv60WHHRNpjFntUvM/TNOo1T2BuoIf
S9nN2krUHNpnuheHf7MHgSebQrdu2p6u4UUaE9W+Qe2rGMZKEa5nrnUcUhM9o74hCgE7BOhNigl6
hXy9pWvjRYqEoDIHYxSg3Xhu0JIXzH3VN3157Ae50iYtduOT7fF6RT26jHTS31CxfqIZ6clcH5r0
VIkjIQXMw9nGmtfwkJyHWeKJhYk2qAELi6y06aTWjyFWacTxKmuwEG03z8boc+taZC9wdFIwWea9
V9jatVWWZrysk+LFIVXdHS6VN2TM4lIdKDU/IhRhm2VtU+ztAVub/SwwYHcQjq323fYJ/vHMw31d
1ihlKS1v1AZasibOj1yiNd60HsiJgfUXU8w9RVjwp0tyVWMyVHHpFDZ1smb/P0YbmFe0YKVBmw08
8sBernag96KmtuJrEOvgqgm5zTpCtr9u0w1pnwGNpoQcIZ6XaW+W69mQWUp+LE5eCZdV+wNnwwY+
n03pM7CbqToBgXx5PeSB2d8Yl58Q9BjtUjOyft/OtYQpKMq0L9o8x5TQPfv4gVnYJIFgww4uFgN/
y0zvEhI3PpwNeJ/kRlvubeuIuI0ow+kMsRFWFL7vLNkWwuqZecyqJ/7c37PgU379GtoL8XJ/Bxgw
OmG6v14AfeH4F1wW/yxVC4UmQe2MIP6fAyhFVikYXqYTJTPKZ/bSbWpOrcOpdjy1heAc9kR+0dRj
DuEvtB4sDaa9+FSTrjU6B+fEgQ/l0JHQgGAGk3uyENGOdIjdAfOPrX0Tc40M90trb2Am4hIcV/SS
/oFxIscBmT6TnJMOkKDg9Fa4ztbw2Xtna6g+SzT3XpNDEfKmK9dDZMsR8bCJVl9eEFBHjL30Joha
JvWBO8PLICt8pW0rdcSYniuzuRu5VskIlIkKJVkc9RQHGqrKyPZpFuQIqUaBgw45mYb/m2JWxP1S
+/H4TQSRnbxONrSKP0JvKhjPAtpsmZTnvSsQwqNY6b/ggPbmwqbSQTlrtMmzYIxsLeFsKxmoKrUJ
cEzH4yllU5vOvV4XovvqYhBrlOlPWV1I2uB2d+gGhVvJpSdRBC+5V0LzOIJchHH1NkTopHKNxQ2B
QfrTYun3iXecc5F55qKR42bP+Q8m9+uoiZWFD/7Hf8OCJiSX5VHFihUn02sxylNdtP18DYzuRDRm
XIYX3vauUFYF8MWOhAq/XyvPIspUhR8ZCZC1sypY8ZeZqYWe7rAyBKpfAVoNMpPjUimlSne69ZDZ
175ifWm9dIcDw5OuKmoZZCjJOcyzyjun6IkRIP2oj0zYj0cO7Ty8zg8YjXcF7zxCShnVU/oMn8GS
nnFYclSJ7sdzGfeEVsO9Rtvq5z9eWjMhfc8vqdCXTSMnyybpjFiQ+t5oQghk4VkmO5jHtSD8JY3D
8WTv0mk37Ced9sljkjoP1ac9AIctDYcSsZgMM3K6/zHmv1YBDtNu51MOv0Gs5R6c7aGRlPuMEg4z
miHIAUHE5NYV6zEsd6299qcERHXos9sfHC9quGf4u327sNsK6NHUl6fKjOCQP88cXCk/Bn4To6Yf
gS5jcFZKVk7D4NhffBpVVLT4sAL1hn2C/l8aetmMQkXrxj1EGlBZV9cBiUyVrfZAxXraqPJdepLt
RgiQNMQHLe4akrzGq0FYpJMJ9k6E408S/O5K31ExlpEwFO95ypVFKKbFh2ieliHIbDq1jbU3ldAe
Olb19NpleEdv5PP2jBZeLMZJlTZDQrWXR7oXlFa+psDJvDJKaSfEX3MQN2Ci5/SVgDFyI0chRswl
rPYctjfY4Nzmdl+Hkfc8BW8HvnchgkMHL9t3923l265CpUyTCLAwT8RDQmm8MmCqt6nOMe+JpIQi
S9UKePSTcmghb0HSn1qh0F/R/zTBny8Gln1B8+sb1aR8ceKee3AF15NZKCMav2pz9D4Uf0OaZr4T
EXcfTQp/nAH24eR4fKPzuvcR2gOnSQ3dyJBW6jRgJAQ6m01rHlvdoU+/FiuQDKFQl2VVcfIr6Uu+
g8CszmWkOqjf7UP9EX7hdNrDQQWu0bD1HKHL7NKRXdjkv1F/PUa6D0V9yMvqBIaRXED8z+T/BJhh
kR68nrT7tMlvp5AcEWqnWwPtSOQNDe7JHtvXnkWkH5Vj3Hm/KsrLQweg6wM2PtGiTcPAZn+ahA8g
NC6E6k/RKodgaBGZ6IP1792KahGymrZaKslj0dSaI5PdizT23KUH7SowMrOCMMXYa0NM7ckh/IUt
9t73Bwkq4IHR05kvaLvgpZGVoiw0nrW0gnghttuG+b9iz5mn61ZNashmR0rHZ3U0G+cvusy2Bh4E
/ij/iLj7BsABuCTEKnvKfZt2LVRyRQxBLLlUKAFw5y2UH/JuyCUfvQNs0mgbSI+ywPrwGwkLMSvg
WKyjjByZrS81Na/kmKnRF2BmwWwOAXUfMH1+9OLCBiPfcVJP2yRnEYvEvuHtBEgdX2Bw4lgystKr
25Ppu92xuJgRWm75+oljpw2ceL77dT4r7X+WlFE+onGmoYUfI/gv4RbnkjqKFQ4/u9kdUs2yFatO
2vcUb8tKhDTUa1PZiotuHjxK82M9l6jgMRtYmA/Z2nxd17WNsurURwCA3bRDZQFW83E2YciPzq2y
MW8yJyQ7XEqO+4IN98FVmFoTGSkfqAgS++kv2f8I2eNSHoErwbfb6VbXO0HgAJrZ1/kvXL558Dco
ihwr1e81xkCEyXpXS10D6ZfWbZz7sxEZV9/BjNp3BteQCFzO0h4hL769A/aY8wZhHMCJpJ6SnhHj
XyJ3BLDMqvf+qcop7k+wl0BPjr276/OJTanVXXqkhT+YjxACbwAGs1DQxsXUW+kBSFhirgbqUulk
CIcNViGOs8ERmqc+rV/9QZFYNv4R4MftxinVZQOg9y9MzQlUDJjDjG4zy4r5zVqL5EAisjRO3i/Z
OzAVLs5bJvP+XOS4J0CjZ9w21CaFAFogEUIwU9iJAKSJL1eLiZBdntGkW4QIQqzvE5hsxneanBIJ
TI4wR9shE2UjHieOzp1CngYdimCzedcUHVLlrw4miUzjrLlUdKdbQ7Env5UFMpsuU9Y2wrH94oEJ
M9OYcJe75O3R5GPvaQcTbs20qacQB4v79raJSqezpRlhKLHZqe0HgYLX8Ar5IR+xCTNS2y6ZqDSS
9xtIU8eOgGj4jBL8pE4LlHTj08VO22SO323cVq1DyGcQNThPpsqzE4i9O31by9tf6quaYNLzcP/w
xHbqVqS2MVcHXBkDSYgtf+RXtmN8iJt2fk9WOP5bItt6Kny9m6ENbRj2O3xHHloCsQWWYUd+i5h7
uRPaH2zUwTCKcbWzBqh2d5nUOU4+JS369Vfw+De7PoPuDdUbz15SGFnyAhxxfbWGv0QagWup2M5e
vLQFHSV3Ackcx2x0pOhIuBnzc0iO9972BAPJx2oS0N4wgHSRADXxdm/2Y4jHiIsTTsUXJHWGYZvc
LH3I5VKEA+izyis3Ea/QT95RjZ0U1Ov/mcUXINhkZFS/FLL9sbrRrwRNq0EwgHlXcUpIozWgJER2
1auCONITEpjAgpT2Ut/JjBg6NnfU4iVx3aRAcgaXEyP0Y4HnnhEsZ/FshpOyc72iIuOU15MZ+O1S
isnjR8/aoUDU98XEopQANk5j1gO0FU+oPaXMmrgG65se8F/Adx+tEJ0VD4fvA9ktKfxWDRV/2/Bx
5w3GAY04VdOoOIEgCwYt4aU80Bbh5BBF+KibMn7lroC0cNDqL+QgUFKsAcVRQlJXmI4cdGZFrDFB
2DuYVM3tNDzaspyyMtGGEVTXbPBeEwE9Yp00lB7/u5rE3YQXAG8VlwbnLsSV3p9K7nTlgUYozJPN
Ct12N5Nmb9v5x+TfN+Vg+nHBWJuMwJ684YaTVwbMIJQD9tor+ke0pbCnzc+A8Q4V5GfbIYRWGgRZ
nEbbEljuXLdn/gOCG1Yxjl9DyALgDiy4vs2uWJcXlgvhNtYftacOtwo8CV29eD9o27xK2TDdtVDr
/p/EyRN4SAtjNMvZneD4s7tKNUouAzFb+NkTue+4ycDpbuZ+eFYiIptWyZu9n4rcpp+3x5iRcRDR
bGg43QHr8qnTe2oNzyUJ5F2cMZLNQ+XI2nIpELH/PpoySua8HAMa/7opQEJ7TfnST66PttAtpX5e
V64VjDvbsngGYy7lWfZr3gPV3B09I8HHlfvD6cx2JCAdpjpyCe3ibS5U7R3pciZvzBtPRMHbGQi2
Dbm9Vx+Sa/UUQqm0EhCgHAy+TPdEMJUKQUg6GIUsuuPpo78mFo+Z2aiMt/az/L/QIJTlM207aGMl
INpZY/2iYoXCA4BEKM6uAJEiHw+96ZHFpADu/4d3qmt2GENyZMXjn3zph1tZOO/PXe0BPFN9jlIp
3FTfZQj7j12FI41UTLRucKm7rhloeVLM9qZoUpxZNamqU6dnx3iHWnJ+QQQzBmVYgyNTeSlkC/zE
OZSwknyhkwhjIEenaOQsMmdhfTXq/t3UYFCyfgARcfdBmrdQi+zsxcC6MHiTlLXybxJcfxRvebCe
GZ05Cb6CqL9D1006tF7sAY5btYymWwS5Iu9YAtUXy+la7mXKq1X7usfhj1IUSG/3WnPD8OOFJ++r
zXEbPm/PbT6ClqsLKxnjZcYxMB0oG5gl/m36pY2tQfxhM67IAHC0bnkoBHQav3x4wF0wH/l61QxS
RJIasAUpqOd2Eo1TM+35gEQkhrseJtHquxrwCOZjE+pikjAPjbzJItOof/JyybyJ4SMet3BIVTdp
DCIes3FOFJxT1XX7cbhc93KsrlwqZc+46ZxAMQFzewzVtZi9CEEMSv/9Zq2B5bvreT176s7boGZg
L7qT+ug2bWFhfcSGmXiIUoqLXrk1V3upcqO3EfA89Q67WaF+GhSHoT3wd0fNUeaSsk3dZRx3fUiU
XI7bdJ2+nZKH1Hp0419VTU4StCc9TQ5WkivSDWcYPyH4IDVbgUOfEi236aeD5Q+cV6e5T+db7ha6
82mrYA1MgEddgLCEl/nOxVjtjYApzBSCpPfvI4XAfB2HxZ2hTOey5/kUWBOLlLwXYa1uIkQCPB19
0ecyRi7bgp/zXMnR54514ozlYPDlFS2hHfAr454tSXEkiy+fsJVHIORYBjOdNhTGWdaejfGrb5DT
I6H6z/O5y/1JsOrBs4s+MyE0z3n7D5F2Tz8e+gsXMtRnILYbQ69F57r8+zbVMVc3ONgnu/j3xnvE
DoMm9gid1qpJBB3sCDXI9w3fkQcCzeNeR576OUWPxWvg6ZFiMOgi0osDprxNh2i1j8+vKymY9u6y
02H24pbI9Iqtc/1/W1GSaTUH/kpOm6yfblakhHunCZ87SI3jEuRekD7GLce9w3/DxOQQiJmvcbB5
y9pis5Ru0GJHRQRmHGn0CfnBNjhFjZp7SJQt0s89eAmIb28iCpooMHbPPAbCF4LYnuTLMmtlp1aN
Lx+YB7W4f+WdGyzb2JO6WWRWecIJKh7YkbzKDi9RF6fcC6Vv2Fo0HLEFQDicltzuhrxR7y0PxaA2
2HeA9OaBOAHp0v+XBmeCH9acAtTQw2klpuFIxLG5Nge0E/Z7EGKFq2Rf3IPa6T/3iyNingXkqkn4
MawRgQrYLP/0mEyQAdbXfx8zqKZLmknyBh7wSplXQV/veu5oiAi5dRRwInE/q+HRKpJoculk0wK2
O9EizYjXhEnjJXoMlTFtl/neTaR17fMgfm3bZUlr6cs355WeugKHpOCgOatjDEUj78xuYqq6FDQr
zYuV+Dr2SbwVmBxaLfGrxOMtPT5vKOTS+gLN5q+/GEiMLi7tnLcjNy3AUhEeNlnKNihTttXWzmTk
u4pQofEnAnw53re/j4F/pRoU8lPMwgrP5Cd2hZYF6o8YrdAwgTM97+I5RKtmD4Fo8B7K3rf2AY5A
x12EGfmnuCwjjB4exPST6+qnEVEWXcAsiAXDdteStmuiy6DZJMeb5dUxGKb+jT4jMZrUCzDgFFdP
LanxoD05tXJWc4vF8ei1FzRIV10ip7kz6Aytm7HasuS+qPWgZovIk8vMqHmvZGGBhgqqHEDxqRFY
9+4WCmyY40GiBkD5F8EbV/VSDwP7Dzn7p0+oy2ap95K/qGt/hhHF7XIUD2OjiO56lJyDLHYaPEGO
yl0NIm/mF4jurZMoJbdDnEz14wAljEMvbQVro4wp5RZjHrZvJzHsRQkxfYx6zQ7cz7j1v67gvZYu
dT4HTzTFnLhpYio+SIHxwOxwyB/X6bA/3S8aAiRCDcC/+MSA7DWUBAIhvD6xImIW1aYTavHyTBAK
FsHReQLptl6E4i1FJwuDv3uXKSthAVBnKtSzGfDeWV9m2uyABEJTxoxEPowufBPwYlVmw2bqGeRG
AsWGOaJGeyMGtYJbhm/le/hiwyC037U5oh/gs0kLC6MVeJVH+ywrRDXQdaTKLvmYWvUEhbuch3md
PY7tEtsh/Pa+ya/XcrArw6zDb/+qFgD4wPKpOBUQMmxmAP5RCN8FfS0wduV4D1SRSNJebcSMnZnK
uY/obQLBwVn44rKW/F5z9x4e43Sv2A/WpaHj1wYNXonQdYnpUWXfigMeSGrRJwOMeN81/K2WnwLr
K+9rQM/8KC4tBMtBNwDcQB7PuvfY7daP4rqwrtGM5eM2UPQSNNc/zpAEwj9G+7mSV1tVvQkY5fpT
6+hn4TWIk+ISTWfRNYHxBfUAOHBYlL4Amzm2H1LtafPC18itwbNFJso4TNrDTNOyV8nnN4VZV156
kQUkbuiJA1CqssttBHDbWe8+fP3IMz6E4Zw4vx3tutQ5nY5VmhucVL3kfRG/gXLMyD+91kWm2svJ
26xd08e6ENzGtGwY+Ign3Wt4kAR/B7DCrkTq7HT0yhbRax4GUIvJ2UGymW3hGfJm1k8s28iCox0N
v3zh9B5nzCdoCxYmVXuoMauaNqAhpZosfrItR1DTrdsEH1bXamW8nJLX379nFobNJMYCIZC+yCUQ
HOH5mBe4WOWWXnpz2TOPbINFERt/oOLfDG4vx7DELFOmA2Ws01e85SDejispzZzs/QLwrWZjltsU
v2mWvuDHyapDMFg8XDJ010FiaS3Bi++h9z306L0Mv6zTu+UfUDkpwKB/AzDxbHpriy8efnQyJ3fZ
rek0UKRPmk27VZsjN+TkffriwM9R6LgJhmAD7haOLRNS0mH6oxOIebgmd/1ve5TvSQsO22rL/LRN
nQ4S4uR5NErPYwx2iknQ0twq8mVKr9qkAtPy2TWf5S9qZtI6/QfYmOp1xxoJ+5s1JxiXAG+ZDbI/
VSn3qhXoiQqa4S1IAwigPwflshyMEmRe0j13D+GWHU1inNchF8JfThSMYoCYzTvrJK2vU2FvBiGv
dH7/AnT64+TKp3UHNHTnZk1kxc+1Y04h20vlqAxz8Ik6TFViUzPs93GAKS0maEjFHIV8CRREYmmu
TNg3uC++kkYq4f8C7AN6W5u/8BnHrItMWuus3RW0YDQFinrlGat7AMb/iOkGKKjLwUaHnoPatz9X
R+hhq7hcoy6I3Ti7XeyPKT2ktzZbdjUfq3iw4SyhBoV2AmXBEwtR2/2F2myXL7zXKfde3PtH6VL/
ofP710kAuuPwwjpoMRyycPV1BhXkvg/+pXa3sOchE7WC73tCn57frj6UZ50KSpBswA6vnUzWpmZY
oV20wF+h3/1CpgLtYV6jNZMDrGWExhkhr4g4NrAXP1Ldyztwo1dunc6TO6wisyMZ36L1GEw4ij6L
vtwfAoJu9td2d3335ZY6mI6RlTx6VMOsgV4XR/XPKwMeJCMtlbCr1HiYcWBEcWTAh32tqA9tyo7/
15x1uoIhF/b8w/1EIOXz9g8ZAcv3L3BNH9umd1Ap1TR15UuBQBxhs/LAu8zGwcb+M76ZQlsj46p1
KAq9YkrltNwA2RXH0cBFdzw0mkB+sQgAylPynv/nPafFXjMAYviIEzDqFCdO5GpgdjmpDMMAXVrg
3eB1ALwkwC/ubuCMnbOhLYni3wDNSPEPFwLtbBnlgvrux+t4/DPOT7fhWDYCBCni0LRYOt6ZAvyb
Sihf1NsnC57G8yFcCrweLXsFy0qrRAdA13RDH+qMmb9A1IFFKBeOdb+/Ou+6XwcXaxiM7XvTMtnm
C8sMGx+7A4SSaixkuakgJugL5/I2o57B3w08L5HqRxwrCcWvqeCJzp7NBWXe+PkETcLWKkNXff8S
eneUJNmzZGS9+1lfmD3B4CQ9JGk4FILe2lrpWi/2j7mXkuR/zS82B6jY/LqKJiJdfxfWeHJLLk/L
jEbeUIVGWj2fMfxMK/ZuqxpfNYxWRVyUUD1+RZ4crmMshuOYtmv7LTZdE690baTKQNf77ZrH1ZYp
1QvFUpQila8TjeCYtSFxTxDULNz/apO+r5keA7fKT4CbNY8qNxy1Y1afpubxt9un2XwU7R6idYOM
nqSez7u56TcAAUT3xRUBYtDY77rpNE/Ft7Cw9rawKUUHrNNHktCWAA1EJLnwUw9DczrS/ukex2eL
0u6VuB/qPkNxJYVJr2Q5MhRdPkxzpd8ix+l4v6C6BNRDDZmgjWpI6fA7g1poT7zSyqAkHUtGtjmw
Sqfw6+rboR6TY11wxkHzj2xMqnur4iid9AwWbJUW9Zloxd3sLx7fiz71DWJytEgVJAwScVDFFxL6
6TvLAy2zqPEMAfxJ/NcydMZ5gLhmz+nekxjjr8DQrRwC00nJLUlxL33ZjJ46D8jkDAFtTnZStMrM
ASTeNhRyIda9a2qX6Thjg0Qwa+FvlfsokqebndOGWWvxJzf6fB3A7S/TY6A5ALbN7uXe8rOK5uGf
Jd/ugLWot7EY/1fR4cgrg0zls+TuLOb9Nl9UfMKXV4Wl8iQKrt4e+914CwnelnrQF4VoU2HbRVZC
M3x6u9kMFL6JXtvrB8g4r1+T93c86sileoUC/JUSyMwwmQ4Dl0g7y3O3RAwzLcCcNP/txxWPXpMv
z0v/hSWRjxrAt/gmLoWWnpIumRn/vfmYO+FbnLaXgQmXZvJ8rxLXOmWLkYELwN5fQeKmkG9GmsKz
PoYWc+OmcN6390axKO7wTNahkkqmWVxxc2j7sksbjU2YtZrwh46fEBJXWNVLnqZ4KMqEonHuhVzw
ZGqYCTcrzwRtUcYcxde2ZY6bdUtMhUVKAbVcGVA2yLjfj5VfS0NnaRyVNLbX+ltQcHz9YcMJBYju
dx9IPooY8BglmpN/Tn82pOt6Cnq/Xu8LmmOGpyOVtKZ59Jr/YIzJs3upwYHFTlQzUAmFCz76gEpq
Fctt5eDIZ3ROYuYuz6VrhcyMKuZS9tiX/xO+Yt9G1bZc0RHr/0rGrXc8CodvP7cM0els8yJ/2yyl
USa/Dleroe3G96rNwLfEVfHBFO7yvlFKciKc7XD6EQX39J5BCH67D0/FCNno4cEvPESKTyr/c/9X
XzqnIoosodxpHYH+wPs3MwOhFrSMATBPTU0CuvQrNNNMlkF7uEL4u964n5HZc1MOz4C8rfm0j5LJ
fJw4nO5/QI7vySW3Nhdb2VdeHMkZCNejm+0EvH4tOsQFX0l58R4y6wJ73CIgPtQXtoY5W4rxPhNL
S0+tF3IMjEbofsNhwlblsVjo/jm10YpxRF7+alBKQoB6aNN7aH0lFGg5Is9ItIG3pTaPNJqmviP/
m/2DvAk+Ejq4H+M4dbDigDO+zbp8q8yj/eEeewBxGNJg8y0p8UMIAUndikM8PXX4YvqMO5PH51jz
Bli/zVxBnXyOAruzwC2PmxM7/OwI8MzC4TwPYyfW30XgRuPu7tl4T9453ZSdkMZcymVAsS+dow5j
g/jShB1SWdOQLkb75fUVM6w+SXsZ2fIrsvd/2J+KG0HnjtqKyugnswmDccg594dkpyz4XTDP5Gof
yArNdZEJ4WeTaaP6iIlYRlZUNcrs0VF2h94BH1nsYATEU/fso9Hj0o4rLoSZa3yAC+a3dTD1b6ZU
PBtOkpfSVYYB/qphjTR79HKBc8b1T783VqCYF4y2T5ir898RIIPxgFsfOq7KAI4XpbQ9HEjozJ9J
xAuF9hc4fOQuVmeoyb95qpPk+YRBv0++mPcwk57Pb1IkMqmOxy0jIoZXFaXlOSjRW/GoEh8QO9kQ
uZndI9TgcyQqloRK80fuqPr69w/hGbimWScQp1TzKWmjEle+WY1k6/eYmxCHj561n9DvTGZJAC+m
BoPY9HAQdMAi49Ly3z400B17ShGq5ojB5kbPVbmhLv14K81+pk5l82W54gXSCUnAjy/0Dh6b6Bax
fvsDhyt+9PxjagRgwPSjGlN7Bt7qHPivnWnxX5U2M7N/NqWiLObix3ciDA62BgIxaewT6HTIeCJK
4kXAXh83XNVqS1TyB6VqHWKkMbIvHfIFHRU05vfUxWCLxcTYEYPANqB+o1piXgzuJMTi8mn4t2zi
hAbj0iyRKGw5J4N2aB9gS1vc2OsOkWrNXaRQt022ln4/GaytEf+0jPLw3CZWkegZygpFZdaIQoz3
t8ZZhls7AgO/viLaIaSv6p8wNg12NmZe3SJNXAF3Q/LrGEO/449nQNIu+9UU/BkBcADajXM32rDQ
gPNTfrvEbktajl2yFhGB0L8f8yifLW961WUAWWIsdEf6b//wT/1SVJCxeRZ7/wlI8rXiiAWNmxcG
EnHwUYD7mnUwPtnRvUbvzUMTlsrk/ezLjVSQq7bt3/a3LPJsUmXyZ/uExJ4eAygWAJM7PGP+VjvJ
aPLn/AKAnpOxBwibQI8PbRTF/mWzCoL0DvSKrAHtmi0YThGQosJW9KzyGTaSNGDWrAnlqP8XZHch
0+ijTLVjZ3vioNseGoexPGLEwS49LrmVC/3SXNrYb4VSI+LS+FKI9FPo/n3rwbdu+SJ/8SyzloRl
ioX7fsaMMSBtJnT4L4WdDVpsH+izdqpK3Q5CR3DdRineyDmrrXZyJD1KQtdnMzFV0e5OvMb5ZFDP
IUeh7C1OlF/xwyifJUVEQY3l/ZceW+TQiLY1ph0vRJCjoEyxD0+95xSZOMkYnoSE8Jyy8PBPz74E
6xosenVFPVRWRYTOxdmle0AurDd9dERxdgq1pNyfNjykzg5BJYOD83U35GUxzzy7HlYRf3sztjin
s9w49Z6+yUw0paHN6UtcIGHkw1x3bhwoU6FcTRswU/AZpuhea8fX+MU+H9iwUwNaSLgww+LNXrnp
qgpBiWKB5ETllgJQT8hRvQ4q+NNMHvjEiwLnFurNtFMhvKSi9fM8/gg2l0eNDRvrytLXxI8e5fuw
nra3JV4tHfqDaRqamvrjba8I0wH1DH9SkSEWRozXgNNNLg4f2JIeMGkFp8UV88rjqJYUv5pWuvvb
vZVsnE3+Z+PUfqmO9qVwCfVz2YWDYJEGt74u1uLFrslErjKb8ZXOseD8PSQt2E19dllfMlCrLPLN
adSGFrIi7IbVTjVCiJXvmJ6/e5n7rC8qbRyExw6ZXfJ924b8Q8IDz9JfStkPGnnpdmciIISIF/Zh
KVK/nOM908A+GHFquHbHkMIzf7bySzLsE9VTdl1UP8qbpjW471IE6VP1gDx6w+Ra8x1lViITT5b0
NA3DTHzpCLb3aQJUd+bVpkcYsm/SUebcBnMwMJxydmb+Sa56KodT99PGha3D470a3wFsV5Th694S
PflY+HUZsOHrcTcQObMaZ6NAJEnnSR6O8nQ99IPMQ3/rUulBTawubO1PFN4yDtjhRpCjL/W3s9q6
iMmfDpN4USnZLKPaOeRsMA8UeYN5qs4HzywUJfPU+QpLCqmHoebTJ1lU55zV6e8cv+h+QA7bM5gj
l+mNxCHjez215vlmwHasRaipL/X7SmKzpVkE1NZUINOeimimHKJaErbfHrRN7IIQD7bXimiHnXjE
bReG38caQ8GT946tt2bEizufzLhF8kB05k3QrxbclAcz7aO6cQN+rcysCYUO9l2ICOUOCPMM6zTK
dn99ujQk7R+le9aCTSpm6jdkxcXQWrWy4fcinoUc939Sn1TE7jMSgCz32i33tSoqU8woLVx4P2Wo
beLq13nn/cO2UIrzd6MJYknR8bYWu7n3YuCBQpHygERd1+txbLZaQZY7YZzf9AWyqfn7HLhDYXBm
KGMLrHq1XziNohh85bOgtLQ5wK5fbHrIkWsKfSZve70W9QSa6G8DyfrDQac8sZNGodraspUrjEOA
wrDN2y6fjUWY8qpkAe7uy0EGrst7rIwLdLAYcVjdlM7eEC2pcKeZRbAOZ1xxPdpSKiKZarMBiImh
zj9c36O3QCxoi4ZRKgKTEhGwcpN9vAfcHE9ufLlZfhYtGl5/3l7frjl0FYAEBNjgMqxjGoh/CCaJ
JK2rbL2NxCSdk8jFZu0dE91PIUhYiAN55RJ6mUShRm3CwpGiogBfzS1TMad+iUk3cpKVpvAqca1p
XWhVBHKHNk5td8kVXu9+aKun5y3rVvIQKl4ykrrrIcP83r7UWi/SSmXEB5D9Qs2aD1Ho+S9rkk5y
8xKSFvN/d7c6I3NBXy888jPS72dRpwnhyx30wFn+Qd2Y/cwJT/qcYiplfzrlZVY/ZIk2RB56oIc8
3TTX8QVD6OuH2kRh803F3joQeq6gVyadLCDvooz1awLA5gs68revXRhRhfC/kh0zZ/TdNiOgs7Yx
/ZzwO6T41pPMALSP6vfc+y2gPCLVL82UMrw4hwdIJ6V5xJvis0JOzY/lxKQPIU+6T9lUdDoa1IsH
O4AqCJHuQ9nsHjRkVb9mAqMCFGjndHIAFnuAF1yvgixacz+4GLh8czIn6yBXQWVRvDV3eMmkwxNr
jOGgHjiMLcznKVVlwkxUui2hr5iE+LtCMaXVlfqmdObsm/k0+fwWVhvqj9BH9xcXBRbkQw1eMPVe
V3iqFBHU+A/cqh7LpErZYPVLyWMJtear02+0kNqAO4psa3V4OW/kjdNG3i/pl1BKbReCbwbXMzWa
JpzxL+wdOiyGZMN3GYKM6zo2Wg4XmIrbHXWn7PZrsMYWoKnVL1kSHJ1PrqiMH5Dm82MPUVYA+0dN
91KSzKrIX7PB4LUWAOeR8K2V+xyROJTLV25JQdaDBM+zqhPwjAL6IEYS/HsPuUe5mIAWklEJY4qG
YGUTyUc7CDOInNJHa8LQfKuFGQwKUgOfPi4bNpUkHypGieoJBMp9YgVR6Gh9Js0+DC84g1dsIrhj
/XYp2LumBWI/AblQFPHm0g5Q6me0RYA766bHkXPANGYx2Wx31H8nl5G7yhvwa0vDkLxTtcPjW0H2
NGxao6AyUEdLopHP2N7Ax6L1cwrkFJZTOjj8BTr5vNbIuwXAqOhvVuvvvKliwnevT8jd5zVhE64X
n0k6+RVOXz0yFhqDAThJ+MBKGvRF235P6qaKNMedHfPS8as+oVkg1gmHQyWfY5O/DMAR2MCKtOT3
0G2jRI383Fvs3Y7/Jnfve18zv7QRTpi6boZiAwgsHd7HIkYzMOxwiQ9V1NDwgqfbncB28/AXTpWf
OWOpiGPQRRNyQkMB0oeluAOyySVO6Qw0rG0c2B7sv7USdXmZhr3tmnzBKBldCaPz6OHgdCF4qEvl
7JOdgh2K0slcy3Q6UV4NDOsbtzR4++hhWEKfcjK8hfybxsU43Hn6HjzKdHpemwY0/9rV+ZynRtkR
J0vt+qkNit4DjYFuBpQnXr/S/ou8CU8pRzbY1tD9QMe8qTnoEGvGpy3HCFREgCTC7km5D8gCb+47
tE0sJU7xhBKjON5EmOuozzNCfe9WKIPM5/4DS/YvZM9xilQtiB8yq2URrhuUmJukdA8j1sFKrCYG
Y3Zc0GK6j7pzIpFVELoBgGyQrh9BICLIScsOarvtB7yyGt4Js96L1PDKPHPhVluxAsphVjz2N03Z
Tr6y/RAnIrhXif7fwXWl39M7XS8QUKz2RRz9W6XTGudEU55nAMtL4MfZ5QnRK4jrgEJhmDVq+Nj5
K4eDpIB3tiPC/grTiRPn5nQJT8zXD3R+olNPmwC0vZY5N/DX2PkuXY4EY6cCxAt1AowPExjNbJFK
IeGEqAf7MXg2+zdTi69PCm7nXjkWHTkbyN9ep+8w9ru0RtkHowuPGMl7vA5BQHZpi2q8zcSJ361r
nmaDW9NAAuFtLDi3DjJNwz9I4LG1VFaroguXSLkAsiC92ojbhmqViSW+s6xW4vEcf25kElQvSY6F
xjiGv5JDIKwyv6xq951GpQVCVVPq5jKP8fls3WQDt7oXuR5gvtDVvyHXFmEVQaR6fe0PICLfQZfk
kexE/HPyV61PiC5HiXZkk9x9R18FWD59oTfgImWyIv6WztygyQfUX4YpXCCY/4WNrlPV8HjRZO7A
vQRjMvcobNLMPdup73mcG2MlKQjlCX68YLMbw4Gtzwb1d8ZS+229M1QTqKS3tPZZQ7diI2WJqMi/
J1mkvDKqLrg10G89/MLhEtbFWRg3DSd9xIpaqAOG9ldPRWyauQfjJSI9gNRZzlFpH6ebNMg29iUy
kgEzuAoNObl1j+nOkbZz42OUdUv0vgXcqOie3NK59Yl2UCy10YOIESoLNnPSUserQCIWyg/YEkDh
dz5W6knr29B9/fCi7ACHWOFi+AKBUz0/+zD2cubD1SEasCblBYp6AVC/p77sUKUtDNKuntycj1Ob
VkuRKJfw4t0n/P3WyfPvUex3ajNwmNg2aR761Cbi03RmlONHKpwx+7rGCCS4V/RsSQrjtBR/+GSL
L+j5ShIzMSF2gcnBMky43nq0BkLoMc+N3LI7IGfTzz4P4uTuLo1DvXts28g7SMoJgb9ZjbzaZATs
trGUk8WJTaHsGxlncOznb9YTut8+CWlWJVYVfk450Z6e4eHS5o4pZ+va23Do936WCm8dyUcTw6kP
ZZxnNOu1mI4WKvbIwfkc71JPcQ4UGwOOLg83Ck0ao8uiSsu6wPd3NZ4zVjhFS0ZRQY4TLqu6OMSt
LWBfjqFYha88UO94Upa7yhBgmWwgS/l3VG4rOfsn7O6P9VTgQ0Lh9DSjS4t9/3XNdPvm/+8KqBkd
lCP634WPvOoGZk00TMxUF+Aitq95gKCrsN/ArB/gsGscOPO1L6ytvkoHJbm+STTvUDJ2+ggGr+s6
4320ybZuK9l5CaGhLFQ83FHbypW/Q75aUWFhUy2t4HFcByOVEerQZz7g6ycZbAQUBFN5wVEL5w6Z
MatgogECtoMHqw6ZSqPUKTD+efpKhfKS7hDAoiGU1ImA8eZJ4W4pv4bcfBvScpWu2JdLMVLmCMPl
VEP/IPjKXLnX0fdZmm9BJMxkh0ugur4TkQENOPFviVFS6pDNoxFE4gOGn06AfpIZllek1ahoGrCY
6jrO0Wg9OlVjc3BykrWo8ww9A74xbI0kyFsdPPa7Wd1XajlnrdqUI7bp2M4rTwTawuDhNDGdZeKZ
3RnYrgowKAZ6u+tsoF/8aZvxHDY3/KwDyaFX3x8JzEJzDWfHv85w42xPclVwyZWPlYjtI79nxK+L
K5i1KAr27G2oA1YSWuHBlR3SZYJkPzimEECgPLxmVfBFDgLp/b8Q5ix1LjUtQpydXNL4uLBEUi3a
VuWfFqt9wKlNuegHpqZzbyo+VE8+HPYhbOy77V4/Qg1p+2HXtTgtyrrh539RMOrHxzfr8t3rrDlq
MhoOxBRGXg2tAl5D9NIwVAJhqIyr86thXMKyzvt9aGb3+/YmQvtdsoSB4bUl9tMnewqHDpZP0Vy1
KgaRTWDZ44u7Izb6D7ZCGBRhNeWEYgcZiP/C1yTDzQcvyQZUqmstEPIA/n5KoGehPHjWTUoZxUcb
8yWbyFBG4a2dGOlB02aOeq97UP5EkjstjTr/b7RPC/57OtpApfUfBfCORAhQDYYzpTu2YcWmRktT
VTXpWhg0dNA3opfJNUogojOtL13PVPG7z7ar3Tti5mzRbyWa6oLhqJjUSRfZNfcKDIwCul08bxlI
QKT0byhnV5TJ+8LH1fm2FgrTvNUBj3xJCkY+t8T4H/MSKuIxkT7DL1HyWa1KAp+IkCbX9WQ/yvmb
OhNnTTPTSNJ7ci1fk/w82NTEAS+v8xF/6jyr31E9Zp13AFhAECabkl1mnEtmKhms8Epjm0dhzJ0h
OHkEQMwI2nN/RMYcZSYh3xSOUFkb6+ybZ2CEV6QTX8cCpzA1nUiBUjm+2k3Q+htRXV20HhSl4G4J
uOBoPA0IR0oANFYAcyRvZq+dxggMs6FiQpTtOEORavmF+ZaV0fmhjNu7l4dQ+xEDwINlYzClHRFw
X0LmpvTVeRQ9U/usgiaplYhFra/8DX5l5EizbW524mSScJ25cHShTZWlk82oXNPTZcYlTEAoE17Y
3Sa8UjznI+GQlrJ3BHjyLyrRVedK15YCtt7niutdVbokhV4ldWNFzNkYVYni3ouVmk62jVRFAkFg
wb8XP2exvWsoBacMlWNI1uYLUYUBi58Z2svaGAI9pgIkY+d9jDPJwODOSfLMDlMpsQdf6TGgvfRj
7xNkmi/518oEbGT5EZh+ae9GQ7B9zJwfD21YhKmjArv2WEUuNkRKjb/Qj4D2PtgKtGcHI17C6bKO
nHhZ5yubK9GHkBuzvbm907MPZCffTyyXFiulPHgQxgYFZVprNwmYr/wbLfme76Kmw4ntJ6Jid9cL
uA6ZRoq/lwi1AImtrWxP0nUCbOUl8CoEyQvcLa1+HoT3LtdIBnk7gGK2g7toeKUesuXJD2GrDcO7
OkXDMEYjDmhbIfzLod9oNNbYeOE73gliK+MtrPV9G0uNeU0+eJ5Gz5rCYj73Nr7bUT9OPwSptNZG
q9V0pIZDDh2SSDU4CeQF5Sa4b9gjY9IDoyfUl2CYG2WoEIgxAGiIybV7JAuDXxawjUAGcTksU4UC
p/9MeVLrZYxVrG9tGSmnjWIjJCCM5KCQ05lk+FB21XZUknf52sfeDselYra6BBs6HLJeB0caupSy
U0mglq5gyD0D0jcOSKDJCoWG0FvhTmVsIaOXf5nnD+rnOs4yipu/z/NfDJsAoSCUc9tgUGuuLNWt
2nvaDr9wsjFfhYEvaGhpAnqS4RcyUbG817KBWtpPdxrbJGTdswl57xOXijPaLvWdDczv9mUC5xbm
U6bnjXZ95VpRJbnb2FXJorDwGvt9aAKWTwth5Mqa1VH2fV1JvOrLPZ6prZUF5oriiEGL8HpV7boK
kUVCxHEEn8vd4wkpz1pUkcN0idF9Lt8dzVgyCdrnHUVs7kggTRGLL6frtbuYz/tjPqUduvjA5dis
1o0W5A8meki7tubYj1BQaobNmAv/G+S5n73stgg2BQjDPWAjrnv/w9v/zvQr+pAH9/WD5lVV13id
u4PMJz2ZGvwN8uRnPbM7+HV3sZSDno38ZeaU7Xd5GIFByV5Da6JiXi9zRt1VjXQyiysQfqtBKuxL
1MFaKIzLuHKIOvd2PKQyA8+c4BLLxQMuSRZwxmiatVf+tGGZo1suTHw0I6aIeZawaHWti8+tKVdl
tIV8KfVpkIg8yCRzjeqzx55Hh0Gu+FnyzLnmGF06aXb6GO3Dy1VhgxPcKWl//6ujJQJq+9+ns+e3
0/dcVuuoKSJjq8wxw2w6H+dwFmIlVHMxfrKtaP3yGxcAR5ciQ5L1vGScbyIZR1WIwNABWsKzMJmn
7HMeRvyQDUhdU66wADDc0hxmvLXcxIXy8CsVEAwwla54+l1Qt9Jl1KnUkj0A6jqX58wr5ijt03i0
lLYsJwRs976Qu9tWhtcG1I1PC0H3L7h9+jPG/nXtld2g+3pTiZCcnHmPq83IQApYk0ZDOH6UmDFX
3P744ikHMmq1VcKfxQRqMDDIqFmB+zK2LDF16dC0zQEcBs2ew2DLZzjsSjmSjsXiw1mB7fm5f8WL
MpKlT7qFP7bRw945yRUmd+yBdRFqy8a+K8CSvlOlf4AI9/Fww5LOsCoe4d3PYejyLICb4lZL0Scm
Wd8P63O5MyLT4IDQ8/42+MvbRVg10DNrBDdMm6fMjptySpVKfknak7klLrOY6VscxDIOs0RQL5Ro
fw9KjluzlSBAgqCoU+IyzykywJvOQOtKBYIO56uzvEIpP/hKsC1uEtNJ6+5gSP33br9IbeYTMWWs
hiiMZTKSk4OgN8JC5Wvo4MQLkaLj83DE88RwzKgvnrQI9iK5HFDfmLzdLVxkgB9TbLBHqAhjlRYG
tR/poqAOr+gZSs2yTadglcmWuIbWetmi1t+vRMlWfX+57WT1hQrAH2JKbOio90aXBCnKwpeT8/x1
1BVl4JgEOeQhAKqKzYJOYZKO7DJ7HVxDdF54LNPJ36IeOvR6uMR7M4Mk5XPsTOnjBrIQ0KdCQEBv
uV0sHkkbV0N2Cv+mYCTUDkNfYbhvTP36np6m9caXD/5wt2NWej0RZlmEGC501SQtIUzQRCynHtzI
ilq6xWWHrdBl3WBpUox8lPxNZU8RD7OCC09YzSJRbJaj1qlFqrQQggMcdD17daakT1KDON5oou1Y
EmwS/bLTgVFtmVDnDZSQ1V9PF5CzmHOfFMQCN6pCCJvE+bHd9sGmqSMsF4knltL5qJcUPNfLgDhy
n7krtu9wrXQdHB7CLHTSjs2U6VnRLIzHWLU+Cm+n+rFjLGbeR2wtMr254bAyuVeZ5yWNWJ4yiEm0
/T7iovKwhYdZ+QgVzF5SBnZ4Ehbz2QNot4PDZDVscHOFcWD7v1XZy6s55ofG5igFPk7x/MpM8q7Z
j6RTFp7uXcqNO0BzgVVfbwVxRHD1ZUNJRjMqa3dpogvVvupgb1xp6IlkpsDQArch6NhGjPLXMJ8w
j3h1q96dQJB+8WMpwrvmcftfWAnWyF6BVPyddJ0A8QcqzDOqX7Cu0fjOERf7LjcrNY7JWHrRUZp3
Kj3MXGq2GdCpTOH1kXNnSSLqwHFw6R7wpTTZq0C/anzRaKGkI3N/80jDlP1dZ2Mb93CjsKuyAqFm
5yVLIwMwz646QKv8ZWyZaJfCGhBYFt0eRjQVVo4Cdfb0UZ9d66FX1chZQA1qtgwQHKn+u+K1LeXe
MIrJ3vCDbIf/G2za7IimAymbILqVWzLsNEVuLmG6sXBK+xIq9Ewj93XLKGVWmTA+u6ljwmXHqjcF
E9M1QpoEG3H0XzVhiZzh5FpHPF3poWw6+tQjLVTmZm14XI39jmtW558tle5w2UHycdAvQo4l8zM1
SnB0t72iGEgpteRwQ5iUFnuq1j6/u8MeFnChnB3pIkPJTKwAfQ+FN2cSQopZbSIaPAN55UUPnD4S
WHEVgAeEEa3QjuS9tp+/pAlwsQXtnYy0tpzc3df/ZBcDN9ycPceKz6lhZ5WdHHLieTtaViARVhib
0XYXaIIIVSRhjCaWW4QGy5I2vrmzuBiZefqXpDkfDg3Gaz5W26OkrC8GoXrjBM3iy0/SymfUt2uO
DBlxgJwPhxJQx5HbBW1FFHIokrb64y42IK3qPaXIz/sl42SdEuKBxUkkvVzmuKWFSogcPGDUzEKl
sIGP5L5J2wvswSrDMlUcRMmnpb7vzE2ZJ8fjiZSGwMOYRn+fPJZsuJWZGhrBgAp9oD0odj4WVoiq
T4Z1M4Q/MbukvoQp3XSY0AFPy0MnkjckCfW7Ld9OuxApaC1OCNhamCfMFHa0VegzKJJG0vZqd7mJ
sexcxTgB3nuiUEtz7hyYIcgQGKB7LWrRED0rFVeIMqScHAQhky9KVLPE3/YAu74D1AQBuYdxiLq3
wx10PaJkTxfpkK62zQk7mBIRbDGQyKSBYch+WrVJSmp8Nt5/R3Ib3nw0I/RoQJcmzTqLXCmVVlaW
as+uxr/C2x9yZ4weMse5zdCGKLLRtUBLe0t8JAx3CedHCMHhNrmZ2Bcz7pCr27hy0LItTl2douH3
dkYTj5ZIZ9+X0I7fg0+aHCM0RTkjn5XtMpQ0wK+d1WLbm0arXu2WlghvAiBSqopzJ9xHfT5EyM70
2HiEWvWeSU6Ixepw4yjCVSkOaQj88q+GSTTUwv3el5xeoOYLesTrwTIAdoUcjiccN92d5xh5ySC2
HmNzlYp/7ofHi8ysyxkDS1tBbNGgBuQ9dz6YQrtotRUUNhzOzC8SL6NJWCrs32KpQtP4n9CJp09a
U0Y9zm+qnjCpoZKDu5sUSfo0EAPUj9ksE0nlGfVTGKIjkq8Yx/LnUfZp3vEHNE1Doizhr7+XozWO
XQ6+ACAtuJW6lHqSfrC/iX/f605oQBMuSX5/5lKioEt+mi2ORe3CrcGbgWKEzEzVMrPvEF5kG/hQ
P3/AIAPr0fKcJQSGdNF5HSnqjqz2usE2koAEp9CGGKjAHfcqQ6eBwyWHwEnizR6NkZWmqjxWkNIm
OlGJ64I9xPXtDaASb5nRN4KAVKWbx2X69UM1vxVIhv+xU0a2CEbysbwqDwidFOJqoYejAJ+zAZmm
fFaJp+d8qetBCQLBqaAE2iDw0M3VjFcOaJDC4jOvyGaQ93L8N0IgPayR8XTfbTlBUwJGqsWWaIAq
dWiKZI1o3f/ytk37Jh0PMCO+66GjFvN+yBZwXLpkRZD4TTakhnD8/fKM3yQXbJXiTATY1VQH6v57
BXYvZcdP6/7jubDmoQc8kQTLC+72IUX6lo6ByThZrGUJGy3naNVYr7MqNKPQhfF1/nsEotW95k+j
EB65ONJvOZNkaKAsH54g6WTDrKqmiAMUh/jfdLImgLjGUkJnlczS9NGRQrxp8G4tL5X1JHEe6NAT
94h3/jLu8vvdNA6BPVkfi5LxG6abbP9KsPsedQJ0IAOa8g9Rjjxvxjdc6yi/9wE6o+iXrxnDaDsj
UWVDGE46cjXTh/WPMXUMyWN14jz7nEQMQw8yN0UO32TMkmoMzLtrp/KPGqWvSvzXlRVSCVxUQm6b
7k421/HzvZKiTZjmzAmAd3vi/+3te8Ed3UWMFGi+zPfXf1xCP8DC2ctnAdrUfbq1HL6vFtT4Xsja
yQqMkRvpjUC6vsdg9ImnCmvB8gGGpv6S39vID2r0hWazdYXjvy5l/P7abgdDe4bnRw9LKsSiFmg2
lrHl4M/pXJmmGRZC6yBshxBAOU/c+5CQF4kq1tBD2laAjUeo5HhEkimRPmtJ7kx88x9PGf7LpEzf
yS6X9d/alaUHupEnyMXkLvLtd1At/SNSqhBCgdBb599GoXw4xWqm+D6TU3C3B5jv8uy+cX11FPua
xLbbvZ8v2PwGKRUK/pIzTppQN0oPXMtXau0Jp3xeJwn/5upQcN1anFGz9fmCqGc/WtMmT/a+Ahg7
bYtsfW49hQkgaOkpaIOMueuSJcYLM8AOhiE2DHR+CNPhG4VzkWnU45/A3BaxEtR6n3v1yQqSYTXZ
k+zRiT/fH/T63Bqr8itPW9MiEFIhCb2PifrCyeLtFnWlhZV28NnFDQ5bEr9YyLNSLTwVtOq2A5bm
QBX37hVKttLG/Cz12HNFPxBGx+5SX3TjBPC/Yc+JCakmocqTViQ8b+/7PHRrCfhjLzXLH2vVXYTz
xd3WQxoeKropGZuroSk+R1kSIW/KckeNp2Ws05hL/exT6LP/emNKJrCxkdeNNycwQDv1XPj1j7S3
1hZEvYA6fGwfMRmWpdQlJCv6FcEsfdv/pmb4UxrB1y4PxCkhDVJ6ZbILYyITBH9VwCqN9BB1IaEC
mt8SBWtglaQDHwHfSAx8gTjgyPR06NxeOjvxoqJujmK1Pi1XzDeIzZIPjfOAliPjzY0eJ+MB2ZXd
UxXVV7bxDq7U+K5fOHVyh2gw02Hy4+6VAmdefRe7WeoxDjg6bnk9npK4W0n3Q0LIR/GUYGC0vhi4
HdmvHkquMxF1DCzXERUQy8EWS4A2dol7K7x3bZJ7mNDtuQ/N62q7xpxNdZ4JAvMn/upsL4xDWuoh
XpHR0SzcmQ5aOBaUOaLZzlfvjy6/TMmJ9FF7OV62lQfUGXjNowPVQTDPORPmtVoXcz9yReQYDQST
hGD3N/5GatYUPTo9EBXgdw91n/clNFHANMFFGNHGFF8m94V7DdUvhAuFBeCqAa6TrHVkShSTVE9y
bCLY/KpvqoaMaWU8yrIuKtretezMRItQmTyIHZ200hb/WE28GfENMyzDlRqLccP40mDcAwnjxVNG
+F6xKw3MeNzvN/5pSRBEkaVwZ0BVyDGrDB6evise0JPPf9yn1U27ZMKq2yD3xho6/wkWxlsmpGHC
CXBkw4lOJq54UaIVzUGE6zT9H2MQtosAKXOGHnCsYV+FGsxvI8T8fjCeVnLXMaP7a/ihfQuBf5MP
YfXr75LVgxwIM41W+xCO+AyAp02k4nXE6t3f6XMxe4ij1IUJjB4IJSyl8kGIxlhJ0FPmvoRVcLrn
r8GX+n8lhkYJYKth0DKTCVmtyfxB9qI56gcvSIhHn/QFo/lZfydJatVkPUsTvgZYOdvo6vzOqbC9
2uPuwec0bbzpRv76dknMpKDiMBSILMR5RtKCUlLSnPIgbhSS/o+icWFC7c+idpZVJ6Xps3yiX7+C
0KUD1tbw8NuwTmPS81QAoKBw8x1+FPOp1Z8Rd/mgsIkanZQNvlMVKYc6eTdRZoFOH70fr6eSjjdY
z2FywLmEjf+5OTiKAYf+5P5kNAdGD+ctKyPTWZzHpJroTB4LR/RmyESiqovzD6xSPStPSk8louBl
foRx+S3VJfn/P8tb1qqqPZtMb3hI5QTlo8EpyCrFwPFIvaBhtYVqNZstDJm7opJJH5fcP2w9jh6k
dp5SuzsCLg5X3TdAcPJDJvzGomhJrOFtcqf9RBFgIEP0YxqbprtKbq6KCApesFOekJ8in6BT05Yu
92K6Ky/Qyof2zBNwCiWC/8bFxOIAJ7KP6KtssmY6+JZ6ZsTiQ+ZgXsF4FRyi7s0ECHihmQaImzZl
QD3X8nKqF4piv1EYoPt4wH/4KDppXFinQVvrIgUooJ1AZiwMV7AmmMbWLk1niVeMrtpoKKFNUrU2
ptw5Ogvm8QVZo7epB9fJenFtMug3UhD0JD00UDFgX+gbDiKWg4DRRvxss7vHSr62wyaeyxbtrCT1
fvrOqZA4eCt5EWle1uSzpqwY7i1vb4Su1ewyerDN8mrklDSkFxyR+ggl6fe0CLJul7H+1IYcO0Fa
rMJY1GpVY+xjoTgtBYYVj8+Z9EDNzfmajIU0CW6KkmC1PXSFemJV+Q4sXF5bwqEFd90xZpdCiItS
3xoH5N76phh2NA/ESzST02OSTJK+nd3jHS2GbBc6u4qBA/b5gzRNB+uPQDTX/8awvXTnQ8s2H/LF
R8YBVriJUQ+OND4WWtbzB7RFCGWew9RdAeiFfL4CDDRZmVDrfjORakbAvMXTvfrrLKJZoaIXnGN/
o77vnUzspLvp2DuI2XEYvScJUKRGZwDsy3RSGgx5hesJbFPZAU34WPmKfAjcaCR2RQ1H6K/MP1WH
KZyFI1/u4B3NHKRMsAlm4QoFD4scvtHASv60NZ/aazhu1wh1SFO/3S0LOzePA/0rxNllUv61Mg9z
aSIijHbERuC6znrL+fgC/RlVggho+Yo38uBRhaDKlo2hnrtvVGP1B8hnsgr3iWf0AgYQjOo2jHA7
uiKzA/qy3X5B+q0haxi/ngwH/rHHgNaDpe2ZP7yfP6X6RX/SsS8+2IGxEwySPYONMz7nbqVXWidP
dkVc3V87ngcQG/bmsoI6LpN969isNdO3N1mqhsfgzknnRMccOs3QoC051+VakfBBsTubwf31rZ/C
FApj0rp1vNhDiFRKTWJ1XrOIeKpuzs+9NqTnbDXUcILcUO0m7HbPeuh0hTmMIn4r4xvn9EXlqoi0
g0F8zrxwTBh6tWQp3/27MptlYaCNGZM/ET2wbUPEok4pHiah6M5gmO2DX/ZTexZug1RrivtxulzP
7hX+5iPpM2b8Bed8vDUQZtUz+jXDcYugOW4GDlZ1RewnOoklUjLLd2rfySnHckjOorieIJ8bPcQK
h8I7roYiPWPAWgU605ZdHFh08FnSf0M8ysQEqyweI7JN4+jsXpI6RZcDA//M/vbf04gsREeNFuTI
GhstflqbMOh9/k1qV/Ay4R/2YqAnjByjSttUIXHi5L55pzcB0ZD6bpzYZg30h8wSZW1VnElrSnBU
FJuV9QzbEattzUDLrud/AfBd4QIrguXSVOR23odAks6DL3aeWAV+yi++4BSRJLoOqn3UMKO3X9vQ
mLp96Qz3736ms9NC5Kil1Q4PMa08Bsl94wsbQnlTW2wBGTgDTNBb2URyUlQJ1ibt9MCbg4l74MTO
VST/LRV0guVXLqy3Rqb+i6YQRg3WrPgSjdxhsukA5z+RiYerIfPqQ/nP+2yNgMXxXh0dhzwE2NEj
5GtNyDg7xzwrkGm7ivqOn8wu8JObehbO12cGSnZ/N9Tu0kbk8RcB14gcqcQFq6NDu/VabT1vwaf2
xPCB+4ac6OX7uDz7C5NsmvbHbbPAq2PHdmksekhkxdDs4DujtdXDyTExDo4Jeme7Z9cU5Sfr0fvT
2x5V0hvmOoBamK6a3kHL+4qPToDp4rUOstHky+3Kju/aZ1/FPp/Odo4AeNqx+mtYdZ9mAAiKvNmI
tRSFRR83JLqnPPzGK/iNU+n1aF+RC5TvVUKUboG1WYA4rCJs7mj93jfYo+rHvwe3F2DKIlAvjZhl
JlsrPqHvBj5JYW/Zo7ylqenN8lTqFU6wzm2BjenQGdCkiuM2P6qlbOlPOGlxAkDjcsqpy/6VvXJV
bDnXvRystI1J3/LNDEJcC5VIDNDToTVVefnFJCoevZOs5keBrUQI1QEmGS3srlK6tlHmVYSoa08u
3wZIuct7R9n9mRLdwkvxljQYMTjAFsO9vtnjL53/kMD3mZTAeb0+OlzhRs58S2aYEr4Xw/OcJUTd
/YcsRGEvk4iTedNR/pYRQfjBwA5wRjw/TK+8nmD+W6FO9AOeL3pllubaTgJCQGKlRYzBAHzeIxKq
Qpx452LC5PE/IayxKzZtLrrn3RkODrYpjO0SaI4ZJzp33F6tdMVbl/wIKciNB+d/kda47vDK2S7f
4bpiFRQqjZOr2U2rIyMiTKr+kDLL4wsqbaaOcTuOIIF2wzDHcgxaLGySnRsiZXZzcvJABLKfWKXp
RXJuEpK5rgtYvzXkiZuFSRYrENL/NFsKbFG8sTXcgcWzm0ZhkCmfumgIxhkZDKCnGF5he+H/wsCW
TmRVDqM24mGQYcfePiYfX8UlVKHudwUN58ueg02SayoK1TZ6BSDQO4fN+JYkdgxu5tFMWKM71Cd2
ur5NodxVlIdAjMN0b3EQcfVl41gwYgHCaXlMMQZEua50FkXd4AWbFgqfqlVCyT81mrKfW54vZp3B
hQtcGt5YOhzoUhIe0b38+rvkZN16rBK4gwrl9/C34aVCZX1tScjheQ8wPR5wDlPRXw1o7rKnf1t/
DhzWv++A2E4uE7PoeBZW2tjNhgrEO7RmfNrE0OF9TSHb9P67c5Zgsm35d1Ycvbs4me3NQQnT0LNd
dqk2XN8eLQeMJVxsoQIW29iyaIE7EwBbtr03suTmYYlXhCzNVBmlUVFba2qy2m9MzajB6buM7HgM
WF/oiwPUu14DwLdbZsvEFvrZODFFcx/muuArEv5RpRHmJW2TsSJMTrdIkHAWBSwamgnK6yBV3bGj
5gPGlmeuHg35L1sCKyX1MMjDKuYSlEs4iOEOrUznGPgaZZcT7izqlbxTlVXvk33cGojxP0raVc+C
7OYKixQYKLy8jJ+iijCGhNTh/x2XeM61FCWfJzhmFOIhKNvbtJgFKaGnZ2a4LCKuYtbnMMBzaFlr
2jJrmRGP4dlr4h4lRVBwTxcURaOL45oJmFD4TjeXGWeClmcdW1I3JBf+OKHtdoPKEoRSz5QzI9hc
YH2f/jr/VIpyJ6i+RnlUx/yr3J06t+WXH/w7m5bglz8jm8n0U+jHlk6gR+WyBqL2BG2YNn9UOnq8
+GwtSNvqysE93/LxfS876tatIKTtvVDTC+sOW5d/pgj+1DlTgoUm67wSQIfa/lgO6dxCkZChxSy5
VyLAz0P8fEFO9Y8abNazLcx+Kpcq913H9jYYq1KP4Kqi/rbl6XFwO7XGCSzbjaNYrD3TBRBW9ddf
/3Kn/fmIt6WJiQ35tVs0X4teSMi1MEQGHXM9DFMkOi7F1wz7YnENGI3HaRAFHMfJ7Vb3U32S0DyC
ah9a8ltXSuNDDW/hR+yQxNLs6+586XK9NNQ+MftuO48bezgf0F/Zb4C/ppzlKeLIispnGgCofeNW
cMiFXH9uMfiVf3xFVeVVUkjVRMg7iwKEVoJJUWkXtBMYnZb24+Fd70XRryc+fHwgxkuiLmzjtt/t
QDPr/dy5gna1KqHAtcvkVwtFW8fdtgEBH0QYkwQa/ggS2NmIWYsyZvscXzFIxRpfszWVbn2L6UvB
A/ELKeneFLeKp2mzlWazKsgVAOAVtFQEVAXBFrU5ZbLeY2+Pcsb+Qqrteaz48zOlvdUEv8bJdu8t
vY7v36ZS8agH3Bfb8eakhhCDemYWhiStkxxUkoU1D85CQ2qfxdK+qgkD+YvkmIz9x0rAUDejm4iO
6aGeTpVy032+qRw+ifOQP29ooWbTip1PnFw/6Hk2OUgucxhS8GSEOd/x6kWK6wXHaYs6UG9uGlcv
lHbeExj7zl2lE0+rb9kwsWGnOrgs+o0LTIz4JzgxRPoDP1E+e5SjuQxl280zJJ211KbLGww5sPdg
ofc3aY43yXCSatyLXUROqRHRFrgqTLpmseSOw6BcuIs9s/ONILt0CBQreS71G5gZRrKGKgcK8qVH
GyVm+YbYoGFmW5jV4c/nWFvXPE1p4KwtD+/HJ1TuMYtttzYQBWbTGCOMcDMvHwIGy+wSFBwJKI4A
die5u8UKpRzFfdwpJi35hhc70DIuCgB3gPtLs6s3kbA6I2YGbWNlT5No0HwJEt0T7dxWZu0znrO4
En2MRaJX65ugLYaH/PdO2VghKtXoWUi1mE/4hZ8MSR/m4NprIf8g915hpOVuyE3BGXqVmPb6F0SI
02G/Qal/NIjGe+VX5mQhnKkrPfpVQVpSe8htttJgJq2N4dTvLJcjuxWsxu8iuh0xEGRosydhVY/U
1t2QjETihqv5ebNJZbSWQZGtLAQ0lYf1rKUvaoiJ2NXCnqO5A8yWsRn1uLRgQURgmKsS4y9CTh8p
NG8/eqOhoBGNojUtH2QD+uPuHfLIFjYVvTAyHs/nGJtkJd/BKM4Pa15hoe9Z8oINq+6VNfQWSP1y
SAS/ggBzvd3yUY7cX9jfp4eOWWUQgnNkAsEtKHHiLNoXsPJCmkt16m+GxfeGTOI7knVID7w6oD11
8d02DlGUzMg8SX/k3q7AD0i4q9KjjQq8Rsd5PdDtTGfIc1RiH4CS9Bw66sMKiL3jk6T3YgAJnmp+
UPHzhLwehCXQBwXmxPpFWo0boy+1wKjsgJnYAyRrJYdS/ySkba3ZSCCFhYj0hto0T9UxafVXguPJ
7Kzigkek6HGM9Ypwq3ww1ZofdZKcg6AzEz1nd8sXkUgeBlGNENb467XHVSny/xmcCbs67YB6uIYU
U9QInfnFVGigjkd9gYHkHMoC6/PxXPB2gfljw6UGd5JmMVE0XR9kXoyyIeT8/9ysMAlWebI9tSip
d/MRvqxfUFQn44uzakW5NM5vPo1sj90jXldi+4rZNzepq4rfbjNP7KWPwhG+LRU37HqadGAtQKa0
N8ANo5AnEsJFaPfbNRUdQcmU/dyfTRTDp240vT8mjTG8ez7jPDO6zIPfao+kdUTBS8BdErXQM+zY
tW36HmeAaiv/d9ZycJ34YYpAXdSy4Pk9j/i0Ff2fNh7Gz7lvgdmQBPfElM073RBEK/bLHNsbG9do
p/e79XHUMP6NEnh8qashFXXcAHBjTMWumVU5fy/x6y7nZ/u4skPu1Oh6rwSmwKf9IOWZX4+FuNpJ
CkMnY/txCOWz40UGpr9SAzIRf9/eHVL2MI5ZRtY9TCzPNxAL0awSqzY8NI2ufXkaCEh9DnfvoE8w
QBOCtOKCnbw5zUZYkNRgbGIvFtYFo3IwzzpcfdojGXO6v2T5MCahmzC2O3edo0A1Vrv1FdFmGzAq
gKv+aomWQDcDS7vPuHb2G7KPm4yh0RienkXXzp6TnabsWMMwUKF1YdovDNbGUyr4yfNIf/VaGO/F
Ml8y5I/SHmmhnkUlAQy4O+chPVrirJCsT+L6prE8OcywebCTFqNIBQmWuCargH5A3Z5iSoK/2Fof
D9AAFYY6cpEhuTqZts2zmQ/JCfKrwqIvQjUCVjRBFVKlpDU3lysLyNeapKgw1St0+Ffi4WUUWBWm
vOiA25lBL3XU3Oo38NZ6QD/2zLbIt1AD3yWUXfx1ulhK0jpbfH4b3qk8k32NAaaUVfktCDeCGLRW
OfUR4+sm+yk+FTYVjEE65j8nNxT47pFrCDwAFDjwqFYnb/wl5sJUEoX4LZRYzOakBKj3cknAMKz2
U9fCXvfaI9HlaCYwIg50ItJWdqFgwI5RNwGHhMbpcFjNxbX69oHp4w+h16qHNfRgGkn3/FX1j7BX
O4My37uf/UVdPpQjvFsg+ca9n7t0dk6LutSJdOboHyh4wToGLBJq+RZ9GtG5NPQwLNk6HInlpWBS
rarG+9HYwWNKEk4gByEOcQURmKx8iqe3+JtgDkZtQNy1e2aOMBUziqvv36ExvygkFrDzikUks7OW
3VFlTzOY4YiMV3AsKovLtfdRrC7wYzDh7gxLNuBPQ2rFxr65ari2qxnvNJdoEx2lMIhIUeDMWL4B
omTAUmLbjl8zyL/+TDW12BR9WIV8VYzKefTVfoiiPIu1+R4pwa4tIqh1uSXMPLQxx824NGSwkDSr
084uF32GbOFP0HdIRhdhQyxEUAK7CUDFJUB8f/JgxlU3gzvQoVsbJXXWpyY5296JiFL/EZYckme4
uCj7YL8GdOZJRcZAl0+HrUYwL0e79X2444tYKI5XBaLcl7FwYLNZiJ1te9fx1vNfaMBcrUPa60PR
rNYalaAqKw1BNE8yVCaBQY4TEqM2XwNuc2Q4nIB+y50Y+HYH+/UlXZyPqQqsLrUN9naZjgmZrZcD
WWffPFjx+wdrMrjuLZ30PnobqVNSmpZ/YCB1h+W78orLMKpHE7ZD4JvyjdIG0e55uFqvKx2wM3q+
opeCtIzlb0YUbRvhDF7nI9nIvKfTiQizwyF2r9McoRvrI4N/KlVO7N27rne1m9CozkqAD41r9zzw
DuGFY0hNUAV2BgyST3X/sQRFXQ9ytE7x++Gw0bk0AgfBaeA+2BU4DfjTrix8rTM6HOweHLhQQYoW
tAkp8Cy6brioMPChbyaXWpdsnMl3+rV5Sy1Xky+wS7tnkoeohSDWCnp3ljWXM37OIqDTL10NL5AU
Z4jOaoWe2dQ/7SKjhSpyA155ouSRMBOdSDzjLo64pUVlcqVmqgIS0Ti3f3JP/ioviDywimJDU7b1
h1ht1ouw8sBp2LT2RK9B/6L6/zd8ShH7rm1M4KncNNrWLxdWLHzF4evczrjcKMDdVqiNlO+JRwvY
gvfeRB0cTS8WMCPtUruySpDn42MJmk35WBcDr8stEB8whOizTGPCiq+umUB9YapFWy4Ln6Tn39wg
L/zwsaIq8/Nl8aDVrq+wBQcwhfBRZHFPT3zwZ/WLm2u/D6dtqTrTNziNq56xZxSooSvGkIHZhile
3YFG2ZIVY9l+rkDwEOSX5tLyXz6v3W53Q7cgI/EEvPBz2w8qHgAq9EM2ShDX2Lb5eCIQo+yNEDl8
T/q5En3cXOWixyF9/ijpmN0WNHv5OsSr48YnSK0I2qG8WLPyLl+teH+OpDVKPczYTxpMHq2i8N8i
W9gSISFKm7W5QbcuLVKZkdhILtDDGK4qLJKxJuMt2/eOxlv5/9jIR4CVG7P+t4+Y83/Akm+6m7bA
VgKwhAykXfWZ6g6nt07+xfx3J/rw3zFhg0fid6OAtDrvvqjYFoTK9Aks1FrI/T3NlX/8gND12Wi+
mD2uhHKnwinWZRgMy+KI8PAj+yXe6ucHZ9xXE4Lz9nMwwk7z6uRz/WCE4E5g4HYZNAK380AnTEpk
dO/y1mOhOB/nf2nD3A8/mGdJBbcj/od7BlAVjkZmmC4R0czGUXmQl2AJZj6Idr9w4FN+luDIo0Fa
dzS4zcFCQNyRl79QVYAUg4AlzI5Tz9ByHG4gvi0ntQEGjA9kiguzul8rGsaAngc52SVlQqBM6Vk5
+oclDGukY/sZ6r90HaOUXK9vPU8PP5cxoNlxhLC3lxdPrQnLvzJ3n8P8HIn/CcMbr19RCUV5bzBU
P3n5+g1cL6rMvX0yMmHKU0gHcaYyrQpgE4fgs9CfdBOx8+bnVHQBFAkC2RgL4w24pA4ZW+/fYrkG
g7BJiH7svTjRJIdYNWPWJish8DOuSAvdj4ndnEIO5kiRhP4I+TFiky3mci0iy1JRjquSo3/+ZyQI
wXNvtDQQ8bCBBu3sfT9wLKq99elvxO4XbMSMprcyJYpI9unozrSF0cBoCMDJsCYxRhxgHh55ebfB
m5JlAQ0RqOSEysYoFFpGNJAjqZX5lEpH4qS36VGEd8t/PGP81BvUhgXcD54ZgCgn+TUcNA3f97nl
G8EwwSPFSzWpM9802bPnv1S0hlBJNdxkKWWFcNzSZUCebO1WjSTlPeUYd8YypdYHMmsjfdOs9vEU
2QCMNmAwegp7+d7GwmtI3SR1xEemU3YCR+sgbvi1Qxk10C39po12OZfd59O9V3tme3YmYc/DXdRL
sn7cRAguivas7w/UNgzaarxdsuTgv4yFRmRARkDq4SSanSESbaszLbpUtYoos872jYntVSaxAlKG
kG4gj0rpYUAPntP68PSJy94riPdU8UW10vIRlAwd108keHtoBv122vSm+l1ilxQkrGx6o2jR7Jge
ouMeP0/GKJDGiLVPduf3U1FqtWy9N2B+Ct+9StuJ4Ny0+0EheDYEAECtKleeSHLCaCsA0rAuN2ve
O8pgPFfgzHK2pM9sJ4klh82o4buGHLrk575NsmrUBnePkBdEcaGEIynZYt2LAvbKEVBqWTJJV1VG
mBfkakU8mz7/pNKzbRjM+b59F307JM47Nobfl34alC1iB8n32NAfpJ7r9i4lcSwbgthm3zFchVNl
h4ZACgdfgWO9P+hiyWM190eezgqvStF6fxIRJRr7xZjFV4rpJG0uOVrPHGLDE2Z/zd+jk0Gv2YLm
Ug3BE/8lDma2+63RO3rWVkpRdBEK3LVqPm13xFxFzcCZaO2TW1op0x+1+rasLqy3qauASA4CrPZ3
o8h09fttu1k4fzDl/kjbOaxcCmFWA/UKhe3IvQHnMJsFF1xZW3Ynz6XFfEUVlIfNs+mz8X6uH4dv
roHBmoOmlQLYm4M0V/b+zMflruNj/lkRpOoypvcu4hwNGKjybGofdn0cda4eKnWFVd4/cTAD3aZK
FY68CiN+5zfT16Q9WLBK6rfqIurbJkRlep0s5P4kO6jYH0TWkF9eIqRrSFVP3Eq/D0s0WrRRI6Vy
EGOBOpDThSo3PY/k7djmsIl2VAOgg9bv5fsRGPFK20X0EyLffRB1jAG9ubAkQuQg+VPPYlRIKaHy
NO3JTiOPn7TSyAdgbJO/RmdJNip8ZVNs7CpPDycGs4kCr/+dq2/L+EzmiqWpPRsSHHK6D/d/hT/+
rEBbmq5N0zTo3kDQfFDf6RjU/gnblKJ9caut46N70BEOmQCIIPGpw3vCSv7wlb+SYoy97HYvB/Lt
2so6micu7R11Opu0fJrtYYiWvcRzQkDg/vdZBAeS3CKg0T8RCv8u7ME6CZrnMIfDc74v3ZEAZmvL
xp4dU/y976lx0uh5ljRkaDm3nqy8vYv3Wm1PPS1vrs41edjtfkDMt5s3QOMBFZh4plgOolbf7IKk
3osKnr+ww3T9OaiErbGxClX8+6xKmNr3WX4uTgFTxEZmGIYQggWIZ6qG9khMvkJR0ZPNOxcWpyAA
wYYwo0kXPMYSc0iu0PVxu1gAvH4QCQ0lmQRfGgcB3bgFSEZeCGpqC/S5tfVHN/y7Zs36bE/EAkhb
n0nPmExcsn8uzEY1T4RWCyfjlladPvI1fzSpHmMPjERw2xdnNntOYhAexhkTqwXktzdC62fDuEKP
+wy6a0OMX9IV7UKuKIazlNxenkSJZYG6Jg2dpCBNM9px6u91QoHDHiXg8ICmtCbrkerCEzuMSPce
aCE0H8fdXnfV0TxbY3yXGLoVJn521s4skp9WTwktBSQgxbeBbOVzNlxpgCvurPITa3BDpbFhmvZO
5fPOZMtWu1HWfBxo4zYSo5M0xZRM51/4ihKvox68LnoLvtwNKyOuhdQR0+FRZeJ63eFVCflVbYnm
8fxvK4/DInib+MyxCAjf7n+ZSajJ1oQ6BGO529+PjuRYrAwx2TE4og6kE/AaWWxfWJKR/oTiOceT
9xsNlzYgpXHpKgufGwrWQP30SlT5Njc0gAMJm1QwPJ6NHY8zMx42WLL+WgWaSK+CX1Mrfie3UGOw
lhE41A6a0p/reg0qXsfvfaRx4sdVOsC94gFKvdfFJrdVIRwxRG/nB0hidKtr8zuXl936ZmqdpHN3
QSXlJ90nIB7kJOo6HMoOezETNCSmewETWEuOR6kneKLPmaTfBn0YaypTjwxIpsjx4UoduNm+iMcA
KRTZ4BrKRxzJoe01FA3XEYm0HWfi2G/eFbED8dW9OBnSw5s++N8rCB8OEYQHMkaLjOSCYJ7bi4qi
s1fx3ZdioVnVw7P7FQlheg4sMlIBwuKMepmbaRvj9oGnmOt2UiZ5Y/rEW+Ec2BsX1+t6K/A3lNd8
PZBP/WdInxvua7OLn2GVLVbapxxDbENaXqnC/slXlAXmzCfW2bEPI9NhFpg+/rtfb7uwKFnNNM5b
p8+jJKC4o0LDVEaaKaRedJFKZ8VJZBu4kuSVcXyVzo5CVYVto00avTGn/zUcC1w+1iuxBhp4Pr4R
1Jtn/yzb2Sibdz2edeAxK1vagPKH2lw3t7sEKiGFG2a4hEmjdnLiMaWhRyQHIyCnudvxyefwFsDN
+vJipLVNxfBlKNoynt04LBd+P1x+cn4oJ0IyWpe5QNEbbvpoIoREYMgS9IulUShrLaF5KUdkGHgO
7TY3+wmeqP13le0JlvE0cIpFOZEuVMu5nXrvj+zIWwG84T/RlFfDn/U6vGEdWW9L9/imgskLdwFj
Ehu2UvA9CWLG6xQ26i9sztmpyeK+G2qynlTetlb+mSWD02UYWJbKU8L0RTxYDekJp4iD/EJriubN
61PWZ3qbqAfVqwwrGEQ0+P4B6Lq42W+CVDFyXnzZRFW2dKtR5NIqOUkKDocUjalODuZVIO0KvseY
gthZq1Zqc4sKU0Jb5qrB980dcxemOon2EaQUmuEf3q+lXwCNN4UgP7OS17uUTGmbduU9C/apT1KS
De0rY/XVHQioeg3ycvfp1296InrXQ5tMFJ0Wh3R1byWUCszeFNMqnwJyaozmQNQwjiXXgxkMN4Jy
mpOGpb5DrzUgun4fKWx0/HFBVsfd+EORffgpsuWr+GyjzUcncSpWJd72mhsco2TbYi/R9gfqfQid
vnzV4DYp9Xy37/7GeM2LP5tUm9LEAMaGbCszo1wtPeb27G5PiPklS1ki/D2GmqpxsXk+K/9ajYg+
A3kILG3MKtr6EWEWcwKbqEEjciXQHP1pEVRXbg0tMKh1WpE5SFhaj4Oko4oJp5gy4r3c/ewXZYvd
jLiN1MTnvd1WP7BUz0KcpGZ80Jx4N+h3abl5/U2TtUuucmoOfbJHq6PdX/a4kHPhg4jL18BkOFtk
VbvLSr0PTmr6zJ4XCWS+m++CFglV8G+crvFNpLLN5upgg7Hv+x/vdmW7z8R3BnY79lPeOxo08/Xy
UZDvcXqvqXiFt1eRnSsiyI4Bp0RO5PGoOXy+mUY/ZtFQvg2ZVUx3MXfJQ4Nl+K5vtbKjqzcwwgUw
NX4iyLjVAmYh2Qnide/cDtcSrFEu3lxDeVslGXxPmmDT3vTscLOl2yc4QdfHcN3pSsuBSc+nDucu
caL98AgY6XZfjxMuxbnIwwlJGUptiG1XVAyoYeE8OyiiiKaHQo1bXQBp0SJYk4unMU68ZY+Y+SgZ
9YwsRdHCbti3WskjCfK+SMarz3Pu7PeEUZjnOJW5AO+LrSgty2dGdEcorK4l7M+0DD68z0+BaBgK
zDPx67htkNo7XHVD0C46LFr30KS2IcRfax7onRwRTZIWZ8NxRe0RlhHl6YVqe7RgXdNrUfjnshjU
tQTUWqsu3exqtRGFgj/FgQfRR2OoH8IyeW+Vnb8sqmtxTdH3OkIdwPXxKwy4A0uVJ83LH37NrsXg
7scsss0s893bI6CjksnBKlJ6IWWXQZgsZGm1K8EZwmOHQll0+nEUiUuRgi8tRMZDpuDbHHnkp4pe
HJeMKFJq1USc5KwftCTavze/ZNO2X0rMZJ5fHalW3YUWwM3f39Ffc8GCo13LacYhhfC19NQXh9a6
6qHi+Ia0kOhuwmkasHLSto90HwwDNpHpTyvdtl9WoobVUCLM2FhUU4BhL6dQ4olrlb8ZaCb1s71t
G4SeJXRZyDfE1+/WtH4wai0pzcIe/vvAU9cdwSv2qILE+M6tayYO75swBMCQe4gToGzUYiC78yrM
yOeTZoh+4SDICO97SWAC6CT+wgZ5ObOWTxdkLUP/x8JqxdNUkj9j6MjlX/Lnhgkpbmg9dJYguHrr
UWAbUBCEFgIokLIwttNLa7ss5HVy8oDB0umONzBmb46J1DvmeNIV9lYsqAHt/MP/dOT1MzfrOC+y
t1UecyF36Ma3tk3vdwAk7SN+Bw/UEXobtFWzwyqek1ThH6sk5KK5RxWZuiYJKy71WrQTgxhUITUN
ivP657GmqC4oYkwosOQtBOyVhe4BpJdfVPRqi9xmb8Foths2PAJXhJYx+L4RPuFOi/W/DGPz5uYl
7U8treq0sgNqHvcymEmDvLjU/4fXyf7JFFctZfGIyRYNJ5qn+plkldMMRZiMxeEPBiGD4R9c5vf0
5ZnUqfUGYY21Lu07iN8LCpBVtPateq28/id/KnBYwFQAfs5Ng2U6L7NM4BLPCXf3y00fDMAQjXiT
lkeuaQ/EZ1YnyR/11bun2t2J+ASxgf51Sn3bFRizU7bQL7dliYZ656GQE70P3cC/mQFH0lHkXUl7
t0Vvq9b3wjlDgpg71weyxy83XCNsG5hSfqpMH89va0ZtfNn/talFzZSeoiXWHqR50k4jHs8oMNHN
s3z2CvZ2cB5KiSy5hhqUhibPQ36t2BljsAqHG+1WlMt6WpEsjaGf+VtBdLCONUygaMAqXwkARF+b
p6o2nvvu26nv3kG8ssLWinBDlsmhKKOs3X5uq8+mCnJ8ieA5I+d5CHZKjHVqv10v2lmAsuZI4gjO
54fUzrh1KI6j1Z+uOAo2zxfHBrvGa8rcCdEB6xOU6V03u0l0wb8v9xY4zYIid+P6W0oP9OA1QTT/
PmeZrFZOGXOlFEqleOKp+JA1LjcLhBLHz9YMdCLJXq2ZmJh/LFPiCUgL/EjV8vPmLaqUvMz/glZ6
npaRwz1LGz/dmDX3iP/A8D7ItpOl1zEymR1cMmabGIQOWeGOA98yMQ61osJbYjxapG1RWubl4aBQ
szET9qsr4d7ZzZ5COFqEuZWeSB50uYkHP+6jrQucpn3EpMQoohoakfKnr1rADwY72bqWalzYaL/r
PdSkcZX7Hq94UExzzSZ76WgTN56HojJRd52Vs4NarfT9LG/ZlOOppagfHdToQgVp4DraSeIchezP
kpgDyrzUt6jZNg7lrbKpmEHmUrsnsYtpLHwiG3O0vv6v8OtgifBaiwRIW4aCm7S3pbojbaLnvjAB
s62gb21wFC4ZG18rXHIytSxQGK4VKfbDHJu68YaAId5jORMBjVtWiw68YhUrlGTf11xguKP9N6fk
5y0b0no9r/27N9OMyhiB+Bh+3igNeK1kpno//Lm31sVrS+hFYuMngXT+ZurHTDmEPQggtTs46HQn
fsW1HVfg+zXZLaCnHifTuqDnBpOX+BHRmVKFyJ9QJjvYE3EHh5u/4/h5CtHKE8eOGsgzuFPpXY7S
PCdCG6OlcIFpOa8BN2eo6RyzMacP4/moIRsMPnXi1xsQLnem0/gnhttd5OY4Jf+5HnqQRq2UWyGD
tPth5UETMpZ+UGr8kFgtEGULRPOWlV+uNM1TO9xxLVRN9EFRc+BkJBx/Q64mWbwpDEo/DpkESdD9
l59fSe17mdb0ODtLO1AwNIU9uIApCE6Vrhlvm3V3mWOHDqJHn1Ze0dnYt+c3bogbt436R1Y5SByy
P8Q6JR+shAs+M11VDTgqFoqYNUpkT1/hH83ALWrfTNpDTHCaqhGeB9B6qCEnRGK0iGpF1eJKf++Q
lvkWH683p2YtHqJjrBCWn5RZPwWUPujOuga+94qpQnO3cwdeu43zgXxMrJAYrXw0L3M/nT5tfdhu
hcIuJFf1OG++KwrUMzAI8WzgE66N8Cb+NA87A6Kqu30DIdr50pppJ/r6yc70xRy4cwvUxe+75kjF
kl2V+u1JMkT8Ish3uSagZVdtfbFIR/JJlSNz1v3FXw/kjXgITjeujya4h6TpYrc8E7sbR2/PS0SN
AC0e9/q1G8GnHgE+TQWTVl2qCoaSANYsDGmNLn3WmQMvS6V131yOETaPIF5zBB65HKNlfZ88LniB
PV5OlcPLjwQqQ/81eM1UI5MFkHQQeiq4q40CIUdb9RuLnDdcQJ6NMBG8iSRrUzsrJfwz62W8oVaa
8xdB+CfUrZJlWaMo0xuTJ9VPxv891Ce1XAcKm7p23ByimAmTeC+SQF289e/LsO+/fd4Eu8Z7/KQ7
IAu0UcTTYlhH5ZimuCrC+/WbOENB/Qlou4vSGUN/s8bERUGH7X29LOsRYYeuSX69Bn+hek9N7g8m
/C7EMayUgaNW3CimiW7DCcublEVOOKxV7XJnJB7PD5t4Q09GosZyn9dG79DFDDlWqnq9RfJlEdwR
VZpvGsit+bvn57GPLrbuU4H2JlbUdDsb+8wXggGMlvbFcz7lZxdxRGMA7+0VRxh0E9GwkEo2fg3E
URAF+Sp2lMQbBioC4i401dbLKiswlGDc1rOlSB3krvRMzKaol/EkS6lM3aJBlpX+zZsN1Nl7P5VR
Hd0Z59Cql96HixtGJqNDNswW+tqK4txBPyOl1chm5Z0xFz5ZKljDIeQ9TtkgZyfUH25/Fct565zW
bFb4yz96Yyjg4Aona0XnZ7cw4CRISEiFhJuRDThUStAKxnzBeOqZpgqxKtS1xRwzWGAk5T2w+BOY
IjcQq0loHGrWrfoY2TH8w7+PxUu34CRVOlAYRX7fPIJ39+DQ7tBK4KamKSY51WYCrLl5LZ5ymXhb
HrdpZaQxOIVeMGZbstng8Rz5e0brTqRhOpNdWS8NYY348LAMsKAzjvLG2NYJVXbUbDdMIya7CubN
Vs0z3kTHENelkruD0aO8jwb2eALG811APZDEkrsuUD7+qT+4Sp4H8tY/7hnK+aHaHmczNMl7C1T8
h/KWAwLyfC+rhG8ASN9cH2EbHrGJHhU+QVCzMjInPRueHwE5F4ZzOkFOmhdwfTQFBP19apRqW6MS
hx2sThOVU5IUWRZiFmNNepcRzGDuDJhLnpGmJRrxmoudAalX7OacZhyO5XxvER8r/LHXlhEoYvpb
/X1Nu6SPVN0KVgfRp/KKtBjyxmejybiLBvPpV0RXp5VwUA68VLlIJRDhmrE0qU/p7ZtL/FCd+LV3
pocjlIR721ZgyiRdVOPqiHX6R26xf73g737UGc8iTdFga3PpCEgr9gPIqxLqveWXqUJWyR2cCkKz
+0iwAWBY2eJ6dvHpTG4DcjlXTcGLf98zJD0naNxhwnZdxSg7pLAO/eiPK0TjCr3JCkkEhFMXXt2j
a1HBW7YdB+NYtMoCkELjh+jUhYUyhNMa+xlXSzK2qz/K1UG8bma++h9AwSpuUsB+8h0RWEQ1woof
k1JBIpcDzwKfou15dG7EM5VE3U5bY1+Tf0d1Z9ox1KQtgTxaLIyh+sZkejksVzB+C4jVoH5H65kb
rKLYvxkvS+eghlDvpOGZdf4rJWp90b1WmCvwHCSv79EVm6zXv0IiMTEoeJGAjG6/PYKDok8AKQWX
cpaGtLhA1TFXv4L4hgCSHx4xQVjJiqC+KV+6KXQ43tHWmJ8WYL/1VP9uIxDSMi7zeqzNrOjxZXv0
nKJuioa6uSAF1UvEZ+DbKiJzxONsLiHPCPNOXB/WINkDwuR2dCG5yJ+VeBotkEFzXGcFdmj8EC15
sS6hQ6KBkmDlP0cFNqRXM1+0HONGoV6rtrnpTLjhdAhi8KbX4Jyr/k6Xoq03KKvwHQrDJ2Ugig3Z
8my55RWKrwR2ty0KQdMKf2LrRub6NNGDSSSKqo3S/LxydyLq1rwp1XpmeZapTlCvFebVoXaHTfhN
WTaK1PVtDHGI+iUGnnBsbtYbQQaFxAywZIOOo9dFEieq19dhDXDtTluP4rupshBfbtvFkZ5ICD/7
TwIv30+u7Oo93VYaEbCqOamALeV+5HcZqq4RcVg5Zd5nZvUmB6ncLPoEelCbqU29zf8VUckUQom9
wffvJXxi5xcpFbHDHldMAcwOgrJcOOBLKV5VrBWwVd2fB6UVpTYvzCqreBCFyq7ztPVOoPbqHwPG
9wW+zBqmrvslTeg+0MIzWnx/R1/ZWOJwg7kV8oFnM4cHjaQKQwBwoimyICRs0/oOONDGEVYbSvft
MjjlVOwKEIxbQh/hE6Pu9GKqlLkp2Gra6/pSeXYGgLaQKwcVtdUd76E77YOpRGsldq5d+PhFXosW
OJ5gxRqtNv8GTeS+Fpz0G/Vt4jQJb4nFB+ttkyso3ACyX0vy+6/UXU3XSA2toPSaj/jti7f8EUhP
RYhIFuvfNCf9Y/i700s2OXQ7tNhc8w+9udDwhXdngApiCbaSxpSIecS86SNjaXeTLWQ3u10LlIP4
TjASaFLBxgwWEk7/3tOyTxLpcdNdbQQtRrVX33Z2j9rA4N8JhfVnkS4eFE/Oah3aML6seSDhAywT
s9RZqgnevP8zmBddu8fBDQp18skjNfy0G4gC0//pKW6iRwdkix/ibTiSJ3gTQOxM38jTp1157AP/
I+gFxMcjTJIPbU3hvJIZwIPYLWBjN/KgmbOA9jd9i2GjkS+5HjPWy/J5pyIc74oQH7Ia2iqhVZLv
d5CPj7j8sufIgWFG/F8nRB7xE6wRdN+kD93wkals+3oQJ5smkT+ErZhSFksdvcVkC/WlxJRkPDRo
hy20jr7oPxiH23EUheMB6MC6pv3WXn9uk/7AE6TZ1Cm7kz00ZAGy9ThYLStc7EGYBPQZdD965mSJ
MgAt835pLt7FJf89/MChlmgBYETwtqeFQ2SzdExejqod1IqM9i21fjfpQQ3xiXwAAzsDByyHJDDu
3oTRqIdOsubwktvC3nlHoskSvhYz9r03dL4aRdlylIwV4lS5FvlQbGqLUWxuiHuKjmFar9AsEUkp
8CxXyBeTNPgLtiLNeFzXuHqDYkfKN7YuP6gJR1/Agb7DAUsiEIKrdZxUkAiz3AzkG5c//a6UwBqj
EmQUOj8VL4vFVpj2zy9SQ0ceLaSughiRsM1vxlEugw5m/KbNv/ZkZgeKhma/40gCUcQ0FHOh8XwI
6VNNMjQKZpQn7r4cdARKzqCYa52t7x7S7DUN9o/TWzFyTw6cwHcmpsyz9s4nhcoAxxOa8f51QWHy
8+PqHzziHoxoEhCvB3jiOKPi5CPOhc0cHowx17CsIsJkDgcwk+tGlHFHFPB8zBKygr6ztyjc9+mZ
roKcjr697ErhH4xcqNTbLP7tz5xKsuZ20zlD6WFhyynSEyIgW3SnRGMu8Jzo5qUVWjBnlyUc8hFZ
XyDyUIYiMuaZxbMzpyOUhog+2jPC0Vp28LXP1VbmgK7uydzi9Wr+6HL9KdnNkkjNrDbxKtAEMnVl
joSqEngifx1dglTyM6fg346BOH7T00dI22xQXUc0NHafUKODlblJ+1uuCJudqxXKYhdFIZkA9aMG
UMyEmcQANGhWsK1AQIWkASOf0pLWe69pw3LiOQIyli+N9/fM7E3A0DwUJrWL1nPKmY/1z8dGQT53
IFNlPmdPt2tiKAzwC/3O1VqBdffnVDiB3luLqWTU/sGflJ1aulsXyJlJ4UWB2R54ZTKSsGxuO3yl
6ysdrh3/pUe2Pkfp/W9bvGeaAvvwfzC/anUR8esD3rqUPcL/Z9VYPJwQLUsMjEJl9AcAJZDDDBUs
nJwLkj39qhQYwa+8zA9f6DY3PScHV+4M+T9ecrcSwsRRArGXD+m8McavTc2+JJCU/5znt8w/A5xf
5xC+73zwe31K/wMts73bLRJ14KRgCQ1hPPE2ZsJBw2+jbpTDlrJn9KFtoNWXN3kjKbaw0LGu0WHX
1H6/65XWXOE1Jg5PT/c6IAb4+eNHy7CXJ1pSnI0gUjey4sKH5c+DHn2pY/fuRZ8dStqHkUsJTFWb
XclUQRrTP9ui/3XGbNBTx+rWvEBjMR9rf55+u+3bHnYoJSyKHuCQZhQj99VYLZVEy8N+1+1KdhPk
t7KEDOO8RBGIPyLK+d0f3sb8LUZE4/CXwUjcfk1SE36tedLWIZbQxynwNC9CfxEHr1YRjrVZBm9Y
XPJQVVUYQYnoBgO1jduPQ0mmV4kd/qFXfZSg8VAulXFwAJr9aRfLH8BmNCsqVpRXZzo0gS/OLGSr
/hWqlqCXQ79HgsG/P5K0lU8uuH8UJUTNrVYmoqwePHXP6n25zZjOXrpuaHRGFmu7X33dmDa08oJP
xRbgk4p/vHdtOuJFGDtx7Jj+p7BDNGgKbWNKZYcLKbbFKVGyPcsPWrqbdeVx00//hzS2yH+s7u0o
yrugJpVFD+KzFaEkjYFEdmNJNcQ0cinSbcBddnwNAFQ4E+J8bj45pUdk8nza2XkujYqCeGlXOIoM
AK7p1RkHJmMm06eqF7nlB7DMlHaCWTO58BIME76O3Za217hJn7c/hKkfV1alYbvjpJra6JppRDsv
LR1MVclT0svD8E6lcn7YLqg1zl348zIBKXk7X6cZ+5T/7b4iMvTeoVTTMLvE+YrZE75YUSupvmNP
McZEhIfJsx2tq1gdDGs/kF32Pvbv1cLp4DGOw53HOJ08Z1oVeGpVWHvWqM9u3PS5YmmTHjSPLSP/
520aTaV7R4h8wwsoB+8RJa5dpr+kQmyCWezMLEiFrNF9U9Fq+b/3T/2VgVG5k9kySgCD9b3nk44g
5nWWkSKji8vcxVEeA8xW3VmzjXKWE5lYD1yVK7YLCx8zyx+LhzQNiMMHONq0o/zgSl4DzfaUgnkL
vOfB8iOw3wKHDsCg4AQgb5NS/4NjXOWViQ7gPgpjVuBmq9J9mbTphNGo2s3hRjoQ68hR3da4kLij
/aDO3/SU4Gh63Z4MUBq+7lIbferrhIrbpINhPNA+ws88wTADO88GtR+xwQ5r8TE+aiXFrm7oraD1
dldHA0e+m5LMn77BsSPEBdo3bknrl1CIVC9ogL/QFhyH1gcyQNA5XhyDDlyxwPYWX21jFd2iNd7c
A3odVA0HEC3AX2LENa5a0lXE9XMu4kesN4K9krjiIGv73CmDy2ILmu7CmxUFpaJGGReL+X1OzLCB
VOsL4UqSx/tuYmwhjvQsry4yBEx0vBZXbpUWeDtNMaE30dQ3184lphp6AnhlCpN0dYQQ8LUtxOGm
3ICu44qBpawVOI5BxQttLHglJXXMMVRHgkIIYzwU0YoPaq5mEBCegiJAqlSEauqmteWuN/6lC6hA
XylVBjwQZjyVNoEgQTMQUozkwohjc6yHDg3vJVciqm227EHl9K3vraRiHGgHjrzHtAVQPw3ZK2FC
ipR+KY17SiafxvJAuDAUZyJd+f6Z8BViQFrubKTWtHbI+db3mUtjhfBBFhlW8H7jPlZirvq144Gk
Bcg+DRF9UA4CMu5QmHg1nrMj0XcQNtkoK3Y4CD9KFgVrXCHIQEY/vGXIQ8zwKNfcC0BvR/8/Pd8r
miG/SgildOYHS9cIO9FBvWRLvzi2Ks/Q9dgP5lnY7xgH23l5jj2hyd2qCup2457Dq8w9tz38Gp+g
vNc7tgdBRKjaarMyHPdpqTr7U5WqPV1mu/N9zHnOG7WOGqxtghNzVLJVWXENt+3SgfKJbUy2nIUm
myvnED3oysy+sR9DObHk4auNSxKlzPReZXRo+JSvaxVSHDAQpF6PUr2HAuQiBHOMD0uF7LU9VYAr
jW0NQvEjerRojZL3TSHaGtJKa4AeYvpWfa0DQ1BvHJGfVs+t7nvnjrBPJDqq8a4CVTAYmBeZPVkA
3yXaLLGw7MHkNMVwpsL05n6DesuTofQDxQnQ72i0mp5LTQM84DnaR7r6uK80qIRbms/stCUSkA6w
l38m5o07nYKZQuxfgwWzsnF1lMoVUBHIgurw1GzSjO4cOGQB64f2VEwNuIgzwesa1/2BQrTlzK1C
e4E3vF49BIhr+g9nQP7gVCTKPkZoBy+SFg+NY5YTTlYRi4AGanqUcI8OPg+Nq+W3X9biFc0F9DD3
qJGDu5eFKnD3Nu2H4L5t+yvYRSIUWCcayakgdEcjYxavjYL6nF4NBfOqCE6HhVGszCE+R2Q2x+5D
VQS5Wi5gbqEp/mX6+Jdha2NuwgT0iKIsQirHbt8G82B0vP2CPRdCQEMihnnyRI8E3x1FRJDoDshy
fN0Me0QNmSY5jDgsTOQJWicV3sroq2g8yNOKNa1NJdjj/ZQUnQApDYwFAbW0SpNly+E8+m6PfPi8
B6yYm5Z3B7TX6OkHUrDDPWjE3rasXid8hOBUaCmvXk6sK9t8E0qzh5sh1LNorDpz+lreaT8sNHjL
oAL/SqcWpEOhCfpTAP+B6e/IXrfO6BKZjwAdVLQlAAiISvzlUB9Q4z9LrYdDwLuebV/4XdZOFCS4
5bFuEQ1NxJchR2OsD11KrbXl1sDhB8pYxpLy3/v/gPFk400QoKhlRFMzcmOaOkqX3P7Zjw3urfHG
sun3sien+/H9klEpM34rvi/b4gAhUcfiqxkn/VQZMNYBc1R2SG0SEZl8w9MlsqPVkc8wdk7qQloB
0qvifRSMHUpU3ZQKaUgBFx6PAcEKMYqvqd8GS2NytcYARhoXqzGpEytF08f5Il1aCoaAVwVUv4zG
xR0ByNiV6hOVu8YdGcZKO7UJ0ok4T701eHHh4PSPYKuCa+iaTVlCFT34nupd7L7ZR/TlgretaOLA
mLku9mRqdftKS//v1XNOyJduQAc3B7eQvmCrDHaangt4QHwjjhJeY//kphS0IAx8D51AnTbNbNg5
JZ77T/QE6xcRkILLMe2J8ug/I8Ul++tSBeuzzyndYlhSylGa3t/7OZVIkSvUxrNtKFecC6wD6+1D
i1e76nXiRcgdHJLLFAOdC49flz/uZd2kB6OBK0ueFFdkWJBx7eGC823+wfGNpiHj3Ic/uvsLNVrR
oHNksBtlnC2B7qYusSCC16U52cVKjOhkaXqBQcG8fG9+4silMc7UlHbWTR6LJYQyR7VvRWsc4zVT
LONLHuN+dsZ/mpXmKrWGW68TprQvSWcszyQuUK6MKw03O0Zj/BDBAlEriDBe80HrgXcZT49oQyzX
QrVK1QyHtaRh8vsYWDgPV/SIuki9D8TeT6OjAq+T1WaOkVDYlNUpnB1Q+avBHsFyrYZ4Ndb1HFWO
L9WM+/DHZDVLVjH6jhOG98esqJsOZ8Pllme8+PkyhKREC3Oar0gkrxpGwQH4CPbsdaUn6/i1BaLZ
J0hx0afcZKc67oI4u4jxUYptFoyyxzYK/niGhXjcUTqG1/rRo6I5rr1kvzFNZH95p1Y9xcWN0Op0
jF+LpT1sMECtUVtzcH2wp7l4WYldOOavcrO25jDpS5zYs9fae/vG/H/2GSygw2FZ9yjDeHbVs54l
x0sqXb4ciyQquhyqEXvgY1w1dWM0zbHK/TzBrWJVv0m4p/hGF1Vxy9+qtcg40NCmtwrngU/QndPO
f4dh+nJ1nBhQpeJyxs66lqkiolKT99pCgoZ+J3YLygxMtpZdRwAkwLw8Zz5zXi29sXCBZwlLggWP
Ycv/lOA9zutbMPX1RPJ4sCbw7iTX+jPNtUHuEfd+JmHUpR0hIUPSfW4XSEfLT6vECzeRc9OPvkQQ
Wo54oyXybHtmOokGjH9JeGO5vjyJEnnY4pMgoziApD4osfMf3+PXnOuszCC7XVHXvElOayDrFAHh
gnVCv66mO19f0esYJOX+/cbX5djIctLh3DvKKToY3TQndPoLCfpQq1+WGuOq2nQPn60RilGlpKeK
UxTCEa14P4amoz+Oi7X+dnNjKXrCWld66Ho+pxd+b85UeoeWIfrssRPFNc8qGgAOgiU2lu2cbttO
Qiy2cXfv+cCWQpfY1mUqokm7cX+nJh33HEhFB7MPQAb4r/ss976QWPE5poYKVlmjiH9RACQOacok
3V8Ue0cpMqDghxZcrb/5tyeHWRCip9eqsHaC/EtVacZC5/H0c8L23/Z+QEFydo5bxJTCPOvaWny2
ZR0SnCyjzuhXydA5L57EZ4S3kRNjPjs5H5esXoD34WcJmLn0sPpeoA9RESGPUmHF7SpyDc/Kuy1C
x2W0KesIOyUjxlfiIlGfBXeHIev2qLrkYnQz4L4jyfT1zNiMlHMjvvYPeC6m1ZdcHJQDShGTR/DC
jB31mvReluG2nycXW0aymIVYK1KfdeudxYL7qp0IV5aD78IpznwX+pNZxkWI7IpKJsKEdrJWtmqF
yl8W3c3ZP7cAucv1K/RPNWu+N1poHmYJYL5+0906TwGax3Gpy+23CxDs/NODeS2q5sUKynmjqGv/
4mnCokkUY6IYyHEvJaT6Ae+QfexL38qrXrEqF8ZWo1iUN57ij9I0ED7kpxRUXSmbCDliLYueSgi0
1Bo4N0yykZcpwFf/ZNmlYmFLPClANHff1xThEXzF2FkZaUCEVpAOdUlYEAj3lR2avjEPusR4hcEG
aNQyIyazsV8WQoBiSPt6CE5j7YK5q1B3gkz3D8XZtJ8T1mJ0RtrMpY/u+ua65p9m9za0CSRBRt23
KzFfz/l6t/CfW/u92zYgTnIXtgiheu4TtSCRKXbMEC9Tnn8dBLv5RBX/2EKrFZO8QSItI3d91F/q
Inl/I5/9VjJ4tyZtMqpZTrMdFFOh2vLK2hdfxcDEaHj+Y8YcrE9/KmaSw5coBww8goKqzfhO5qc6
FW0s1h58r++rzhFjS/mNE8jNnUYQ7gzx7EOi47E3aiPfca6pznIhfTFrqNulL+RYEWRmYkDZ9ks4
wWvIPAb2ISGHBRcmc8lx90ruBhM7OOn7TbNnsD1zkyAzgJDuuWGK3LibwfZ1OVO3P/h4/6DcQfjj
HagrI2OkIIkWtRg+Rfr1aApqiDblRWrd50urufHuV2J7HEVzweTwZfOUkWVeoudH9iHSOLskST5X
c6x/Dir5rKk77xLnKsye3uhdjcgjOPNPy9C3eeuofHJrCJo56XeDgvp8Mx47DZDvwh86e+SNl2AG
1Eq8bWuEGdeAGV/xHUUb9BvpeeQCvHCJ08F2leaLEym1APblk3KZX3N1OEr86zdRrKe9KOGWOG3E
uwAzJAb7TbgmV2oddbqdxGM21bTRL0OKrtm2Q/hUH/O3b9ZE9ka4961wXxNFrkGeNsCcn+IBEaXn
LMQNJdDsPtIpQG+W7lKPqdVjVRvLx/PoO6SRun6moV3Tln2+X2qhgSinzCH7BKhRBD4MD05SYI0c
SpePhlxoMHxj5cJEyLKVwSx0PuWi+zoXI/u8RKvYdCVaBp8rOuBRk2NUNfWKUFwbzDIEKXbm8T3u
12uT4QAiJyZY9LC6lCJFlOZYYSeE4Y6EnaUEwxfVnFCxyewb81g98gMpPZNb+HPSBo/StIZA98pb
2DCdQ95hWeVUvMFrfGYlLicq+zJ25xIwDU3wBol4l30pyjXKENuxz32MRrU0i/rgIQ8A1lNTZF3u
mX5dx1G5lRHYK804nR7VszwdisUuk9gmXDfnq2eS6DxouHjs6tG6aEz1mZ+pzZYfWltBwN+goVWO
BtuOV7RuBQPQEvxDGLkhk2dLwhMjFE1+By6IwPtRXfEaR7VGND2HvWYkBB5/G/9YvnPWOLh4c852
K+2zvteS9xvA8GOK5lPap/UdsFVx5Kc82AaxAMPPRGhsSZrt3XRJt9FxT0yAhqEBqk7ZRaKRCAXZ
5m5C6rI8hFPQKWnTrHF32ki665IS1jX6ACMhGziMg4zvvYLyye+2X4HEyI/dzySuXiIWGcenYxtl
/dNLoXY4RSF4ObbR87KXfIDHuZEtfEOG/JnPaqre0JF5LS1z2Th+3gQZ0Tpzsbsr4baDwBQDobDO
FkvMCWt9ISgUocfAj5aoW9okoUs1sBfXQMdR2pOOxgc51RLm3E/iLyeRHLFZ4r43HvEh5X77P8Hc
IMwJRSXeBukbduWoTcLNuVaHScDzH7nFP/dVzLUFcYPcsZwwH57YBXdgJ6jB0vwHuuqxW5Ynp/bP
dRgmXjxAuR+LpDanZI7mRr9qjLL2n1SYPcu48wQdgnLBk21buWitVMeTvra3lB1Li3+g4S4EM20U
S9k4iRUm4Hp400YS68+OrXwhRxbD5axNNY3PBRJ3Ib60aDeTYKAER+9ZtiMy4pC+tXQ5xA6DO43Y
y3WfxgmW3NEs5vxH4UHo8oltxlJfyXA4YjMbpoNQ5vAkcQR8MQEm4TLyK4YzPj4WFmPrCkrTw7b6
Xg0ayOkje1a2t6v/4hZxf/J/fOFXqcifBSM2C8INhrrLwHKoxPTeb8GVYKwu4Rdbvt8cJ/Biw/DL
C6YExoZyaIsA4qBjUQu+Z8p0EU5puqjqfqX8ueNWm8UV4jxugFsMgrpW3QLMMG4gNvaBl+lle9RZ
8WXke/Or/QEHy38jkW2YS0wJKYOKTj/62MXOLnVWsJ0b3SLtDxb8uOjqZrppOMvEMP/S8KnMITiH
QkSi3HQaHfT6m1ITJDap38he3Hgv6s+egbeHaxG0SbWcTFDYEqY7CA723AZJRMZEAencjxC1xoe9
8sIYm8Hp0r8joert4tTsBQUMuasx52hGG9NgYp6GD4vI12aIiBqeTrPdbQQEMekQ1TDBYwEEY118
R/1x6ffG9bG63MfumheIcM3XGH+e6xnBXq80XAqQ5gbmKQmcy/K/dbHsMNOjxa9Sp41Enp0N+2NT
2ePQMpCZ/PPhbPKije8KX/wWkr6+h6M9ckhD0eSZ1cb0KWpgeu2aS3plfTzk+ZJOULNt5gdxfESz
8030GOFQkvljwcDzvo+cuchbsy2xl82V1w4KW9NoSTFLjU+OwqEwqJTBucHLniQuXdCIVdhW47TS
6BgTx4ZiI0+9yNNSrbuDr7ZfRQmXDhoMw6RyqEgpCGVrRK3f/0pVvnia6sLDJ2z0j/uf52l1Npm3
fykfjApq/YTo50QZTMkU9oHQrAIO9yo5UuA3ilhgWbcJoXaXYZprlJInsBbVb8ujeCrN2GWSChmn
naU969afG3+cEeExbiAEnI+savIwV46T2nb6jIZaBAaqcHwhw9klxuyq5gUzrxaeWdIeNiELoROZ
D6Ywv0+Hh2mQpEHtqJCGUPDzUpDWgPtpmXgqSz55p3VNoCnZaOiEbcMT/PAPi+FadBA61QKI2Spa
GLmTXPTxRrOB9v37tWJjsOXXSlP3QzO0p10QqxmtwZjRgpC9fU1kzg0oQRrZ/WqkSGdgDSkD0PKx
tRqI5TekonWN43f3O9X/CxPICeAOUldPk62nzMyORs3aSZMgtFF63G2CBqDBnwqBUnwEbkYXW9PU
2mvW+UqoKs1P8j7XQ7+eK/6YsviTU8U7GOgxerJhFJ0bSBlitQb27bbhqO/8Hl7Afdz8fyuTeBbU
w+V91oEPFDzsMJ/J9EcHMqIxRlJbLKKk0E1rX46HLByR0WohBzBGtYkzCrqMrnb62EUT4WMXVrv5
qiQaA/7BFjYpvycFAqRG/vhDDeyJXVsp99uRjyPD2NVZkE0DiSSSBks6FdT0uLhlueHCc+I8bja0
QHoSt2Bu6r9jhq0v/9o0imB1Z13UTNsKM+D9UTcNxFpCrtdrKcuNfJ7QtjTnCSo5yEgUr1EK9mC5
ltx9PgHgGywe75aQ9QD3y9kI+TbfHl5CSFS4DagM78gg1/6LuxY2ZR74TeMYCeW9IxVV/9GE/O+V
fLWskvhCqvFhkaqbKUX8tvjPpmIR/XSaAufaW4UPbmP6Fmin4DCHYclqYMugWSC0PfCCt3mh4PMe
V7j8daZUN0qiOz5p1ZpHWGkqQtaHuGjgOz1Hp8CaO4A4RlL8LeYHoveIbIyshHHXCx+DBS5kvAa4
vnq3WQYQPt/1AwUYbJndZZlMUJNf+/14Jv0iK38qv2EANTrLlfupkAxDQ99kOHOBaLYa0i69NSB8
ZfdfGJDJ1HRk4wHMnqmW8+rAqcOqQspImywtOusJB6VoE4rvtBuJipbSx/TTV1Sbm0FoaLy+aC85
uIgjP1WFAx3r7ljgaDXVTLoygq380o9+0ZUxKChKEWerbD0TLFUWmNJVb3z9rvA1wjGjNg+VvzUo
Tp2Ph/B8l3J7ycywQjG8lmM9XLsVkEmpzZvfinWYFUYNraWFsJ4CJ4oclmUyPWJ9rNuuFlV3OiPg
k8iACTDmyl+5rC9q6NrIZetbpUx85y4bz/K3q4VmvqrhKdJSzznWC6qhV0Gh1Sto44gYIu4JDU10
h/AAWAcdHhuRQsdNgfW5CPM87K/EmlHcP56X/eYoCZLUD7GFwCpWK2EPFWN+yeDxW5ncYMQSWVKG
/hKHYcre02Ky5k+AoJQmv57CL7Pn4Ag97hXGbn8wGTdNudnncUrz7C6sshiEOVsCYJKJzgZs/q7j
af0NMgoYMiAoq5QCRvAj5yumwjgJk0Jl0VWlXoS7pGjUZni6RIZUmadVysRKkYsud80WsxzWQq4a
7i98f1jkOpqW04t3P8RI/BxbCSR35tr8BOYbk4mptDLlCAlmss1eykkWSuLMoG/m1ZPjBqxDAZ/T
aBbOCUfC+wrchBINUIGzIBRFREsTXT3oGMf3fte4seU+oVB2KCaVaADTj63S3RvsVScjO+vDpApM
A35Z7DFj6ScCu1w0Kj3MszqaG0/ZdNIkMHA0U2aj/KGubvzTd2eR69A0bg6vBiRTPHgzciMPgaoJ
b9XHKYtEUdz5JyDdG3Zu79g4itG6xBbi1+W2LffXQjcX0ynENKZj3q9lrqCtHq1H0ERs5ONaAP25
LzUFC+9cbLKUf2/wlTmyRSZtMcJeFw81nBpzizOmFpn2e3ji6HyBtXbb/UWd6VUYo2O+Qnm9R9zL
F5wWFQQbkPL4wE30InDDRXIX7EIBfMT1SugY5GdkYJ3ZPQtlXlZfwUpzPsyyqFmcw9HBczzI3k+w
i2VBUgBNX8zzANSS5Xw8gR/2x5ICsTzrJHAHziC/kiiNGmLlTwPfyudA/j/nWFJN8J+FozgZ31ky
Yf8fyovl1niRmIBMFTs1fqopykN9Y86bIx97aiLwiE3uI+KCNfmtxExsfzFmskH1WkhLF0yBnUKi
jM2oujtltQ26S/jmL2wq/uOgIZTixuYa0voVXNCzu76ElA1hWsIvJeQuacM5kIYXWotVCzQOyAHj
arzMbO5gr66yfYCFUI00Mr2s8kWV54EnSHRjOUDmQM6NfNRxkQ4wA+72VlFuS6mVmTiH26m0pHer
zqfDb9XLJg379bxTmUxj2tcrliU80ezv70jwFx3xixEGXEltX0c3R074xtLZfQH4mpCB8jMQn2LT
0UmLNmFXkkWk8jyepNaVzucFguutdQ3RwPubNYytafQd+8UZdFdCg/SQbsgsUzx8Qbsm6KtdFtdQ
T4BSnkwe16ekcJwk21qnxBJcrBZVtdWGMSqEXtKpI6SGX1Rj/6hru0BXt+mVUWcuLTM5g7igGjcx
JF2dd1JC310OWBdWjHdfpLWyyAkGTDA+D+LgTvw21HvrCblFuLq2+KBYjm4+BBKGb4aNJ45rQkHX
GvCGm/OXp+H1rqZJdsfnpiaePscQdyot295Pouv0lYwi6ng7SrzvcKF564l9FDd30kSW+BZJkMsA
YEI/Lkss8YNMAHdyMKJ04wUJ1XzW6GkJEeZWX7ttymjJr2R0YFwTnwiJv7P8PS4snvockq9Q+VCh
rDfDa+2J5DRUylp0eUZFEXio54MXEJ1k+1ndn4JR3h2FQpaDfb/jY91uIPppOOXR4d68tzXd/7fo
uZn/gGtaSkixptIxTIzu8QROswkBLCiI/57QIr6EaJdyPs6t4lobq/n+V5fSlt+4lIGDBjxDd5Gh
tLNLMSoQJUAkoQc2Pxhqf9QntVD5i0FrEKh2pcVnNoWgDCVThYeJvns3DW9w9UDEXnDqFQD8ZVdD
Klkf9mut7maDSfm5+0zLN9diLAVDxIpQ1cBYaFWfjZCThXqPjp4W2KF6EzEMnma6obpuxqgXhXG2
pOfYTkgCxxt3FxQL+s16WzgSILPRuMFXK9puixpa+QmkY48t8O3mecQADgj0Cw8Th2hGz+WRsC+R
SW2uj+mQybX2YFWAOVPe9io410XjeWm1ld3H6EWle5O8Krceh5VDWWONRasNb16J10qdt/Pytw9W
72FAJyII5JKLBvPc8ZRuuVc/Y3maFjtw6hQlVV3vkXH7SNis1vn6ngQL2fP3jFlDXhZXM3KEQUG+
vkqwsPddgThIzJLep2NeLDfVRP5p1xZHbF/PEvH3YAx2Ata5jz7AQFtuC58x0oUg2ibx4VxG0SbE
7K621A+kSa3wiizeqjlpW6DTWjfqyql3fVFThx/2CFHrDKLd9S5X2huWnENqykP+4UMt9IFfomCQ
jCEtqiiHO04aLjQKqj4kMCLmXDLzpEypYonKeNnKuRXRKi9gmjXkvcq98a8pgbxBoqIcuxgR4M4I
/CzfTTAW5QgOcW4/wMdgzJnro97DQ2aWsqHGQMFqILE2HInUcgH3HBPlwXednpUEDIjC1iMbCqqo
mQToVYbgDBOdlNbJyhZeIf7afRYKX7wfQPz65ecP/gzQs7nmlWx/QkM0Tbs9nQAsLRCz16HhiV6J
zVTa33qcOxO8vSq0OrF5QvTMX8W8Ek7y9sq+O7zUzzWABMZsgXYp4CVs1rqhIdteVoyjtHVIEFcP
aIKXOq2/qPL0mxVvCBqr6Y+Zgx32QO1gdQueYQec0sSWzbJ3cR/2o/Dgug5L4TJVv+Ujbrarnom8
NhOPnXOnjjbp5EvzruqQ7K8XWVGjV1XYncw8DtY+5FC3spgS5X+V73QTCk1QAQqVLrtBskXJhX0T
zLD41wTybJdSPBpFgmTQAZPvOcaEGzVAhARBzi+LKWKJmk0V4saXOzNe049LmAcberS/j7KQkyal
xOBy4/L3EVP8wu43buatxsPrIA1d7uM8p/r8tS46qDejcDNiqjK5HRBkCsY0gaxtcxraFLhVKifT
TYNbVDwNgONLIgNf220fjoOx17KyhY6yEhlvocO1k+DhKX3M6T9xrA7JgXmgnHq2chunooKpLJC3
V53OX+LQmPO/W7JNkTnANtLzz5cpdJVTqlynOV//iWabkyJ9R9QcjhvM3g3gV/B04a7qc1zlc4FM
L8xX9NOXn6h8/GldDLMZ94wbUG/dIP3kyxaX+jS09iVt4WHVXEM7uABgcep1CL5qS80qF3avgWjx
kVEE7Xe+R2+dQSyFA+Q4Sm9CPV80rvcjRmmLQQ6KhKBLJNB3IexqWgwqpiX4qwu0mo//GJLK//2h
WGv6U53q4Xj8NGo8RMOpT5CfudDyZ+bP22SiewoBYyfc79e+b+ZmiYWkyBbCwAfef2jHs6jCnD1G
QvEcqjlTIBR2/wWy70hq0n0YhFFVkV5C6NOh3iz+416GtT1RQ9bOQVpKi+8WjoM0adGinxQkW5xE
AnT6FsaScb2uIEDyiyEUroQSY3/FNdMJDaLcdQi9/BAIhKffnqFlpzrgJRShRWQ3WNQDOIJV0gCN
OIg6q26pngrMJ93C7t36ms5MHzTXCyBCgLfmnUqkprqMOICPKCmyBl1cXk2vYBhWmJZDpZAOOm4s
9jCWqj4zPumxgFdoEP33PJoL1o9Z/brTkuvfXC8T4VbsKiOG6t0M18kORlNEGUt6TBbHVGRkAkrE
UBVMBNfY7UkxuqJkpnbDWNu+vApiDbVIuS2fihun5/W4Ppl3batbnwFUndgJf88ODd6uFDrFwV7Y
0S2HUj6IXDZihshuy0r23qG85q1l8nhbirVl4G8I91/WBb266AbC/Hg8KXwX7AxNu8pHlLeR801s
aEP2WNdB70yUQf9t6HhAusp46rzZq23JMnzJZguedgrlS8eoB6zCU/+ref/moOihvnLVUDgCkge9
Ks/eGOCtIKv2gFpMVQL4q7hTpj+zGlGXntfnP9EGFs/j/gnLhqi3NaOassGVmqwNwdcGOcucIbEG
rEOKrQvbUuK/8Wx5Mf0h5J/fhPoB/2m87t1kOuZZrCUEtPOMLtmUB3VKZpsCG+rEQWRABn2Eh9HJ
Uy9QCe9w6q+zN0lSNsxoVg3TCQJgnTv5dCuQZ/y8z7rmcHbiw3F4pm1yjb7U65KcgHHE0z8nJGAZ
KGqV5V3VA8z+G/j8kBSobGfVBv8lKwYaJXcRpSSMNu+DVmAdC/vXm+J77kM8zPZYGW/WOe+PhZJO
YwkpB9KqI0UB3SbsQ7V5zZvEr+BlNzvVEj9Aywgnalv9hmkjtmdLbttuaLPpHGKSBUgsOfBPDQy4
hkvH9wvzf+rTJspEU9htQwoMj8us9owl6ISm/Ip//5qAWexAPaac0mZUCNOhUdAvAM2/CKtCckl4
x8g8U/r2gA7RS4HSUKOahUry1OoshHEtQc/uZfEvjHoNbuZXhQvLj9fQ+CWmgteuC6DOZ7G0R3hQ
7gbI5yPc1lG1wR3aT38OD9ruFCoYTCc4zWYIirQjXKR1dX2ophn9sELGdlf/Xras0dxadHPViqtH
xG6VDCO/3PhEQmLFba207UQvDvh1GIwgatW44/+CsHZZt5m72DxzaG/U0KZUtSyvYtjgewmAeaII
PtlrUH8oju0OSS1bZlyeGzEzHNuAVpus8TApkLcoUGTZFeIxp89RiGSaSorMKREatdiSQJ7EWKHg
rgxKTeW14pa15d5DRlZh0V2f3Z2kQnUg+vMTMOObRMIiAbClA3fMKd7xLUXUgkw4cv6+nRWp6D7v
K/CbtTQac3Ff0RmG9DkkiM+yruBvJb2cBBR49ZpfXmYULpe2G5djsV89Z1qo+WX+eS7WsxlWzPIs
qhQEzUY4r1zW1g/7FRl8fduq+U9gJmOmA1bQ77C43JUFgH5eDhn2pIkIsYOzrr5mzrZZyIzvzmLB
dY3IKlJyc4nX/GfYtbkKoKcf5jO+2cgbTIyQIXCa0NXj4LH7mutW3M7xR8jl+cwdO68PtUciGrJK
NF1swU8MdaA9N+kJxoVynvDpbb52IhukgvSAoRCITitcmSkcrjCPb957YJz6abbunUaAeKAq9sR+
pnfPOerUDzGIoT5y3t+ouJgiXPiDDBFqgjC4izHgmz/5xzlK7FHk1/X/Tgt5AfNauIv6l0rnPC0M
6zSV+UDr6vYeMVEWEVslu1kokA6z5oISTPnTSpTUBlRty7h9Vy8k2isZ4x8Kh2Tl7MqK4sziGvg4
qFeG/tuMbabF+WygIvY6EM6o8wzy/+SFRfCv+o6WcKFPFGpf1d+Bspj+qpLkm7E5lvOuXsx0eLDJ
dWA0TmpbyRrlVi93M5nkqU76zfdzk33hWgBD4YNCQ+Gq6l8rsP1bpmCBEtJ1pLXvUBz5ISaMLGJT
Wn6MsX+MGhq1Pv28t2HmbefYBk0RfbTF2Vg9gPrzh7NRqeF517xbphWd8efgE+Dtl8oVOL06lyja
QAaIQy4fNwr+MWlup1RBQICxUU2psOXyy/C38yZlwGY+gxVRTZG7rkIyM7ksRd6aQ8h+RfYJDJ9L
jNanx5rI4vMLRW2lPBew/xUq1/Qf+6C1YfsyHousXVZ3i7GrkydSJK1JRqYL4tsLwLnrcBz9EULE
f1e/NQyy+l89AOybCIwkwvMAEtE2wNj0y8qIoAVMuHwmnBCg+YP3O4Po52tdkGLexNmLV8ojZ2Oh
wyCNuJP7QXgjtLaedqXumshZbJcxZys3//86iavS+Iab2DOd9BzCvM3/o5McmN2haS11BAu80JZT
OdE8W24zy/1aXppJ4bf+4tCDd/r2bRM0Yy9plXZqDC8ECi1d06lYF057YyAOrvLu2FKL+FG33eJM
RaSynz0o9HrTfhDWNw4w6ipmde7gqljoBDIS4+z3GvuRQe7M+B1pS6ySyGDt7B06znOw3gjE9hKP
N1QSQuxbfMCj7BrWAD4Hs2jHVr76lN+latU1I2KWjaq5b818QEzQjVkh3K2LvReih4TM8Etkxlzr
IAqFOuV/ImNlvZV8hiweQiYteFj2V/NXnxV0I2AZI2wvC+NzGiSH+rWeo3SKod3PFsS5FapLjvaI
R8pCGCdnAIRbLp8Ft40G2FtPCa3HdbmtLOqvVi0/6g6ROiuovX2gDst6UCUeggvvsQg1hpcozey6
XBHGWTwtG3GSzAH4wHw/ISjE12GyxKHZqRMrIv4MG5TcEIQw3o2rtu/iJKjzBsonJ3JMN2Wk7ueP
QFk6K4FoDFjhdOhSOq7Y94D2HrXPLOa2Ae5oh/Skt4x95OAobHb/qW/RF3kMM88ZmADjyyBVSv3V
vn0TexNPEgb8cD5LL9aBalXL434KS5PXTDZ4TtWvh8EdU7u8PFl4WuvtL4RI0Mau/Xeezhd8JKwr
oZJ7+UszSSZxiQk6DUd73e7OLCR3y27hgPhUeuLFy12xKfBZmqm8qyUTyDwwGJPrJ/kFvAm8tvci
AfBv/Gxp6afkjeznRWOWbtTRAoBID2PJVwMCg44L6hXOTsyrHikm172riQ70SECCp1uPfUIA1IAv
AiZoLmJbsy/knhzeQfpaoAEi8+hBwpzbU4hBdsr7D1cm+26+FSqtWKej0e6QyU7psDEARwww3Y1n
qmeLAF+C2ZCW7DpO13hR9LdUB/iMwWDvKCbPyPaSf6U2tIgxVVOfe7Ax0Vbm0F687WomSNMKmmcL
YiVmuUgQs3Cxt+9I82i2z8z1nYXeHApatKWV8MA0+tONIeStxKmVWtTi14zDMC37O6lhM7F6EMK8
UCy196Eh1XaJmewhVQZjbaiNthGEoTr2C6wE/z77VcNxpjHAZH0sEgZVv8Y7epweYuLZgDbb32Ry
uXVNb4RT63ATylJUnRxafBwdEcsB8MbeC0wanPphE5SLtZ57ueDysa/2z+P1QMq6H8k6TQWuJ1Eu
TzslpXdfhSDMqyS/DJpvnJ1fICm0amE/kiPygBTCEmx12Fw1u8Cy9b+rvkqUWUpakh8x0Ceg/owJ
8Si2pRYx+u0hFwpUNdxFMYpM/Hm9bV5ysUsVC41jpIc22tX2xsQL1S/IWcY+xGdqOf386bEHHvIX
HR4cZXpyPqCOTUWRFVsQeZ6iHnLiC35KtIgW9oTKu2ZAAyuK9gMF9OrmtWYxugMpPc/CtQUwpq/I
yJiYBwrS77+CXFSQT8tAa2gBNSnPT0Si4a31UrwnTL3nE1hP01QZby2Zy7trBnhBrt8GzStkpjJW
xmQTAoi5HGPU+I2U5mZhtfp9gWcVHVmdO+ZirWIUjAMu0daEfF8ZF15VVbhdD3/cO1O9OnL0iFD+
guwo5arkMzF5U1Fb9CBNQwjERNlzEBJ8fsNMMozBzK9cXtu0xXfJ/3Iy8NU2zKSL2rLnhR05GA+t
w+jrFqt97YLioWdjlg7MFGyfYYJfzMdleGF851leXkeSW0tMzcVwKJQ5EMSCNKnfLHh4fLBx2Ilw
/b1hrSDsv0n7oCz38Uhl9JimY30M7CGYzabS5tyt1fiGsvu80L+7Ioq6e9XHvb6u180e7DlECsqW
XJBIj/Iy3x0mGXgFAveVaF9Ui5QUNwNtNNCEU37fvhi/0DaEXdhtkKKVTbRpmarHb9ooWl7E/fME
ZHg04t8sAdY0Sd/NzsKzBSTBao1cm+GnsnzlzvCywUkxWEHi9AmY2hI9cmDnpwoz1WnTLfQoOqBK
PZmpoM+AybaCixU2leiL3ZNgXiPT+ggKymXzTMyo7tQbjbfDuB5a7RU8lMWFmsBWsLZThgIXlulZ
3Z0mPiU6Xl3K2pvGTpPnpTylhQhHVPAv96hJ7PUNKlT24vZLXtKGw6KtJNhgSExG9+R8J5CjFnNW
RDH7FprJ3CZSpUTtGhowVNIzIEz4/7ZrlM07YFeIxLjz7swV6wzgzoaVXMWNd+sSUOLJ2OeKV3n7
bswtqC6VW4NDXSUm5Zjc3NCO8v21KjQ+zTOTrBCVGlqm9BZsTay+f7I2Z18P0CTzZPKyUCrvotsL
aPidt3q04bpRKsSaIgaKgjt0qKXo/h2aqAYKP0giIoCNS/GGeeJDb93xhn/i9G4ZIRDT4Nj5aI8w
JmtsExJkzaKmgCnW0W/jhMQx/avR6wnifFjlj1JUNjQKYIax6ZnouLHqGp2nlVWihu8Z/hmjcpCw
2g2EPNvw27sRGIDWbmyD3c7mqhRbatawJUHE50c2XVGNK0ta8eqB7EMkxkq3OnFnVGyE8KKEfqbh
CaIZ92GjcenZTs/OmqOH9w8oH+rtbe6r5VuzV8OmEM59ePIt+8/j6I4a5ecyrnHsomzEZMpvH3kX
sdYAZv0RjjmiO+zKo27TIBw5IwsXXbeZVGw6jLOj0HN5kpGhQz0e1NZ24BVyHubXu6sc43/0zlYw
Qws9bTTS1dM0oA4hnLkYnsRLoCPNkIRCxI60sY7OfB6keYuk4mdBISF/3exF2eUuRhgRyY+NSu4G
EtW3xQ09yjyZiOSfpx3V9UdM1FEQnb2RYiQ4wsD2+tr5PrJq9MimT5t4LZnqDxb6YFlxRmJEqqG+
a7zoFwuDoxOU8VgnaT3cMhAIQ93ba8E7PHIRKT8eDKkbv7ICHTIiPaN49ODVKC1PU9cBqErgo5L8
/2tYhVQKR4kymcNLy25vMRGyow0gR5PTwJ3fHMfYd5TLNWhGCJ7340/jd6Afi/1rwrB07v7t7m/k
pgF3OhpmF85cJjIBaNnzVQraHCsHRD0mQWU/W+x0LtXMW+Ki3ogl0aOcxQgfMgjofy1YSPIal4hn
gKmNgaATCHwDfgF2NAZomxm6Lfis/0EW2MF+kxpD7Co8BIdWr3Dgzlw3tQ2E7OwNQ8N3xuH4wave
P/IOjmJ9QDzlwxYpPD35tN+QEzN+pYhzH2nkCQAAmRBP0CDRnw/DTI/XPFAacFhyIsR6A44NA7VO
szBex0937iu7zGP8ZFdkS/8GZfnmaPTQJvH2DRpbXBeZQvxosXir0dN8VrGxXYCND8HAP/mfh2Ep
L6qHTCALdCzHRL+1YQN5qkwHVqf1EniXzBAK7AdX3QzvBQA6BeCUDBAmo5qiQYzvOqkCe/+jWUO+
k5DTuetdrfoesqBIi6wa9GGuAF7Z665vq4uikjybcrK/yO/ZUNJLPzrf3tTgUIpiBHzLZTYox3lo
MWiHpqpKKAEogwxBJsZoiFK/+/sskzCI1pshCV5bW8HuUYcL93QuMLZTK3e2XuqA/7PsqdwDyjGc
SV/w7v/K8f9thYsfLZn3SE1+lAegbSEltIStP+i5jFpllmK8kt7vCWgALqoRorYCJcFBG/ueJ2AY
l00m99z8uiRO9T5QmKKB6LV61Xc76anYUCDlayZ8Fw7HszPQqN1mWnp+cKNj8Uox4zs7MMsWW9cX
1a7NaReoSnXd5c7NJPJtRV2ebj6LFVhIfkOqIm0p3PwC57aCB6wDiqioqCHnoPjKgkAyI4gkVqo2
CpxaWl1S7q62WRVCy0W4de40iFt8TXnw7U2T5k2jibXcJf0/VCOXBySxKyd2ASLldW4yiBzWwrON
0g9f5okw8WDHwQetciTngsTGr2IE54y2E8PtioWcuPrpz1qK7JiY2NOArjLGrJEZ74+OK+uEAcg0
090iov2uSXayZ/kAUcJvh0SjJgkrHvKQVd8tXcSFLTs76RDrTjip5UCt80YtfLzXnSEfhdWTaTh2
nYo9faph1Vpi9f3rG/ajenLP9dgwzmA/VmMSbQaS8Y+Cj/6p9+QHWUi6LOuSqFDTXAFjF/h7YIBE
5RK3lyDxhZjAqSVtca0H29UKV8+mjfXE28xqECdbJQx5GDl0g43RaXzXDjchy+4/GStCTpkSPvAl
zvPmFTAv6oiygafj/3yn5GL/qWDbunUxlGNA5V477A+b2gWWAKasaoQZatxG47NXlQmkYeZbU+aS
5rCHmh3tpr+STh4Y6J/4pUopbq33sm7jXFr5IBIqLC+l3PlTqiIcPeEnGsDsZruW0+jbNLVzNqlk
QOoWfe6ArgOveEIi9qnu2371UzE1W634Oqg2ViyJyCy38D23uutzEip0iz7YsHz9VeOP7E0GrjDH
p3E2YrDsI3IUSAaLC4bQqj+xEr9CH50xNj8WtSB2HmXc3AYx3/XynIBM4QTOtpnQdYxxYH5dj3jN
bkhxNe55xEqjxa9RWREXDA1PNPRV7ZeT3iInxzOW9vBlbdHCC+uFrcafajj+S8yx/KXAgGhLVGC8
AVRE50nrSdFijf/zPpBKBnCtsnFQYymGKc7hAYmB7qPt68rOV6zL07NhRFuVTWbFq0U4u1VyJyJJ
zHek6W3DzctWGf05NZVNn6/YxaZXbia/vonH9vZzaWh/Bfwsvwni3TjDEkfNyLOGUcq8CC+B8a0C
F1knzzyrLkUlQMrN/mpPeemL1o3q7SaOi2YwfIjZzk3cjVoV1vwiMhtbYXaLH50Rys5hkPWcUryL
REEXZbdFmFjbgSMo7gtNDRpOGDQM9D7G1HpHMwZs9LB6Ux7mMsj7PUnwx8vQbzHPPbxQ92eClhTd
b+SZrU6/Bs3I13gK8ygzwCeN31nRMLAMK16RxIZ1YLbG9FdJrp8jn0EdBdicp2iQ7nxpewaQl3HT
psIqHjolQyIs4jmlJHdVftU5Zdvv4dyTKoOJlhLQ4Y4kQp1HZTA1S3fTuvnl1DurVeBkXxcdS2K7
zL6tz6iN0j/5GXq0kHnbb0S3S5Na3Fu2N7JqQLG4P/UBhcxO32kT3grN7xDlew+CTKJRlGiL+TxE
yWSyDuBx5KPPEpmPqklxEXYZ2TS63OXfeKCvFXWmOFJapacmViSyw3cyKVFKtDVvt5N+FrU8AvA4
OEdlR1m3vgQQwO+PQY1+2qwIuzMPfnJ+lovZ7HkyA6SuTNLFTwfan6xeWIDH5oLhL+XxhAUdOP6v
jwkeTriNt4Ax4vRuPwR3gwG/9FF6rxvFvIWHc/QrcHceH1g+Y5A3tUFBF4dIOMVNkProPfsRIzKn
zx9uXPsNTjhSVz8sf50noOvdmuUVyEPdoFbODD13Sr16FtmHZKpTWfC075emLEPn+veuEt8YoSHy
z9KP8ZVAtLtBBMMWJZOsa/nMtuqQdLU/lUiTIgwmLD9eWrMaOWXSmk8N4dN1EET2nrbh6ifCwLWM
wZuvsetK5EeJA+Va1uog8P+jCav04jLvVqy5M1i4aRStfiNH3aPqJBOC7jP5JkMwglkWZU55nexl
HVjsWtAcm+5HrBNS4NX+gfbXe1dv9Qdxi78zLZTCo01X/FAiKNmA1jN4qIB5thfarm0QKcat6ySN
+OxwDqqU1YtRjeNR7+ivyhKjTIGBM17N61L0da5N/pJmJnwJqC4BHGm/isteh6R0rOe7nCT/bEId
7vDNDTJ5OF3hAn038bccQSMLiE43FI+Th6eDosbX+C7+DZvKBcyqSiIyd9Q1ZgsmqqkZFAuoVvk3
m3yXJKEcE6SHMtBP3et1+XTstLFcYs9fo2s13OkPRMBFzSHuFiBD1IqyPg4gYhonaj94RztJf5O6
0KG9sXJRd77CtgDebqYQn5Bn5xXn69vN8XhbqBgu4PupYk+3OzZAQFJteZj/0CvkeHpprxjTMYWa
0QU0W0zC/lg6AouPTwYqMVWFsYmlc1QDMkZAseeST3WEQUIjef+X2N1Zz27sHaN/+2qTtyDUrqV4
OSnqWqaajk66OkRXZazvy4TvcZMF7Qv47sQhOrphLZpHLtjHko72iv+lL05LBgzWsrOaZ9U7ADgw
iK/TPGKBJvWlm67jbfb1zCnunqwIe4FHaNYX1KrpSD8+i6WnFSLltikphLLEVDtzV7IKxqo1VrDO
6IcB+vtC1P3GmSM1GZCIw7v34/LodErknZJXrXbnSJYeUldnnQolMegVpZsX+2myP+sM2wu8MnbA
j6Er+3xPjt1s0R7C4ipqRoOt7wOU2SoScG8pX06ecvfvghkXR41y20HLnC3o6jSkFi35aNqV8M1t
p9+vnsQM9wDwXukGQa2qFMprllZ7KM/Bpwy9Y2ztTV8L7Hv6ng0D5GtqZZFPzS+UKd2jE7ZjH7Yg
pcR7zmYBntJ08KIeFnd/9ILU0Z9PJ8AmUyzjM//nt8AHa9IRwMONuaDhBh5inHNOuC6nTZLyx/fM
vZqiki4y5SSncSzUga3YEyo3Y10HqVYUAmYpxoJyC49wQ7ak/p2+hiiP8MVEZA0iY9t5hDGdPtMg
Dw3onVLW3GP+umORDNFfx0Li41W7ZDiJFsDDgNhVGDWZNtuEt1Ssx57kGAMZ+sQc4+kINlr6U3K4
oG4F0Ee6DYOZQIm7ez+D5V967okLHzdIo8WjU58RjPBCU2wsE765Ynxkuc21hWbAHc56fJiLySYa
/P8iYxoI38Edw/NsOAtZoyvtNUsXLlMBsXsGY7ZSfLpPEHZxvUqmhC9g1Kyua7obTUCklCb+xwGS
qgkvVSzsSlH2BOGyGrV6DH6xbigNqVS3VIAv+xvjrEjqDn1RtKe+G6aLSSUi5pi0EsHzT6NKcByB
qo1qmHeBVftz/ecGYh9OShsREO+8ulr95XlrdKQqaC9URiieHS2o5kUVsiNT0+vDWl7r1pSYTVk8
MibVmOJBx3DOvkwBOCHw1UvvuR2e5VVMTTX46nuE8gAnf4nhGK4E0bQl8syABK2BOuBevMva9TlA
IYyePbabhC72TCKSlnvYIAMP76lcaP/axdD/HiEbZbk3691tYcg4VbpGMlP2AdMQIlCyXPN7UfED
F6l3MlcU/eJeeyo7YTaMzGNqUEjaCbEIfMgEjtkuSf7/7ZCfim6lHzntqn/4tqVJIDxl+81lRNct
9m+0fcqXPYLrWCbOcUjhoZ3ROvJnRbkCKo/AWtKAogknhiqPU4vE8yGhYjtjKAnBtsJdsG4e/xUo
aZIesDLrIjK9yneSXO1GJ5dxOiIx7xiIfsPat1PcP9Q1mLjLLi77cKd9dBSt7dfKfob9FIFwpfeT
mWfNM4MRT+lJ9zpGdqU9RlZsjxHUO4iRPdzxeYaaL4LZjGPXokCQWKoOe3o8Pd5vgso72xQt0n14
lykbNpSB1KnjVsTS/BGDOPag6HlR521GOgfRjzthmJFB1tl7Cd9rEkOoMtFT/y76/kfu6Pu09kx3
bWS5hSK0m4KeFQ6GhHzca19FOhr/fhuwJov/9tW30bkjslYc5Mlfq5mJcPJ/0FGebgngaN0bq1l0
g9whf8Mt+WIPktw5q6ifq+2rpEh5mB5KYedpFlLyeteAnl+bJi2mXOPt5S35nRVhP96Yydcu5Nfe
XSYIxSza505UuJR0Rra/0UQjDlyMtE0dSy1YdIZCq8pylmPDfuTk9U+LNIbtK6iRCWQ02LQ8F0dE
fAmWuSipyVy5KvypaYIulzB2Gfb9Pb9w0mxH04EQxQOprK1MLJ6MnKudgamUFSaMRKEJeuFICHGK
jdWelgbgLukC12LJcLM+PxZRpCG1bnEjPnEXAJZ/zeWuqHIiigb8RJAWz9lz9qhVYIdXzumD/m0M
8DuNuWZBk8hoCgHsGn/ir7CpL6NO1j68daBPuTd6LeeiUQS72oPYN1G5cNdJ/e189aWJd+c9gB5j
YqEt9oLlRbr79hf7QWZ/ji/6REVKLceUnSpksySmYWOVeqyrRRTnAtJCtXjEn2/8/D6Td/JKqzTA
drILeozxPrY17TCsqZVFnYLGaSZoY0uxc0AxXAqUPJ4UnXwXCZjtGseN93Rw7K4veRUYyy5SRjB8
HhTLHdsXvglD/gotOo76b131xBlbchnuStlRKtfRhhaJK7U7M+T9JeRDK0HtB0x5OYd4/oVaP/nZ
7tv2fbVF1ggwBJuZ19zSHBiD3IXMsnOyv8Fiuit4oys6bCpV879+rTrd32ptVdWeDrrOCeDDDuo+
vE6910tkueHX7MXAovfljC4LG5qsneY72kSDkwfboAupWYFURyTSITmCmdqSigyv48PvuFpSLwEq
p3mpBDE4XKRMkDGMkp7DIdGmpErGA6ZPUKm8KT3H0KVN0qsDyRudqOz7c6SfTUSDY/Y8KnAMIWaX
1P1/WMtxrAs2vFCqGf0HF0wFcqOxIqHmlTE5LwCqAYofw7pw8vn+At/Wbr95gppoB9VvOePAcjyU
cIOTt+5h5e/bbWwVGHY91FpyoAOybcYIryZEKlrPO77AVxrTe7SR1m3Ng0eufNrR/hb+AraRC6o6
xXgF/61BQ7v7yAUc2FHPDYBWCxoWKRVbHBQwfN6vqL+JFt/5pfG3ZPZmbvUknGKaSxvLNH+PDxkh
Ypm9AWINgPkYOdLkdXXbILexkqs0yQ4KCWEneeAMFziCxqA4TI0CFFaAej18/6fbOTsDe0UaTFjB
Ky+nQTccRU64DYH1xEvU8ZeSZlj+Vr/Fllutj+ovEzkH1vYSwLNB2hh+562YUAx8N2XZGJX0B8bv
NyvUviTTqOP0icG9nFzzLZWJ6E9zMWrda9alLBj5axrwxs1YVtByzVsu31XamTaX0l0tldLXJ2/G
MBOvMVb0vp2ZSvhMA3UmsctnrESNJe5uIVsnJaFLWsl2PpNWQEQSBc3VCCkGK2wqzSHpPibm8UgF
0RNdezc3B66/vBV2YtWMHwOdHyy9CPoxK2kLwsh5ia8B+je1YxmQ1LQ3cEbQQZqmWGiSWjaitDMm
+RJ9dUAwnppbYIeImAngeyad9e2BUXWV3l61eLHWD1dgbCdXih523JqcrJPn1fNmvkHmPna55bhT
nvHCI1TPwQnA5hFuZMDLONZnuInhYWSOSq9JrL/vMkuwA0SinPNMFyQnzsJnt+ug9jiBufDYG6t5
w4u+kKxY9V7Et2/XuVyK+OkQhrfLhBVi/V+CbjosIH1osZ1XUpGZvvYale1wdS3IZxSbuxa+KC0W
qASoS2AfZ1mdDQpqhNUzKP+9aecOkoGtCDBQaN4S+BTIuQ3bnjWYUqh0Xdwz2+xkFaEhJ3mKSgg0
zM1hFE+byM4fDwWzXnttbDCF4EpiDywNyGt6AwRPhprESOV1UgIJ210v7cGyTEYqOHlWct6LhB6D
xfnnnUkXxEg9vRno5lz0XwE1m4PpLOJmNPhsTZCT915Yd9Sx4ye7s/+WeXh2pzK8Pj4wwVEROu4u
EmZOXHBff2HsU8lVZq5YHrXAWkywfMi9Gb2375/uoRaYUYF1JvGwNwC43Cq2Vcp/ox/4CvL6/hSU
+FuFzN0FT1t1m19U0oJwHObQCVYdoXlhKfO17K7SnH++e1qKpLLogePrx/56cKtDPFySp9ywi704
irFxK/Tu7AuxEF8AKPfVnGl+jUNGpJsUCphvA20tZEqIuRTPkq/uk6UUI7vy4/gV9+xZpd/CAY70
5pNEO7g1kmcQG6hKcGnUPIOzo864AktEBlGCeCbIso6vFlG6+WRsR+y/njOoUvL1KWwIhQ85r95M
RTTYl/ESIQq5BO07pwigHnxKtlr59khTG3OfL7woEJJVYKQbnX5ZG5wpl7RQJ2Makojc9dUmUNNQ
TwL7n7oZ/R7st4UnekDpZljUSRV/B744YBdqnQu90uIDQdzjN7WjOvq91Of3IrNpdsonPvAawYhy
Y5a1EH41EKZg6mz8sBUJMwxDWyUZbPQ6xyoKCZELSen9hZDo4+LOiNNiO2CYB/97VeCVe5A2Fpb9
ub3ebePtPt6Pamkp//y31rKSNN+0wA7kwAPw/kgH1h1mbrren92PX6krlY9BXuGoIsGR2IUYsqu6
38SpLUQQk1se1dEyn1zi4UhSXAePfb41WZFVE1/8KlJN3knCbYJp1MB4hU8O/3cUdp1cIOpovXw/
RHjWmR2eW4C+4pE0LDe694xkcY+/5OkH/IEpxUoc1qbXsQif4fHLoG42Lpl/ZeujEjrn43pvqN77
OcK/rWJYOEsc99fDv33sabJBqIgafxn+a/SMKsFGUQ4DNPkxF0nRU42vV9rZPyZNHlB39lJa0vVc
yPMA3OXoxZmQBa+WbmI6pBpHCUBy1U/LKb+fOQCS0jIiagtNrDTjpbpSpeW9vn/++Z84h30ow8j1
CncIM+3KHiMNZLnd+x5qtbmRStWDGPblfZi/h46RFTMCwImCchgq5YWTYz5Owiyt727cXmNATo+0
gjqh8dhn0guG73UbqBBd6NQutlxvmj6dYNxbcSvi3tfTM2WqBYnbNph5Vo+0uBtUeuZoq+t3f5fa
lQ8e/NOhPbiYjsG44nlgVdCItmDaqRmCOt34RWK5ufFSNp40E52SGujKfSI0CHH5nzJXk/0W6iIR
tOdrY0sJcdkt1XiBRWz40TUtxJSW7lsC7QuCZ14SB5jSrYyrWsohwKt80NvVZV6nXfRZCumHMh22
OtweJ7iyyqsBt32Trk27/Hy5hkO4/GbDabGf/gYNFexQ0iuj0wVrribgjQPfq8QYPR6dVFuoDgvL
mypQTC4MpQgWg/Sbelp2YSfqD+9MCQ+jq0GdANF16nVH3RWwiAXdb2dHUZea0UMOsK3+u6hCu1Xi
FgRcU8Dv5cT83B6/ZBa0gl+LqkXIssq4cUR/7fanlz+eoUKAywKTsMbjaqFCfNsK5RYjYW7IvERh
1/nmggW4eM2KkFY5zl4+VhJB6HKLFBBT6INHc8I1LKqU4ktXfNZXptiJ1wn+x5ztRxY8kcqZclaa
nmc8vdxHhzFRYey2pMzgR5gnDiulNWe6glmeeyLzmBPOo90+sLdMNPuHzAJNQgt1OKJ2qwOYTO2k
TX1/qlHbxZdXWSb/q7MU+HGJvzvWUSejJjpNKe39MOdkKFnYqtyaISqOwLOnNXOMvM+76p1Exnap
vqGwVn8LvabGFqjytJ8Ad6RY+bcqxbugkSaZesEzSxuHZFsbq2W4BL5dp2KhPcFNPDQ2MvoPmP5N
iStmN0oILSyua9EI1sdeHZEv57Y61qjth+xyBuB9OV2cB5e496f+nwcd+wxgMQ1WfpT7yE1nyVIB
ajyIYNG3Ocl2QNPM2/RgNvb/Wq0Df/KvilrQmvOyMh5ocsxV8Sy11mGP8am4AYCeZ+cKiE4Cwx0C
vT2mF7XEwTQ5tG2QwECBZ/JcXvQTtazBCptX+LOPZx910vXNfT2yhAOIpRoUWc2pcHAoh5L6cCXj
dON9iJmbqfbhjWhXf7bcqIto7D1lQdy27NZ1LNkELaJKgPlH1stvKbivTlRn/pYtbwekpNcChUt2
CMCR/mjolxLmp3xtXVnF06IANzUoCFmHiqQsN1Yyv6SFMGuR7GQZkCMh0JCyDZH5rplYAI4HBSHS
foICsv7La+kDWTLEkgxW24uN5nyfWdnmpF1gR7SgOROXnd+fJOMUiO5CWupg3fdA31pcHuMlFJ/e
JFx6Qp6qpWCYbO3pdTgf8YbAzS3ebXHta/gaZFqcWDEnsMGcxEXSgA9KP9hBPD/FW33UFkC4AYVt
sevyd2O2vPl+jULIGb6G319WszeXYKV2Eo4qZG25VitI1tjZJWyRtFGHVzhMKJnr0ZGOHT60nuKG
7Kcc6493KMofnmtUK2ei1OSJOe0W26OvIr9U8qWfdzKYgtTtPTRN7slGeD0shC8wzaQ7YslUb5rX
f9Nj2XEVNlJOFs2fIVkevfhf4m4wERA2OQm8ci5DexqB6zl11I4vlF5fhV8ePI0r0EfdNtjDHQJi
kgLDK474ZHK9RTkOHWj4IZaT+iZqMChxTX9/ts3ZVh21FVg8H5ZoYvCnDDyLAGsJhj2eoty87M7j
86vFmmfk+YNEVkz8w9ZxRwhapyp2w1k5ERHTdyai+KSJ09MQHpofSfnQymupwxTCg4d8JDtmTqon
SmRlAMQkcp+/T1LQ/d0rznSOcGDjCLuWOvkYO3DzuPG8/UO5jkycqi/RUlPLScl24QHqW0AeCjDs
Q84nVrapqOBgCn3Ndi4KEFWoJntXymKWRM1YbXhWoLaJKfgse94Zql0Rxl77oeULqRU8ymzNYNfo
04XaxMlhWnNSDf+bSOHJSjkGp95bGa6Y+5GHeD+QY91mL2V17BLyAoPwaNXWPbDy0AeO2Vw5I/eX
tVmnxm93LD2BslEGXANNdlbLo/RmaYhruuNj2tsUUD5R8Yy5vHEmfxTzf2Rmcqh1iN0VfBCbizZw
4wGzuh4vTijLEvjiwnZvZC+HvT2wZhTO8gIGbfx100x01b0qudirTgSLRvLqLwcQ61qLqQzLVhtp
ytdy3NDfy8IvUiveiwJ/VjwkHZdGAnGRXnBdubsdD3AnrQQQQ9MNpclvX7NIbUeejywDgNnh8Ajp
3y9PIwnabW6ZPmQtAPBk7d3ezPmxNnf5YX3ngy9AGqCyJ3/px9Q2OidoInup3lPKWfqgvpc8RCf2
zvo0v+AeXe6cE4Fzgx26j60bg1d33lyw4svREREjUs8oZSwaYzKy0DDztUqciV8wUgQ9g/t0K58I
XGPq/o4vLWFuEI+MV+xjBfFa6sP0MVQqTs1ifLwc9z1Kg4QAwg42uPL2fkSWWJ1VrRiYrY+TT1Ec
8XTMdcA1DwcWNLBOJ4GywhfdLBFXu48+jwom+X+KRZRI6Zr3VcIG3hyukjnymwfgdlwkgYlcDQU6
nmT+zXbP0tc2zUdubvW7oXaRcurrqV/znTdpdhigevKR+OLalDL84jiIrnv4Vxkz8PrKMFrHSRH/
GjSmbgjztkcJsdVgegHrJrMt1K57hcepvfmc2uaaMK0rkoMdkYo5KvrJgISCOMm4QUqv/DDzrfw0
Ft9uqgN1KGsW4zr9UT8/fLC+ywWTpQzmQYjTWnFFOyndrSE2+jbCOINWf4p1LWwnW3hJr9xQKQV5
CW48WnuG8KLY2kKIssBMCmVK7yXv+pJjTTNcONWoqfVu6+UeXYLfD8fEZ+mMMgzlM1S6vUDhKW4E
4okIEmY8NXoiNPADAkoUnLzxPv5NMa3CGJ+XXBYFMN2Hk/G+iW8PBag2xUO27HfmvGwRYWxET931
tFf0hnWqQzZ5INpIBgWq1MfwEL66hdpegrwLXhzgpzwOuw9mm9rB7QxgXLNLyQ4711I9nnVN7JT/
nimSz20pLXtSlJSbojICdD3PvQjnPm5Dkbz3uEXU5R0kBk9ZmfVVmKwbUMl5vRji7r2yENE5btkf
Weg5zRwdzUhrl2GODIz1/XGFUGJa67LTw/8HPQO5C3BjhmT/+o2rjKq8uqPpD9+5x8ImwIteoFb0
DiJwFvpsgWeAKcqJsznlu2qa85bEH2Wy2DsvjFCpxel77uWzdLkQILjq6yXE162dV+TrUhwTp9gt
Ru3F32vGU+53vTe/CNgX78Qk4yjxKOOWOSrWH6JQ4JuuNTZboujsEQTe48lD24WBD7sdvaIVNeBN
Qv0tu1JLPffyrZNIFNGFFITScraHnMmCba6JnQzfxAdIbP26CcgBfyqrReGjIm9a+MZsf17SI/cz
Z64/R4yZJ+7jhNXp5R301xEGZHYGJ2xhsvKGn/cFiDAg3pn6K8tvb85cIlqJBeyqvv2mes4ZPcyZ
XvyvDa4cJewX7a4uUTHSEChxvDXKqjSzKCrA3rLh1lMjW3MiWLHLAz9c0gJTPAxASqfP5DMmt+PJ
/Y+pOYR9LWx2kgCTQyfyzmN2yfx4T5YizFaobjN52gwLvDxbsVFnt5V4L6DTC15psFPNQXSEhYJS
qdE5v+PGR9cAgQ5K0fXCzwHI83tOYexJxmkBOtI+C9WemZzsmJ1nNqyvMhN0cr0h/NNGviPs4H32
c4xne6wsHzpJw4DLEIpWL78pwri5vz+GJrUaIlV4y+2JzUDI+BpjB+kjsoxc9HTVuDGzyqKDqxpe
Rf0/PSfVvPuY1pUEscebRGQc+e1ASkXzliW+o5Qfan5EP/Klmse8Tmn2xaG+mEOmjqVRSMlh0Xqw
4C9nkvanJBG/dKNuOXsr4FijkGmf9LIqR27XHcWL/FzRlnUWViT9cTA08/a+uex986eG3HeaZvrU
Dzn8fb5GcWJSzgC+WRuE08D0T+utpWZOR45LUhP7GENfWb/G6jG/MczDd6q99gGAerx4V/bP4TkY
dSmjROXkq62GD5R/6v2cdLrci8dXIpZhzR7jhG7fE4HNhsytz2IBOx6k8WThf9sODcZ8ckoJ4SrO
1Ay/y7vCdZtFILONCINun0RiVZS+GfxUZiQt4dwdEL+fm3CnnYDgSI1bOrH1mbobF69yHDdmS0qb
7F7I4oOiOwyHX3xdv+HT4kKooGn7UTwzNvzSSlBn7aD8aCFNcnzOMpjph0xASgiV9GSBFEH8pvNO
IJDVTQFH/5W67b6qDy69k6h6b85lYTu8RTrnTRSGqPzn5LlWp/crG0cab+khJdTugj7XsBb4Hbv6
SmBMHNCC8uIVYxiRWHEJSNpT0Dh/utfUhBpRoN7E6z2jrl38bau5btW7bUejDK6XcCS0pBz4gfy0
6oxz+0a4cY95lPrjsglONbnEDIfj/3Mm+cU00+6toq+kBQNPE7ys+jKXgK4HDFqOVleaYa8txmaE
ENm1+5UMyrHd4f+FEly6QNGwI3/vaDMymt2A66YcFB8EeawKcLCY3q2joaJDV8XhugvP7aVWfg1e
V7B7SO2ht1YYE7MMgJz9qP5Z9MurF96NaShvVojKKOj3ARrEdvIPBs5FZQMweHGJaku20OJB7fa5
/j4mI9LsP55yoEfC8YH4AaQXcuC5l2riBzHxOO0siiM/QLvoW7NjWS9qoPcQIpgl2XfqjJssFVil
lmfnzGYnObHHz0Vg3SWqOjs8jsFM0k+yfu+5oCc9UuwRfqt/l9yhmKH1v7gws20k+6hOJVJScbT5
oFHfsaNesBpDDkMdxFk5M0wQd3uuxTIEW1Xa6RTfiSEE1CAR0oroVuYeJWmINPDmu6tWW+o90Ks9
gN/7Ybnot95JXh1QNw0j3sROfeIbPKpvPXdT8cq0CWy9cM4hsNDhzJP5XX53KmyFVDBNUGLYJO7G
0RhlhjBhaDD+JaTDVzG1NQpan5CLPV/eP+25lKhkQYsDJGRVvzETXtoROPccQV2dLEUL6Uk30Vv9
sfuncYpuxx6CSRsB2gc2gocVcyzLsbtLP5Ogi2bGi1gUEhAcnxqFamqXpKvMV8gl7jNXIjM5jImZ
4KchHa5E1tFaXio52IcRrO9QBCyzDirS+0n+j3PqTgMCHCJuCdJB7V5Wh03DTJbvGBLl/IGyUBCG
FNOkAs9pdNPvDhDKRfuI9ABPpjegwi/8dWJMYgtB2R1b8q5Ssjz6Wx0y5+Mdwtkq2BA09qk+WYvE
68vlUdi6UZVz1BcUyi3BgIzhZVlsBDoFYdEfIUPGeOqzLhSfBsroo2lmmar0McAFzoQndVOTrl9z
wYzNz2iTSgrhN0cPWwzAMCYUYYgHlikq0ceOlCykeSUhM5SNx5WE73OU39R0S1pqKfIfuOZUYnvO
AH89fpaFii/4VrFTT86Hsf0GSrSu4v6ZDkTHBR9amwvN0dvlSWrzdVxRorwwO8bbyBcZ082Fgac9
6ZumY8RTirtDqdt2hEuslYrf/2wmIQJ8ji7thoEfCy4luVJuES84zSoXkGwOjLRCaiNipF4/yekx
KUJC1JZLAaw92qooeI+V6f6xQhS9U2DuAtM6EfoST96qt7+TJZ5b0eoIvfirHSQB54erncYP/+1q
lFURcQTKAb3gGD9hncnpHT3Yfv82Z2/7wm5SmwUwpG5pkJIV/l06FaG/kmp7jmv8LVhjlIGRFcv1
T7tJY8FRLXBkkS/i829FsRwk1BnD4yvF3LabOLrbuiNeHMcYsEZ6vCCJC3Md+DXYAqNVCkhyXJgC
PBhoGncjBEW9lwuPv+QwHgTc/8GTUZ5DBX/eOg+0bR23mLZBqRULyGtjssWu4JRWJEC8VsVSmJW2
AiM+KNLA9LU5EPh5KX2Uotpj7N1fcCO7EOpg5EzVlXuyiwytAHV1GEXYVJjPtdODf4l9Xk46sn5q
ASt1Nt1rB7k78xfgWAlRFGAtBMmQJ5uf8ZuzhXPK3CQPAMg5FT1/F5ATlndXEPQv4Li1sT9cuhfl
SmcTFrAVB+YmN0doWtsbRQ0z3Vk/kX12OANmxoFTLvFKtmWjkErhfUPiva3m9z5P/Aj2ulpZyBR7
NlBgc3XgyuDTxMfmMUmWM0gdcpL1YVJtsikLy0a7kJKSDnqldNhP+M4jR3VvmPYJsZpy+c4hVMeV
RDln4I6Jl3rGfVCXUqLgomdhb/juHGdgdAm+yLyKs1yM3FlPgElCXDdHSZ1Z+cJX8iT3e8mA32RG
l4AE67Dki0ufb0UUdkQ7s6LI6qIh9bWbkWx6BDWNmoVbkM8G5oVAvD9NaFdlsvCRP0Vj0Rlc0kmj
2jReoFYKCbIzxrKuz2y2xG3eRKdeFqYwc7rhaG3yPB+wJL9Iw96/yJfxF6ENhLjmkXicI8XPa1pQ
bDO4LtJLfTtbQtlT2YNX4SQOii99g9t+Mx1MwE7f7FoTsApPFHmqG+JUAQCLe4T8AhdGVjLqbcj1
qn32obA9OlAwhR8jN2Yr0LNcDJTCpPa7/ujWySVmSoDLsFZSaFu+OjJzUuMfPKo1XuTqyoD53lU2
Tviebrtt0OCImJaR0/uJeY1XK85RGmgyjtakusPkfB0ASCMVEqz2BQ42LUa/Myft2xJXC3sJuLvs
1UH6NjC/4plVmkYvggviJ1WaRXAe/lREA0YL+JQuVN63YSBrnnF0aNqXCxK98mttNIRpwmmn6XCv
Lcy4xP+L1Qr8c8qM315tE/3WuWom6HK8EE3qhRliRFesLxUAexZW8wF6ugfhe2mNTh5wC1+2i0e0
kQHa/LE1vSZwhjAvgeqHefyLXkHltAGky5bvIvYBkO1xUD6wzfWvQI57Ov7RaDJmadbDjLU8SAJN
/kohDfugxHc2a+plsXDaWYOjjdHh3o0OHX8zzXohgwaCRqH0Ebb3+ZJZ/i1X3WABmavCjbBVgCO5
3+aQKmrB38SMaMKodkS9cBr9AxmUal2rJdjQkxgTctglYIKk4CPqhmcQzwpTkkuYcivtYzuMVej7
OYda0guzV7QCVdk1craTU0jNinqgjyVFA3f2klv0NtWq7udaLMbIrOeeWRePW+htAgE3g5HgCgEG
VFEeyZfxvb4m72RXIt0L37p5HhxszFdEDHKwWq0iXHoN2wEGv3OWcGqSBplOY9DSBzAhNGFHjMaS
YqnYTKlBLublZt9zuGW3xs7wiqoOoPbbzIz8bcNbqT4RC/pV1rbnEjz1IRcZRI0IU/eM8oV8vP/i
udKxOPd9TqcmBafhVup+Iu7DPg5CaOzxTJ2u/nJeMbKhUQtIAxADCe3Ve63GqO2zm6NMtn7YluMF
PpohWJisgevqLaBKJF/9PINnbU8+94Kxy5KWvb1Yq/QXnypXnUNio8KNuPOyZy8d7lLNKvQY6mEq
1H4VU4e4NNxjQlvRrhoM2srUQzlLLaEGg+3kUUoJpOqNU9yLgAn4TkWf7r9dvVj837H4A7mCeAmU
oiRyVgR5zQPG80MbrvH1Uvtc30N6qzXWQrwFTZgdvDobxY03oQukTd/CGUya81bYPspX6/hzAKuu
xopRu5OFrL/4t6iShjl3oUEyjt5CBAJ2kBWU2o5wfhYnrH04WZHAEc8jWXxcYYfkUWJI7QvWAjW4
QDGVQUJLvioXUtQlEdAEVTpeUZrsggSY3GwVts78SelGK4/vxEyQTO/MpUs8uwvH2vJugN8QgznG
ywhk6MnJqB1GYPNomWlGQf9HmdlfKheeX4Ae50fsUnWk73ZUtCOvR7OCwi8PYB6I7cgIrOQ15/47
lzTV7ah5RCcBevTpAGD8dnyv39+hxkm25b9Ih2U0aYNvjTIFnZ50nsbkywTeIL8AofcWYJXEqicX
mM3t91TPY0oPXf6KP8THPFZqh5VSLH3P4zr7QJgfimSxhbyl9NLdE0T/EJrxbucw3VnFkpH7l5lq
N4gFgf9c88wUo/QnLM3P+zhOjxPHYXoS2TMFTHI93aoyrzSPvZfgukybsMk47P8pwrDB4sC5n7nl
oGvyks8lScBQSLpkhA5nar7GLeVbCl2navdmEVOpCic/1D92z4C8yfhPleZMx0KTVxibIO+ybdsx
WCuaIzRgtqUX7bOzzqV5ALnGARi9vA632tYMdybPSyz76gjOORFywBFTdowNw3zVz+BvFnOvrN7J
DyF/itLJK29foeftYyo+Ouz0SmjjWOQfsNLjRGjf1wAX50jNDODppEXktijIf/v5wszUemU5ZvDe
ngYGIZ93A8VS+mnj7tRA7j5iegRF8viBSWAs1+s0l2g6TE0kCk09sTUXwYpA8XsB5ArFpKVA2c0j
myikDl5qKkxqyx39UmeHdbXfd4iKMHjgrYuXd30rN6mC2JpdE7h2sXqTr0V5YVKpqNw8FX7Gc3cL
GZ05XD5qK5cyD0sQ/0Y1uVX5ItUDbh2Hs9B+OWL0yTgQcCSBDj2RhwvM/7Q2ByoYsXhHQdG5k7tP
9kAPGg7AtBSDo0CVdFfyY6gPGx5AnSnaY8CvBoFMdfVUVCjoibq03J2suViV4NLRkt/NRhhlgjJH
EkgfYR7HZKaPgyWpHAr4mSufbQ64sNNgZw71I6O/rNt50rgb04QskSqtHj6iUsSwYohzvj1FO8JW
TK7PEVINUTW0IxpgTCq0mNBqaOi/N2l8zJSvaIS+U46i2LVoMuwC7yh/wM1Rxa50fNf5Y65Kicpl
ucD1dypc2SQQB/47JebkqF9w4K8k1GROoOdQgXrTp428ARfYXlCH+BI8Gx///XMZEdRapNOlfWCM
1ZRns8UqZ+hePtAPty5EGa+AHOEuUZnCuto7rQV/vW/rMdy81X42tS5lyMadpSvjy3LrVEig9aR/
izAZq49K4VEfC7lZmqnhQqXPlxOlYUZRcJKhF0kvs1JpaRNbut2xKcEBDH4s/385tT9wU23IJO8n
TxbvYytp4O1gIE7DpfIvCAe2YatzzDzPmyUXHmMM0ecFVmQo82RKy0oRCTxAZP3pPscjUykrxlA4
qNvGas95rEmXP1ZkcE0Y7RurBjDbNArDztj2Aoq4Ha2QEioo9rgVKNLIPkh6RpN5tJQPcv+zZFv9
OBVZxzuupsGDlJkUDySvb8nQ8HsStCcSgiTy8wmwMIjpjKXJhCe/+cwqucX20x/zbMcJJMPyIh0P
gCs7iH91UNe5phNbw09sEdARyV9q+BZYoZaHkpPVLYQKuH4fUmEK5u6JNPjauVYFTW9A1/AnY38G
lSBc2l805OH4PAlC6dSDpkUlvj7m/7U29UBFU8dQ+vcX4Vi07RDAxrvlHUt4d2p/YPm/LpjgXCHw
wbBBspfXB0Uhf3bEgI0A+v8iWXF4P8n+qwZqpDvoKCF2DVJTliPoXw2lqefdjde79SAZ0fpJKj4G
3GCy2lCZBUyedJP/mf8ywB9vwwzlRyiO/gUG5C4Rj5kHwxeDhPyCzFoJ2uTwfL0py/zcsFkHzh63
zxKTTuNef7kS3cGa2fsMvuByY2RSSKlrcBJ9OudPSJrNCKRNaLAHKWClKiXRTIULis532ibEtHQz
UQsDG4scotFslNwiZ23VbmFAyDoGVolT2IsOeKf5/EeFINKIRIwMkwG32lndlG+tSD53yVhY65Ew
l5Esu09x49k4Xgfhbsbn2mom8u1St6/fI00/9SGdqEYsFoJeeAT3spXxzJl759OZbgYqxRwWZuDj
U91+yW+uvKfhw08ndpBtylpdpZa7ihxD/ENxRB8SylDxaH0B8NfzGGn3EeaUro5XngWOgPXPLIWc
17QpRgogrQb1Uz7nDVyoRMrv6LwCcJntd7KYMYVgPP4Z/BesozlIkkXxzr+XKt3fhvkzPrKqodN4
p4DTKzvhvaAqtbKBD25M3huIgHhKlJJfRtNC2RjzWMOl4LfcsJ3PoaDjJlE67ejapu+gcJlKj4l4
CM3+3NTLpaAo7l8uNcw52VhoP84StJKIyoImCo7AfRx3R51NxBrgiwMaSDUMuCLo/nT/L6L6oxhT
TUBdHlGY0bHczhcbbCX4QS2dJEeF1HRAEcKe0P4lJ+pi4Axlb4WD/Hje9Os5/iAhjSScCVIED94a
O+RckpBFg74rd+ua1oAw6ZbdCyO6oHzamXfrHUf3oWylfb9WC9mo3kAcPvmowz6qKvxxYJ2C1Jie
YNS3CubBvzRxpcyn4ghT5OOTZuVuqBkPw6ZZMtyX77nle650mJqfCE6zpSQYog6pS/JBfoOoQsnf
nYiWAnrG4rdm6BJhBC9lH19HSPDYPcSxnH8RIrGbgWEfB1c6/U3Lic3oa2wzPz8bTvoq/FCm920D
t+aGy5lwyLpANqH9qAWSkbvMisNkxIGRvwA6REGRzGliU5R92GQ+N//8YlR+7KREYi54y+CyLEHL
Fd5mLwy/cTHsPSMZklsEM3eyd551AznAFHESRFfwyNIj9Z3ILgJv3yjUHX0o7jPynfvjlGPD4FmY
CasPXgy0azgncaWRdJqFfxrISOWEsbyU7+fVw9UtVDNUmXfqrksI5hBu2bS26pHsyq4N0TPqQESM
f12j08VraO50kcwctJqcHGSIuLsry9/B38yMi1sjbzHcyg8fz8RYgXfn+FJUjRXK0vGdF4ELNmsl
Akf+VMn75LsQlGYvEQPkvU/6l6qdAR0eVGEiPNjo5AqT6HvoTEeNtz2XF6vdlZQfWZ9tcBGporUW
T5zP0nHqhY10hAIZYJXaDPFr/ggNpq1o4ZJPun+pC0hjh1YMr0i7dxBattFiHdELllzpYIlM6uag
H5y/hdD2lD+40C5m46a1evQjEQhhUb6IE2HdQYCZsW1tDd/vWWfTzQo4Xq2I2D+Gf7udcVVghzji
NcR8ny/vqKni0xWvM8cEKBU2XXBO/GS0nW/2tI+cMoq0EsgrAz5JM1Oou32Cdp8Oo11CC3MbgOm7
BERt2lfKsSCrPcsfRMblks/hki+mEcjI5+FGvDgkvBOS2wvpaOXw2AplSKrR/1KUsreooajpgss8
GNx5XAUyFZBG4yGyiu12JRRONbJejcPiXrWS8pg9RCWzXjL5twWn9NefVvftRjedortNwsoV/sP4
pQPbFH5nVTCYp/ITiOnHS0gExGCLy2lCvyIhB6Cov/aukkf0oxEbyGpyHYYNxitKg1q+KV0RZiZg
laPDO6ocgPVFwCuvON+Pw2whk7DhyuOfBfUH9e/YHSePzGYS8N5ROTbGB7S6BBLv/LpigxuEMrOx
43aJj1Mu7XeV9JRbdHE4FdyXEGX2efd7unb1fWLtUgxxab/D1N6nM/gA0v899bzsZ6MTUom/QLDV
9XzcdYWjZscXXbmUOKJABXqn+PBGGee7qlIaXxKyBhsADdQJp0M1wuMjT7993VAuGg6n7MhfGcbk
fWfiOur91r4ecP9qNsP/oqjfSEudpomtqt+i3QQcfOhCAeuu7vENPB/Bogypa82GH5O0tnUPU7U+
Lf94ueISRINArgiNF3L+KFEnvFMvzJ39qOXDIQwTI8iGX7u0xMPKWJyxNEMyyFAAlvsnO2t/7/8G
9GevVyrG9mKLfyQtCSqautqCw/OEJMD7pLAvFf7kBCnhI59AFx/vvqdmP2dGK9Aa1+4LeXMAxz66
UnnHt213zDif/bg21blcS/UqnDEn9UKFb1vsIAPemBNiWF85/GGYXL4Pgx4kaKQwvIuVm20zD5LP
PvI8uVDmS6OAGU4m5p6tKZWsSJhfzlFhvxAIao4pmb6Tnnia03BvcEYkBzuAwjdWRnLUYSXmTa7B
CnRdt4NxwYGgCcksTjGDhIX7RYQp/9VaT12A/fcZNK5NkJTKONZY4kJ/HTz7yZHiqNMLE349r3W+
7qBr3vBJfSIyK8u4xe6C0msZYHSFz1kJ2tq8GTYP5u6tzy0JkReevLN+2Z9iTh9Y/GkSW6HYxc/E
apcDiy3xAAd7PpkRhiyncvKO/tlZ4wZUIS7aQtsgIW0xrCs23uk/QgBks4DZtpw+TH6Yx7c4BiFS
CKYFPJFGzKXDmz9ji56E8WaWVT/Om8hLJM6dArpzRoE58cpu3vsbgwloXe1BW0gDtxU4nWoZyy9E
WTitGew4pTAuXxMYH942XsyDy8Om5gfeqdO6Wp9p1OKXBAVnlTQ2tGIXdn2RFTXHdcYlYDLV2UlZ
pOuld+cw6PJKAMTVs+jE7XmokSsU/6NyGlFigjXxZbQ8cuIdR5zXifugy3p8yj2E5fbnXqJFJMzt
ngRrMwcTVQk2kzXrwN3MqW8DH9xd9m/FrPSUIPEUwfcoVRSib7lStYpx4VpE8B6Ga4J+z9hoOAnL
9qKoMzPpmPNSfanrslHY4SKKihr3xm8TXIrscTrF1uswOra442zptDlqr6GnNKRP8/C7woAeEaCt
gMPX47sUk7bRGVm6hxY07FGkh0wn6XmlFmURkE4s17VjkDtb6VZEZkmBSFNAihEuNjSA1sDdoo6+
mFdoDPkB+plu5nT5KqKS0cNwrmEnqQxWWTtFGdxtSaVPrbPYrN1llUepgWRdWGGQixjhdJCKS84l
y1fSSkL8GU8Fmr6EVMVaBq1NVU6VMs2OEFHmL5CJWgKn1c/0ys+QLyui7uOf1IlhM6jGH54ocn5L
j0X+WXGXqvUTfDX21mmSAjXO2PR1fGSbD7TNTm43YacMq+Yht0iwlyTFjeYa/S6LqX2VpO2smunH
8gx1Boy6q7ifIBTdc3Ob+d3sLDzsfA7LcWs9twte0XMCbOdPzgrEVXV7v+rYiSjPJSCu7jAZFies
G3S44Yy1XvVlNhtbR7+xO2L3RgYXGh1oIRZ8dth2LhgZPbYfAS8ixupnuNDWVJfGZXPPNz8T18Lu
V0qu2vKn1RvrKsiYcuKwIL3+7HRJUtiRCTtO3/4klNsDMAREEUvQzqr4iLUQu/1ySqo0uVgP/Ly9
L/B0SPaBLn/NSHzS2a7f+/zS40B8WxLNq/1cHP5B+XO8XPz+xgc468mAs3wMAcdcSksf5qifw2bc
NUC8ZgDbtE8nyqlqayglGTm6T8PJWg2yR3xDf4KjS1Q058FjPQheTEIh/D+ceD5RbM2YdMDMwO8F
J9+stf9rTCFWos68l1JMfDTMtbplemXY4ZSVUrKcS5f8dJoLP0Mrhc2/70w4idoG6nAPulgip8Ev
b2Di8SKTww4Pct+tDpkhPRrZEeRaZgmpf85GKuZY6DmeLmzreb7jYiUN5GmGtVJcfctMAsmOIVRY
324Rly9ZLTwAEHgknIROb4zdKmnkyRUmWLYVuyx0CL1VAtV8AxqJO+LtChtZ5gIUX7Z5i3Y6TmdT
HC4znBXK+X8QiGIKR53de/vWpQfUcfR0LOU4DqxN9M7+5VImO7orXSIpgkTWpabj2XFVlIXTTNuQ
+gmimN2j9tasx0r9ZJJVyRsKzDDnevdSqIqPJTZHI5N+HI0qxfd6MB9tXPuThdC3/elbNp8ZAeWW
2aeF8dcm1jlN2IoevoANBUXbJT2yr7e7LPgMp7JIZ6kWrdFFQ70KRI75AWfm4G1xoNkV9/LF2Eno
VLwzf2RL4iT9O5tYUOSvyzOpkfawsmVXEaf85cJZcrCefVr3IjCV0k0NA0sX44r4NyGGSQcMrdXh
whJfTcE6y3O8Y78iZfPgXIusQd6aBq7jTWV3T+xQxMiovcysLduVcmHK7E+mu6lkCMtxbXMMI+8U
eGUFT0jfUdbaAkF+LQK26lFqbjoVu1u0e7ZTEDP+3Ci0qQAGQ5Bf0sm6g9TedkCimEukzW6+PsJG
f5Y/CY7BT0Q5qxuHtZkTaFG8f/Hr9ly1C3KEncnMuQ923Sq3R8fceE0q7S91Se+XOgRtbzDQZdbY
DYQIL6D34l+0PKPxD1fhMSAjELin+ZUP8W1sAPHPLH45QiXRAF9eaxJl8wPl1sdoFhTzPamsbtiZ
Q40r4kaEeRtmiiSYWEs0ELbNZS2LmYyXBi8LfH0l3PWKEHubPzcIbYvxfwnZBJzqijp4kOQGayMK
AhNF0FHvz69XJiNbvRVwCFcqoK8brPGuNWSTF0tToWym8bX2z/pOOoDCqBh2xdpHQPARZLUa/4LQ
BxNtElF04jW2CEBl/OOsyxv0AUbYhWHIXnoK5r9Ow5upMt+JFc1VQH8iX2h/Lo2mzom6idr5SxX9
YY9aMJqo0PNnDbpMHAmETUBjqyHbLAhH4VT8OcJT4TJBSc7/W8SLO0s377kMaKcLUrX/oITa8IWw
deXWQfzwDwB9EpMSGNc8/rPLhebcTqMhy8ye8QmHriJ2aSzfaZ4zl6vBDXbXu7JoJmuEFAtk14Sk
K8Uro1m8m5a4hlodcTLg/dpsN+xvntwAtSpILFRzQsBmS64sKJSzgODZA1go+0B5fs87TPNgKsCV
2KfMR4zw5CIr0KPEKRd0uyPojYzJa78spctcTXSvMQSCzrjeqmMH3xu5rzNRwY5MD0aXv3bWwykO
IEziePyHwOjFbky2p3QZEuGPoB80ZRKOJTgLhzT7IwCIlOnppxK71iNquOiQN4I1GxCAHc//i7Ez
lP00EDSzQuBCULDDtMQXLp+ZK8tMLcUKKTMukqTdpeV941qarIt0g91WT8djdh2VlvxpWWloBvdS
XeYeCc2QOWrtnyRSb8eSiOF8NYoftlv0HsH1r9O6qti8QqQdex+Zu3fXidDjZ34sEDrhwtcqwjjs
OfhPzjAkH98KfiewZBu1CRPezsbyXVJR3+2K+lKYTBx/de7qn1p2acUY7VVXI8JymOgstGJs3etP
HvBhu0aQtOsen/H4OdOd0PmMpWer0R9MXtKSt0EtSG7q53rqGeCHqhu8CC9HF5vcB5H9LG3dK4oC
TbiP0WgffjDvMe+7sgVSuiwY7hTugPrEsGnlrWNZKMQaGMEMYiIVqNsruIo0rp8IQ2yA0tLUPu3Q
MHqGjIjd1u3cgliVRnTy7QfSEKoejotnzC6XVQ7+p19+ESjn9osqff2p6vWyWh0dW9aKdR2ftLcE
E/snKSHdUzG75c/HN141EyHNPTF5WjLvbJoGIMXpAG/GGVp5BpDslh6j30jlUau6ZuFJjGwsRgMq
FS0GNzqFAYf+XzXE5a8jFulS6fQGn6/B/H22vv2VkhpMmmNisd0w74u/4VdH9TeMv+Im9RZsGD7P
Xq2qpItzr8OiW3D+n76IJxBjUiTguYZTHWMbJGvzboBceOfHZ+BEoUCBuelrrs/Q7QUghPXnNPOF
rB3tpGmSneiwE0052OMa940SkK7EsIH096xd7xRxLCcE9ahuE3i8/8a7thVBZCCpjGDPtNzfa0Bm
2NC4Ljp2NvEdIWlrmonuScjRigNqLDQhh0VyDOBB3A7OskBmQDr25lCX3jkimsEwl9ndeiUrp5CA
BILA+QyNSHpylu46dqP65q3yf4jRFx/rQrtxkp9zf3x22Q/dtQYiPEgRAHgEW8PoLLn0KgRf/YK8
Irc+q8faCk5IymVFBL5e9PAsgFgzeHjLsHP6G8/K1dOYSz5MuABm+N9Pu/MRSN5t/kpbnIDp6OQo
nTSyEVehfRl/KvDLPApU6zH/L8e1EL50x+LQYDvS1BNjs5WFAI28m/7qdMV78lrD0ZbjSKYOtn/o
90oimwemogLsFIfvBDwDgVAHDskfYp73Z95E67NH2z31v5BjUApySf2zWRNzcjGi48m3AEwx7tKF
j/ffRMGSsA4JA2Lqyw781qKqe900uHVgdD+rxBpsH7egtDqDdPd5hTnaLpXSNRkY8uI36A3zEIag
184H0+H36Gq+OeLm/IAqXAnQ9O4d1AfOPqH6F3szcuGCoFSyWqy+nIpRjYU/mjJYP2S64SJMVPKc
oaxxaCEWVfZMMFwcQciwt6pgu7HR0HLmp8LLkE6HnGii/qyYxJYpf1AAcJbAbEWtBy7ZVptuGfIS
xi5jIKtkX+J9pY/yFG0jIHsHpo0fACyPjHLOjq081/m5GR7oQ7P1SxbX6v1FtyiGYXzfE+hEFjyi
aCnef5+hte32F+NXya095uuJnKQYlJ1AwEY53my87jQelRMO4HqJdRScAnXATn+k/K/HSMy1/Iwk
BS8qNe5El2Wa/raVE93whko3keBR4DnHTzwwuSOdcE95JfC7Rce9HnnWqop7nqRO12BQyITELjTD
p7Kc6qmlHhWTz+kuy8+uVd40fwmFOXZ6XtRgc4dx16lxmMObzJf+LOF+MggGJNzqhQ/FdLCkoqH6
ScNHb58kd3DhwjBO6GJ3XH0tmu4whNg2oaQweNy6NALXtjgcN/5bDs6kLkFd+9gxrw+ZHNvSKsuz
8kKmB6Ejqx8zQrAAD6JlPYUsAKb0qVfAHqW3VLublyJl2dL01sLkDfIGiXnWjp7X83x8bIsDYeuA
2idlbJP28e0rmWhnxISz83FXtN/gOUzofzw9RkBtYSHlwPA1wuRlEWXdthxKETvEMBTtydhzQAqE
8wtv/6K/5lsnuT3++My3814+/IEPwwuvAwD3z+s5cRrGjgnVze5Cst/cBRtWHBB7++uMPcdzWbDu
zevt3uQLIoTlZH0DE7Rmc0wBKE4Fo10ZZXMVcz4av2s93/geMfn05gdsapNPIagBGQZ5CVdnH6m3
3C9/dFv7iK4rm090ux0HiZOOp4O2AToKxeg+P02+ih8+SMJ3NefFYTJwvdbCNGTmWm/reJ1NkmWC
FsxO+N57JgWFsqWkxnJDE2ebIKISHfyVk2PJqBAloYqU4BLbTvakQQ1JpXiQHZ4onNOBY4KdkimR
aX0Wo9ukcFAkEQOBrsmIOV/8zvJGTnPTtKyPntGmdJEU7QzoppjKt3VN5Q6l1+h+ryYXVkN3IRcB
TRyQMcMYrM0G6J+hoiW+d9KO4B8kMUAIqkeD0pPe3qlo6BeYJ/e2iojZB9kdLD1184nkMaqpvTY3
LkHw+j2ru0EKT4nYzsEjtnLgxpDbK6IgEM1eLDoL6HtUl7rG/NspUyrPwwfnY/IjRLDlUg/+JZQd
cydHJG8siFhLELwHKz2nGfhXxUri50oIfGO6gkj+HneCO1qzhkaTKvuzV+Yj3t9ylbV4000Cvnug
3vh1YGzx0YV/tQQM1N7me28UtU+tT4Mbyl5mHFSIRnwHxCzwTmmaEd6x1EiOwxrjBbc3uB6WaWw2
/5YKfu2FcIH5i/PZMVY8KMFQBgZTYQB92+QABUmcvXsR8a7vn9+FsGGEmM3dM4wcJ8ItugBBv38I
U7Z0UlREQ48rmbCmmHEtYb7EmKk/cOWVZtF/UjngMGdmMtcTcn/edoNEkXkwsgkvFNOb3fzFzVU5
yNOFMZkiZJKKL2e5bQTG+6gbL3UmKF5tf5Budf+X+iwNipY5L48bJrKaPJnZjDCXxiCdnJmlj5PD
PeWAGcO/R3lTEB+FNbq3b4YVF/6WogUjZ7T9QJm+TkjnkiEpkQ1/SZ3TTMm2UWdrIygKdBe3zoka
xXPMtk60ZYYilIiYNp1HtQxIvE9Hyg/msWu8Ueukbyf/aqF1OLENtBKUTJLoLbda0v1L9PMDIRaC
TvO95JUrUvrXVTrLhcl8aDqCYA5VHBSNGRkOCNo7n1hTS0X6oE0fU+oPE65CJdtOA9ihpaDR4HCl
cK5I+2uM1KDq5UgMuhla7Ye6zUsMO+1tn7ouUJuRPj5X7amy9mD1MqYE7U8F/kUB8v5B0Bm5X2GR
rYhEv3AAUMyeeMyeqHk5fSYQ5660EW4S9bTpQzJUPsuR7nppOHIAbU0DR5etUA6zDCB84dtqNJrK
27U4XA0NmzOx2/nHx3uGc3aQzAZ9MOO6HBGMDC3V94KaLGujQSugDZxJeej8lqVbJK/Y/ZKshWSM
z9T4EGU7N7DIIqFMnNCBdsXixNXJm5raEh1HY+4N/6szTz8rPmmnHJ6Sz2++werm0JIcs0PaHRvG
eKq2hW6D/27a3XVrsI7kFpbyqpnadxDRCIFgE0WR8LpWHmJ6yX0/Y71abNjo8ARUipOygxPnb7h8
rWendm7iX8AvkzfLOQU/T452v7dPFXLELbisJ/I/7LimMJw7uRMEGD3ns5aKyc5h9wGamkpkzgXF
c3GjDURXj0XOzrzj+sFJ9MQNAEyrUMSEb5FwdTfWigJPTHJqXqSE4CQMFHiakAKE/rYKYFzZbYFK
aGFb6jwe1JIsmGTApNTtln3lcixncVysbphEl39uZykco0jEXj0RJq8M9U3X8qVY1vi7ObFMcv8Q
I5EmNcujuf+d8k/IKhnxuezSdpWSDgl2EGMTz0h1bScZmBUN2wliFTSItQgS69BPFSpzx3NZpo1K
7LK9IzVOhF2tkO20WvTTSe1fKVjKPhSso8JrJN/kKiFdCTe0M00tFK4axBz8DrPr/O7uDa6xBduW
ZLl/+TiysLSxX4gwY1vkbr3EL4qssX2uiNv29xYkIIkVScQQVzyOvijtuyMFSP4md3d3uZVORX2o
wKNyfHmt4tF4KFOlKng93aO1I5Mn+tbxBVGpWy8X7C54WVlZpn0qZawL9cX9eKs7ikpxPUvHKt1e
Kuhoo687iNHrFnhUExi2PTGFIWx/sZJJC+vZBt6d/kQmvWGdmWN84eUw+l8fA+YRg/o379/CLWoi
XnZXleC1iSmoGpUuHd1537g2TqY/new+odLorIJBVrRWWvzeSacocysjId4xXBYdu0HehR3ZIv/d
keR8lw6Eu9NfvWeWoA5djTNHMRtW+SvOG/eMC1uvNuZU1/Mw1nMFAb5/NC75V3HylCe67Zn/H8yK
tjSzLszS+EM2wfPjXXSROlarbvtX2j6qzZFvKRbr86DEtWsSsz/Z6DZzFn1z5vphRyQmDN4m1xYb
/EzHMXLei6jIEDruUe4+VyNHDOci/F2tFnTlcHxzusJph0ZIf6Gs1QGTz0GzJVrMFK5FEmSzMDFx
M4czlF7PgTHCJeJwXl6M8EpzezYQDNTNlpmhvNliyvmvF4pCCeQNeu5i1SPa3OWnfIBshM4j22km
1uyCyIwjmB9SJeDlQFAx7/1nxRvJ2DjDND2Vx+rDtnxt7IqKLQwq4JUuz0NTh/cp+fcJuVat7AFT
6hCHlBcqYckzOjtrWnulR0Nm0bB3GfD3K0E63isuBB8zgLjYi4BdsTzpT+20zhouGipcYJDKKp9N
8Bh8hFO25NGO00M0SghXck31hbnQpNFZX4hHnLEr2dBRQ09dxtTp/B9zf4ZYNRHwj8FQ1oLT2bhT
G8lBSCWAR6QTxLY3KNXK1hFuULBxch7QpNXnoG6vSTouqUov19MDLLHly5T0YzvFopGzzhBvtXSD
YP63N5AuskXK0BxUJH090ZewnRRlH7PbK+Gq5WpBMLTv0EgljQIfH0WuM0EvW7+/qxltzMsfqQKL
h/yJuX8WGAj9pFlHyfIPHBhnrJUbrklRVPrwvHePk26lVtp7udp6U18YF1HOs2RzIQvkfEHu4KXG
fv6Ul7Ff7Sp61nP5MUu4SbicH8fd+CbPYTe4i2eVkR3QwFkTEr0hJy5qRvB/J7Tsy4ppYOBwKHFl
bzMkcwVXUB7MmTL7gfr6strLdCK8jNk668QDMfGlWIQ+E+WnHVsZweR/MEzhHiZkkmbwHnQleJwt
jL3qWQzkT28FRSSWZV/C+Y79xLpSRZAIqFqOQ59pA1qQF/ELo2UmkUxtCMdE6OXLUAahCnSGZyYq
7C2FoBO6X/IuNvhbgrbuxuDCJ4Nc7HIoj0H0wTGs2o+49TB2MrSs6EZtaVo22cRWsJbATQQDaJ1s
r7cxsC0hFfPMsB9/FSPR9AuoHKx9NNHK7RLLIZBSU+RokjlUlQIbfkzdWiZvGf3iH0Qrt3WX/w+N
2m5nC5vvo3WrKnJd0rznLe0Xi4O3IFE8/ZTyWEzY8Cv/a0pdrONHJknB+17dYcqfNapX649OkrwZ
zdPZVO5rSZNv0IIFueyOvfwxWBR2/Q0d77ZFk+febySXfbIZ4jy5aoQFCvBrd+dSTc2hPPSfB6us
/Dx8JyeZm7Q3nREi6wCLaj0/MxjgZYQiPRs+9gBMmzMWPQCzzGGQZxGc7PrKP+IVIT29eGkG8u/f
j1XNm+IMcED25Hi8XZ++xGDjYZI3ir6mSJ3/tAWyWL0qsLJ8FuxSJeus0I6ot/Rfh77xwm5YxXRO
M6Wvnwmcc15N2TfQ71VyS6iIMzpm9QslLOH7L1dvRvkH6Pk5UHW9d4RFWQbTVqAiLzpNdGMQZmnl
myr6h2+hNWCO5zuGzJtRwJF0mQ/LuSrk41mlwXja6WvbIIAW61usgcBwjrgaDjOdbIQQbakCs4gX
nDbA/WjbWqLKlvtIneDdWG9/1F03vErKSKcstHZa4JAAM7ub1oorDrgPhFKdHys9sKERHeceFwz0
OxRXBLU0Sp3I6Piw/7rq4CTxgc1zJp1DIpDRVVSqr6n4otMSHDZLqW841PZ+Q/krCvKcJ6U7EN8J
3dV6+JYPmpDjFR2cbo/eVZBHRLh5p6NVEQpPcYdo4xs00qkrMBGikRkxAcwu8D24CtoYrcOqy+CD
9YAxApakZ3r3lJb7MpyUogUUOS6oqAOyH4MgQdzzA6JUvQF7oPkLtv+Q9BnR9Qk2sMa5c9woeg0R
jvomEDjF+vRi9xWqD2zrz3Et9EW/l7fyZ22VYoDcP2LtCY4+is83dLM/b0U7DRyl5V2V2aswU6P7
hK/3UZkfySKiexToBTnEzlshHg1fINUIwMcWofMtHInTZeMwkWZdh5x+a7iNdkIcz45qVdKenlzp
mz8tDsHdrxBwSvbqczhMkGOTCyMixxF5Vd0x7MUd2hopiVwRb6vk7auzEdKURnxcaGlWh2CYNQIw
cMx0ZqPYnpSyE1zBz6FOzCuLB840TOahrs0j9UMAmmmeHUPPWvBNccyLUQ095IyP6QoTSpEHcvNw
H+R+PesRGRrnVHMpjmDfKoiCeb3hFyft9jn5NgzGK+k7sxgYNelxdCIzZSjSFbEqgnPa/61ZOyMD
Jf1iywCrOd4a0SfqPw6WqrDvIesO7Wg2dB4AJh7BKeGbWlutgAggwHYxqz8qfjeUQ9+6vrJs3f1f
0y2QyLB69pLocCffjDwS7IsSTqQAOWmNIiD/S5c6pD1g35TKQViCgQ2pO8lNcjaWTPRPp5d5N/05
R38hqv/qL8Uo9tm6MlEupc3xfRso691X0r44Rd/7xhk42XLfJJNgZY2CCQqVlaGG5ItV2x4VNTz0
f0Mu2NDWkL84vvMN1ks5piLf7ZSnTOCFcqL2ljsTZIjWOQDgcKARfifC3ibbnWeFE5jV9PGTQ1M6
F9gsUUz/TS4LTq/RJCJkTUyxbXI802fJuXvGTiJiOCI+HT3sjwycJVOZItqG3FJ7B2xkOcAHkUEQ
iv+MknxBsjJSRcgawKhWoe0FDQ1BGSmu1R9ppZFmjpypAIj0IJxG08+0qrxCKd/9Tz3npGqZJeGj
15Fwa29zRpM4LQzajYlP3OuuIoKYUiiSHwDjMCqr6Wl7QCnFWM7Qh+PChQ8N/Wx9uGY+RSJE3gt3
2MGTATt+dvOIQAJl4vhiinxNL+jzA12DR+Fr1EWsrtfqVgHnLYqWikMcw3/O/S5bNsWqIpPKno/w
NQMyhG4EdO2VHCQUIIfNA+hKWmlXsirDrVcRNeMujF1MhTcd99zyYZF++2pdfrTyH0ZiMh9QuuSn
+8480mlnIMJGPyIpt8O4exDA0NGtAZlJLnwxfo3g3sDE1aAAoVH1ypAC0WEOoTptiXLwWh0uwNRU
q03FA/znG90tlqO5LtVZCOfR7l4Ohx4110DwP0flqW2Sijn+SUt/ZSDQ1HgjQW1vv1VlzZOnlW1r
moib8dEhdNWlQLR14z5J/u/9hRiSWIs9Oo9Gj3h7pSNd5p+Aef2RMpRKaoYmEJCE/U9OwxiT9MxA
pXhqkiyZsQvDOtZlsWpbwugTqLSo48iX4nAhQyqggXfCTG89U7ck+6cfdpwc5Vv8WaddPXWi7Qoz
OhWVu/HWDpNl+8TVm6L3Zl/fw9nBn74TZXLUnto9akvepWtRZPhtJ3ZyLmKbdLcYPXQjHLI+xi1W
o/u2CMqt7U+wxmVBNYgFkysJZn0vMh5JT63NNI/4hOVzNu44iSYSzSwaeaDsQ+2DVn9/kYka4byT
v+SfNTyc+Am8uq/idKN/QWTKUeyUjgnDWyo0rU6SYB7Ru2269Hta/kopEejAsuj5TGIFKcpAQ4/w
kH2U93Lfx3EgGtr1OH/rOwTOnfYwaCxBWMnk7tP6tQQ/TZUPUzDEf0Cjo4pj1v5UEKRZrGhOkjCB
BMxCvArvtD+LRLCIvOarfvoz0ZT+CKgNL1kvwk1tiVGQ3hWyrgbYkuOE/puS4fg6xlapXqtivPpN
Z9FhRtOqNowWVYpMR/2EMcdmdwGaG21J0+JaWB8ssCUfIEcJ26Xe1N8zWMhX+ldOFvaDIa8JgVxW
+woi93ZCrlCOWzocGDKB/B2FquEaVGRopAYuwE/C8PHpEYvwQ+ac0s5j1z/II7DZ+PgEwZN29UZo
7UyRiEQDtMsYXz4IcH8nPb+rb8LBy6kK+VxPy7KYbou68knNh+ENNDp1Jyq4luIzczbsesBsNPUj
V31PD7vBlzg0jfAyNWfco4pUTkAGtlMts4B4jo3S5o8S3Z4l2rPvWshmFamVyRfU0eHlQNJiAt0n
rT42dJqofUCXuLfQ5T5lqIvxFq++9Fvl7w3c6pCE4YHM6E+4NCt9KBwGzrGl+veg/k9pxho/5INe
1K8gKo4zYu0rtGjMzdUMzcvkhcLxo3bGo54hSUTqWbrMeSZQKG6MvkS9SOhdYFZZV4bg5itcv1UF
EFkw0+VAfJyODceNSIWg4oXrH/tFBo4Z8LMVvI+2xArqKFhsry9qZu2Mpi6CNNz5N1zBUvzDFc5Z
5jAT6x8kojD+GFZArjbtTSvQ3RTjZ1JvnJ/AAsNmoTHN8spWShv1iKQ0a38Y9jdv0FcTxEUxPWlg
rwGc8WzLT1Hk9bl7KhKDlI9o4MDFT59MLLI7U4E8/3Ni+gho+adS21vMIFb4wWETt1r+GddwoiD1
fIzdHSoDmTzXKq3Ml1+LxTz27TkKYc+TsgRBAv6lM9L7IFLipdU10c8IWA7q/XNfueJCBPSZM+FW
DOdMQcwFeWuu8E9tAla/1ZzKE1f9wSI8QdtxtHFY12pW5pKONI/XeyVAMAjvpRP6OwP1M1ZxqYWo
LdGIP4mVHSo9qh3PnuPAGbAeh9hCvhIZPSD1lg7h9kW9egW9N+kz2mYPwG/jODJ4Zg6G0j9x4FvB
Q0bwjPet4I9BO/qB8YCqzNPnbi40QtTrvBlBfd6Kqss1zTSltMdFTtFVvgRsZTDA0cowGlKtJuL+
AuThDXLIL2LBmq7HexA1ydaCRKqc/icXl45dPc01Ocvw1hOM7JpEbGnCRNTXsIuoAhpuFQ7HHrZK
8c7+5TsO+zVzOZh1kEjWWSNBXghCphv8BzT0bf02rhjCkiYFG42zctjaCPVtldTj8jP2Ch1EepUd
qhagQ3upcVbnkF9RWHWGlkrPW6IynorWy6nFlsvljutLCyKoM33GTjPOPIlJN5/MKNwvZpOVVg3t
xmJv9k/FIGzLJwLr74FTwi13tRgD0TIT+9tjkMrVm8znSMIGTwwjTb2HNNQHX7xFJvu2lQoGL+vB
FwNApLiqyrgjfY3hfge/qbn+ABwnZ5OeMKBkUIfOGbHqAwPSBP9iXDHhWASUk7afOk6hCAxKbGJS
fn1CJdl75WzZb/YWIMtB++7kVTS44pfvGbxnBHmfAJrddD5RVbzel0Q0yymJ4Di4WHrVvoo/iO1t
fOZRU9Y4p8rw6lN0dbhHdrjgkOCScemaKwlrqh7NJe6ThzeyhADDZ0FkvGKKRc2aDpX374iuBuSH
SCIH3Iu6DAbDrjuCWREAF8C+Hz6xebTj2YauW44mS3CVzF6Ke8b7/AmzDUPQCNrVgHNzeSKC9pGD
csxHJ6hcqGgu6pN+JzpPYjvOpAg6ogjVhuGjOU1QbW2wA+YhI3u+PehHP5wzm8RXtenY2Sdc7twP
BKbGWAoo4wl1Gzt+fsrYAjLB/DupX0oW97OhWeqcI7g3JYDxrd3cbGuiHQ2SHMnHxDEXQ/3H5TSO
8YovOKhpUyIh9d1s9k62PU6j7i5CgffKTtENMh344NbbsTpx4U4KxccLF8FS55FH2LL5VqjG3YtF
rk45kuVV3pOjbFpZ0Qq+SgDaEYspjkAe7DrPKAQERl+pP/VVWsKOgmNKcq8X3+BIFtF1dJARDppa
2OJzShWtooB2iG9sBqsQE4D4CGovdd3hZA5g97sqFPSYX01HzWaYfm65c7yHoaeHkD9mpOd2LB4x
DR7FgylN2pnIiCu+C8VjZIZUbsZDg5nHZjapFIMY9sMpr7w+0NGN0nFTAR4HWmVSq3jtcubUQ1Nl
3Uu8I9ojDmpHiiHCVIPwW+ytNWo3y/82pCNMM1dNhRpZMyA1zJkihvgtX39l0C3Oig5PM07GTa5f
EzWtmPRY+RXS6nlAaYGUftiwzmdpDT/KVF/MUcyiiiBMuURzH1lBkdgM2JAcgqFBzSpfskfhQ53m
95DNSj6I+7ykpuo8N8r3IpFqHSCZnTshzrFaygMyt3jmhbdhTBaN+vfhe54chlH1mE2vmEap9/fd
BG7DNLtyTNtJPD0ttqD4MFdvEuNDtVcyMPNmn/SaIQKCLBcQRThQXwb930/aa8gpiob/mK4ZTNl6
VMk1Nj0PmhOTxpPQt8CzySL1reKGejbJrGdg3p5j8VrBIjNNv7A9mitCXwrKGTcn3+DvdgJuM6fV
IilYufrlvp+A7/PYCOXQv26d5BRqNaFAkMZMC/ihKVzTCzB115x/48ouhWByMBRCz8arcG2ENrv2
sNda7Qch2T/dPQXN4LzQqaMdyH1voNISGe7YQ8g+oci6amdE2srke3gxTBps/jv04QmU9g1saswp
Musk8hl016/wVdTFS5Xu/A9Ce9+EqJ1DkyEoxbkLzn5kCaVWwT+WBTZBzP4LtoJ9fIfeHm/54n5T
zGf2BNSOXF93UNWYmXPuWDYaFfgjO1eKSNhfH3kv2jWk9tVE/ahkTqFbPXho7/c0sMPQrhq3MRqo
neKQd1pJzLZAfyG/1Fke+5kfG41vABd0eJeru3SDHYYiVYtig/boWVUCxvb+B/7eQgAAr7cHRqfk
LxeESZA1LEV0r5ELOo6/6Kvv5ovay/SrLOY47yz4+uvKOcmSLVeb0rGCteBR1UL6LMvWyfZhS9iU
1tAzwUBB2vC8BNCnmL6VeZ4KrdT7TxGAxuN4U2OrCdlRj0xhNDKgaQuSVi5x9ILZtLy/bNP80sZQ
8R4JXCxr2rGhcFfFo4TOqfSDxULceGUotvAlm/iNXYyH5nA1481Wa/N2nSb7uthH1V2UW3wEkTKx
7T3t4Z1a7B5y/8ynADapMS4kzh8PJ2IT14R04mTrQ9CR7c5cD7Bn+ZRt1Oqn6FIlddDxjFYDWLoN
WglTa+KxOlXElMtrniHlvgPyFeY5W2KRJzFGbe2mxGU9bTUfkLZSrHDcNPX+nTxL+M83+2uJpjgp
s+2TzQnmlo0nsBj48mAbxFaLFOAsCxSjJHgDHqLEC0X3mQDl9Pg0jQRd7+NwEGDbHad8Eqh0rY5q
FsxdwR/RVztQzKt+SafpnfasRwIZAxidzdVnLBwDgvIqZeggns7oJz0KjVbHW54Y5i/KumhQYmQg
bykx1Klf3Dvy5qorKJevEVoRrh7zR52wXmds7Ia5NfVOlLCHFaITzRL8qS218sCefY8MQDVxwWgn
ZH5wTEZJ+Z8+k0PJrVRS1bMSRhba1qpIE3eqBxz0jMpRYAtgpU4iAjPaXldKP3VEWLG2qYdG5V5s
2N+bFFCYcKUSLjBo1rMRbaUDdMr8blNWQUkQwr1zYuLao4ffZOdOhmXFMkw+d+t+qfrz3U9oPlZS
G7EkKSnu5nqR3z15BO0Yj38WU6FHqCqs5M1CkN8yBBaBIbBXAhSPJyZ6dDHn513r4/2yP2vFdjI0
mZUdATPQR0DMGSDwFWyI4zYHdZTv41l7aFtUfrx8+BjUr727K96LbNL4Jj8XCQi1tBDZfzBZjJ9U
Ic76CUGAK2Z6cAmMl53PjuUfDEoviqn7cGunYfEwDkxBQEIGn/iYNkowNFqMRBNR/ddR0x5DXdHk
U1edMPF8JSpRRgPG8kcth85ktkTM7Nr0UywVoaS1wrHYp7MB6Zo9tQOA5VHpsq3NkUryGx1vcZCp
Z1wGTFdSUucHAuisjQqFfGV1NAojeLol/KyEkeY/JaUva9qicH/lE7fH3XMgDQPYBzjkg8SrrcAu
dx2Y8wmSVo2EJq7uZi3HYQ5IZCzPBFsKu1mwedDkWmIF/Mo3epGiBIP7cDbbpHUVXJQP3hLqFaop
IjwZAC2dTQokGEXlrGbutYZQrwo6kALV12awz+ATSb/KH7165iqcS4vgkmhshiTYZxPW6zY/NnGJ
AWkXFMDoryPwPDMWijD7Rw4HoFrtDz+1ZlT33ZTvRhGvoDIaaluSlWHahxnKD60F/S0lEUso4wcf
89ipTQFe73wmqvte12r9lGW38xy0Ud8343g5lpYPk9tDgDR4kX5KF/9zlVpRo62MjrEIrDB/weFs
yEUk5ubK2j0Hc/CSWQ4qwEiPqq7SdZRX0Akgylq9NdZK0R2GKjOucClWhKR53sm6c2/IEtUZfI/E
9rRROn5ZL8fREv9gWZNmX6IqbhDPTJL0xFAo6EUeYcyutrgbZ2REOJ0qiOZxMCUAPf0HJh8YexN6
53lw27aFW5XFMPmpjPrDsaGj6mJL2EH5RexRNb/zUilD9ul/Q5Mr+11hOnSzdmMtqk62IyED3lp9
xCMKT6WQe3uqIjShX9hn/W17m4z7wYI6JrmPXGSGWOcL3JKt81gbwKVA8xKgJdqabdmg+bXSTD0k
iAKJbYCCnZdtJWcgKo33P0uWkIxs/TB1dkDuQvMCnHc4o8cYrdToDBofVKyO3sTy68BA2plIY/Ug
L9dXzdvcp7zxb6V4sUxHl9xrkUUaeMbUVgcJY8dn5wqXsRj/mdciwkfzfoA8J2mG45OWP9A1nuhp
2MZvObQdbW3+1nmOTJcsAujsbFli1mdlh2xC2vrhjtGPC08ohsMGwaKG7HrfZl7ANJS0aFXg4nXY
03zDwXwLwBBxLltO9u9HvJ/DBcCkScvZnGufC4iSssD+93z30E3SyUB6zXXf9D+iluXp5O2sH06B
NBSXlpOfhCsqPUtoVAKs7GKZVWZs4RafupnVx5pNbI4yxVgLrcitwxWvRCaaJrieI1Js1M5ZkceA
zlUz2GtfmvNdFd8ZloR9nhFiXPO76ypQO0sh0HrP4x2Ave1RXoX1nLuU1e5hT3uMf/HeMYLffC75
+fRujZj6aA90/uzi2vGeHg0RAhaAlNSTE0jlexrvxBlweVwYoprPE8EoTVhzcht3bJcIkVE/kdWQ
vsMM6L9ICEu9PlEczMek8sZApwcVGHW7+qp6JkVzkORr8S8m/m5jYTswGqBVfgmiCb1T7l4OooV+
AQo+DuhM1PaxCA13UuWGOux+Rare5LJ5r0VlNqcJ0PCxDg5CP5QdIizjvx0rD92+6oitzynjLKA3
rCkYdtQxYseE7GE7ckZhiv+nARAq8UUWqLqtf7N40DZXaVVuuIoLYBNgKU2QrMzHwrYx/E1zbMuB
0Erep/WQUo1Is69xeLo/Qz3xT7yynf0ybKT/KIOO9H7ji16QMl2SfotxlV7zZ5/1lo1qdauwljcQ
YXyWlq5FtQf+XXuzvzLeRX9TKBvh/xYfYF5eGG5ff2r43+zssCCKA6YaAp7xDLbanm2434/4xk/c
v8DrOxDooLVkml0IJMznSbjlINvKR/ViOC4vhzC6dZWJgbvyfww9zzQVM7y0VGiB3+WvbiCl0w0M
L7CRbeWx9AB44hCbjTxo7/eFaYrIW2eLLKVIonZarKRdS++++LsD7Sh4uxGobDWMDiQlcGVah3+R
PDodcC5iyyFE0qx+SxbfhH5F70eHBhbb9aQUGeGlOdgTAElpZetvrrlOovHEgcmp16FpxPxUILJC
3nHGWKo2+BZPjWY4nyG02isNwB7KzgyYZTOgTCSMqkfjgJcFqM9NI1aVuKRpnhcG7IeqogIcGnAo
bf5hpYqI0dtf4G4Nqq4nPV/sWqWb8zPOz0u2YIwEJg5de+PhQ9H9m474EAd0pPNHDZhMHvjoorwW
A990SdmxaxnMKhgcsrSJmaBQMXYfGC8RqhKZ0XalazuYlig3nK9WiEiGoR2uVF9d72vSL3o4J27C
gmD1u37P/wLQQEg1uJmIrM2bMob1N8WJp5698Epvp7wjcVzdIp0tz58e9WN4sdhLGFAJUx/+E5Du
hGZdXAx/nJpaRLc9BM/nwCA9cApNYgl/t0dwzyVQvvBYYkfJqQOBj69MOLlTRLWyYA8JJJ0uIas1
7e3b4LOIYrxqfe5lO8MJcoDQGsYIXVYY6k4WKSnSqzlTQxRDDSglQFw0rLiPWOGJHpwzIhanoAqV
+PIsXdQD2jaCtktdMAWGp0NplaN5Egtl5RWc/Ep+T1a8gCOsdTQMTCHNJQE1+DDBWTzu1XmO5ZyF
LIamt+YTj8LFIfVedzlnswtsUyq/waPamhVlgEurCEGpB0ATip/xJnNQXrmioTNwznnEiu4MYceW
WhLwEP/ZUJHPH2E/INTE7SwEckjoYFdKJ40q203a3GYpXQQ/UG9xL5fBCetAkxwGQlWY3fDwql5y
cXGYR7FsxKXi7M8ISEBq5iXwZdynWH0FKCyH0se/K+tHNXE79vba/rA23PKEfceyu8Pfa7GZJK8C
y981JQnvxcLwVPhOW32WxWqQxDhOOShG4ZWMayxG7LHGkFFpCpNFhpUEQMjbV9vVlYLovjaN17eq
RqZ+4r/F+HRJPs16lFbTMx7kiIvxVRmKOo0VxHGxQH0ftKW/5aPx7UcMWjAWiM1mv+Q0UGOZL4Lz
+NBRG6DgkttToLSpdI8azQ5n+XabnqB1b1UcK3fbOTTj51S1WHIWDdczK4/veEcgYjUEV2BxL2vI
7ltvusw6tN4yo1uzGwJSWVwSOrpmLZdkFj5QflK35IQSj9lFSns+T+HCX912maIN3aF/5m6EHhDJ
g3Df9+bmg5E2wPPJguWGuwFoEbXa7qNAe0aaHC25S8IuPzp1DvcPAAUzlZAfDSWNQmXxpkypEnJ9
XRSWkaVoRiC+9htrbww3p/sx0jIkQDP+CRRakSiIwa9T4IY+DI+pv6WMDdAl3o5sqa5YV9D3w/CH
qX+LXOKLwKam0lti0KWng1XqJA8cK8lgWjRfDdlpqL/fG/r8yOrR8bfyseOtdjfiIfbsn4z7nmS0
8UkgUAiifdNm2TqPMedSCnWHub77PFwCTApHm5yQdzCpsgDrrOJh0i7StNVlVHnEmZ/GwAckZ5k6
oU0/6gkJNNqPGqrpFa7XJFyw58sBeQ2BWEdXvNtV8ZZCifLqELAdg4VAp5mGr07D6YtuK9BgP6yo
NECq2OBB22zS0NU3mPA3Zw18tCU1/JBA0klS0NExxhy8fBol8tCSUwVyAgpwjJpWR0q9Xpwk+vEP
eAGK3/GP422WkSrKSneGZ7yKcPfYmWYqOk4n/f0aaws3kRNSg8jpBzxoRS+1gXZBNpUKQ2FOtXn3
6T17h5DhI6APZbBXyVH3NN0Bx5nrHG2JjSOimGh9bpQkoa4AqggZdDgs9NvlN/IEzMUL5LZbyIAM
9wMUg+ueOWY5cmCoayJ+CODXgdoWcB2LA9flW8n+lvsOM9tBlYKNThdwVPQQ0TJLwpTo634EHv/f
8JmPZLs30plpYcqP2S+Tg9L6yvMCk2Ldc2JwUhwu7btLul/pM2bdN8t5Df1B61bY9ezOBqRBknm1
KdGi3JsTb73h15l03PrAwXJkRxNzBxm0YsZaPoTGVNbLf6cbnhYhOM6GikVeZXhL3FHV1+pa9OLZ
+o41a6TO5Lt1nBDh30fikYUGRjHifqGunqs6/g+73BFmKgICYFjIG90rSZCgGH7+3Xt+cGSCngIx
MdsxbZSv7/N+9ZTbOlqiqtpFHBW597p/Lrer1T3DzvhdoSouRErRkpXF+PIp4GGFK+xyt+LfIUPM
1GcaVykw8dhzVS+HIfhnnKQrbbMSMYUdLiIRs0jAXOIiA7I3h6sYH0pJlV9wr/UstX3EXDtYqX+I
BpD/CWZtfcMAihAWv6xclj8VUKJE7PSeYQFpS8sZk7SMtataciGgppo2Vv3sxiHHcXIUfsNWcm1i
50VifqoF7Y5jbEvnW3g6S6L9FChsM8/uywR5FbxFf4ZXNnYX9vMoSpuL3siAU/UXh0MvHHaj1bMj
GBa6nC8HjfeIvSDhB3gGMTbEaE8o1sNmNHt2dA6w2voa/0Av28rbOXb0S983tzVKy4bdzoqotGdr
+/+L2ExyvZte5WldttI6BCYWGJL6IciKJ76cpKzhtfbRa2iE+KkzWsgwpfp0ILHlUTpm0FxpZJG2
LBSgiafx2dYOPh1M9vBscPYAr8jPe7fOCRfWf6af81qkqkyjLEA33laJobBqW1m9gFN2Vrioxs/4
lJjXt6OdGespx9A7788QXW2f1K7JkJiGvu7NJinCeWr5ygO7Att9eqkUF4fHflJX/ntHmi1GiZ7N
cfh/9KSokyXIsFla8fjGvCaoVpNpYHv4B0szo2eADSJzVQWUhOCw8a6n2L/8xRakDUyKDGq4HSMb
IVUcMG6yDMFSMrMzRXLyEx1sGlDDHjl0x0sWmm0uPHF3RgqlQt1bPm42/Q0G9F1jZYJtrDS8wq3X
SAXwn+rXO8koW5hiOROXQIEynZzgRyEXT1Uv5RzxLc/9FyJV45AOzoGoPJ16WBSWpZXBugFIP68z
TaZSdSA2fgp4+kGsAMNYPt2tyMc6CdRJOv1WgLDZxBr3b1ui0++qSWsqp1tnAmCCFSVAFwrkg7f+
S47kKL+cuYrQhsynuHfMSRgTD96KYYFFtgLaooBlPIQI2cIX0kzXJ6pjYBhytkpmVMSAIJ67vdMx
OGoyzc2wULgle4ik0veBL44IRt74cz94lKVzVH59kiYO6YAQIDcAVvxx72rFS8Z7DMYPhNSedd5J
/xaPZ5QK6KSPP9xgmuVIzGNBEwItyHwZgbJZOx1P7+IhewnulYFljyFhYRv7PKGNxSUd2uWxC7OH
xrCfwtwJbg77ZNyo2PXE0bBnEitDGITh7vIeqJRJmY8vxXbjstH7qw4geK2javwmV7E4OctxhbqS
uNQbVJVIImM6PvfE56Vi7beHod939uvHrWxJlvjgMLe5i8JhIJRydN4IioDnLvz76nzjSYm1d1of
uGSvs3hwilbXqjjK3pvFWW4Df9yHwXhzHNDAQ9Nr/uzGoqEtthxt2Bu1UfujAguinkHui1KA2Tpn
bm4b3VvqjKmbcj6vYqQhyPfrDQpRmfrQ8vJ+NTKlKmlm8+uoXbDh9lTual16UWvM9vbfM2yjquPH
c9cedvCYquEbz38orPxYfoSPRcSbVzNVAQAxWnPc+AxTlvgjtehqvOMIlIMpUhM9mcREq9Dgdh5a
B+eG6D87ImALWWk6gjKa5IfjVtFiQEu0Y+ecQME45+6+QI62EbbA1AndnPcd/EY2onR0FF+qcrVc
n+SmzE7pGlQ2k/esZAqGwKRd8s9YdpjGqgLPbcNlVHmHwr+myrZGVeyI5qggXNkkc24pHT1Dd4N4
1ues8M48H3HnA/qE2fWyKPUYW7MloLri8QXO158iUNYMau4OBu7IkvtAbEqkQ2Xru8QzvvA1adaL
JygUboTcReFNFWikwZXHzXXWFT+yWlCDFc8XN8R+PWaXHG49SFou2Tdc0hQw6UcLIMDeHHwPsgh0
GiuoYo9hUrSc8zf/VwFEbd/xubgJ1+5UdhY3Bh1SOAq2fasshYqNfavio2TB7F5QdQcjy6LxO9RW
FdVq2diI3J4wjsxfdWncFGnbYU99wudXoQsOjm+EydwhBzI6lHXK8uvbaDG/z5dKR/Dr2tqcCG3F
o4ZZau7KLN0htoh5+NJC00M/zNZgoMuuP75qMRUwG9NJKdzgqgnDLBfB6H7fg5C25F45i8pdj2fv
WTUpKfiB1+UD/h4ZmvQY2Pn8sX0iJAWYKgUT3ue1r/Dytv+WwtRNwjs9lD6RNCAkVBr6xC+vUNiH
vEFDDU3TgAdjgdCuoOJHJ+ArNgLBYJ18CSRNV7EXEBMbp4gAxvyvODDK0pRjmwUsUw1VVjxJVMJO
uHa8ACE4LYgjNNVd8AH9ZfJUJrvFvB8ON1sI7gIq5GX4dHo4FyIBYaDaR0InDsQpy9q9smC6/dnG
Xdz6/OCD0KRG5pv3FD8O+boJUdASA083y1wbplOMz/EobOvJDPOPHTghatSO3lTp5Yg1hFLT/Gkt
MrtXMZI231BnyuvgiNKqLSKrXvJmrAzwNRgo+l+cnfmYd5iYSC6MMkGAvqk4FML0nYOY6AVNdeql
NDuN7vLFIgG3XIdnQvt+JntTRvafAJGjSbPjy5l1k3mSy4mZZln4NNk4n6nd76rRKLeZFTJM8dMA
BSe5Bf8HiQ4wMvIhorf/84CviTgsjolOUJrXIjt+noa/+PWQcIIr4Fiy/pU67DmzSf1Y5LR+hjIj
ChMfGBJZrb+fjzcRxbUIFsuffcfsrniJpnJWFlw+/MTBM3Ymm8IvlfOMmMyD746aT9ioVfft1Leb
KBFbPOU29L/dQ3P4IvCObK1TaHgf1wE6kVb1F7tEnzQk6J3OgyV/l2nI2j/5orLGPvOcGKv7bC/D
8nIET4HwAsEYkmKTCZR/mDiKf53zmuNiKgfH44pdOp0Hw1K/G8J6kqOqSHCkKDnq8hgFIqap8v3K
Ofeg/Q02bMz451eta5qUOtEEr19IxeEEkYEmO0uue4W9OPItF51u7c2YM+R82QbqO5mEtIErU4IL
vB0g5tzCSa9NjKzlj/RoC8nLypJR2doGf8t9yZHFvjD5v/Lu8IYntByv+VF3rmzqnE//aHs6c7Rn
Do/xaalzhfEKkdP+hu/xF4K2xpN4PS4qrnPSLfSLl5GOB0K1pIcQ2yDkfJ18689IF6/Qc2kOhGyI
HITua6rLOwxyTnzkNWLOGCHZEYocIm2DH/0Mgpz4gtT/hVlrtFI0F2I375DbjOsUmKr3W5gO7itQ
WeEQA6fEcnojju3xkFAu/BOALmoK7dybwzNP1VR+bjVreV8dzu3zTT62d7/7GfRpCzsAsunsQ1Ku
dR1ZU4Lq+48ApbtNcZxFmt+g/RqFHuLDByLDdRfw+Ac7YNuW8XUMyAy7iAzwaOw0GNmMa1eoPB+Q
lHS7d2tPKiezyaQ6+0YP1zzl3IWFn85uT62MMx6vzjC2QyZ5+0BYITzfoagAPkTinD5WN+T2buam
bnKwA339txYkKO0GQb9wilgs7cPrqmV+etAfReKXZ8oo1olPZYz0PSOkAD7f5+6vlzaaWcuhjA9t
NoPw7meh69CasVL7XgNPq5t6SzR8KZ7vzi0slqMTo6Y9Ve6UXipTU0oJh19hL1Syhuxk+zQZFu9o
e0WwDBc4DRwEEGDIylqtTwCIXZaByqOaBk9/s1OttdtDsg//H0/u+vW8RxBid/R5WPU66mNw0xRM
06RmKOlOHDX5kA0UI6IuEwzgyMjKxB5iJU6uKBFYZOIqU6eKc/oYxxPlx7VK2RrQgn/RyojDxA2/
Eg3JKI39AN61pfLhCT89ZxVAlrflGzWnZJhe7pJ9B4+gfvIwOSv7YmHK999W6S7WYMGQ2AofOwO6
gLuFr7F8tncpOWuOhfwzUE/+e/gDWXKeYQ4g4/axD7kAUZ5XdQmVhtbp2OE93q/NLviXEvbzYzzC
qOP2EhgCcuj8Arf7F2NOm9csOoHfsTzXpxdwtLuACX38yfBGFOzlTx2re0VTSAiS4/iT+mMpoBJS
F/f9Amb4Bj8x+MharMFQZwfw2HW3JENYhBFHGpHKG8EPfLXERknuxMzHuG9pUrJhZaNKbMqZcuw7
rkLnT9RMAz37WJF8hP8Nz/AR4e4V8yGK3u+aXACfMFaDRS4thzqtz9h2a16eRL8ZtKdX7UJzKxJC
ApLVQyF74UytD9gDeGHTn1gfkh/byVmyh2oCOcK56eGqkVXR+CkNdRfD/kSsTyBI2+mRAkfAu42S
4XQUedB+GNoaF49nzR/x9bgpVYbsZz7IzXa5TMyX+sawCi8f/zAfyOIaUXsB8ZWy+7N6BN3012KK
XBp0Eg6m3Md56TF2TKlaX0qftOBwRWno5UR9ZV6/z95xACmzJeKNmoksyjAiko/UiqWghOPOGqJX
wt3sk+Uex1rHtwBoh0dTAA8CaMRY0p5htxVNXvNFBmICYmfEqytj58Jwp9uKBJNQb8RbHvQ3Rwss
23qF4ufH2kQD7BWH6M/OLlTJI5bsMUyNQmrcA5cFk5EF6RfRiD0TvaknLHrqUdSxqrqJ8R5CDXz+
m/VFvIZPco6mmPD8ZJ0+vv9yXAmAOzpYHdruJhzVyG4vhclQGC8qb5KWVwtmnd8mxkRSMNWoBBXZ
CwFpnvD/5AEjraCfW6i6bnZWBzVktT6d7IAQKEJ+Wvgj2AXEluigUe1OtxrmdnpDMWzp1VefPslx
8gnd+eEZdgBNLfWsumrNCkeEvsZ2ZqaYaiAff8Gowog08qC9FlD5xLHD5WG1dETsnytyOQAsktcL
2Clqk2hsMiPDVrU4i23klS2kgviQ3XSKud8ZYSCYO0Xf4stQf3bIic/VenNK5wui5yiJXqYi5Ljr
5N3QE2pTRB+VchoE0cnlDq6GXvwBjHEbAQsMpSb8hUnc/ur8bfdoEUv68ZD56aK+R3ttkxBpo/WZ
gWMLY1xB/BcD6e5jebo3qIfOGoofwx8aDSW7l7sVKaFRJklTZ7btEbtCM0l8ztLrB734IRRQYMvD
F1c3FMHv4+6++witwegKgjJKEFJdgbdrxSXXZ3gjy3P28T/AgV1VBmOBsatHVtKtYi9EAJF0i8VQ
4o6FfzjG9L6vrJAjru0dZtLTpAaSyZdBuGXT5Jp6LbEsbpuhjUQQR2kyjJIEg/wOlSbxRxLN3b+5
x5HQPYTO6r78LmFxr8P3xfH148TX9etjmVfLu/g3v3x5YOOjPFQNqUzMU8wunRf0wa6YIGsD7Kq1
i+9w659AhvJ4YpGzaIYa50elrW+FcbH9AJ0pygdR+G/NXjKYVDAIq/n0HGe1jkIHaKETSlWq6TWc
0RLrd7BxYHGo3nN9ZpP/Qlh3ZEVwrJhGBXFE8LFHjBI8+inoRooxHXjT5ELPVT2WUwWxgW3XXU6e
ULeqRQj9+4WFSNIpPul7mVH+cRNGk3O9QhPfeYQ72EJaxAnWna93i92fPCf++HyFk0T5QkRfVtSW
ZjNu2cSKfzhdL1JNe4tWsB4rcyxTiXvDknAUAiLxxpmNUD3rwRPQkM/UxIPObk4LwCCCTuBKfa+J
V6CLf0L0vj3Zv/BV4iXkj7I3ZsRRxX7MbKfx7N5tSc25kZ1MkKnWSK7cFOscnrSm+A0VpzM+UNxc
sxZSejwPgM0cs296F0/k8qYQrHU9pzTKErB+x75te6jeauytCtlndxXApgSiWM1xphM6F1+F+0fB
3TTKGQuV5d5jm2A91e9dh+qpcvjmID09z9lciIZOox2O3QxlpVFAxCnRlx+lw9FHUTPOfjc/zE6g
fsT7hMLpyVvL6mZYE92VGmbp2BnqzZTKvgGWx2b23WgHleOYA7NiwYzZ+4Z4G0KJx6zIFC2va4SO
A3xdtdSwvDBnpCluVf6LfebJ8D+pioTK0OYigmPJvFg/YqiKTLZAtfCW7SgHK0kNs42MiHJsjhUg
xSIcrd9QHgvqjbQpXuXnuHMLd1EtQGoR3TuDdBuLXt2kODu3T6kQ/6ciAMg4r8yuivoneunZRHp7
Ut+OIbHwxU//qct4rsp3Skq5/I1wZIUpkoA0GAMUAfH3+QNMBSLnmL83crMgCUi6OBwxGyqhzsvz
5/GXO4kqop4Jb0df0Pojvr19nXaPcHN/qE1qxClUdPNw12OBtNl//kBaMLaxoW5T4cATVOQFwCpQ
p8XwC/skOYMwU0EM+FQiJPo3VvoULJ0r6lGw7xNLU5tanpEuGhFcl3KZogD5LwCfpvnVyzdS+Eor
oFD9gdEi2+de+lUbe4/DCF2E1UaaIrpmC+OBN0NynRSxB4jI7Cwd4HujZddccQXBHUKOhlAShWAO
PrxFmrdvNISVPJaDiH5B+MEXiGbQBkbxhMyKviyKesSP8Sbh2gjt1u9ExHv1OzryLVo7q7l86YK8
WHskzYeUzwQTGXWLhLnwWhQVcOakAAULyc+YhqTY9ADnGMlgQ0cvH6f5c4reuwuUQXyD7dTU/NPc
OWhU37gUFKZtAtd7MLCb/WX1PKUFtyhz51RUyV/lSSD4tHYi86Hzl6c6EEhyvUAHZDTDY3mDwEYT
81/jQWrngVKgw22/DjdujMMf0alYvxxipwWMUOFctnGACdkzV7wWlUnGNC7lOoEtEde/EDXjFaGX
UqE8UXk9ERyoOP/A0mVATK3XNL9E+lxq0rUMeLbgr1a0/hICA20uPAFGFaVILbG8lnYmu3rpJzN8
xyFH6H3rzk+cDjYyZ/ZSopNCXlW1u87umGaFRLX+Cs/UmzOt+GJvrw1EPwtsgXS/1IciJWMd+Vt4
EW2uNeenC5HbeBBztQiw6BhxBM8E4cTTLXXY7NmTO+G9wLVAKK7Hy0WYUwlzrIlOULawVdK1xCWi
SrITVkwtd0WULBn87FZb7UAyln3fVZMAnXW9spqXd9hkEI1QXNNLGi/OiV/Mg4r8vhq4JXCuw7yr
BhCFu34ovQ6oFOAmr6h2DvHiAVz9LBQWdQM3mXWTlV/kmju2Lmds+pzLbzhcdxBTSpO28NkDKVkz
J+z0s9WBcJKS8ZsuxuAXkXwUzKr0UuoXipOLsE95FdGzLAET8nlyWJAbcs5SRA2zjpypFV9G2XV1
P8Q7jkLh4EgH2IWKpEeasI/LrHfjlZSpSfQE/Kcv9PGFMcHN37q+dqXl1EjMOgEqULeqsaIC0X06
/ZJnl9Fw/pjmgIlYPJOvrSSJVihNCM1eGfhjPGZF3S9T/pAO3KbRqyGryeuUStPO+pfF2vh/DVPf
741tA8/O/W9mXRM7yqpEjNctOnk/92np4aAkilvSlXimi2tDIR+HDFmkW+IXiKy/+xpIe+DPnfTI
Vnnyl9EGheaZLentw2DTha7WTaVV+Q7bFbeIeeFdsV623/uBSZT5ONRp7lzs33iZBgQTZlf9L6oY
RjmIuQAglgSe73LeVu/lbSvcMhQ50OlYbQI+VKheUbqt7U7vCKZh8XOB51nP6BsS2vFYLY1YiD5V
KAjmhK6eEAi9qixWY3t1eQuEHIdMSWtvMGV5tiNcTf01l5Nd5zvJVhy6xeIpqEWinalXDjVlu2MV
6VS1iyaAZ92zZ/GjQk3H6f6nADtpdXFNVc2nPgcEbdzFqfcpWtfjzSHUZumTfT1K4KONta9+K441
ObGDZK8+nTzqv1BGxAVDhLx2gaOgr4SO+5FCO7MuG6E0g0Sydio+jjgmW+x66QxgGATG05CX9mC0
Qjpr7ZphiAB7JABpeYCIMEBHA2OLfNRr+uUEitXgbhYkXLb0DjIjQUkdwSHXWus787nDmnqCCYPb
gjkTmXv1JYly3SUGYM6H4XYlVnD4e69lEVN6jogbQE5txKo7U+oyBauGOd2WWgGsLKc2w6Vo7eC7
JzKIj/yvphrc9KRXIu4v72JMY7XxKpk6AWpToO6jzNfgfkgR1EtaEqLXnMzSo+dtwd2P5zpRE3Fp
REnpr43dghINInogY6uarGZbAZ3fFDYsqt1hILv8Wv2oSMPTnYHdMt7cz75oo1dlwM5vLQBsrSp9
Z8/F3EmV4kIKvHkOCXTxf/epffb9+iOt9M25n7i6WD6wQO1jg+eT0bTK0LlvLOHCcyz9c90POFwt
3UL0VF7C77kY0EKeFe7w8zpTQ5sVSv1BGD2MdGpnX0Unc0NO7fX2VgCR6AsKbN9VZa+coeeRJ9Xe
9/Ubzczaf8oGjNHxQvwNj2u9unh2WC9CZYqMHxKQHF9vbg+17MujPztEKGMXEn3VrX0dxhck4d3c
Gsfiz7rYPLPLOgatWMiy49CHoRVevBy/DK27357YDHVgB3eWsJPyiVYB9PWnOCITIjuOsWBX5r71
pMmkC9W5iLVentBxfd2BRYntJ4kcDspSBynzCRA30vfpZSRgM++zbev1gEOIx1RwFiJ+pL+ChjfV
koMzoIeBP4HCHMKPFcMsZxxggKegxMI2M70XMcWB08/lLHbWPUZICVSth5vn6lFnR8RJutMOAqF6
Fq5ti9uk2FoXZABHs0D0l/rfx8gumvbMPZU7Hc0gvdU0+L762HZN1/1iZWu+X7CcCOO/ZW4dxAwD
9Nlg/o2WBRCAlkFV3NQvybob6iVxjkBBxVUopSy+0ycpcUeir19ziX05ueU+mj6ZQdBQAWWuiewY
5tAGNK+nrIhgKXygwwfL7d0hw+IAgrdxlvWx65C8bsRfhspY6DC/pj1L0lWZYlGXWGaU+C6KEnxw
rzAD/zG/a9GWC633dm8YPAYhy7Dn7RKOKIREu9dGkbCdACxiHz94QYBoRmFFI/teXLZmV7RdqyDy
XMWLXDvmCJko5Rm1wJuNkK9hGzqAHskkDqobZt0fHtWLh52qMYVSYWIQnhskqu3DxgD8uYCQFG/T
q/QeIrsOf5jC1pX+2jRVfJm0Fd5j3BfdlqBNzqLmffQpkd3vspPQFVJ/BQ8hLpmt2kv7g8FaLwl3
D7KHRiSvLcKe4qZ1poO/6nraUzSbVlP6ZNgXIBql8gFB/2c7Mu6vifoEd/Sr7O4djt1GugJvDeRI
aWYLpZnHftctV0mKKWx3fD073LxnqE2fZaq/NEB4NtPS3Mm0xGvK+KwCuV3e8Wi42tmDaYVCg+ZQ
Z0I/FEAGTUOp2PhHhQ51DQLI7KuW2HUydF9qA048gNJUxqnwPI3ZD3uPBT64wbyGZ1oACN/O+MBk
tOe+BwGS1G1hGdDdGv1+OUP6Zq21moOqcBdfg083P16uQZHBChEQJpiGrOO+bjMZjaN7ZGxwUDSI
Q84AZG+xLj8WmJh4cR47cSeY+oATECCW9ODbhBBQG+KsOi/Ogp1VaPDL0E1lS1xmltAJ1n7QZ4hx
F1KdIYAtJ4qGGVSSH+OwYPnZD9OsfT/lKSL48aUaFGR7ip0D2hmdg7UBUmzN1jZBOrb9iyJ95HHw
CbUYtCE8ChAKuCPHNDrOMHAKGoHalwKQlZz+iewpeL/79Vo4oxexJVcBhVKp7Fn2o4LosyeXt/8l
CY7V6Y6Qnw75M/EWYCUrJ7MSLWJf7S3cjkCBhlrU7fy+NIpbrmp7SJsuho9zjC+q0F3WJFhsmqDm
um8aldJ/hRj0KXq7Aivkhw/335pLEgwstIKN8Krlgc8IHdzYzt+XELlbwXzqBe8BICZKUGAw2NOe
waYdp27Lo2wSNYCva0bDQbeuincBHeQxLd1iPRcCEWft9pWZzDtBGFr70M6N1K68EVtMTxi8qPxU
8rKjLIBLREBmuyFpBifvLDskDWCuUrrXvEvf4ZHXzZ8TIxpUjYVabMuR50YRU1si7LxBHGicjY7R
aud5m5Cphy4VvgjcwowHgKrDVILbEMjm4/WC1Jo7J7JqL2Y26hrpEL63Yk7DJi4lW3eMPlFkwuOp
cqBTa6VDyy162Jf62cIyOOjh+v0o/LOKYrjHq+8Rw/tKdLHgR+YH0heCrhTZUgkkpD+Qa2k4Z1QX
LwXFR71E6KPZMUQROZVA4ULbpTV1zEmJDSZFL+36J2e0K6MmAhCTMviFIkTm2mx4p/AhFekD+QzD
Visu7vlkq4IdK7LTjVxVVkFjuCj60ScQdtmfpBaXPge7o+b8uTtlNeFsiykVwI9ob5gpROiwt5vV
X++dbaR/Zl8Yo3+ivRN2j21byoN1LqB7wLJRWllkUqQaP/p2mQIC0+Je46Zoa/Yh8G3f8ux4MCwL
mdQUEJ4mSCq5YTmEBoaUpFxEPdLzv7eMlAlh0XWB8F7ex2o8/MawfFvqzk6OHWoi6SPJ23HRYtR7
67ql2H4kWa2VWZufWFZNuqYjLb9fKOqA8s5oI/ZRjCNIGqaQtIclI8wK8ofUUY0jl6dtxuj/sYgR
SHYFbV1oxmmre7+fqXYJGb3EMDoWxIGBuY840p3bYfJ0v0yqJIloQ0fYh/7ZkRXPDqLTEoDgjVK2
QKs5FGf+HzzNFQFEQT0Y8kqMBNRjsTmwgOEqgif6sFvsB9n2URLjaTTLOw1vIGdwFyi3LL65/StK
5YhOpdbKKQmhXjTXQwNFLuTgaXf/gPwuOddJyFOnWyP8l05KXUUn09nga5VoSTYh56vnJuscMmiq
lxo2EIw3+nLq9Otmw1rkZEBbRjF5tTrfK6hQvt/ZUOfeCheXouToXlUev+S8O7wb5eotsDEWaqLo
lYKothpuxHLV2MiYUJIoyw0b6fb7Z+YtxheiyebcR0nxGoPcyNP9+jTTg9OpMJd2JI7Sj5E7qLxP
mTJxjWsCwg8NSOg1xovwh/wG2nZtWPWsb+l5onxiIib6ghTXKwjA2QEs8ijrwgYqwa8WC2sWviVl
OqETAmXunxxxJ9LwgT0DhKI+DZez/KS9dlpkcfO3+Kw4TkLQCoGGYKtDhmgn2W6OdZgIIZg/mRPE
m2ktrmrBOd6dBjgr9bqNLHyHO17/7t5p1ofj35gkO7KaLykFaPB8F1ehYsprh/yrpsPqmZWS4yUF
T3ddbJBjoRvIRK+4g+ptdnTE9Lx1OhXnwhk88a0AFehUGgRQbkoeFGMhy0YD/DMYBzQXEug/tvSR
r+XJsv5YjwM1jK96XEZIapP86gXqRpUmoLFxSfk1wyzQaOxvoQ3W9Elv1qcHdI78MxcEsgKyIJnG
4qoGzjEKIi48MPcHpPI01xw7KsBEPjqXI7TGsnUCRPLIjGZQqtgRK+NKGsTa27TRcAQ/o75/duT8
R7ZSbmzPdo81MoSsr3MC+C0YKwtI5S0LzNyES2XE/R8fm7zhUOh0q1vTb62+v22m6fcpW66kXwUX
Np65bRDxgsBGdDKvrDnECWcNpwhzb2Afge7tw/s3iT62QrTiG+ooqSmj78wBO9QSjdlsi+UNknUE
aax3q+cICk+vCpH0PsnxB9FbM1m3u6b6VKkMAE/JzfF7twhhlFcbSo4rM9kqKVAi2grdZqY3xxfg
XsWzAz+ulQCKwLK8TFc5hiB3gEZaUN2mNHBsIWJ8m3hHPH2KGgJFKhCNTxZQxFpWEfFgNy7vZkMX
h0Hk+LYUpOgq8rXHeiiS7WY8thQ8i4A4qm7ILewuEaPvQgH5oBYoX9cBFttsXB3ljmWuPF3Z9ERZ
gHSJVNokJlReK7GiiP7j4VAKJMmiSGZ/Uu+Qa02h/bgoVCOr2cfQx3LyfhV3kkRHXCywaDgV3g7f
i8KlnKCWkxS5bgvBgIv2ApKRDU5GvxEAUhRhtfOXR36h1pHDZGmUC2FODPA1ytEf6DA/q0UmiIg8
FWC5IUednGFgR6jVwzqJIpKj+T/CtA/0zlnYsuQNXMdlp2p2FZk8hJKCH89d4fnbeclkq+SMTpnU
HKEJhYWf8PicRfIqI9uozxmh6koO80SfdWOUQ405BWOYTZDGlWe8U6zngRvHFQeAz/K4uxRkrfl4
ERFTQD+zxdSrnm9/xT6h7ae7gsjkfqVvGBFqtYLx4oOZ1te1B6jKHHet2GVN9/htfS9ksEvmavgP
VbAqK4PtqAQoP8vwF6uC6PvOzOqAbVhZkgdjGFB34v3pWtbj2nRJtFDDeB7XP/CWDeDkTcEGuIDx
VYriO3nRL3EAp2QZCJhtm5oXmtOWpSDpzTP9ejfUN3sEdEZb8IiCFnQpT4BhOgCEL9+WoB3FYSdm
j4R/xR/UDkD1/EItoYaT9QdsoOXFji+KQAl3g7OWHbktA5PtXTgU2+51IOz+ZRNN2iDJLNoKjlIV
Md6ryELWUwbnZfwkKdFc9FEy5xVTnKfle7HCLcVb80sQO+bNFv12rV7JFX0mtcWStO4YIu8s8M8r
QV7T4yOD9efATFDwBe5q7vfB+zFydpkY3tT78oE3S6zMaxw2dQQnGYYNBSI+cpg7DT/O/e3yRuR2
elSas94BtGjQMmavziVcjhBViLpSA35z+ftKnllKMCw2vKc649k05H/PTPtJS1GaUrD8J2wZjVrB
NxtuhEz3XxEHVPHEUhrMUU+wNzXnMgCJh7kcUYw+Ga+jxqXlqxACiAeS722cSTVm01Tp1HcKyAAD
6xofT1EFBc+LhUv2xRFNZGgbvCCl4EdZevJGopPF6P7Y6YpNLorPUGd92FY4UjB27JuOTesk6cX6
CSLIJbcR6KqEFFHQmp5gw8RN+E8Ib2wfjRo4X+uf9SeTEMPogQlMesUN+kiRL3o6ibtO5CJMg8SD
p9xFIWgBPhYp2tWzGIMrDgInf7WSWYwMCJwHpR7+UgN63zD+PfYrThMbFoWUaUp68hfbE9ALEpTz
huF3w+n6Xcwx2BQARvEsIh6YsMmgvhmvGjA2fpZfKftM3x9gS41TL2Gehneh7RhB/4uWhecKxg9C
kxvTmMCZqeyYgA7yaurmMVH1OwAtbUGw4nNl5PWWVrdXzWxILlYqt/wqTay/iIZ0KFD7MJMKMgp0
8sS7AjZJPaE8TB8ih80xh1BDyeD448qZfspDmdgVAj5ySg81WJOhbvoLlweUHnBW0e6R3mIhTjJg
cpzeePTnuNg0ICzuRKhvKpjefyjzclt5kVsc25tG7oAXaWDynzzEpl6h7gPS9CGD2pCZUXoCgg1v
5IPPn5uUJfjn67XKSaPsvbKXEBDzpOBk1+VfUPXD51JRKNfzINXxB00Dz5fvsjPr9NiRcixPJYL4
zz+aDeNS3TjlV/sV/fdeRUGFMNYmqYFAFlTpjn8m6NQHjvFefAVswj9ii+K7Jma5wJiCd9U6v5xj
r0/TsmnrSn6XXrnjFTXcALofG1mavLVbpJ6GKvKVZIoMXrOnWIbbzXuvgY10HGW6lmJJQfURabl/
jG5pvVR+Em8FuKtoToBhixfDF9LVQDWJ5O26TnGP/qYmuwu71uDlcX+xQZXfKcpz/1w4LgbcEmTn
WG113WOeN9tkaTOWyP/YNQi33ohi4koFTrwheSRutrE5le+/7z50JNJy4s3BO+fOD7Oz0pPeDDM+
Yt7tF6NQB1MwwfQ1tEfRH0bsLYuu8BYpmwraEQgGVkXSGhVXhYhnqHTuP1ksbM5N6XAoMYtABfou
vjozcEIgmitlb68Zj22QsZ1Xbn8HDv6l+gN49LR7AwSQe7aKYqj82cmseOolgBOfQHnhgzDx3wnw
Jn9nPnD+Jq9EAL5ur6i84ov/+EisIwewgrJZApbvYyAXWnGdUoVUlbzgM3kfGgbR/Xeepz0+QIYA
31GJss0PqvOeP4uJlQ/8uVl4lp4Q6y3O+TP9DiG2hB7lgt+8T76EsU8CDR1yd5ZToNCEbssxVRrH
FYSwH3RcymWkNHHZlnwjMZdd+EWHHA/S5RVxc+xOhUbRduucKQq2+b/ZWNRH6JQv4Ick1FvaqddF
WcGIiTB4Czu53sjLtlTbbwQs0BJUDqAn2RLTzIQj999KFQpkUMdl0msUV+ZT//U+3/ha6ml2IHKS
zjBR9Wj8V2QsJF/h/DPypQto7mSeyZm/BmIrcNkvG7LnyHpFzHY6jeQZAapYx2tH19f2LPrVvnWR
OLsnqke2X/Mz568/NpkEeJrlVeisrZdvTojS+cbDJIAfDHoAnh/9BbIEg5wp7jQ8FQwW02LHwqZr
sC+Igpb5bR0NstAENrPn8QT5qqyG2zxSmfqGeO8yChsR5LwCArGiTVhx7i4UumQ3fu3ALyVbxdKY
UyF1SEr3JvxBDsY2bwzn0N9UGv8PtZF+ev1c7zy8H4JrAkuaYdWuMcUbXr+w7LU5JJ5TqnIm3mHe
yerLm7u6v/QDr3hQGr2icDD1udV7w1mxiPpkX9pSjZDGrl07+L6qySboNaSvdrSc0glisLAnleBv
2SAMNtUOVJxhdTD+hQKDs9kExicPypCI10RofsvuZkpkT660jepl6W1Cwbq8/JIbzqc3mkiW1hat
lQO8d1AYqJQJx4AljuKLre87X3hAVkF5m4DEUvPkntEn4tLvTfYcXznUxcmnxp9MbyQWCP+h0HFL
/WGROOR4d8QMl/lv12PrwkLnN4s82G7fmzM4Fj49NTxdx3iYltZPNoOFs+9C9j0SHrZnioBwXwhB
IqzVNhk7RJnwzUKmpSezq6Yon3lAPBfsUA5QdrB8lPd8ZBi42b6b9SdHiH9uYP+iYN/PGoj6Y7Ls
gecLAj3V5Y9Z7oZoLya25L662x3l9v07l5+7sf8wGmnW0R8tpDOKgJ+cLNIv6g6qu1ZNqu9SG16h
tCyqvg62c2g+Ch7mGFjf5rwApD2rkrP4cbgIb4493BbiWoYvzDBpdmhRUPXMm3+8KmHaOub+6117
TzzaWSkN6ZAlQKv5c3/W7V5+t36GxdnM+xOecKgy6boETVIbkzASFJWcmJMpaZEsMRL9etaXq5zr
a5CaK1Fps079MWpBOm3OF76r6NEx69fTFSpujfpS3QiBcx7dmYjmLx0vTlG51mb+8BtDK9bu1r5L
ZC81lzJzCnBg7jaNNhVMyw7jcapupCquO4RYeJjG80DnmY/HTZFz5RJQZG2QCbC5EcIMp1E8XxSF
8U7unGVEthisgiL4LyiIEWLl9GYeFzNRcdq+LVWOpqdCeEsxAs4ztNOc5NTEX3NSMahG6BbCxVPf
1+rqNTrAxwk0iQyf0hS5uXa7AboPHFEMn+3/jyuZndA8hH8S84rV3Ujel/wta57+tlI9USXwfMy3
4o0IyIj2SkKV4NxDZZPqgpkIlm8cG+C27KWR0dyO1UC99a+5Hp+lAaJta9j51I0Fs+0vO6aCLpXO
IZAzXabgKPiHh3fO+skcYD8Jj6WdIfmv33I70DXE7MXBIS48gSKYKv+HuBx/5kTCWDLxX8ZihdEM
VJqj6oM0FYPg6+C1/A+KjfUcHFv+JZGyoi6c/LkqTwDN9fNqt/OKciJpsaLv7iK7/hTnJAlK5+pK
wkW5/z+R8VoJhmH0FWvtqiOz7vz4oCQBWxpPXxCooL+YW/6j8RBL4TvEXOTflZQx3zLBAh2rBcQ9
4aYutW/+glGWGVBIoqWRwrjOP/SD3V5WI/5Uj+E/Hv3d8wGJYpHl9G/AnrlvOB5jHiPVuFoDlTLG
BdMJF0RQcBsRBgiUwdlCrawpn8kpYnmFCLdV5G/JFeqvobOVDQYoVnuu8t88kfYcp9WQoojFhDRA
ABRRb5R6gXIMAmzI4GrjO9M1XENn1iP344Nc7P/Y06GR1kwyJVDNsVi26N4ny464vATS4GAby3IP
Utm4cH9vSZQp3Xy9YNNMrPuZh6Y5v08i64BIPT0U0p5HssPIEOuT94PAdSPuR+w8/AekurkZpFIs
8+g8xWfvs9ScTN673QbjF3UKLKcq2xy7jkLWDwmRSJ+hihIN44Il0lmx88PM6EwvzOwRTbMyEowu
7VqXQkZVaoGeaQaiaxaHx1g/DMFjxwdoewiY10u7QxAEmg9iYDr3cYCLuN+JMR93dGg+lMr7eZFQ
9wNBMQs6B6ZGrYr9mX3VW/lieAXBKHgSHRm0x8TZ5y5eVekTUEM6VkSPiOyp/A7P264gxgT5Uepe
tLEVVK1ngNs786jhNvdn98UI+o6scilX2sHE0gpLMQLbblRAWOL9nm3udBkXOp9CwVBd5BW9gFuT
PVg98yw/GsbxHpWt8IAcaVHPwBzl7XOq5+vCFEA2AL3lc+Gr7lKc8Ko2xHWqRZ90myM67BUKOloJ
G9hT0KkkCrmSGfgOfa7ZzIILwcjpRByxQY9q4Mx7ARZqEXrPkvhSZbe+Ot1VxPtukHQrGsZQhrQH
GJlxV4SWLGxrfLacDEct65xSyPoqjMQBBKph2ZIYqTvxMNuppNvt8ZPRhJG1PKPb3WfOnX7e2vjq
DZXQfcSjQb4tXlhLYhl11SeLLFPDJVd1s9uyE58WeLva/doF2wL1inIxI+U8DPSD57ZMMgaOjmGo
1dVmISTvtRH1xkbLHEmOF5IjB9rQ3IDw+WTTiiWW4kXGD2+ar4irFhMp7KJs80RiZsbpgPlcTb77
Muh+Fd705+JVx+kIXwNpY6wiD9nXrrMMu31J1DlGCldN3eBCpiC24gS5zzqSgV8cV86oOGgDpC4P
i7t+ROdrVspe3TRcz4FV4o325mICrM18m1+9+6c5o5Qmqcc3y8kaKJdfbhf1YluGu9Z2udE6iA2w
lf49f+p7AokRbJ+Jnl2taC062QPiondyHjybD1vBGYC+xod7DRlwJTwb46hgtPB/CxUNkqcYJ3rx
RmNeUFpe7xnvx3tz8GNL/eWh4SyMi7yElmFvXq/k65GMpYyRqgVdgiJY8G0D98wJPDcO8+t/gE2w
Nj7gwkyasidmYfRhbhV/IsP42lDFy96bs9xhyVYtk165he1VOB51yQcT4+ZhHH3U9m45FOX1+nBt
Semvcdq/hxzR0mQRM9nqzrlScpl04rFHJhDaeFFTyJi/piS1D8scEIUF9t63Jum0xtp+0KEw+ZWE
F7MX0X+Mt0FhT33qoc8Vt96OcsHdrJyH1ji8/1kQiSlfGT01MknPHJ66OYFknAwOkNEXBRLdHSyd
qf3ktQK9li6/oXdIq6byhM90gofLC6C7i/w+RjrY5U90AoxKC8ztdq173hkJaG3Q7LOBO3hbRrhJ
GeCeKBXQyykqy8ZkkSzDTjJOKrBlUm/Cqx2HbWUlPP7O6+uAqqmD1hD0KaAa7XwNw/9mN96h/3x5
z2kcazIvL6/pVM3Zk1guP9YwJqgbmN0dPhkdgf7sn9Jqqeu6ECEWG42yAWiFgjKccL23pVfXiDZI
6PlloXDpMaZFDKJ4rc23ajY7UUG77uA2XvlyT0iTwx4tziWnBAVWs2ZEw81z3x44spHIdIh6nJur
jzTZ6joqvAKqxB+gbsxyDbkEFkVqZw9gMuqmJEHvkFv8skIY+uiXwfwVfXIDiTv/Q12OyAPVDAa8
VS0H1cE+7UoIxFssJc1NElE813tTSmq68cuOKFxSFFJrR9bL/bgyz+ZZQSVbg1SEmBRqEawX2Urp
Z/nL8wZjFKn/ruky/YWbvUYYEE/oyDtjGBCJTRCo91urIDul+48wAG2O2G7rCoaCg2StuYW/38id
BTCnhc9A8Z88LkWLYoAkYEfTQmDQ0T1xX6U66ZPFNs7DXLhxl5qG6V3oRDEAA/h752U2r9GN+y4P
uzwcX+nrtuRTMk/aYqRD/hq+oKigUn+fSHL+WA264zV8H6Zi7DzNgHPxCXEY+8ScXA6diCTZq5kw
5DK9pYDMl2FveochmQRURvan0iRRl8G+o98uJRVkqcmUDp7W0SU2dbOOaSSsT4D5VpMZb9LnJ5GQ
PV1XndFWxIJ8MJBoW2V/ssm/FXJkULim5Mo7uXUqjdeE2TmzeWLJKyDvur241eJuLG4/mRFhWQne
AVvSIVZic9bIm6WA34dkksTYYviqDzDwpiVSquocqd/hwCR7laTJpMKjkYOGysHjMBvfxdWeLhbs
dWwGSwkzXHKi6er4zsSopnaykg0yCj7NutMjL7db/MC0JHSxvd9JY0GY+KDecmUmPy1wRLghoLrl
0wZL7WDBcZIecDYtezQfOuQXRun+1uBjHIeCDWL/Z9HThTx/rkAQoWyUJoSyB+f6EVDAjyyU/1y+
C9sa8+Jc8Juh5uNpG82+BuCV75N493eHwoiICRPoAH6PmgDw4Jx5fXxhD7rB4IBrGGgdm2wJNliz
VCioVJEEQ+kXjjuWmtYKiKOmMKFsqFMmdpzUhPX/y1unpNczhqpIV87D6WibuuT/wJ2B2NaWoT/p
+Anis1uaofNt8crhkAeep065sWITQXjOdnetEmYCbTmwurfRao75n72ADjZxbN5HkdQbTheJp0hR
Ky9pWEivGcTopL3g19TF3ux8iv5RYQNtJZJf6mCFwGYUW9CugD/MxcPI6+OPwk6Mkpfahl27w+yr
mpoJOryV7xE6Skxi29pplOujfGubBTsQ5OzIEjQ8/Y4kyHnNOtNP7qKDz2IAcoNKZXd5TkSD5XYc
bMitERqr6MfKIcguK73KgXqKk7KTmyxfXiKvXgDB8T9MG1ytpkjnqQLz68lrY/nNB2+cWeYvGdho
pU9fSVOVbiMymZxB/8apU0BGtQVsZW0U3NEvC74Rh2Rz4FqK6L6x7bzMiefSp31S51XagPZOFkwV
Z0qLCMC6lzw7IByViRSAKcqsh02kDsPKsuXnxE4zur0mf5ZnNEQMlkXvQsFlR5aDxCy9LpkCFUOe
xsG/oUyimMZCrfC9JR26T/R8oReHDK31FI9orFipl7TfOJ8mszHRXBkLd6zXWUDhDPEb52v7Il6o
pOrFby2MaAnxW2+XSUksyjBD8OLbvGpujK/qJhOrhyWztuW5lwqIcesjcObzNn1f1KdMLXY+/Ou0
BJdpQVQbQ1rCjJR+DPVUlD6xhZ5TiI3Jx/gF/3QprYS0JpB+y8cRMlmPmj6+c3TfQhGzhTJ2WeVB
C4HaZd3CswG1WUaSx8gKscB6ssMFyDQVc7gO61xYOiPQlOOjULLm3/Pvmqdm6POKifGZjIwdcjA9
ZVOlbJXF1n8CqY8w7Gh8ExMlFr9DUiJFyMrT1OEXeYHkBpCe0E177yUXiJiul45QvEEPsROWRHF/
AUNnjDp0agvGhnpnd+bnoFdwVQjrBdEm+qEorOxp2RAxywalkwIBH/v1ppd5f5GfnPuk/hFYi08S
llGF/otLmjugK4e/mHMJBxCw53ITedDGHSlml/S8Fqx/Huq1V78QwEuSqVXMh7vePVG/5AHFB4Jr
2+cD28ObdK4j1lcGdL42w9VrTVDzG//K+Cwmn32LccNpzyYINC3ncMtbKkOQZk59tdX7qnxdpggk
4EONqQqk7bafaJ/Bhn+7QqoiAh/Fc8agvy3Kw0zGamT/z3YGLx4aaoi2Aa+CzkUYOQJUHEmGM3dz
uhEBsm6/1XFJQmJPeZPm/bKbnlDLOGxo6NeeAXD6tQzmWxsfULhIAyEI9HsTWcXAM7QoBNrgb7ju
QQn4yQeVZrKV/tSFilgxxr353gn+kI3v1rmJ4Z6tJhvIQC0Z/1TkOkOW5mCSjA3Ya10ZL7bGcpww
3kQkiMunSQ+Qigu7+7xq7/tpoqRGcTOMvPrzIoOYIXnAjqbaQYSCW0LsyRVN5XDNLDzC1Req3wC6
jMDkYE4S1grIJtvnxJxHfyWMmLD68R9a3v4IogBh9V3J+cEsV6NPU9tnx7CyxIu4fJZeeBL11Wp0
7ZeejFA9uTNlG7Zym20kAo0eOdFriopUViR+ypz+/JQZSpz8YocLtC+jLpwG+Y2mITa+SrVGXUI0
J8EX40OPCq34yrSa2zXXIpGzVdbS+wIy2TLMlEsmSKzOdAEmRzvueltRPTVPUQO3rFNU+j80iyKo
U8ZtSUzvztqSur0kOkrWVKT85T4V/qISDaPidvMusaM8ysa4CvSzS/Pn572pL6huBmENra55xmsG
qCnc1PF6EpUl8FuU+humAXllot00buVCXKYiWqhNfLBawVC6L5LCKIKN4Pnvnk1wEszrVR4EnNnV
mBnslU4jCTqJLEcGPRJltXMMgz6ByTol55ONPo+XCwEFpyQZJdG1/V9lS7I1VIXpE7ER/4nChU6e
i+y4+GwJ9xR9AIjsHulkqu0mUi8cmNE0BnUVvI/LEt9wpPitakD+++XCrJDni4H57kDCHh9/xIq2
fOC+ExWT+Dwo/uxbtiLxBcAsbKKy/uUEkpAedGhyhaOB0coTJuTOVwzZ00nX3+UxAFYHA0Wj9lhH
WYveyqifyAqFgg03nLXpA7jgiN13WsXVh9Wh60iFgfLE4uBxz1o1VL9aBDnP9mahHrZdD3d5o16k
baLYGdhrqTKqcUVEVjtRVxb+emqKT4RK/VAh3Kp55tLG/VW7Oo666UOq+ILqaTvsFVRRvU5lOabZ
hVNcPndA4mkz1GkKR0atK6BkGKXmQKaZ2RtsBWZNjD+1x5/k0Hze+LqVbTJNh1GS2zlS9L8ccm/B
jaMQjgrO08Rkxi0jm9ykIv+NTrvE/nnUd7wuQR8bO1oq6m2ffNOn6DoDUhdAyjbkT2RdHQF5cKb+
NnqAUTZoZFD6/cHm0TP1EXgdv0vslyIqqxV4TryRlStiHCNng1zKCgPbVxf7eKLCPL83KUZV/PtK
NqEn/Fg7EGeFJpwpLnMS6PA2q0qEEKv3z4Lbkp9B225Ix2mpBtIoxStYKLw664ZbImDL05rjrvpM
jChFJI83R1v1MpPi10AQQr54TIspVpb24riCi17LxFyfJ+ItkItDbA5k1X3NRiG4YBn7UdGOprli
nlsAPPIxfX4VIMI8B2qrUUR9yl5DaH8BrjT01pdjR4BpahlBnxTc3pZoTS7ikhwEtPedqP4o9FQi
5xC90jBDfOuiC6CergQIc6wDSlpCS2eCVaaG2S5LhSaCiY5yZUKNdOwkY/MfrzaYmBqVfjIKMY/x
+2W/1UXa4mQnEiMGfvwL5gQ7x0lVOH3YOeahYChkcAoh6ZO7uaBAr5AE77Tkr5ziThf3oiBPT+gF
7VgAWhKT9fIh1pRHgxFBZSjSezS8qOVspFi4+JMxLliGqaoOdbft9UFjz2xRA7wHREviB+gG13IQ
+Q8UB+7SI6X+ITG5DQVpD8Oif0A416UKhgdeD3VUz9+CfGmrBKm4ny3EsfDBLheBVB1A7IiN15Hw
ksE3quQKo59hLEb8FrbhLL1PFYhFNJ6maulVFBQnnol9xn+aYchvF6VS1HjwBvAvNTLNw7BHT4Sb
BkcKrj1myIbYtMRZMnb0KX16/iAnjTIxYnfoZ7EFPsjs5fLkUlu3iEoRJzsWE8b65quyhmejEJet
Q8v8KZ994grkl9DNFox63tJSGvd6De9vpOQkRGSNdbZZc6/VffWaKDWlvUlZu3a7AkOrsv1KaXRl
2Ne/rK3pDZz2rBMsZ2Rf2qj8TGxVZzKIJG7VMHYpIKkZarjgcLvgE6cfQNKCGeZ67h0hfoLLfvXR
Uk45zZfBHzp6nebZLg+5PNDTQGW5Y7rNfnxuf1P/wZBrE5ofOzHmKs/hZzFQd0CVPZJuTTuRdMzM
EZAstfTn/qNHnp1NGGoxmuMuX4amONn6/TMsPpyzmnE6EtGyQ+t3lJPy6kzefGSTwL5/tGD2h87N
z2s7iG3gDYEoT1ygRLIPDM1nl64ckk7VQPGBlzr6OeLu6M+AG5xk3dMkAbeGqYLaHEbPbis/kfdh
pJgJCOKOuPl++qAtmtUYr4V7BpHxgb4uHuAxSYM579i+0OghGid19XLhyTusFHZKK//JSsuRnWDY
E0oM0fJR2HKCLR0k7hagLJ9gxUpJPvJ2RcsRzccj+eTtnPt5jWhbNrMk9N4gYUXo4RcDDhLKPdfx
qU4l0BxfaZGn4BKKiSb4lsY/EDMCwTL4P0lBjRTMsw1oIQlcNi7pXyDd102mBJGS7yK+lnTWrRpv
9m5AE4vS/ijyQ2Dgp0W6HAfleeHDrUmc9QVMmnS3OaysBOBXpZ/vj2ZHm/XL43BJDYpgHprM/c2/
H4LQKlDRWdt7kffMgHioxqaK5z+7+spjGdykPzwaO1J3g5ypveyUdE5DbHvKQRK7V27egl+0MrMB
Mr92ePBQLpG6742RmHNyc5rOG8jJDP6QEPvrWnfv/pLh6pPF3mhGSJNRQ805A3q0KqMKW8IlZIds
djd08eRal4NaqSEwHBgUDm1Ql9ZBYjvZ29A2Tuf/tP8XSUsIYycYwz6KU4Stg72hOHg0sRjTqePF
m4aKQbhsrLYWS2Hp6S/6vYIZrVdKmjj/ggg7Mb0kcI+XCR5Ms8p2EoQhsHvh2Rex3f9G4XuSaddl
gbXJPxxiL0Y6iez3gHRL9dz0Ho6M2G3cK2OLwQ4h6uWyxXoB7LfN4MgfMwrbA4hz00syCJOz5RQy
151k6MztI8KEF1SjvLMRUkSAXPJtVgQwNkQx3cYPNhtT6xwz23FEE7qwVIKygKA6zUv96/zcY6BJ
eUKq6taHrZ9LqBGJFRd0Kg+cPVAVOjOKmQmWP5YuhGTSGOeYCxPOFGXLx3oWYQYrPQPK5Pmn8zon
wxz+VcjwZOBoSRgWpQwXCsirFuLjz8meW8Jox36vcSFqFN8nop/r8udrtEbwNf4ZCf8ur4/tfGvW
tsRUo2S8Zszz/DP6wfxiBpFPQ5/OxZPxJpbIKx3eSXKZ3Vkm8dE3S+jaLwdpByZneFCQRk+9QcbK
h5SlfkWo8TbXD27NksJcV8ONxxRGWTeI0NCQeOpxX0eTFZl4VQOG7ZW4hLlTp1hoCoM6stivQaYo
84aVoM1DjqE6AlzgPT5oFxqWnaodV4vUTqjpsVWNWgkMafX9lRYYchUC/Ku8sYFE5FORxJ1E8RKm
/UMhteGK3gIeXsmjNZsm3DavKLpR51/rlV+lTk5xbeF1ssqNs+f0kA7qvjW0dTTCgs203j+jpPqm
M/qJDu/63z5AozZFgGCvaLFeNlZiIdS9+YX8kFxHfcAmpb5kUz2KvVsrnchFyyGCP/DPl2hETaYC
jYn2VRiSS4fGe/+gDW6wBwFhIgbB0JY8IbAgmpAjeMPabMR2v9ebS9yble9nRrGdNSmK0j8KXs4D
4vb5TL/Lz85jHXQZbTdPbGaecSmmbFbdIW14IsmZxAXpVtqpTGSFW/Rc77qIacvBpzptmdbxFJZL
plj16pz16fA8LZT7e0LUegbSklDKzl7DOPlnIEb14pv8u/oTeLnAdBs0LQxisK2sSJhQnf0i2DcS
h9KW2lIFA0j0LbF7DBhe0YfASDvJ8a/pQnaSr8XTWJujT1cS1sUiwblMf4moGhrgixRXMTzibBxt
09UbQU+5C7dvznEmzOpHqhH4UFyw/iYxP/rsJ42dYU6Vf0kNbjUQSvt5omAYKwIkYpheoxKrIS1p
8Iv79C4KI6T/4b5fuyt8rKRhKlczbRJwp0gY28X4BOvs1nyQbXE4xOYuv1RE+gJudJJBIN3CCz0v
2czszpg9iV+uyUh3iqoZUlThGssQuOQ5PHo7R5taMRc9oUfxTxLr+tOyPDUZh+8a8r0wRw7GOyKQ
XTRWnwWffyjK+gj9M9+ecC5P2Nj+OTkKgQHuQ8Nl9RVZfGfH4BGFSSlpp2SoeEtLiFlrUoxFPKc1
7KC0yqcxQWsIF3d61/dWCEjZh/NlBllyzpL3spdBar8+hteyKTnumWUhe6ynafB/5fQSW4VK/4SX
oiGwyOGDcXOWp+41dhhZ9HvjIs6FdvxT8sy2nUYN/5RFRm/RZML5iApgpCjT8y55qhF5w7sVfqNm
M6E2cGU4WVnkGFZunyOCIkhi0T/OQP4T8ZKswmWAVQ/9jhvw2Kq3qXl2mkJMJFRPGi8dX+jcKR1e
CNzOH895fVQJDQ7jLdIKzf3SB58ZpE4EXyEJaOXTYJqyU5N0+78juhqzhcOf0HRKntCLne479Pid
gZzfbKJZoDttjMdC3GQTnmh8UXgTAVDRcyAKJ/+VIuwArgqaXk0lO+oTNyPri7q7MfNI9XVTonMP
vAaW2V3JFTjrtiIiihpTm/uOkTA2y9MosRRRd1BMKApOxPHmqIt0gEpVZ7EvW3+IgcdykA3Fnokd
njUW1lnXH5+sks07aWIJ7njV2lKKoAY9CZzGQgkg+nyBsU4yEfWa0kLoyrEj7Xy8P+aGlV6faaqB
hwRLA71nNyt48rp9E6p/j0KZP0kc+DncP9QCBOOqSujGGv0nisy5nhy0pkqKNRIFBYGW1txm/Q0E
NlbDT43VCGxvLythN7jEe8RwC6H/xk7Q2K8ksl7vQWJXkDX0sglfg+vuysXdXrV6Qsc1GRMqLM++
61i48lljqWAvrocAwNDiKOg5rs9yivRzlIjUFqCAlNEgp3AGAlXTV3XbPg4G6FsCvnKyDg7zMdyn
mv7TZHrZjxUENlehy5DeZurVcLIdIpM56Jx6UWJ/r16NFQgycAQKL4brXk+3HPBCwyc6N6tnT9IS
NWyQNRweZg/qVhF8EwBdfl5ck4TPPcJ6NXeuFejKI72qQamhgLlp555WJEv3+Rtde8GWOPNpNqvN
oYdYhc9zk1pHPpI3kOOrDtD6skms01PMXbrieg4nNW7lmNFRLjgVHz2BqoL8ts75V4ypFRJuSaCT
48/icWoZO/4/DCnYcER+/oFN1veuQHVPjTJ5eJU6x1ByX7eZs80XwNPoS7dgiACw+iiDwa/fQmrT
/TTIP4y1rSY/eTMIQx7E3bXUndDD9oOVe55qFoDhALI9BirNvNijqvtEy48K1YGCN8xNbfac1p+/
bKADNeKK0HdM2LZhKtOR6dla7e/XY6zhy63+m4ijghOJGRSoEoHPKU4c5BO0hdMF3HWrjwTaghwy
vYunVdabq7kUUfYoAP8WzEx5c7pv3X4VhuCeGvRXFN/5dCMQ7CLJEh2OJPWM72kcLFIcpHjNYYFx
LkevQ4c6IgTGs79WtAhnK/0OKx55B45aQ0wEzfDPqBby9g1dHzeOmkdryYe7ZoE9SoYkMjqXPRYX
yL69Z5EfsIN5ouZZX+PrOpKcIv3xMUKJFFT/2xgt74KTsq/JoSntHudY3O121rjy6Npy4j5Tn6oI
0IEvOuvAPZoyWAvwfHADgZuqtMyJyJvewv7QeLZI949QqCSee//99CFFZJJL2DaezGMfBo2JS/1q
UanoTBluSNuq13voDeckR0lrD1/08s8jvPkVyk7uPqxuW3rRouyDU6UuIQlWmrzE6L8cZeyqIl5p
I3SQfVV6rHkY5SbFOGgVbIwhrmdBXoP3Uiew4k82jPx6u4BgbWziZzUY+Yzl+rOnisj4HG11mKQM
M8uG+Sh6OcaQLT0bNTfSVYNVaAAkSBOb83NAjxN77JNUL/V7vC8jGXls8xRSgRRueuDcLzm2LmOI
4h9/NbpbMNXuc4aM0B2EpMWmDKD+GXGpvQX3GvZdYvRfUj9sNsZSNXA2hxrMXTlNFz6tAniwr23x
zw0V/6309EOXShMQidohWhtvUZTg2JAksORC14O1KDQSY4puq2IZkucULEFUGisFuEoE+So6Pi9v
mWgELUQjiXTV4vAbFeYkqjU20tceovO0oq8knWwgEZd+I3wsLjp/rpd6wegPFlKtINsWLUsUxYHG
iD4DTq3250IT+DfRg3krOqUQHyGPVZT5MoshpKsto+LPDvMoNtK9bqqY7mFUlsamEVCZGdh3lVwH
05A3fuJiLvGsUOlFiWZvgW1BCwNAZk0EzRHkOMMo7TNztd3mGfWJSsflouQ6nz5u/LsbT9fSBHCU
RZHc4IF+WPOulErvUM6mid965N6qt4QN6KsZOap7shqEVVH3n7dBMTwiyLeq87c8mIhApTS86gzf
hwPLQGNOLIRmGdeVx01Nzbn7B8GuUW4LEsbPmbkal0angY/fn9ZE3MWut3Ak6bBWZjciTGP6iyBe
U5JeXM2522EQIltQ+dnLArVJbzZG2defDncircF+4xBUaWRh6H2fdeHjzGJLVsD9YYSYH3+h+CHX
ebqip0dkr3Y4wHIVBvnWjYptrOw7V39Eww4DTSUrS2vFtd+zjLUBoj8fe7guclXAQMgppnqxGXHr
PT6wcWzvyv16k5IrNKdyj8PG6PmNpSFDDQ6s8cNhVqbxv8wFOoU/qbr5UXaKD8NkMSqK2jp27P62
/hYtqOvxjhhmcueW99oF2Oy85lXOpeceWGEczq/nOxFSBSwcT8cHm6HyRXZScDWOI1kOENBkfy8I
a1wqaxKccsxppP1uYNWrQPZvF233AimujB2qP2Gykgcxkgh0pwwHXTJWPfabBkDN9vZHk3zFG5Mx
cecO9bt4SX0Hxhjv8Xp36QdNcEEP+HsrStbnpkU6gp+1jHgMgG3QQ2eO+hHm+U6vSC6XJvk8WLDo
F2mn7e5q+SiCRCXPif9e7qr0WirH+n19ytHyeJ+UmXnJ/iM9VAgR18pMUl7Hb0jURsYZuJX6OCZr
Y06oDW/ogAbpt+ZpEk6gQLMii3Vkj7JCCSjmGsHyKAwH/WAaOrVUKixWPneNrPZ90OvzHZA1Ja7f
0xTEnWG6VYvgMhYeBuDWrRrzNKfnYjlENoSJISexg5ONjlbwIiiLo0qGf2uTRDRB6vz49nE5MWgk
EKNZu0sTjGosBs/3ENRABN6cvvZNaa7SsKabmK3uxKIyKkcw3aR/DR6/DQ82HQYgbRhXlQmq//3J
aEEWc7ZAkj1dYfh6mpzBP8mWZW6oHoTewl0+2UDcfZYrF20Lzc3kBZZBz1UCENLFj6eR174Z0sx1
ZdJHsptoZfHwMRkA3lQ6gHxxb7ESlJq4zuBZcY46qFRdV4Hed3f6DQbAmPK+y6fbQ6O0p0abLEVz
dPDi8wnapP4LSQpSM8zQzF+PJvcbN2vgGsLMBZaecJFSZc/97qk05QuW6nEyCHGp9uStRQKu5pys
XNcS5qodUC0OUMs37M7DAF5BWEGICD9oAoLkUmsPk29hvmDU88CJBhxSAOcFugwBGvcFsF68c+GT
SkNsD9roFoS7gvukjbsBMut3fZZ+AWmU/k5jo/dvXDqJhTUl7V2awhjTeInRuqrkH2948WSfHA5K
KM1WbBzrA6u233hPeb+fgWcb4E4Qk/XyWjWqIDlKxKQqMsRst2Gtk+CWElhZXmHDM3/1VGyl5oHg
oo8b5lDM6+nQNw74WSt4cRkybXnXXB7HEfSIJzC00p3BJb5xPJDJDYzEpxS1/9rXAva0LsazyAGM
dax+Y0Pvqkv0g7GVDu2AhbsG+xUnwMREIPh+EPvYCa6KhBlmX1tbfHuARJWtJjq/c4C+AirJdTsL
gb+Me9k2unqgu7jNLEZ1fXBRq0PG5VnSufi8UriIGd2BOKMPo+sQIsIJdnsnX8IPiwNV93wYBqhU
xi9q9fAcCcb/6KgWiH2tLDZvg2uQKnd8as0z7CVQOPastwwz1cquKoLF/MkZBnf6ScGDPVReY8/7
aOKvOyjMjR7OInRIB46g0b42IgcnyGfvepgCcQdmg90ZdF47dgv3/4F0ITZnK4gsbr5494o1eYkL
IiCvOaHKLL+EaaY5hUh+tgL7mbk/yEpCt5CACFaqkQto1+c5aMut9z44pOjuGp+8rv229EtE8H3y
F53ptPVhUzkL2kWwTwBt6bjwUV3sY9Qdbq4G82lQr+i9e5zXET9uUEMterl9cOqRznCvs04qfVsb
WH67VVMh4/fZA5zY/Hgm62EPASGwD6GcNcxhe3vvXNlWTsCVumG/SdQSmCy0xKhwtmEOUI68KxW0
2H7TVEGmIglIyP6yj13fW2Bom95NCP2rXsZRAu53ZX1fMU292iypbFJAY3dmH8F+74AH+8QrMgpe
nW0Ft0a+xYYa4rWMJt0A1qp3+f2HuK+AwAyfOQivqpU4JT55cv/p+SP6MQCDRLs2TsitgqunpFXk
FaRxiAKP8kN6AjYtTHLmG3MXfwjNunVZ5t8eTtC1IfqdZZhriFk9gpxx0+9gkG0fHXpSWHXUS6p9
con8AFHWP4C16NRTfdhQQmCEbItJ+3cO04jPk3l4nqAGoEJZ/hfHwNVJYGRmwwXCMxn13YYWxauY
SIUBvF5tvoi/jsCG4tnl1Iy6d0owhtOH1juYTBHR/tQlkzMIF9fg+bT44naeRs9Wj4HAhIprs/JN
73cymq4JLQ3cqlFaz9G7ou/W839rMaHwWfoGVBLWZeVH/8BTAAvrTbESGXq1CmvzCK4ZXE72uzXL
uuXmRdqSSKlLBHyhWKPHdy+VTDiMhau0xxRFS4tlkR4Ztuh2Gi0TI8wV9l/44wENIEOyzkhHv0EA
YkELx3nq5T7g4Y6VBLVawAi/JMUXs1BTU4lKxxncE/LJbOgeWsUie6Xc7Rd83v/eFwNslWyKalYn
Uc1pFiORbTcOVtc/EbYMXeuPMVieyzlMKJ2hRmLIIepNfCVeTF2O+ZfNYFeY3tFi0OzPjkwso/ex
WTkHwXFohXKKzMJ8kobEXS/BAFqLQUzTNx59szGTnEtdQihwRs2XaqKt8cGtrfa4pK8FcfzVEdPS
dBTeP2kWjdSzQ+MJ8R3UwKCk9KemFjHQ0sFzX7O4rrWT8fJE5oMDGUTBU3zeblBhPkx8+1+NdW+6
usIHmuyB95KxZNJzLAaUqs6QKbioTy3vx6ch3vpA/KhnyvlzTAjB4KeONLNoz7cCtODi9tubSXTz
gnVSM4+4lHK7+E4UMqwYBDf8LRo6IPdkjbSIEZqhns5Xo3eX+7W8/d7OIxQSCjbMSUmzNHcQde2s
PLQ4ma7KyAZm8k+M3COvyuGGLKL1kNvdRpNdP2ZxT79VmLIphOHQGT70qhtU0d3b1/oHoMuvOhXJ
XiMdhJ1iRIONBzZwUt8IBN2+At/I34KSWJCbjVXwotB2TZhZutoTJqDRLQmCu7SCayyvN7C3YBcK
JKS7RbI1LksIHaFJV/DECwUBkJLnPOOfjfyAs1l1oVGtoUNQDWZ49bc8VDgeh8k8Ks6Il6loJhJO
N1XsWsERT7Vj9108IGkAiIoEhUQVK7BbGZfjhcQtxKpLRk62ZJEPyKghutqwAnPszxQVAfiut4AV
+Ij8Teg+Ncji0WjXMWoN4FDNrD3cKB0BjItPED0UJWnNUDk57ug0aVaCyGOUZ9PdA5uTWyH5wWkY
wbxoZ5WhKU8cGICrpm8QnDMVAygFhUUOdBYsdYg6zqFZ13qU8mcagiCiR4FMJUQSWOpM9Yei4mlu
N4PdVKdWmyNJuK936Y2II5cggSFJF38UJYTRDmvsa7cKznv8kwfIlCbEZxnyJPNBCxXsrr+/3C9q
zadigouKqcOB9IXsqIJCFaCQwHK2HrDFeiCwlLgLjECuW4F1ZZBVgftBtbipNJOMRc3fpWx0CRc4
GfNHSkKaqIxE3NCxhPZP+5MuzP5f5crrn5O634c/wh4yJkMXpVh3kH261WBva84MyCnLKVoDPbtL
xC+woIxgGL4Ex5H8+0Xqq5JqSUdCQ7xUwzsfofx8wGqdQYDw+4oda8vLLoGHjDUtjlx0AycJWP3A
RWGq2uDcrFIPzjL32kGxS3SbnTk239D0suBc/LY/xS8dJse+vYCAM+stcB9q9W0nrKYrndbpc2TZ
aTnJLVv3GvFqxdEZlgmFuMuoSs7JXSIPiuYxKjS+jLtQiA7Lu2LY2NY/baYvq3uo12I9jm+YexZo
a38OPw8L3JD45QU/Z35YOWnrqp7NYbDasESFla8xxglgnBkwdcCzwVMNpqnnjHdUH0Pi3RKutdJt
5eWkAcM4LVvSUY4xa6DDRlhiZjcO/l16Q3N7fiaOzWkVjg+vBUge4f9ZR9YyDIVUvPzHqxcQBog9
NS0R4JrxH91Y2lyRtApcbhQaDrXKyqvqu8w3++9cHC0YIjpCAri/SovYE6hv5TWeBTeqyp5hlVVb
twsSqWqkFB8BRjK3W0ytDU4fggAjvW+RLuxE0/IWTcexVZzTFrtCRnCPrXtggdIec7yOXPh9HWcc
Uke0xOZO2yGzOEGoUSYiWlqkG99rMk1jOlegBO8/qEUqfun5PDg/AKRNmA6v28DGZJuSLwkdVYsw
4Ilt1tkuw1nxrKbPyXdHKJCv4035vLNJ9YuI20kasQvazivANLHzyLIFGG6INonf86LxGuty1QTz
v/8Kp+zKAjYYuaTBmzZe142LIHbaNZH/xmhAfIR7NzyLvHQp9lRg/gV6mLjqWga0GLOwWa4CQIQJ
RO98G4uKTFEsVf8U4fLvHKduS4wGwictW7l0wflBOSM5LstiH8YgwIHcAFdmIapzgHHGAPyZtej/
IwN/4+YDrVhSwCD0AQG1h+a4cncre+fIST2O6eT6lEM0zFr6BNy9x2vmI86eOU7tGEhJs58zg6SC
q8NOPCFb8YAcPBfkI7dsGEtAZIrpE8lrGSK5dg/i+4/GwxhS62YtbErF7t5CoIQX1WEBLZ0q3GJv
raHr0Bmj0AneNz1sMhJ32lB0UhUns8ZUejKkEr2Id5EP6AC4gPewf+g3CzX+FeymNl6iW6Jwp1dQ
uTUsqtX1k+DwHXDHgikd7cxlbpeYErs6qKv9Nl/k/8D5nSJe1s+3BxYkHPBBkPQjfo5CHB03sjUE
Hwzi4C5SlCCuVKdEzLgWAUi1UbCkcpQDfFFcEPJYPptUVXBSpqZ7B6grL2pwvTPYSgPgp6tR6OCF
kCjGkVfWy6jNjP0Ntt+MDuxiwthXUWmK+u4re3v+EFM4Jis/3VyKEVRvuEseCZWNnuKZg71fl1xO
NUYdb9n3fAGkWThKYx+VDNlANEzq0uOG/srLLamZ8S04c+W5qMkbXXPtwnM2jOx//hln2SFvOSVO
JnC+oQF/18DeF49WqwhF0Hcm/EznSNpi0vAMwoBhKrG+46zwVPfYjGFfVled+iKxevc+/iOX+CZt
iNpvZnMs76wSOj2R3FaMsYqpIMOHGd7fOyAYBPeBOlG+cr7ZFF+YURSzRUQBbrHZdlQ3rNyL5R1y
wRQJ5ZCpsym9EYj/zsokPhj83avjjsLtYXtJYQkzlckRxyphlTr0Lco2csYlMwsThaa8LAICQXtu
ZjD/y8RvD38ENEapTywdMI9Tl6q7P4xDUcCZsWUzFa+CA+ZJjM1GqJK0RvRlqNECyT/hNij5D/vD
DiwG2fRPfnCfO0L1yIXamOWpQ6PLyZW4vkjSc/dXMmZ/YzSHQztdHpxGHu/Gy5Wqs1P3FcqgPJ8n
xozOayCOzd9+5Nl4NHnVEEMd53eAdANP9EI2M7JM4dqXkQOyGFLiBW8Afwa35NBHC6gUsvb4Z5gR
pVqOfN5V9FyMwcCu/C3fFVg5djS///Y2P6pGduQb3H9Jt2aP44VjPFvewhWWn50eRrkGl8WjODpR
s3BWZYJEZdSSANODUiIWpBjpBWF/MQzCGD4G3qz28tC8bX34vNQuORltPcuxMMvMLTsC3LDnm+vJ
g+IYV5ABAYzwW4egcQjtbV/iqSy/PszmRY27NwC7OYeO4FoP/EIMYtpjUjdNuNppts7s3PoUc7Xc
GZKRQkfPiY549gpHghgQRsMA9qxHS32t0WKYl8LEK5hj3o1WRCgAw9pcitFTmbT8QoZbLae8otfe
R0NHrv91cPOsezxRoQKbbJhkcoCB5Mt0yUlSG14Pb7wvHNNPUjLfTV7FgQHsfPleA7957nvrJ1FG
lgreOC6BOvlQBOsLeI7e+CpKL3U8Yyj1PApvOtCHd17AMZArLgfkwTsBLlwd3x+yB+Jl/UXT4mhS
IE6P2Nyc9ZvZ+LbYIO2h+gX11Oh4+eoPc2L768mFGuC0nhw4zvgjYrFJMJl0Qb2Wqg9zZpE/Kjos
CRL9x9JJ78lt9dTEkT0yNAPOTf3U/vGwgHV5NTI+7GeB3ZeoVjUYbirFxbFaxr6Spmu5CBIJbZji
5i+3jZO3G3sHDk99hiSlC5dre/9RSt3D3UaDM1+zGgfrRBnDS/sBYHpdh6rEOwjSPUfGsSm2c5Lc
7p8ZUYuBMKDJ7bwB2ZPqX8sIVJtQe5nY1eGtSNjxhKNlj7/J2sp33Qgo521KED36/al+e6LwbUgk
yiWQSqRzpuPjgnfDG1eduKlyWuTRdMOBh2zy9NeISaFtRMwTmEN8gPVMa1btelldNo3dbH42ReNo
Q1eMyZYEKOWYuKAqF7mWHZJGdM0DZOXHxy4y7oHoVYrRorcqSbM5daA1YOyymuU8QQQFGpH6n2Nh
uEK9EJeREMVCSlyMlH1Ou5bqGGqXI1Ouvz1OTt2Ue+4cLHZbt3A3pkgYR089BeS5Vtd7V8Drogkd
z9nzxYMSi1W5P/O2sPXov33Lobd/miTpOPAjWAURQy9OcTSwjbdC0dgXs+r9z0ygxGBZUG7duM0a
/naJ5lEu9flE6DyKi+i41pEKQzeVSVoVhz0Kr5QfL4Rf43O6EHe0r5E3s8HvIJUxQbRC3FKLbEJe
f1fIVbmr1Z9SG7Nvo7nxl5mXxbRc8QtSKmAaiQ2fmPcr8ONQVJrhQqfQ24OnYj02de9GmDXibZxm
/hjTHc6OircAgcID6VupQIwd8l23qmSeWBFC79miftjQL51VH8eWfND26667hYHroH/ZBtBAHLb7
HUPu9YV8hpREXQ/ubgd7T+27dQdqkVvyDtwK3DJf4LHYX8vmZlQp21dhlfbkma6Qsj8efUKvsXOj
oodaGo46/djNM3tqVQNLIw34WW3j3j+0u8ra/L6zdMg8/Dal+bs4NZUbm+Z4MhQkK1RCvpdy2285
boD8XSWbdwqqV0mBmpfynGzY8BCx2qFvxRKIfYc1o+UveYnrPm0WVOsmDPXT4IzeB7QChKjvxjKM
KiHkSQPjFDEh3j7odWG3UlqvJtm7wx/KRjlVka3hgIx6jz+Ho1Px0LdHnvUb2gkpsc0NIW57z+oL
PlJbwvxC2JSO8o6Jhz4+L1eDd3E4wXae4dZpIigYqULojMipnmOOkj0ba/lVuwY4c6GqRzW9tnoG
/OpQLraPUl7fAICq2ZsiPovzq7k12Q6ogxso35IJFO6WBcaO3hWAyN39QtgVhOwhdygwLYL8imim
v8kc72x5nWRM1oxRGzF8wVhXKTWrmTsn873TkbdQwJSb3oeIB4EOo15FMo19EtF9nGQ04CW+SfPA
ByBeZRtL3l5WGjWZjOh4urY83B2eQ1jlXoe6TU3zLV28dbdbhu12Lkf+a9SLkGV3VldOtMM+rZVX
qNBJVR+oBAF0AzVmG9GcnJtuh8TdwkyzajONFLgXIr7MbOk0M8EQgrJW987QUZfEPg8PfiacVrlL
zJftRuXJar9MoROl/74BXRud1RAX3jCscLMu5LeW+Tvo+Jcn13Urxd8shdroZlMii4T0Mv+5x63L
RBsaG479R980f/jxh1WZdjC+eno/4u2iaIiwCzRFxi6SoCTJ7JjvouQwCYAICT0bw07fay4BXfHZ
TBMq3CrOzJ6H12efTeMVNfev6xdXdw64bsu0sJMufqYOXPfESSQQj0RQw/NVKfZ2nFZbGkdkketR
hlRU4pDvHOg55bevnV1IZVB4CrrcoMc1i3jFddEi5YrVC4fsockMOr6WsLWiRvfAth0CcW5GNWFK
FF/QN580EX0q251e9dt94ChU/Xi5Z8nPlgy+R64ycQuvVNvzyUhYDkbaPmq6VlLnBs356jMD+5Ss
479Bo5V9IBHn2xCJAPwb7HeZaTLX3dZnC5YC34ZCklqn+DDFziquMNQTgE+AYwwuMLyZ1UrZ0th5
9VIpE6tf/Pypx3uNEgXOV0RnqadAzDhAGFpDuvILet3Ml5nqYZ2hcaQQrXIFtg2rhZfZFktOeUGf
aJmr5x2dJdbIesovu1ZTu9avLv1MsEyUw2Lxq8ykN6i3TIZ+BubEDanvyqCPC7ClBfaeDSaI0kun
ao50uLgpV6XC/C7PE8SxiO1OS70DLqcZXBXBFYb3Jgh0ExOUuxHSIrIzzTxQzgD0EkVVbYYNOIzr
Qy2Ls82Po11CJAx3bYqmniSnsB+o4DxNUP1xNv3+sDzgaUhTKFIT/zknqrfgmHJiNej8EfjE51CO
nWFk3k2KKyllLMJVyDf94NmPLY+J5DmnjAKJ29XD6gMGBegoQgss8vIk19Qe10ev+Q153v3oRglw
IP3/UIUw5dIP9ZfG2lNydf/E00oyFnDoRkOH8h1OvLRQ7NhN7/hJ49pnHcv6H8RZQ5zbKnOWqjjP
lgvh//2t4mQhnBDDoYV266gKIexGXCGwOZRHDXSJX1MPvuT3JRv78mB0IGOiU/dbzzT6ojgf3R58
GQxEeT72RqMLoqnE4s/pXptNHDhA1chPr0rb/qNiymTj8I12uWvGze9TRigdIf7mhAv6sKiSWNCm
q1RNaN15CQVk801d3KDlzxQsXYx3KOJ5grJemXXWKj5VJnRw/cpLYKasoOcAXsLkAGqnzrPMzCA6
wNExa5k8/85xgqRfnbkLGN05cGbEvCZ6SoGD+rDfE2WPFK671NlZjI+/jktYN9prN56GCMBNJgyK
h2DufgraYeDEPXQjby5o6GK1ampemM5ZQA1aOY8PSzIBzzAvSl7qS/Fny0RuokibLCVHRKVzNPOW
ab69W0QeZGdOrlHE0XYyPn83rL67IsimY91nPuWjlg+Vy4fE855QaMOHupguJqBMrPggTDGsRXuW
qy1+n8aRlVY3yfdr7uzAAgguhG9T35ER5hqVixIArZ546o4TaHWZqwltnzrkAMo59iP16RZpJYOd
lmEKKeaCOcM7TBP9rCKVo3m0RUK+DvcMH2tnJ1ZsmP/YjSrJideO41XfISe92gI7bLNrnSLNbbm0
UIoB4yiQAmqpbGOUGkm4/WrmGeHn8KkjGPW2ppeOhSjr40B0Z2ztFNe8J+ZHKf5nnblPML58rXOP
5inP0ompbCgPvStJsu5hY47E3N2IB/vS2Z+/DFUh0uCmFwQzFnftm9AVqlWJ7NN1cYDJFoJibm+X
XLqNGJEaDh+Ol+qYOQFq2So38V/Dkm1t/Lb2abYZ1Z5DRxSV+qE+Bn/EeqKKMn0wWRcnfrFYzpT+
xG0bvZVImX8nUJaxSM3V1lNkHPgeXtlOvL8I5gcNoEBXsELwlz3qpnUZ1mQs9LtY9Dxy2MFKRrPi
l+u0Uy+XBkxK7C/OoE1RX2A689T89lo1UJ5Ab/Rldprtkx7qdq9OIgL1ptrxpBLCWicbCEM9mwci
J016IaGRxFmm9AdXJB7FxfLiPCqaD4X+Xn7D1ayC6d4Nrw1AgE8WxMaU2ugRHprk/XUtGawBPdxP
OQCdgPZ0pkUc0ZWE8JPGHc4rcJaDYiyw1cQxNPGE5LiPOeXbsNRyRl4Xc4mUJwxyVltYvCAcaQSw
UyUGf/I9ynvgRYoIPXQnM/dgwvso/SYgWAXX2yI9kREkwb0lK6y/fbj7v/KhzbNag6eOz0pvqCrx
4KdAEoSQdeqY/BgNlPqxsrXLKSxuRXOm5ybyuMITl4+mnt79Qt8FaBegHsmPcdGnH4fWkxFNqtVw
Egj3/sZvllKiMkycy19K7QP88uU7CcF+y96KaGSsUVhV6zObkCmeUfBsg+ZvrducLsQDyuj1Gnnz
/ODiV/NClsBvLpB81LglkX6vPOGYz0bEv2DY6RET96l/euzw51aGCGDVrP5faWrSlrNuhGCTXvXZ
IcW0FO/PZBaed+Na2BGkCTb47tH5j70b+/piNhWUhWkbAVPZThlwCUoNC/6Xk5kr0F7QVhwheq4L
NexQE6SVINgP/LJPeGlOrNWe6Rgx6prZ5UY5Zw9o3uA1gIpAXFLMrvL2vEy4J1UNRD/13PNNg80M
7agILIAW78D+J9Bp+lNTFvC3YNQWNqx7f93z6fGzji3JhFqVxF19rJEywgNUlzo58666xz2xVbiy
WGV8av/0fmYDfDyz0Cf58d+A6+TTpACndC0GVq/Xf45VEhDL3CadsIkffV5/tBR7jLn4SYJrGOan
4KgMyg1ihd4J3vu3Z1vSRmi3k3bfXmAzPJxuUTtv8T6Ew1OtbXIHzlpMNTE0hjh778ed9MOp9gHg
lA9J5JbM8fFe8zsv8BVF4ADZlAepzUylt3B7w0cfbus7DL6fz5xVZBXtbjiQOg+YaS9w2EZVLbfq
PuXkOoqnfgKoTviwim7Bb6uvNF8mXgcxEgxnV4LzM0v75sWRfnXPb4IO7740EJpDZFgEKLnegp+O
/ObUX3v22qu+bgKVA9l4ENNeL0IUI3kz6g8H18pk3Uzn5mhuywIA3IB3oNShBGLAHTe8FMnqdp0C
qDCE+Otab8eg2d0kr1PJKi0IEy3Ykv4EH5uecN2SNyFG1UNRGmMnSMkcEPGVeyaue+mCU00EmPzC
IKq6p5WkNFvqpLPFu+YyFu6/CnLdvC0ATG1XF+aozxf+CnfHD2d0WGBnm+ycFQhaniSKsrfcT8hA
wZDR4knTBZdkbRy/vI7y5/AYS2TkHMwhSMfp2vtSwF9M3umcOFCcLyVzQt0HiFHaHRs3KX7eqjKU
WHguBoOF5cJ/CKYANVblVNNNAy3MQSdSG53Sxy6/67XIt5HLHRPUPvIbeMEXnoTlQ3P1x+6YUDPk
pWqPu6czq5lAeUeI7zIJU7YGj71gZg9xyjPyS390L4hBhT+PM4uWzmBPZBFI4fmdL4+tFraW9Uk5
jlvurAk1d89fhnzJ/jN7C5Mvzbv9cNAJ40SEGSEnxTwYbFQf7MvydC6/4ebhYOI8yS4y4nw3izTR
wqpKX0h4uX7UphbzuuB3MOHqXXZlcVujQoqyV9wCok6O/NuDx7kgayIEUB4ROs2a51+Sq5kfgpiw
X+zEU3ai3f4vCzH24dwGJxH2Pbo6V2aoCSHZ9Y0Oj9Pu9a4pn1avEj0bir+ryo5ivHWqaEQPzLRe
1KlNt2JLV9xYUuVKIQ5mSbZ5DXkcLBfc6zFz2KafYMQmfNkDXJQ6PODPk8iBD9jMDH/EYggTrK+2
9nDY5X0TvR2N5P1CbA5QUJtAydZOaY1v7ppf8UDPu9rNXbPw4epyhFCdSlCQGkgEnctyAuYVK/JX
5t+X7s9cRMm9GC5rF5YhdDJR24VP2U3/aqd4SPOL4234UHhqsweSj46NEv/b/zWXj7wcwHQiwUUj
uew8bBhLP6jjwAF1ned/faRvJkLthg2+lryEOeOcGbbU4uONriHIlIiAtTV9n5qZmz28UQljbpTQ
MgvjpkTQiORMghppAcvjrpGKcM615zf7P7XLg73/JMqAdtZjdgZAXKrXHeaX682hwKYImqvbSFeK
rXS6XxgMGe+qHwukBpyY94iGpZDoCtayiRSWCIISKqf5dro0Nc2CpjGicHsV3WD+xmGuO8sdj+OB
+3m2Po2PV2JEkXV/4ew5/bDrqLiwqHkrOa+foY+/OcbA71CgMJr2J2gLsFMGlEQ22/jxjb9rkqom
kEfSMNHoOgaVByPd/LKqSlEYnBzJ5B1U0qmQkXj17WoLuLQbzJ7JtquTkrIvTFHQh6XWmhz5GGae
6KkIYHXbjstLdxyJz7w7WFvRkfoF89kSzUwmk19tr8g1TLDUDlX05+6gh4OXbKM39i6WGOqHOli8
jYuJt0RirTqmxZWuXF5U28tOa53NtRAofIxyLfb2bF8AqXkQlmKQM4iFtCoAqs4psY84fuBVzG88
Wohh91vpgevS2T5mh59kQ0EkIxBRrJBwtKke/wu0UrrTxV9X6tGPUeE04ayQAaQ/SNaIR3W+OoSg
Fhh8Xdms6Sw+HHvTSn9hqnEls0FhV/fecernDTN7bYMuOLHgKES8uk6Y7Js5VKm7LGaswtb0ItLw
vO/hVoQ1V48IeDCnEUH3ajMFjREUSELiNdFVj3NSw6HwSt15fSI8OHKGU+U88f9sX9DqNvN9nA0M
m6F4tf7b5Acox1HLB7fGwlmWgtcy2nfePfYYb0X0tSh5fsK4v4oQP4xJjWQ2wCaPRkGTzM0lMeui
bjrjtRrwi7kLdkvzLYQzZy9Lgev3SNs1oRR/FuYSetPLHg6nVEEN9Ws5C2MHlF1MX4UNlxWgQW+E
Dn1EH8Gap+Oiy2qpuUyvOv38QR6Nd1uBjkcNAGzsAXln8V74++GzD06PFgMI/JA1jzT9a5S9FtfF
DvOKbZfNRiPGOpS6wqaCoaVPcstV3N4U6T5dT3QD+KrClBBcYJHso8EO95+QisCZ4FhRXZ6Llrp4
5K/YtROYXmYdjiZS2jlxJhjbLLtB1/dVZ6TCF3AulhQ4fW6FTuJyl1mN54stp6M6+WRD9+T2wqfb
iZJx/HqyavKo1eVpB3MaJNK/GCKGJZxGmhnUEv2k/8sFav6dAcc/HGHmLrFz9wAzLREhCAeCXZRE
C+3/di5l+XQgDdLoZjbJSZa9/9Ck7wv5HQCI7VyoNWPa1Vg9cyLqArC75KhKxjujP7u6VriHldFg
J6z4pT5/KL+VwDYTKgVSueEs/nMjTT+qmcZj6j9zuya72R4XHyWfgiqR7oWh36JmabNWtnw2rFDW
ocKqI13cpAZX+Y3Qsw1AHMWeTUOnIVvcwIgPgLSuAW7eAeGSJxYwnwOOyjAcgv5oKTEdP1ZykSdY
Qvk3WlhJ8ICw9/y7uwWy/fVHd/0Nw4nFxUKWMyBw0lt8ioQJA7JsV24DwXgpF6Ua0FuIkSTYtjVv
Ap+7SdfK1dKw/qOmibq+oCg7daRUlnPemJG5JNMqnnHP/Hjt9vEN5a4+VciA15sFMKXiiHH2ONCW
Y4opkpugY7tshBT8yDFNJzErjYgX9b4XXnNqfmitqulW+f/CTDUuqLUXDwOxdWdGjImZA1VUw/sj
I7MkGGKBgRaHbhwFkrb7nQ+qrUGdetB+4XgXdUgzA5wb0boa/Vd0EXjdXEYvYDqhXIZD+OYHhYnl
nqhUdM57bA0cYbNfWb/e745EDwsS+qCSfQ+TsizXo2EELZYQniEE4GIqDT5EJH4g5Kmgck4WXtsv
L1N0Y/x4ng1FeLf9FKRl8MAYfZbdn+dmyTt1YWPC++3kXcYxnOYAuJDQH5ZWVXZPkrzanofYnHXE
7WwBm03k+0SYLgc7N3PNBIM70DjbsmOA+yjCY8Mq82Ohe+Hz33zln/IjOrYf7kSxTOyuw2/xzF17
5hVLThe0cn/WwOsd1HmVH7MsWlBu5u1He6Z3ZAoihAzxbIra6F/Vc10D0q+D+fuM1ealH5hyXODM
X1j3SnwCPUvwGM/ruWuRSBhoxs2k9w+1pHMt6/Xegsw6emlh2Tnamcy5JwNtQfKex6SnSCERSON8
sIqlS2pjs0NTSddnKIsfkECCAnInfqo5U1NMxLgtz3QFA7pUiR+9p7FfFWkmCaj3C1C/SJQB/+Be
7zjgoqzquxH01UXuqh7aZPu0pm2vzlIQ6Cch02R6uEXzsn0QhhT9MSXo6ugKvSEjpXcbApt3CDn4
qB0vXrcnz+m/y+CQxrI9UMQyEHohrb1gM4X5Bl/wGmb9lgOsNEw2vMRiC3so/JemEwBhez5wj+pv
e7wL7jEmZVOFjYpNKPoyXOvaIBs/G7XQPgRQpZOMP/9M18IwNC3JVwJjDNTWZhzgtKtEpgEyMOVS
V2kF0xLlZ88weSjiFEQcKhhpEdI5euF6/MwC0/qckL0khuoq9WFbEIap7TKYUBlgH4MTIWwEBUZn
5T7N2AbJ5cdjKS0kqNwgnGqOcuY3VqBvo6Gm7nztSg3sHbs9cRb4d76CyDaSFcJde5cyRNEhBNgk
NA69Nz1wlU/pohed7lJowXOZDGl5sPPUQXEly5ZvOSgLm6GCWRlzBbOMVXd03Ez7CgJbwlOtYnNE
+x9PUKqYrHgJxoE7iemzIfKHXfYvPpr+gSFThK8ln+e6OYlhLoKEkIeYdTk26rmpsdBq1A6HQAkM
cT6vloeTJfUiGuSMXoSHBV6G0UK3xR8sUBQeyhlwd/K1n2RiqnlcCxatwKDPGONHo4bBPTCRgzYC
drVMu1+VU98im+6YBDlDuuA0ov3tttuyeAtomzNqVqL4e2LTSbo/+UuPRD7zqNY29tcN4OqIgcI/
Ka/kL5dKa+hzu+q+Z0ngFXiJTOi6JnvwClSVaLmYKUq0sIe+MUkKes0nBUjXZBEfKMLus6SWxDG9
6rvoHjBlB0EipMpL/glSs2Jy691OyduucVtsrHZSIT3eONSIV4y3CG2s2Y0G7jMLPYyJZUKJUTTc
SBUdhz6E+9vRU5fa4Bc1NPxM3tq3MPjiTE8Nc1w+6Gi1GOdEglk4o7FAmUkEOlsWU+3J9Ouz9Rp7
Y2ox1npV5JHNkuEInIwSuiAFrT+devFy6oHCZi3BT/qE4HIZUj38HgnANNZwNDAliUUyPkl8injg
KvhTeJWlkUuwtno0Nt3X/jpqm7ZoPD7DhvUCL+JDk0/amFQK/8F/jszIFyy4vzmZ2SkrgRg4++68
ErkjZX4S/1ylY8d5OCkPSUNOnWPbQDffpCRaMdp8lRKsZvuUumdbdB/UDlig8TlE6KbAlsa6cU3W
ji3/U+hCwLwx0pFNQjfDWaFdLXydeC0edkpFesxs5EPBgjbB9plquhmiAcT5+qdaWoTNkFC/T3E+
BM+XiO6h7SdK6dfJjMnJXbmGVkPyXUAldDLkTxYo3armSgcb7U8m/oVK9tztClWF0n0V6xQOpZoc
/O+sj+oSqYBLYn9tuLzEGbMiyu0gy6uxcN0FYtF+uNC6q/WBsHxa0xW1AKa0vzRy09xs2xNUSa3j
jlTVXtO8fowkjBOLGfA6Z1+BKcJ5sef3+krXz4gm/mblqgnRfLbb7HnpbYAodz2xPrySOYH0m8dy
xkk/uMPGmqDaeIK07Nz7s8/GD0m7D/XpRXcBKf8Efh0VBHmQkg+dW32P45R/+NWY4HUGXTaLZeS2
Om1w/AGVfxwcBpFMuDjttlxcq3EoXWxNSTPPVny0gbAbnZpCPIvwt8gjbrcF+AIo6NxkGcp9io5l
jqgkH/bYTYWFnJaZ4qZ8IcWGH1+rmads5N/e74sZlxZ1B9SS1Rni6sVewctky1rs5QFvnLgu/+9h
9wP4kMn3ktprc9QY3VSKOeHAMD2G90VJwZS643GesWBvkvYYW+pwJcaZvtkJBlBVqsipjbSq3Eqw
STo4s5S/IOc70ZTBRdhu3lB+N6qd7ckN6ZAfOq+T7O+6rknEKIdt9N5cxQQUA8RxIRRBML4es6/K
jrkqg2WTJ6m4UC9Ddjuooax1PAmNAt1L721JTvJjsfvyP7UKHeYSsxYl8Zeh4Ldy4nETmgr3voIo
dZoxGiEIktQBODlWTM84ndvvLVfWtP4CECIBOHjWLglQsczfKbzoGRvjctS2EaTI2HGtD3lHYpDl
e/LWSdxR3YLhB69wUseLcqEffAfDVff8FEAPbQHv+Co58BNIBeJpBsKE62iG6/YSPrwZ95qv5/pA
UTC/y5UMhgOWQcjmOzl6BrIWYQRAdrwVF6d1c8+efpg+jz/fhpC8/vIRKPTDpAIPJMRsUiK57net
IghjWHPG17ha4GFk5IoFJSVgaDXk03yQBOwTe1fqgPbSi36lUQkyUdMZd36ABf/hMnMVp0MFxMLJ
XCjcAFTJ3PizxM2jHcK51TExCOq2UCs7J0s1Lgiau9RpSrNSo8NlH3SCNbMHHS+xAOuzkSXHzAu7
Uu4ZQBZfHUpkf2b0j+28o+HocrP4T+lABmdTopv33GdINkOMi4ntH53NwD9k7gwCq5oE6I5sghSi
5ZvTcW+MZN9XYRtGhHR/FcFiR/n79Gde7slvvP7pwa7wg2G00kwgRUCV6v2CtOeFf2CyLc6sWuuh
RZFtjmNAI8wOEdvONsOcwDxdq0ucKkpZGGtMZPmOK9R9zqEPf1aiVq7b9nD7M0AtkpBHpJ3iOItz
iG7W3A2eEmCMJ/jZvJQsS/YGKOVKWNAPnYgVvzEmgzWHQ0ljkZrGdBfc1wG9va+x58FtVnvlLER1
NE5hQcY2ytaxb8RdJSqIHsuT+k6JEIRfAaD6NskOaOKoMT6LmYJOBhqXGPDlE0IM8DXzw12JR634
A8YPjp4PfqWs/JfxYUtJA8OzzMbw8Poh8zby8T0g1GJPXdY/t5DQjPMNVSk8mThuGEEkYccbc6KO
hLV1AsvD18JeFnUDO77IEpuIA6b0p48dk318EwOki6dMnwKPjYX5lfcDoPbdWD04jdtQDEk7f+gu
z91P+bzVQeK0m+JooALPIx1IEEUazYuKoEd8zpzvYrSuRp9g72BXpSiZoH/MOSw0S+QZxyvWOljL
G1jXUmS5ZU0vS/zsnhPLCpEiiLtF6JmklGaG0u/xht3u1JOUcIRt9hp4ONlA8A+wkYzCo0z2MW+C
+V8CfrLRKX72C7VmkGrYRkgskD344BFQOIbckhfqzNhZs+UupBK6A5wRcLfmnI0YuU+4nDfa5QUb
lNGXScLvfKeYxNE6TWCBq/s1MkictIcu4ASgx2FzHm4zvkYsuQVoIn2fYxpi30Wh36302XaIM5zW
mdQ4XUZFT4tirxy5bdqDlr8YfXCHTtw8LD5O/cjwWXrT5US7fkIO4wkGAki5ivJS1ArTL4m2u1aU
uIb9RxwypjZ/gdjf8ZAnIGiFF0CEH5IW+zqMVhxihfeE0FT/HN9B03L4csJ6435K0LigEQXLFyPK
SPO4HSExloxtBO4jJzByqzvkVLd1GT5txRoSCh3OGgLhogsmaGG8W43s+iPl4jlTe3UJdnaffjBF
LyqKFTzSoHpEcuTAos6XZarmdc/I5wU5Mwq/IBcaNaHfQyI1qlT2mrWDd3DKmMd1CJFlTWw3fDvl
ZBvODmIw/MBY0v0LSKt2VFUMb1VUVjEBONPTlwefIW3tdmNpMOFlF60CyywNRxk6eNnLiZeOD5ZG
zy2nRvCAvnhMoXNxcUErIOpT57qWknYmT9LioLB2WM8uJi2cEIQKWWM1/JogCR2YivOUVwKqDvmZ
eu170cK0MqVRGsf506GEmgJddbL5gsJE7JbqcBUqQXP8bpq4+gZMuiNGEzak2uC0VEa0lkjK/i45
OO/WEEcwkVjJIzBqrlSPRTINqiq7/oU17y6WiQkcA74AEPc78eGIE19WzwfiljkIxnEaKH6ysYFj
uItKoggM/OWoSozz5nKlTI53XwEABBS0jCmGiXRl+E3zZuZJ2n1C6zfkSKIBuJfvlPpbUzYz2IRO
UjoYc5LQHIor5LRM3ucFAx9nffefNs6OsHHD4dp4srduY0guZg7LiJOdbkpLTGBiEefT4DE3SRJK
pK6SYzXB4o0RCDEmcC8EXycVC7Xi4gdNylfuCFBp+uXE8MkSMVXYXYY2OEZbujONwJvsZevqclYr
Ajsn5DNmdtOhF6SgonVTe22lqgey3okXGgxvJPJwNCV0CWVTI9e9BDIGKfVSjoE/+79YPrr3J/cO
Wn9P8iNHpsYJizkv/SNWx0U2QEM/oUUeGWjoDOJRn4eULCBPPnXMFJoDdTVvYFgchxJIRxLSTfeA
gp3aujA1pKBPpCuI2eqd3MtRb4uYu8EIvkumLkjpczqoHFQh270SIH2djiJ6xO7mfuQQPhBOtQQc
nPx7ymUbjp0l+pycHjrEWzfHajUeYspMJ+zGCKpIZ70Muiw/RoWs9vJ5UAxar7GuJ2CmjL/Ce9XO
9AK4dQ4ClVKUzY1sNvydJ4S/BKz+C6hS19unkupzECu8AIHjYmDOayCeNtTXIu6JXbPwFgLSSdLc
5V2oLcdKmWccwjx3JJ7PjXkwhqEoD/GPxRnl9nnrFt03pSG/5rf7o+O4oN0Cn0vLRomSGyGmdfO/
g+Czzc/9g4BeZlNHh7q80LL86IBC3BdtZlRug5N5z/qlMfqea11VW0uvz8+rg+VOIzf9vntrc79K
kKthY9Wc8dbKe8YFQAjmkSnGu9a/5Er6YHpmjgc8iXTG/pJsBuj+JYrHEWzebLCK8xAzPKsNGeRi
NPv2ZrkFTlSgrWIVoL33IhHCJYKpNRJZbrL8p79CS0BqRj/ntOOrZiOGVmq4fbNtrejYj8SGSwR5
O2aPrFXJlLnJzOpiRgjzs/K4xSuJ0Vw/LVGsSFzMJKdryse96JAJhwVXQIIasjJYaEHx2/U1C7io
gML3d3K28hiWcoC7F2HYSvZ2Gdi0PWsnTMSylRde1s2qvoi3ZjjS9enUTTCMb8cqJBrIOCK9/WcC
Clx3089EA33WnAR2TVpZAABEjYUVBLqX6njEIpFnaZUT10p9uhLEsJ6EQjIJ67+moxC01Rr/g2YU
QsHCu0sNNETtMedW/k5rgdu8r3yHX/HoQWDpqQenuyxJvxPQFAv+zf53MNeQfXe3OGVAlVI1J1Ya
+sy7rfVWDMcsKo2eWPpLQ1C6JnCDHEbaHDMzNd84bx8IvbAdQJ4VikaQjXqQ2DP0Q2UyYRfzRuHX
u1tBuH+In0M+2R7y4u4lx3ObOLkInxbe+3RsbA7RkhZ/g2L4a5R6Yyy/BPzgS07WUWG/+5sCVtTt
qreISgXht5VKnLnJgDcNgxxj/YYxlVEDkylKHsjORhHx40OudWfKPxqnae9TNRmWKqdNdBdrzg3e
SjJwFNSINkmXPzBjqL3JD+X9DCSAwdyS+ojoDW0aDs7oep7l+zAm8n7IHwql6t+mza5gKH4+d4rL
ToAKz4C2QqdrF+cn9FRuVLLj2g0nvPDQSM5E/AtjutIIX0Q8x8z6ACJ5LsoA1MvwxRt1/1mNx7o5
7YYFBphdkIlRtKai/rCq4qn4b+DdPnoHsqu8FAvDX9xLJfbKP2Wi0VeNVXibVlZTnb+pd+ED/PEI
+ezT9L8yZ9BEkqRIFOpIDYdewgUV3Kp7HDZS0dA8X4no54rSFa3aW4BveosnfaQZvwUywdEIJqEn
kObbOLP6qy9lHBQ0I2DkXNv66l+0MJRstdhNWW+IMiWo5QelAA1K4jlqUvLe7i/nstDLR+O80Wsc
mP8h324W/AC3XtFiiIFYPX2f3e3LJuExXU4UNAJh1wTtXRJlp9OfG+6FJdGbP/JMa/IG4GjVuzwn
cfN6wrDva9s0OlFTTfmNFcrX4DbeJTmNzWTT2kgtky3+pCfeOwnq0KNvBS4dE5tapTmLoydTIOEl
ggINRBTqztQJoYhaAkzrLIzNODANtsFGZA+VnYi4qd+LnaFl6be0AdFpADdsyOSutFxiBWDG6RXn
rUBhTdcb5+e3to5fF4HnVcwSVD3zG2Np3oeN5LiEV9kC4fXA0PgF/juKK3Tnj8aFa2+55mLKQoGY
JV4yMRzNM5iTwGGCfsat/3dGHji54QcVS4ldyaumMEq60UtYT+coiYBhfrcRdeeTkgvC0Xul3xyE
D896mt5Iz/bZ2C5cPNsjPtLSB1aRgTytVFdKiTRnGAQPDp60cjjY6P2WJBq+G2c9jHbNClYaiX+7
B66eNcN7GUpneZOEHNCixhWALB92/Likwa5vl4b1NLYMoFMlMTG6XJptLztXpXn2rnQ2DAC5pE6H
Do0FcmpHgARi8UaEKDFwOotF9bxd1lzLAAZIC2MLnWONQZq6P3pNmFBtpmbUn4uGcJ6Pvbe7wgaD
6a9dyu58ohqVnotCi9TgHZSjqNHCQVXPrT/IpMkkAgNNH+fO5Bvh/8SNNZRDyLw4CfmVwXji7LID
Ls5W1a1RP1hzQeY22FYSW6U9tUEZ/FMf9yQtVwnJZVcUjrFJMpWJdLqMAxDw9yU5Lmv4oz7n5R7I
ZN8Hx/1oDs6fZ2seHuPlH0/vyl6JzrmnPC5fzvNjsvPzJ+Ck105I6zJ4J1GStvAN6TTRi9lZ03aN
OsLoi1KpX09Qe95/qA0wk4spISewpDwgp4NfLC71k0efWyW6nmHrVKblF5c2S+svln8T1N+QGjHz
1yaPogu/i69JO5fnOq/HfDlskX4PZRMPibQnRTUPVNgKrKt4W4Z0844hrbwe2VDFm3d/anzjqz7W
rr4uwrwVoJm3QXsF845L0CUbsh6BIDM1y0FiMxkFDeVGJRAHsxFJh9amtHLCd/RnMTdWVpHBGGkE
6NYiJoql/AJ26RarSUjDIsvEmNvQJtXYs1+giiiE5P+5wwTcbo5zc7GD4ddPIWy8ZL/4BnrJ15Kn
5P/zVEoSY1krVY6nZunGICise3bx49MGpt7igRTD7+rr8gsjTN8jrO/kzj63E8mAVeOhEjKIXMcQ
OynyibhSBN6jJApU6jAziwTzoG72hG5ndVYY4aEnfCoeO3WDBpBAj7Ve68/rAM95gx26JxMW6f5t
v5no/Bp0ir+76rK35AzMGq3scNyQNldsAZe60z0t7KW94WGPCC9QTjzgu3ze3fPZJRgjBCrl+XH2
gHEY67HUSWcJ4xylSbwF4eziwsn81BPBrboyZiZb+s796p/nORjbyH4AYZHyEy3gQVmuh5YgBBLV
7rwHWp4nH44Q+FxNgQ8nl0TdNB9zdEhBz7YPOp+rDTTXTVguptS7ttZVXpVZpM24yPNwlaXjxrM3
hUrVAY9nQ+J6U+TWsigPGBkQFwZ8cFyirk9OIzqn03nc0SKYxI2XIiX53h+4MyuECc6EE5TbrzYp
H73rWgfIEdaHfoUNU76CfWM2rDWXIDAl5tnGLeRIaVYl55e3B9HDzDrmZa8kKWtGkEpmqtczWn1n
Iz4qexdJ8SGK3cHPqvUzrfhYAfcVfzDGfNyOEbUC+X1zia3m2K+dxplcrgiPYTQRPuUaVEo/kNwh
99LEtzG7OiN9M1vuIMTTFWPAC3j6UnwAJCkc38irXYjnFsat6nXJp2OBreKc+84ec97VOeVk34ir
MjzAnOY60Rj+uxS1YX+huetjour/zBHByc3Rg+cY2reRCtB2xbp78TJEtc5Bp/xOdTPGIZrY2olr
A1ha2eVQsUFAjAjVwKh4iKR4rHKcccCzb7pL3EoEqH5in6X4Nj/pF277zSfVkSbUIEn7r7Mi1/oH
7a0L8ktA/rY9k2e60lkg77uJ6mwOTwZkC+H0tPo2inb4P80/Rf0aAow9WhWxg5i7y2P2gns68Q4d
yr6mR+U2z7sJTpSYJLBcvfulxVmGUlNScwbG/08rkzN/E6RJ96UmYAfIJSBOyQrPxGHln/m6Xuqa
zvOL/yF13/X4s7eIpvxGE+oiLjTU3rrhNF6dtGgSYtRhMjt3vh0866dQb87phCrOgc+PEOv4vOSb
F6saP4xhiAy5WGoyC4QWVAljrpKAAX51qVru/Qb+x0Np313Fgt8lR3urY1scXCnQ90msiJcLxw9t
KUNo6r4KC0Trt1q42gMAJrMilylWUy7Pa6QNueO3vBWC8UzPk6uPjWvfbg7qXtw/FTl9+oPEzvkn
g3/JhC99UJaKgADIEzsPCIJ+43gNRJjTx+HzrvK7s9lsp8tx+hkfmVDOs82U8Oxo8lqy4l6hKZPT
leEc4/9llGn3GYLBxc9BRzGLq8+QIJVKwfdgQ4M0F1u7HYM0kxATN+HFIVNvAs6baZwpy35ltTX5
8c/C8MN/IQeg7w27o8t+eOFK2zrxxRRnnyBxFyxxmkzW9kiIDujdRw6mytVSwJNPrHNZGpkEi1aT
Er+h6kuTFuLnVXKImdNvCY8Cudbbe/QUcpSfeEMF54AN/AIpMyBpwn6li5U/yl9wOglUEVanAcIG
BRMCxJOjK+CJtkPA7ZU92x8QNb8lYa00+0Zu0Y37tIgoEKUvxIZJM4sphR3svhps9NENQJX+Un1i
phRN/uE3wAg+lD6BWR97N2hctXAStXN7qicaMhbyIjyg69g3T+nAHm0/4o/ZJ+LCBilVpNWYjbQV
ySAn40RiCwylBmf1q74VH2HBT9EeUyyPeriLSJbbwu92hl49YE/CMVdKFZx/2ECyEgMaLCJjYJLF
x4/MyvRrVVAv9yPtZ+ZuE6HVs+HNSCOY6050WjdxRYYrNful2CehvM5WDLufFVaADNmlbGMQu11b
3rUZpl4MO2kctUimtYyCdW5U4OxMXHKBks8sztXR95QXOzUsuFMIiMR+r/Qh9E/tiMp4AbBh7q96
S/IsuSKeW17lmuFkiCUUEGIdBDKi27I38yp9Nv2dnHYqkblD8UtqTi18TDrUSv8rxvz0UZDX+eUJ
g9G0n4vryn/sWFPZjRzysXCiRQLTOML8P8UTH1wqa80Q96w8JgsCZDnKyPZEHcLEmMdO473s01Zr
FeV/qlwCKz8M7lU6sEIb8VCm8kALYVO5a13lSL9FrIT81DeGN1N7cMpGu+ULny1RbuEi0hd/PSkO
qWPB87spDpu2/FoMJtwuD8NSumJMcLWQR5YoijULhRMJZgrHYpdhJlbN679j4Ibxk8zXuYYshsSB
8sMtWnr/SHF20x5wAW8Au53Ge5mPz8Gkt89943iLaVkjVYhqxroDzPCO1FHgnvnjtDkq+WnaoHV3
ecZW9JNejT6lPEktV3+44Cybn1JSGV1EFt1OErUbHfxh7qK8xPs5aCPt2CMcJMZnoJvAzsZ+pVJ3
JXWXz4zvttlCs5UnqjEpWjUwNeVaIE6kikA7A/Cu3k7MPvKcW/YhGORbQPOpKQlDoZch9K9HUxCO
U4pVVkWF0DhVEa5UW4YIgBp64fpqZrAOSgPqMz2NIccLw6mN3g1rNQbKRVOWPkbGcYZ/myj3daBI
hs+MeuHeY3VXmWBhFCyZemKHJnn1/GFxjrKaWsGVFlKvyrAHiUXiVSKj18DK3JOj75nCWDb5pkfm
abwKiMEDPxjYB3mLgFNZoTQ0u/8AEmJnlBkBnrBMicwY9FS2H6muW5KeDZbhqdTsn130EEnj/X9d
fuhm9Nh5f0zzDsnbTx5ivAHpX0M+5Ks0TTATMT76sjXMNDBlSpR4OEWO7y6kl0Yk+FJUqSWe0HGl
JOyyRVMRf1RKEBgzbRQyLdm9axXLQ0EfRqtwASXYZZtoX027B4p2FOtbu0owofwm0JaroocIOGKu
3bDbDhYLz4/2N6+hYm6npK/TVymcxf87pAGP380IZtffdjwRJ7j4In1pY3KfsuOzweaB3K3YvwAw
2L3/D8jDZnj2iag5fUl4sjPS7sBNHz3SOcFAnP9EE552EJEEp/PRTyrrkeMCoV8X1y+ezEBHNbdU
U4a+axBZRX68AJv/TEtfwZN4Js0oBvam9KF5q4E1PI/Y129bh6vSgeMGyrfcCjMVP/I6WOG/kz2M
C3qrgclTX5v0HOdNC1MPaCzc+daKqb8cwh/GPnOrezvjuDA+kuyMnvEAtI+C5CDsDvOCYPKf/Nwv
hmCkrYCT9We1IMeQlGgxk3mshOuIu2FjM3rtwi9TjaGrbASpoUMBgTxVoNEF4W9s9XGp4Ki4sOqx
pZ1vQPE+amMwgtGuazMwJC65MTkh1Ci9gHo8mGI/Jc2Mb4bDt6OaD0pKhQfkCdA1LE3qXz8dAk37
3E/nqcJR0JCO8q3IBCswcomWJDdO7OVYvfAeijxemdrSxXQIKziHhY2taXOZVm+mUHFXpJ7B0yhU
zP0nbsQfvk6iuH2EscR+CZbFpMQBP01n+rwme9VXcRzJXYoIc8EQwySpzXd3AIT3YT9WRcLrPAue
OA0SrtKeHTfrs3VbQ/OSxCC4jVLiXEw2cz8HFv4+BWCFVLGBAcLNRK9omGuoQ3qRs1PAXg+wM7TU
R7RJB3tMn545K45EJAmH6uVogxInBAeeGvLB5scDxHd1Sg+7iNAQRM4CfvwXBTby9zQSmsqxnyNG
NGLEJ0v/G10lu0SUFnHPISZKKZQypj4Tf/3gAqfhN9gRDIKGmkI8leWyDHFzhiJ7Z+I3qpqKsTZ+
StOT8FsPLS7KfxlCZuxK38n9vz23iOZrmFPlOL/XsfAoTgNO/ydT3qPbJrZU/89DTb8KoDXwjgLT
fCwQeLav3Fjr3SP1uy3SVVqMB69Ix1dRt+8ZjWy3OE2ukQ5budsefri9JHvyAze51CBck7V8HXs3
WcgpDQ486njyDip8qoPTTsuCl0xUQDNPK/RXcenBeVdBXuHSdvwwL2JhlvRWZ4qa3xijti7WI2Nx
x00OLudFjYgdq/Vd4RQO9Y6j8PcuLEWyLadg/QcZrFsOcgrMI3kIvLB30g5fkz+kaDmP5TQ2a57v
6bG/4I3vs3txBJ+isUrPXnf2eIeQ6nJ/JBPIykWsC/KEvPbLMAp/VPCgg5H0dw/TpCLNALIRlcfO
nFLTI3m48xkP3b8OExJtmZpEBAwkJfCtPy6P4O9anTKwRWnDgrNnjOjzdAuHr3a+ZCJcI3S1Dl0w
98LD/diMi3CHqZYeY2US41bTLjTUA+m/yBpg/FjpgFgH2lRsYH8rfmhO3AA5T5q3ZMYNSD7NWw7U
uRTZGnjJRXcwSaBrcCjVQHI6MFQWhVKgClooB1xDdziTC1QaTNZF7XVVFzWU5nSivw2NnEzFsrxN
3gfjESiXRxukEPedEDTve9DpEuWSt07qk+4C1KQRDt9NxWepVqqWdRpn0D9scw2o0ZRQVNNCtqYn
jXEnXm6CVuhh+t5U8VrcD4N7Gjcc9bNt3JmqlqQigfWa1WPkl4CzAUyIK0ITtpzvVAFZyibU5ybf
GUF7pP6NMQfNt2udLYSbrdoOQaLJ9Y+xgCgH/rsxcMWqBGfsc/sk7w/NXLayjBGKZMPG8jr4OyFe
rSWpOOMEyDhRNzMMfSqikUAnfE/iZD/ppofe4Yth5epSjsxwqjewN87wCp0ZlpL5KffQIPH4gQdj
MN3QOUZlWhPaM/UeftpJjDnp8HOaUHQkxi03+P9pwzYU0fakkqUIaURGuhwkxjzsLrap6lsMFEZ8
RwjiMyNhBP55rSX6zLsz4HwF74aRVL0IjlT6u/yezvs/IGtaBSpu7FlmSjXOM2rtSnUAWF+KN3md
+bvbm307yc2B0S+4asbepwwl/OJFAwFjkPWv5uh5qzkTvEtHeTMias5QxP+wimlptyHmJ/glyTBx
023cbsGFyViCblg9xErm0PWQi1QbmT5ZjNVpNTeFJb1dBPhwYMc0L1LWZjARkN+c9/+X9BVJ+QRV
dhbtoHzy7/EjgT4oRXBu2uoaOdezIAZrH7v3Pf40buSPMz/JCKDUTR/9R/W8woWPVzvkR1y6eLAk
FR1zQR+U4lmfdGQHkJZ2hiAcviCUKpPs8WCP96SWMMG7+iMoD9YNgF7MXTssjvkaXrNFHtvXzYel
xoYKODu43H6hbnD5KCx+R1FYhF4MjxvIAvkkNs1RysK0YygG2ZMXLWxpY/qBZp3Q0HHEyfKFzITI
iK0sgsyoS2KCk2EJyuyr9rBP+MLH2b5BmsxtjNqv2GzxEsKOf7H4Um1sQ0GdW8p7gDUSha6gbTuY
89PZHHN7m8uAcIzGbzqdLlJDUz8ETtPTxRcXTOxdVvEvK0kgvUYOSkDIiZb1j6NhLUyKdrNtBGTn
MAFmqbTq5LoFq4jjyg88bTS36q8Zb971uPalVT7ZE+mAloAqSEPdZyvr0bpTIXfTwsMLtJvCT8nZ
TMptFW15b946K8wQ4xu0+Urp5CFmPVjUXzUlRDauw9OzY3D5TTQGs7bkB8vDfYudgWa3vTs7HJVz
kc+2TEfavdWEBL/K/PBhgzT6UqkPg2ltBxauNO/g6qkGfeJ60gfkO1FMk4mQa5RqLneD24j1qaKP
tI9YWIobC0qUVGCQxxlGu9Msqmz3yyNXq1aVIKdEtjhKOCpsDFSWTgOlBlV//OMdqWvFln9jeXrw
kP9ui1jJEbykZmarTzOOms1OOC+bEUe9vZGudJEIPL7MTpMvkMiOvkUw644PArcvfXirmyDvB9+Y
zDR+FnCypVXXlga4/ONEVbjBUqe3P0TwkVFHF1VbIdkD1IfKDewrj2CAZvaNUPdarKjvt0D7B3DU
FRRFejx0Wjf3om0Fl2mqlW4xaA0sTSOKrclR/kOGCOIB5JBjlb17McY0/bzeZ4lcxyB0HtcYiruK
jwDCqTcnF+Dz6gI+azPUpCYkUoHkqWzSXctZNtF6X9yvBICmh24Roc9zB8da+azJqpefpgX8OJVs
xjA1OfWvwuQQ1/i2RTekyN3jMncDpp/+gq0RsAo5ZLuQovQJT6WdAt7Y++9FhaZApBVxrnW3wERb
nhZu1Mz/UqkKEusoFQ34fIZNYycyKknS32oCo+nMElnHYqG/lSTNobubw7CE2+rFbeDN4W6w8P9F
K/rtuHc1xINzaBAX4hXCjBiqz+kgx0Co3ue7e1jMNARY0R0xDd2Mp3oH2EjR+hK6k+uAJSUT2r05
J91ElnLwPzsnehOhhyfLv0aFsgA/blLHZD9bq2ZbHYRMF/76pPWovoPhKmzw4VMveWFyDonaKspf
/D9w0ILMIZdXG9Mf/qMSXVbLBnAxiewn2xbqbgBQKzvnPVeJO+EL1fGqOiCD0rvT7W80ajnfvNkT
ZhfMajkcfPcCkCocuO3SFFjr2FCWktg5P8mKaXcS05iWUgeWND6w7MKvB5I6UCgH56NTJrC43nYa
wCf8cBAgUfxqZf6Reo7bORBg5T/rmDSae7Y0MKrdJkHTWoEZQciQJleHhdHzParHOxqCgcoEM04x
KPNCW83ms6JvWMbvDYPym/r97OceL24kV5wiscXz4g99VbhLqapKcRw+DJSTbTveM+G6zp/ZOD6J
7H+gFft+nKHLWM1hXgfzMnk2RsOSLU6bq8pjs3OSCBfsXohRFfDWLkxN6vaxQhmwqgKl2QS14vOD
rF6D5QoQ96lVYG0pChhKsKArUNQ/H8qCYlmu9O7gozKIgH7kxqw+zY6M4t/DjKp4F4c4ifS51nmg
W60uueOmW0qFpf4XQTkDb9qMiCA7Cxo6qtl06LVnbNKhqXXxpVroGMx1+d65viFwzN6EyXg0E8Yw
gQ3ICNStpk/eA0hGUVCmh260xpMj11kel53mUAJq4qIy53+xQNCPVrlOnAzJk9zKVBsD7jU3H60i
OZSMd8J2phifU9nqWlhbxojqPL8bmrNWkDGSk9O3n0UMxFz7Stj+n9nawoqeS5Hn/rIdChJtoL64
47Z5cwuzMcpSKpXGn6Eu1cxDB2O2GmUJBMicBvBkEXF4LitXYQ7rjQE2o4E7WfJLxjKdE2+W97hL
wlEDWnmcFerOhcNx+iHQ/X8ZCBYe6fFgomgHmxzJ/FVP3xefm9EXf/PqDy71onBNIgdq/KgyiHa5
Y8SaXaUduG9rILxA+ZPJdhdvDnG34p7IklpxBFypSWvjEURXvQmuOXNshZC4MUuLbYIKP/WET+Gp
VuDvjO8JDa5SfbkEKBXOzpI0nis8A4xUA7+pReiZKvX/f1YdDoC8C4Qo6v1ZxKuINZJLj6qGWyYN
nGMtzrMeIAje3dUGPUdat2/PMCZjol7gZqwBV5YFQeRf73xoEq6rrOEqtm0MBYAsD8AeDyVHwNbD
9sRbQf8+JlIaf27BGpPIHh24Rgb/JmPUv5t5/VyfKQpwB1Jnf+wbvmzhIFB2muZ5/JfDKIGIGRWB
zV4/ErHdaOFcSpgkUdGzUd/+aK8N1PKh8IWWkFl3DtDPYHSV183dOAjn9s+9SV//Zx7nRiszDgo1
5iopDgwfrxgHyJdKtGc07+nmvg+R/qr3j6Z3/1nzUFI5Sdj28VsmfVd4an+rEffa95mBaLbxMnCo
E/dZVmIGSKt8GFYXb489ryKk5Fy+YEu1ALiH+0EqFg17apoujm5bR6Hq0xcSCrMdJBpggx2ixQdI
GmHGJpuACOo75s0MDt8dCSdrdLZjPGAggeoJmSVZhs6RavqUpXWRl6v4xoWxf/Iya3lMbuLZiDwb
ai1YWh7tGZplNwdI4TXT3W7tXGLXsJhmNFZqGDR/A7eIlLOVplbh+6snhTpiqvG81EpjrTt9mEVq
atdUoi40a1jl1F/t3wE0yCbeKWKGIgTcl6Zb3AWOlPWR99ezd/yqVQZZ9tzMKav4PPblmECYynnP
6nWd/q/c3/7oKxj9X7N5EKJkMD00CjD0RQWZWmw0S9RnaRSR6pLARdSeGxVUj0e+iKwP9uZKAz9t
JBIHpo8jk6x01vUbIUALVABexVPwWgxVu9Gl9hbzKrppToyxdo1IGsLYyRYTLkrx61Cu9XaKfI65
7Mzfd7B6QqZ7W/X///1ZNRTEvjMTKK+MGJP7RRd2SO+0QuC9mZqLtD0g7FI+BmncFAIyTEXEY9Ny
mZqt5sfsw4I7pZr4Xd35CrTj5tlPe6q5784gYUtUKGTQeR3uIobrETecPtKRfSNrpFRH6fA5VWa5
LPYPd1rcCm0tjih2+pru8w5NUxyPiKQPUZNwKGAa+oqPhnWcJlfLe2hJnb5P+ZojCIGpEuQC8CB2
evG6Z2jbl//Yif6X8HU628mSLm+xd3Tr9PsNYkB/ciFqHwYoooVw8bIewQknJ1gjMXvepNt5qw68
auvABCbcVCjnKPPGdz/pyyO5nrDICaLQJI7z+yfrvQO3CTJE/Z1O/vkOGCGLFcYxWfuIQtnvhqRR
x75NxWQgwySh1fpE5yzWdXaVHM9A7iaVy0hDdFxVdSrtD2TPxLeMNR3m+2dSVVYKpAvZjn6yutt1
6oYeQhIcQdA8jzBXKzXLw/TWP7gUnSYWIuvpmp2QZQ39fCVnc9gRIDLBCeAbUuWK0WmpeXuwdwv/
teKxUJT3Nyhr2vJmaskDzyOEzuJ/+xygi7JHSfMNmnZDzpvmlqGYkViZinIbjjAuNTJ630oLj//6
WFCKTRaFcmxZXzHByhyIpTvUmeejcYYAHswV5/iVesoTK3vcI5JBWEZthBEJae8NUW/yHLg9SXGH
FUroWfnWb0ivs7Mt1lCv7kcxMF5T6qvbHVhbnwiA2hWORfDlk1T/62nWpWtAvfxqBlofWBOS7FeK
E0raScwq3a277WxjZ/BJtKuHvDL21Bz4j6zcitWpCX9HwbjwHhC2GZnNAYOdIRNRRYfUft90Lkmc
xV5QZLcnUN6X0C3vKis4NRAWsL3WqAJkFYKWD+dcuYg+P+B8vBuwHsMW3/Xq4KU1Sa/8072IzRH8
tGW9fE0n3t2ZGiIXCM3OMLxCVenBwwn7B7WB3Gg4H2TNyKhruVQzroqtwtY39U9n2eSaASE+ltkZ
HYfusnl30cWdkLvmfsvrIEOKzXLL0t2UoJRppPBaEIwVwcZggeYLMhVgWW1ikkzxOKFkoDSFMNyx
va3zdvY0ZQDLtJDgzOBowwjrj0wgs80pk2Th2Qi3MJW2+1/mwKe82789IrzkD+8/mcdp5gLIVuL6
4HiGSxWqJRWXiKaIf7N6WDQOp9t8vWS/JxWfqfl0z3JxgDcnFxjiNTiMo4IaKAjfz2MtXLil0bol
RY35gEWDrk4tR14N0y5a5sMyD+TV8rAr9k0xS50D+dtjXoXcVaI61YpDu8N1tMAHZ7ifhE9jhmuj
Jcu5wlqh7ieKzZMBxnfqDjGeQEEAvrB4JIWKUqRdb2zFrjymSP8dnpM/XIWFV0lAR8jMzDuHfR2N
S6jJRpkos2gA29mFmmsPW0t9BxNSiiFlFaFhfa1iGkjSOAVJDIfPhGqNT0F5dwKkM66m7Wn386sV
9dBkkXqNqqwuVgkDeEdhRQoddX0+G2Lg9GLSiM4W/FaiSJDvHODa2e4S/Wc89pq2fFY1bTjlCVKt
O9/LYEyFwAG0QTZGfA9hCKKcyA+u/dkca9dQNKaMLGuQCEhA/2Uw38Vlpj2FW4a3uW+ltZghgsLa
Z8GaN5xU7palfCIXhO3JN5Nm+Nq0Fl5a53GrX2sCsdfGd8K0jNaQjAHTGaCXIySCGVfzJYZ0zjzj
at1iNAzVUSwtImRi0xrKykwBLmIm1dxBIt9Zu4OxLqRV9GJ7a5h4AY/d8OvJXYI0vy8PkIl7gDZ3
b6r4CGUTFG9/TRQuCaDng8P+O21C3FPfvwQcgEZZ7z1NCsbT7xXpieyXdzeo4r3YW1pPvelibll6
ZQ5ESw+UhbYl9+mOXYfGX6WCo2fmtDkBaQQp2ILIANDdaxoz9e+ZfZKLr25ASWQKCkYcGbSmhcua
cusBMEe7daFPCKr4c1MxXXtystu4UWpiCEgSWc60Z6ls1+DLsRRD2yION/hOM5bEeoW0OO8uLkol
qM1Dm9vCjZDHfDOW4/H9uQeNg/kcRY50JVv24IzunxGB72Qb0i4DckAh/Le57RPgVat6Gie+8Jxg
KkuFEme0DDLrOJr1cUJDK2PGO95vkpnMJuOM65kf0ojs+kdvRHkFklAJJaFUid4hZZerF/uu2Fn3
TE1+DVvgbpFkpXNgLF30rzm0II5wJdLWHPfp8Rclo/31yt1QfyqfVi+vaXdCei6Z7TF+Cc0svnBB
vuM3GkTaQequaqZUmTu1mEnwcyJmsLlIbsNS62KR/0s++w8Ybu7dOoAqhPIgNVGJCkbDBR5kWv+B
SQAcQUw9+zUYcXk3YiUy7lrbNz4eqjWvnuJDy59fCfddBIJjiYN1410xV+49pnJ2qbFD9AyR/QyK
jmgZQBxhDqK2z7PIuRzJTMwy0+xf0p+aivpG5TsRthvZXgg5xl4W8JtFuCCxBpR9NhtZzBEu/kDk
ue5iUkJn7Gd9GmBSVQR8Jh7tLBgbZuT0aaLDekeIuJ3LDPkeQ9woszMH6EgTtLfxxzwmJqcvEEB8
C7C5b9zmJ193aI37ULsIthUkjBdVmd/LkFdatmN97jTY+6iA9Nm7HKIdR5Lw1nHuHkcBRk/DZxoe
KZqeiOE5ZIKiwMte/HsfTrTbUO2rHvxEa2PEgVilhSCKnyDxzInEWYjt6deYsTJ6urQo+rkWy9ac
+hwKFn4deINEEXYqMM1vN2K95EYuTfF53SBxgBD+KphoSsxLyU66Esq0PIspEVKhR8OiWvX7TQ15
5ETWtZSXDHY7sByg4tGb8rSN1Ozi5diA4kuK8+JBXLmemiA97VvsKs9KFpnisiGq27iAxhduX1hZ
RA3NbpiiM2PpRug/XxPtupdwrCJzHvVVa3KYkO4UOjSYjQMqpdkQL2OixnjxHYchU+rTfJD0tTrM
du0iBcq0HfHEQ4G3dMIx5N6FElQjlpMA6tmDijLtOpmRnQlseLqBiQ3JXjPNz9AEFwG+M5ZzWhnX
Kg88cV856DFm6BIY+Fag+z+laLmJ0xwdKam05IjY+UYiZZ7IXiqDzHk2WIKLpn2+hh2VCw4zo9BO
NC9ZfpvNiRNFZeu77Nd4HopZ1SoOkcmBdyW6q4sKWTJxo58J0t33nBssCaVleFE3OFyRbEHQ7suV
/IXBeHKD+qUA2np2wg49s4O3vDFmBy6mzb4jk22x/sWRx69yBkYBuVr+mOUgED518PCl1FAprO3u
/bIqpmb9Ebb/B1dP/bwjqAkaM4mV0sclg4kYQMHYp+vzX/r18jlLRstMwTAmBjpD2t8lUo3iosDn
0zjqO+5sFpTZRxcLkDLi8Nm7qrPsJhDKXhCcYB1NsxXPpfmgoXhTRdGoeOl1Aw4mXxo/i1VkZbPL
vij2G6f4ICqHJby4sKZUX+UaMyRPhUKoyGL/q3biADyzpJauLIGOSbmkDqgw8pN5RCbcSfMQJWx4
N8O65uO3W7fOfPdo7pnhItcSfQWPX6HGX6f+Fty7SPWNWlcREmIQBd/Z/9V+123I0CyLf2WYd0nK
laCm7Qjm9ZTkf9v8DMr7QQJirnhghFemyZczHOn7q300hHqZkAGBXGiKlMIawGAesaF6nqLgpsl0
c4O2jEi+d4dUbT22MXblPS0oztlNyHwlXFwAZs9j5yLY+BZVPBMvygysHp6tmjRVOnMQnW750ToK
AfpG1lPPtgrGzmVTd3Z8WeNodDIfNnuGh+8EY1AlXUYBomKF4XeUOKS6WtAqfK8hl9URBo3kL2Pw
63ipFTVpehFSwX5sK5VCwK6kTzJIaCRTtctZHwzNw9oN+ww3hzsbAxiy0n4oADihCGaYMI7fAfwM
aUP4rncz4mEq6HAheBhvh5B8njqze8NjUs4I+YmxtMBavqWenu5fVPGiJ+WNKU19SoOg7sL7wxeX
b2B6OGHr+Na73HcHogaqdtuN/3X2UnnLMlKRPAlhoiC7JjhGgN8i3t3BN1WU2jiyp/Im/VvIudd3
xKzQptvDDSXy1j6uazZBey/BYDQZgtf6vIU/m7wGysDkX83EwrtYroDBYnmB8OPyJcvwTxUhorXe
Dg6TOcBRe4ogLEFSVVo1NqG+EIjviXkOBFuA8Xs6j2xYPNh6MAaszx0Dx8urz3fdHLQTAPvJNGAz
jqyTs+9A9ifUR/zjagXzsqsf8SSqmoJa0DMDHaD0MWHjb58ULWHZf28Xpop1OKscONARzs5ry3Fp
C0oP/YAvBLTk1b51n1tSg2EV6LblWQr1Pnfh0oOPgtTU95DsINBK5ZiAQaiQYHykT92PrxqNqUPQ
ZfWhabLDyNI8/fZAHyRtNO1hj7tgAsmd8jyITXELgfbQbavAtmVDUYqyFoEKl5WQ25meSN51fAel
RZmHgmVt9LIQzK2XNC5pA9MUn8k2S39adxQgkaX43fG/muFFj2TBPcHuUWWOTLKOxUp8VoAglDeA
wYWSOgGo1MtsFDkNAO9xMf8GFxUHDyR7YMQV0Fd4aTbw7HkAUcimn2/B+peqc0F5qJHpqqhthKRP
AS0AG0ehyniy5Bxi5xdyetLNN7SyB5aJyD9888hrLeGa7+wb48bstDlOaPIX1pTIRetyyhdDP9gl
7ZCNQLV6WKtu0qzyr8pavpdHiB8EdrubLFS7KNQIt3/a8S1+YQTx6Tv3qhM3fuvR9G9KG3QBPw82
veXxfsDhAYeEonYDlUkUd05eprYz0cHnFlfCVCgNVzQI/kJi0UOmpCFDvyLedLBupIt6uuvcR1Ea
r4JJlmXMonp2UVEzzBk1qZG20sD+PBC+sWk3Vg0z+LOpYSlQ/mvxCSVk8Vhazo7upU9X0RcZ6Lqd
hylc069AJn3FskatoSLqY9PoX6UH69NZiZXRP4BBqSodxR62Gl6wq5pkAbdelmfjKxwEGkY0Lplw
ArUwaG+CGvnRxQbRiRXCEPTTvpBpaXy0hQ6LeWMyAXwM6OqVEiLKIukyzRo6yypX6T/IMOVQPVz3
YnhrSDiNttMY3uh2DGeR5d/dPKPSy0PU5D+05Qgt0iH2acAbZD924e9WJo7y+MO4qI8UrLi7bTfo
7Q3eg6wl/ZUkiXpS+i9bsQCAsUFEWfoN9pS1pTtwJcrv6Zg5An9NBPWCS3yzGyvnCazEhfmQiwyi
7sWxawoaCZKOmr1yUt4f0rumTlWdE0YGwiiFCAQHXrLi7WFvTXEFv7eIU65vrCiLD4+2R0d3+kyV
NTWyk0QKZBISCpTzFTfTkzwAg5xGvOS5qJQuzWNdTpwmU5xCo7BhFnJ2un8LdVhU9bIvPjo5DD28
BZyU9LYuk+p8t0VxgDJX28FXPxysj3if8aWl6zgx0CeEJlP43xuAZmPwRbRNqFriIe/jm/qPC93P
4b1gpLNDMMRfB0PhoEV71Xp6TMUHNDMhy1isvQk2AV+jdPSI5EU56cBCvL8vaoESCUOuOAO7jQ2n
rmib+XVLMe4S2wAkvuBWy2WWqX0Zms92iAmTJucKueHV5ROYwSjUIRXfL2FWoHILGghgDxhCU8iE
9n0oET9QX5WwMbAPkDIZAvlbs47Z9buRBr/7aNPEk2EPGKB/HsmvG4Eg8riaxANpdflmUjJdIJRL
zJKYvclGHjNbQ10vufwf/KsroiEHa7vQFpg52VKVLseQWbZS5p5XkMA7YTsyvX8T1IXUAXNHeu/n
4TnU/SX7GOijJzqBJwuD8VNzlHEZUNeyb94Opi2YNy393rO8v18zzcBd/1Fjp0fO5/5PGf6DiBjE
bg7rw1VF6zevoQPCj8Y3tIrMX72Zg63GVVlNu1QH3ghMc4MkBZKY+jHFFabHswPClnSlQRCPh5M4
UeeHyApnoPN6RZ59kU7TsmL1Z+rdgOER7/ZIEDtpJsedBU33dWaH3YFGkq+df/YReb7A5uPUS76f
P1M5pLCq18D+7TiKl3Uq1Cr2j5cyC5MF4h02RtPEfkU9yy+QbMKWJgyWwJQXPjnMkSnUvoSWWAnU
kfx3RyyRzVRjd6Pk5vJlwzzDyw4FdV22Q5p8ETEbEP4nAXz6WFCxoDC30ZsPuMAh236y2K7vhb1Y
XbVEnd2L01wtHAwZlJuF0UQ6FpKq78O7T4YDdIsn1yD7gd7NZLs03FgNYQRLj67yIVK0gdZYM1dg
ZZCtHKDLj8ooprExqwr9bVmOMi9jCktGHMcmflE0j+P7jthGANlOESdWyRI+d1G7JGeMfXZtWofC
Shypdaoz5Erm8PbXSTR94VaPTtLc3K6QDhEOdcZ/VSlYb5N7TI+V8EHc2hc3bXrxWsR8JZ2Xm/MF
NBRF0mUbiE9ZxsTqT8QEiRGbfK5dBfiKB5JqEj/MthXzovtvUNwcTkLvFRRjq+3oHI1o2exCZ3uL
vfOjOPoX5j/W51Svsi8V5LVS6heu1s6eotInkdvVt+qjMxOUpvynNFfx8CPM6Gn5O6ltcO4Evtqu
bAhMRHeX5AVZb2ujQKDKAExJQQ6bSCu84EFcn0ttJlN9zrhPUr2pJPiwhtQygZ/88X4zgkbAaXnj
FsDabm2SD1eX2/RboqBt+JOKcGOKnUJkIEuhtjU046hg/YXTho8HgPvgzcKF9qn1mJzfRJ/z4tv6
qjyu/T2dc80HpplsnkJto4EUjpLWtcPEagxMBbapb4BdeJcBI+KSD/vScEo+Yin8Ts634cfGwvGJ
GryExVcmjmDCCVr+lrWHXD3UtrE+IMNULm51zKV/CVuObwGYdYW8VPhrM8iARCKWBSsnUDfCKoWU
0wjqTNwC4Na9FM8dIZjnIpNuzbiXbwjt8px30IhBupC0A6A1jzOah3LcP8sxw7OdJ4uTS0wAB5Nz
nWxhGalzfNYBVmPrwXC4LSo/t6PGdvVBPz3A0UcM6s+DRSmKGp7fKU/4QihEDa1OmmKXNTq1nntZ
pBwzfEQmOsAZVIjES8oLMwP/iJHEVOtvuCqCE3dXiybYgAB+gWpAwziv0uvvHOfhCH/O8wStud7D
WSw/NMp966MkHAXkE5pW3BJs452SDGykUx6dRDFLsl9BUogCOBwJ4tm8L+eGjvsWYyBppj5AGx7C
nTWa11xDR9s1aMYwRA8V7WYUtFLM+JpM8qu1vxdZ4M4d269LlsoGCHUIC2CJov4usY0mM0pyagml
vGHiLqZGMszGcIOspyu6YzTX5linwvJJIA3xz0b1p+lVJnPWnZNSsv1tM5KHR2E/V5XTLScRwgC2
VG6MKCLPRp7tfwolBVVOZ3aTsLQUr3FasBKhpYofRv2CfiP6v2qeR1RpiNeAIxCU81W5ePEvcuL1
VdvbOjUZkP+y1tfSPmBBH0Kdslg6B5qHfYsQadilg4Kj//Ez9JnkyNpTWPvCZKJ9rd22S34AidMi
GMSnozo3sL7/exzlOwXVeYotobdkfvKUAhEfCZSmC+O3/mlsGXVOA5T2cDRmhSuwyGuTMakAFQyW
uZoOX6PUo1nr8KBJ+VpE20efwncwRKWJuUmIBIs1+2cn4336PW1k/z8aXhjcVbQR6xPy/v39fJpS
ZhnNfHbDmvbvfhC3QQul5Uq9qz+xaCTRUbhJE2/aYXZn2yCt1jqmxCsKdeD/vgP+429jfzDwvbfp
owhqES4uyr5eMhiW+K721xl8ATDeZiONCR6aWeQniOVdttmf2RDpxLCtgoQmDUE1/2RC42iMrr/t
TbAaRSXBna5cTP6oWJjxqbXueWtK4JjUk70ZAqCSH8PrkzDMPsK53tuTMDK18kUjtZ8DeySvaufV
0EchavqaEoFTd915YpXUKZp8iZRBw2Vzx7O+HFBA5HNr9u6fP6iLMJfnex8QWmAUPtyfO51tTyQO
SRl6WzMg9b0afTY8tOGQ3/wlPlk2j257rWAlHCZXatP+B+9Q18Hc3UbS203kedo9qRg2J80sCtLJ
ojdNYNqAb57m2RQAEvr4uYjC9HFvyG1L2UI1nhVJoYn8oKGkMOTKBKEHNmNhn/qlpbtFeByJJclD
29RKWhdHKjkdklWMgYT4D+8EDpcVhY0nx5XErQoZerMJYSMMwDjai6tXd8YuopjR03PNZwFFTtOn
r+WalSqmiY/FFHCT35GCjO/+n8csWxPEbrQges7BrXmoiII4g351lud+P9bRnIef7dKN83yBWr9V
LDdc4yYeCHtYxhvh6ck/B++hD5w46Xz4aDEvzQu/timRWINZCV/Ea3MMRYACiHBt+36An8vrvDYJ
509Jl5fP/oGXduM2IpHfF5NC0AzVDB2u1r82iOwmbE76KQhhs3cCEZJAq+nxDi7vMOkj4R6nO7Oi
7hMVLp2ZWchD5bJCUeHtPyLNVHylPXpgMd0Mw146w2rpmqyHyU8zIJmqAzsXJlgPVvVlhOhyTW8T
/UFSid6aJsVyZIGGWVbX6Rhna+W8vlJ4XLKNWhBLvpVN4y5twK8wT0/R4Wc64mh1Axx1fU7cLvHJ
o9fEJN2rQ600CE6DKWsMIilViMiruTv70EmIYBHIIybOmwqC9RIgH74SD5Kn9nvHSAW9QU1NaGZ3
6Ca0H9FyNddIw8PAXoz1LchhNOhtNSkq/D/YIxlxO3ltkpMIlH+NZ8kVrNqY8TdvZojGNd6OHnck
kzps3lAgrubb1ZpNtmAmRXLYdT6MSBxM+sHieDiwByqxhxWR6uv39vKUt2iEd7BcLRUsWtXh2Y86
7mPH4qeSQwDV7KnFw/r871qlJj+4l8RQ+SsjImwQ+iRVJXgzOLoS6KdDC07wLJ8s6bT7AM7pf1BQ
nu/K/GMkQY5TuTFdliyBSXlwJ+erK6Qn6Uz1lRAGBAUKuisVklZbppGgrPAHc2oYh1nKiYBrM6AU
W+S671JxPRD2pJv6i2jj5GOtgFHufelQON3GjkjTUIbEcDSdzfYkaIlXHl/UHKd2378Ly6CeS2m1
CBx3b/tKas/6Zym7scCIIUx916xdBsFOAnQ/kXGt/wK3BhKwr8SFvvV+auKbLrtGAh3oy61shzz8
pO6heaLbUDS/s+3ZCB9nlx8+pmbGwIQu4N9/ITOk1Az0GnhuUYZAazX8b44IEeZB75S73afsWopM
qKrJvNnCfETQKHaAth8RhTrn9u7AvRfEHHuDDSv2F5bPHdziEfmCikakSEMdJXm82i3UL3HGczh/
EUNpaaSEo5z9aPePUJEHetfGrpHABcsgBsPyKrvhPZtx7ZQPZHiahIteJKinnlrkFXcg2D2Odfsp
/9i0ZcRlJXVrOBbdhf5DQlhENtQCO1S6pwuW83/pWXOh3SxS5Bflnz4MZTAG/PqMShFhqJ0Cls+i
iqe8cDrP2gqL7hV1HIP0t9zdjd7ywteYoPt9y/sTfQ2ajKvN92PuysR5bGwMz4sAkkSBkkSDPJpp
BMo7SygvsWu8Q3LeKFt+6GqSUKxhuJI7V8o+iJkn4EpPbCWXgSeaANTHvfJlTMQcfahwHCWmqAkY
vWBEADc5MOWDmqnhSCo3BkoKIO8s6Q1Iev1yfkymaZ+LcG1Zmyu0jZPIxhrb6/WgA6QjJD1OFux6
Vhrljg2bQzQ3uI2FRHtXUgY7GuIA8FhmwiDG8ANlYEx7+7ER3c050BPBGNXuyxVzqIQEttvgw98q
b+xdtBcTuIA1LaShQlw+m8sTv8qIKKJoY3FRr2hx99b8/yOl59/zFxihF0XxH3EeEUBLxuz5xNQJ
xXYKeSBaXqE+m1nWOQOUet5U06qRDPgHiHG0qtRIJ1WSKLhhTezSoItMWQDJ21XfPUvHiaw5sV/U
SJfZiciQpKyg2Tk63pONEY1CclpQGNGhWB7YaaRjtDncfdydRmNztn5iN2oZ/L4dICWv752fIH6W
SEaa1BByv64zKLO4L/FRw9qUzDQW9hgvgLPc5R6vYFoWvOEeltjs2xXh3FP+k+z/Y1zrvxRC3U5L
oligdV6cI2IYShcJWllYFXN/TbOjvHfLqCql/6J2/bQV25d+duSUqvW86slly/6Su9slVjfhCcYG
FPtsN6ILMqdUehrWP0liRsHSd8TnsiJo9Agl8rnJkHCSKk34nVKXC4DLmHio4bJsNqMH4v6OK4Qf
2Idwcoagoy8SXg2VGy9MXvYmu3OmM+Scx/R3n4FJ1MW0KTtDVzK6+fcK5KBAeIiy2r9Xp8ZNI0iR
7i6FBT8iYX0bK163nThxuUoPDt8J7gUow0w+uAbf8fRJ861PB6wA1l0TvcthgiuHt8SShetGm01P
bA1WXS0qgoP/p4h0VCJdkx6Io4mSfawpN0k7E9wUlRCYBtAbM+t6FPTRj5D8yiikB/B/WclRkcms
ukeOLiAvlTQuMK18HeE+JfdrR8SmkYWBbJPEYJ7UQZsnmDcH2uyHoYTy+dv7c4qRDJxKvtOMEiCk
b8pHp88+Ma414Som+e2ooRUqU3RLwGOVSDiUL1r1hnSNL+Sd/ESNQIXklCSK6I4jP+fzqJY+u643
gHLdtaG3wcnMeuLcmUb0Xe9VLnt92hBgbeA9ixTXfw5El1M2f5hHJFVcD/I5jc0DrPOi4ZqowiQi
yCtJg9CCmxiEXcJ37IVQAqrNyQtGUeaI+ZHZL3HPcTBtzAly7MYzTlCU1VGbFlH2SkH2SkwJfcJ/
SUsDOCPfwfne8MJUfx15iHGjnM22AyP/wVm/dkydJPTwU5E6f6yPguGp95wbQewPVd/AABmCpfIY
nwMVX5Y2xP85+n1tY1bRgX2FoLKyVJkEwBlLtq8rXT560PBYJ8T68fwzQfjsq3fFiJzs3IbpRKo4
XtqsTFglFw8XUgw6/yjlkSDOuE3BGSfQQ9Ey54oPrALmO/BLricUg5STGV/y1hHtLern4/eFT7EE
O8LfOAyFD9DFpMtZN/U7uJnwl3glrjAOAxmMPvm4OjyaNC66W99ChZbldvvxDRqJ0/3nT+9TJOYz
D+k1gnd1JmqCAz6bulKw3znWISgfizu4B2MdQ2ZiLeraSOCq1gj4YLp5Ix2UiiHSBnV2ROggZznY
JJp+BkG8u8C4ViIumvfSYYFFh3OmG4IrDZRmyF9lrPxYtrXnkqk+9VNCW/89Azcr8eIcGmBPkZz8
uYgDwz72KoIroVhiq2ll7dXdJ3J3V8RY1BHmGzgCKcDmtxeghESASczrg2666HQVO5V1Q+bo/WQ3
j16sUxT4KER9dsP41oKJtsAlKbXaq1cIykFaE9NxHMyw5DZx4pSG/bfPX/Bu+cfrpOBKBPMTcjJ/
W3pPyu80tCRh6i8qza1bbNIwPb7zNlnZ2SEduUEKdKkjZMkluyDePtlP0uK6/qIlFISpahihxSVc
I8DoloMrlzE9FBOfe9CsKkxSrY/GTsf8KEAJi+Ctvu0152534dNAeUC1dYJRMAHgTyRKmqSumSfD
geWoNvoT8DxL+9aNU4x/yzvVlmpRBdzt2A9Fbzll/u1tKL8FK2ae8NLrofxmGfPIkJmA2/6VZl9J
o33n1IMaWFd1nzuoNEOL6DqxIcAI+VpkMwPbFeeBEc9zlyIRHeFOJKZWBbCn+yHPUoZz0Vaqs0Up
SMdQBMFnHYDZY+SwMjySRBIGg6vuPgWvIMGLbB4/5EsB9llXd0eZY0TZ4R4EzMqVUFVU/39DB3XT
gOBHTgLjgJqWud3Kqb0/BM9hIOyed0CVLc1DriimSDvZ02bFhxGIzknOrYV2RTCQPeXcpM6U5QfJ
vbEGJEEERt0HZqm4GAmIyYgKFAMHkgB/uojj5iZT7qQA/KCMwUYpY1ROjCInPvVijFnnZsFKN9q2
KZFV1KK+zzM5jEqB+AjFeoAUtXYP/VKTeux43g+PKaxOnIRxOv+cVD7F19KKtzyBegJi3pq33m9r
CIZCESb0VcWASCtJdKV5mulsprxsl5XUsr19XnBjo193kDzBhiTq7FEZ6R11x0CxvZnQwvZVdbVn
gdrF1CLYIRQTPkW65QYMynB8mrNiKVrZSDFZjDQITuheoGs5DWH1NXgJKPD6VH/21XiBu+5mRE/r
ZRxCd0PuLD0p5iur19s7n6ZbaH5/Q5GQArpxaqiYdsM62nBe153KFm9qIbGbc0p7pceU8zPEDewb
bksIj6NkFoBlPV/NuJB5kx+cy6K4mAuR73ZH2dZDAiDsRvnvP477uTV2yHmt7mzAqyP6RNY2CIan
d5058m55NWd5Tj5/0naDJaUDiTnonvCNcqw1wDder88kkfDQR9iKKHsEmLGb5lwn/7jP04JrjFuA
YPNm6aFuVfhPCHp4+OgYyGrfr/wRAwFdKfUzwiwfRC536EzqU6X0fv7lgY8GrmwlOT464BE3elQa
vAiE5Iq2unfL61+YPUDCloOqKLIXRw5uvaiRrAkdlCDV0MQr1e+G2FW/+h5ytEWTWdz7zMwXgGpQ
Gs2BIfRKzJmnRO+1umD/mdYfUjPWG3rM/D66G9uBNzHUsh0Bje8V84GtjqpgWxM666cJhmezkjx+
7BvK0M4h4ns380MVQewYjYgQAqYr/7Rx417Fqn0Id64gcWtiKMdmR0ziehsS7nqAmXBduGUQv1PW
icyn+Ly2jRYzjZpTRqg1viB72tAvurp7FZN1Tjkwe09vhpgrGmo44Kbv3mXzWVf1kG16JuyCpn4D
M/4IjIbvN4VH//OCnrYeVD5R5Z6Chk5lSJicmZ208rpa9/pEklciOODp/4l7h3iknFrRSy4sBDKa
WWdUIkg6O16YwcKrsOSYR3gbnCUGK1+6yJXUba0VkgHhJag8V69VhM8jbJd4ONTtcbqJjoBS6EDv
laXM2biNBcSBgPnJO2uK+ufu31NHV7pXkWxL1cjuta/3IROtzUJu6/goRHiGDlKcJbXRRrZuhenq
zEO1/g4FMHr9Sov66tSjKGyx6Rd6Ce7I/YJ1zw0fFAnJtP+ai8z5ufpQQ/0nUTQFKLv7C2ZhiKbH
nKLM1oE3sOLHmOBP39mbFx8VqLDTk09qXFW1OcFwCOYA9lp697/pOMGcDmUnyqZ17Gl+rvS96O4O
y2r7nVpyglTsmZKUaBR9ZustQGc7VHPg61qYY/SZ/J5nacF5iRJIuQbmHoWqeTx8e5Mkh31GVafM
qj8nhoaspft1Ps4ffhgNGHjRV8CKadjnC+cFKT/IqXUG5HV5MNgoYOSMvA0YNc1J1/Y2oUzbWfL7
oyGh+WEx7sABibFuieoCn8wTiZyL3iYRqA5ruUi5sOz1QRhFoG7wJmhP1uz3oEZv9+7VDGk5Xm+P
KEuGwB8OXblxO0OIhPpGHjSIXiE99cUye8L7+YlQnnry5kyZK1OBNBu9K/9WFIq/0/j0uqxZC70u
9yGU+CEBNZqam5Hrkf+FW3x6Is5+PEROeAS5XQpUTLsfp0noBMBE/F+A/hPKlZNOek/0QM6cBJJJ
dADs97BECnP0evKhOliTiGGtu97/ZXmubFwNjOfr2Gf32/2l8omwumWRbIdXiT3GrI0pk/57k4kY
xqvbnKMA2FCjfc/6L65JZH/C/+frzKA6YWFauItR4qVJ4h+1ahOW/37WqmT6x7fE//EZ8u6tYnt4
W3qN5mU7Rn/QfG0xzLWhgu1UHpxWeJ06WdlN5QdYC0A1NgTTRXLK53StqIrNo/TMP3i6OpFus5vJ
82byddlJDAdgMkp9szoHmJ0lX8KMknNcn+Aj7T/FnJL7QhZvexdJAhKxARYPjd7VQMb3ka7g8qJj
e3FeBZV7lfwbDXE4km38RoRs8GWKmpXlx8u1FMXeR904KL/lADTQqIZLazkLmGK4ozQdHK9cHgW5
Iwayqe0+/HXRACEsREwYRhzuBK9cPovpLU+o2sFVwSW60ULgat7PQaTIkpr8n5cTiY3wQNKsAvRF
bo9Fz+HiJM1qPbH0euflmXtkpjLaU8mlv9MMXuuh+sQH+vra8NQy6rFiVP6zSP12D8HUjBAbJotb
r1uWNO9yKpOTCYacywadbmoeZL8G82+j/A4CkxWqKc0pOEUlt6er+41XWXz5r9r9jBSYfxi8dV0i
BMlK3ZWm/sNlmQuHspW1XIpxbFHjtVDWOoSJ5MSDUMY/Q5GQYZXvbcYqvMboDcVV1wDhJ+jjSVwV
DXeNH/ClVMxhdq8HqALJKGrCMfRll1DRdQxDhXfjEPhO7kcdczCPVl0n+mGGlOINZV50A66QOAup
5m4qMIa0PAew4vAe7o16qzISBOQTGG8nyYbAW9cKfGcEH7NdViJW0jWX8WQt0Yusyks8T1yUbYND
hlvNlxWG0qCwsaumVrU2Cph6KfRE0j6BvJu8dnC01ANajuPH1OSPsEZ8pB6587ZUWNkesGBp03yF
WhUPerNXHWjXoKoer+RRjdCwir8i1HMWQm8ev2nn3ARjh+KXKrq58D/HFZ8iTMdf2KXSVJdMi0w8
0NA8y5pLSGcoAb9i0VzmdY5NJsR1xvmTORzaDjJoQCVzMNiWnbO18d7a5WxVnEMRqi1DDjgkhG5R
fHHeVyqA/VcmXisWPgyX/8XFmtdQPjlrPmvxDhsmZA9MxV9jOBeqyhz1nzzfq7r3yRezwwsw7ojG
gCbWlesZtSTx3K5XunhEcnjVGAUKti2+IZ6bdafbKmgWHQtv9VCiH4JGTHUJGpgZ+LTuZUDLAv0P
ayxsW1UJHKsoSStjM/IVexzkefYrVrvx/OqYF8Ju2bH3dq6TrJTtqeOQCYu0tBCixdCAFY/O0L0k
IjFahMsE399oKq5Uq4K3Qoda483blDd/sjE1d2hFwBoNUu7hPaLvvaBNaSsLVmwMhSRA2ZJKqDMj
rDdbqY5xuiW8QnAGMVlCT7HOhW+jPX6Ftgq/wfrqu6dVQqaXz4uuIc0H25CvsejQ/umjfN4W3mgD
qPvYm7z/POfsyl42VrljNu17KIPG3nxzo1dMiMYx+utjau59a1rWIT7PrexjUT5J4jNhysAkoxKH
Xl9PVJFx2T8RwuyssgplFM0FuFJbEmfQ2K63iGArsRmv1XaD4TIYcbls6cAbw2fP478ldgVElbhC
KSYYCJNEOhqEpIoud/lhwj1Bw404480FA9TvqC8xTiWzMx3mj6VX+dIFJ3NYj84BV7lkNqzQ/f5f
eqjeOUzlRZWErlGo4dE6fDa3jLiHd8o6Vboh2ucG7c1Yi0DxKToP5AYPC8nROeHhP3c9pjReFemp
OfA5lVNwqDqYyBglvjisJDAUnEWG2rInCkojjDqY8LPzllipOtBL5jM8CEd4LEZx8+qZmxleg2Zn
WKooz/02WwsveJMN+CE1rM1tP1ZuhbqNw2Daxs8R4MB//+Gj+PRItETaEbhjJxaqIWWyeok/ax6N
5Zn5i6/T0BXTijx1SSdN9h+Q92Npc4xI35alNk6n7RStifXXQMBn7Dp7JejVeANG3nyfYLdwK8rL
FTHQMGCJL64eZhxJV/KZNqIl/5MzqsX9eqwYb9Ey41DHeBwLDU4mpZQN7rrO5RCkJUjcN0AukAmF
DeXp6gg+ynQmyHaSQmjVfcVgvOfq84QjWp4T7UqS3pCPmiNRjQngCYUzB0Wi1mOdgL0gaR/A2z8i
2UWTQizIBZQ9FOt2K14hxAPHwGzSFRKT6+7Ii7KQkWmHIfD3kQakFJzGJHdlb/L/ei1yJR7GcNuS
V1N0YL0rhhXcd7RqPf+CBkeKd28OyQ4INHER+YXBikiaManuM72/fAqSwm0K2FdhklZ0ZF8yJC+Q
h3kfUxIhFihW6D5DCooSBdDeqVYiqbOXV/dYPFMkyD1Pj3hfDujXQNSngzFpSP8j81G6Npm1QW3I
yHigQssz+oOxqKDCtcFJ2/roSH+yMOdO2PQAuLrOUH0sIhGTiTYgiaZAtbbury0uBVmajqB5QhY+
vaehpJkZBszeRWCUN23RiDdkNmrttYea39cgj1CEFkH3gSPUBihaZKT9OZVYx9W+MgsIPK0oCnaJ
zRWRX4Vjm4aTnVClUKLBdGJTHnJ1c3jVkEnln8L/PmAKEj83biND6TeMRRC61Uhs9RZV14jKZGqO
WzB7PNWSSKoCdHXmtBqyy5Lrrn02Eauf4vo0RvtpEq3zxWdfpoLg8D/AB5xYjLa8QrtuQZ5/FX/3
vp08cRY7EHZP0TTNZxcgxMGZzfP1mySYHsX6fJbhRx5m9rG5d2tOsyQv4UOXorWpDn8+X/cSPRKw
yOsGhgiIeHRhb/Xw2POJ3FRjMtbIzr0oRQj/TJZtSrNlAbFwH/BDPbes6RdzwAaCwVB0T7UrLY3x
Y2DIwqeg7I9Mr0mTpGTQQXGfxK3LEXz8EzckdUnqB5+ENgrQEnB02zfHctOen+bXMcmgvqiCAnrM
MyV2qOzty4sgL6T+RgCxvD55AQ52hD52MYYBXNPV8cWlw0LE1AmgXlvckbHtTCv8yWWvteidvllE
BNDT1z/g5XM6nqfyQQr/OmvCtDX2eAOWVdZa57iGT+We4INmJW/i20cW1KK1ycZCdFD77QjN6H6f
e5oLA252ht+leF4yH4n5wzoljXPNEehL2g99R764QinR7DxCzzkbKXW6PZ3/Q7THTUvmuafyGDqV
4LxhX+gJx8RHgpVEkyI8bZ8IvuKU6z0D3+m2LmWJAjRY7uW9Xgo+2H6otL6z+hJBWooFVzv5zFEk
BGvW1/PGpl3FqJZapOwipQBagSMRDWrIT9vXckmzI1rMUXQtkzYH89YhYHEpj02wzOxA4orSKwzX
T2ZGwoBauPl+iRc23yQLOV70TDNThCIg5ClsihFukSyni6pvKCXh90cX33fjh7oA0KNilWFqzAnO
hVHty6abe9Gzzf2h8QQTJ4oKVwBxbEwA7C+VTzvzH1NStS67f5wSyfaNWXvBKq4ghG0cosaRdzmT
+zFPrr+MTNPZ3IMEYHrKOn+ZqHvESmhRpKEMEh+ta8uFBRVf8jLOt0YzGoLQJ9lLJYZoogu+zdfw
UoHhqfs4Ltbv3SU4O++R3Q5pcXMik99AK483SxgFC0aLrB/2mlSz5cATfuUmxRhuXYCut0Ur7Vqq
hnk+4HEq3HR5YR2pEhM6wrGJKebRXfCkhaPxdbjdLYeq1i1+oeTrtd73jHRhzSrQx5JoEJg0FBjT
s6IBnSKjsECqEoAgFd2/85ARKbW3YhQJ4MSoSFkasyujy4Qc7ur+bz3Id3AbDG/PHhrq430Fdz3b
Qgo0h6gt2JDHdX8vozHGE+6AY/F0sSw3Tvw7Edag9BQLaK2gy0wF8gvRC5osQcvZUXn4DiDTfUes
CQTsXaBVSkgy0+ktC39pDprNmFy0/5hHucRl2qA2+wIkJTY+CGTpMLkq1F37DneZw8yfIKfxGX0F
ULAWHgdim9UsNu1wzqvZTzslGI8UdwkJlTW4Hou55CXpiksS0P5mOF4A5n6po02gy6e53SkxKWpi
9ReflyNzmG3s6Sv6YkQPy7prye+8+Hr3KnBsFHdxaca/64YK5x9pLldocEtiEMDTmgdOpNLBTHNk
5xLTSw1goZYQMtWE6s7OeF+oCh5mNIzSlWs1Jxw0KETMerihTWs/k223qxFImBrOrB6xyztqkk4J
D+WAPxpTpIMLySjmLbfWxUn5gc/CM7/XmHcYAxaYACw8D1/hXLGinNfpqwv/gM/sjXP80eobh2ic
NHoaTnwMN7Oz8sg0IIfcnWWRTIoaN912mkCy5SxzcxU2jjUuSu5P0u33ebJ1qBMo5MpHUH/r6d4l
YtwU5ox3TRzRPL8diX0g1/VVHopFQxTqjW66CpgaXZEs+ujQ3JXKYkIZeaJgqxPt7o0VDOLiNnaf
kxhJ+R5Fd1Llxkb36mJtLA2qETt0P895kqua7r2jFBMPhXeM0lPNwkBGKLKhC8qgojTcjI76Muhy
laPsVbEYq3dG6VH5ugeIK/KV/XYmR7eZLEwPR0Y3zD+IKeoil3Pt42iNVUoVad6O9zcSf8r+Q32G
ZkZi0vZbk13uSd4h9ci9YzZUCP6tSSR7CcN4FQ+KNWURZxhTPiH2JNLXU1JdsLY/vK2jmaKFDR9M
Jq7RTMOw8BjDrZIBktJt9CP9YFO5iBU4dXgygGqzGCWo2+4fCZ099Ay6VlJMCKbBa/08hvEg650d
aBjMiI0fVTT1LBqhCJSFXfHzhb2Z8AHYlN7wJoNTs4zNYhVab1lPOArzbPOGGHRChlOVDHvsjNCo
Tb9DziDvTJCoZrzdfDu2xpfWjX2XW8uQuFXoBc+5D2oY21udXQ7VXXTH/hVifRPTZGIjhWvjrfnO
SjrnezseDSp+tMBosqTsAneC4w/XABiaecpqrr1Rjq/2ERH+wkL7jP0lyxtzWiZMZCzv6YO198rj
FxahjLHNPzlFIaZMAjGbsHJwe+U+JoQkbLcMg21o5G5POhXEKw8th5OlTV4UYeooGEx/OO1cXBA5
hsQAh7TCiH5fTFnkC8hO3AlW7w2NGo5dk7+Hu5MGjcZqxKH8qcM86JLaTh1mg0uklcrg4xkQ+15T
GRHN3PdDhlYnI5encbiWX4Cu/JFmVtW7BPUlTpb4rT6a0loFFiqtxP75yCMLeyPtVA2UrjlBklMA
0QLm3SUaYec1z6QfPlA5teMTVWiQCN8RDo6ZY9Y+XlOxEK9IXDvzsNIuasrJJSO4AhsDiZ7K3kB0
1xXxGRtHMSlPaKA25tH75BBlUVNVKp1EPcvuCu+vah7BB7BG0fkuol6WRaIu8NCOWQMIzMq2e2AT
LqeCglBQ2N9os7OP0fGUsXJKINq5RAjQcqD4I9IXAUfi5IluWmbrKallONBypTV+R3k7zHmzWjl7
B1qGEHzkw1HF+zFkzTBe62C+kuBq9c3f2ousS42q11gcoxssN7UyUhmMQ7SrBETN/Hc9Yw0MEdjw
OS4FTn2Lh7tBI2zmI23Zv1qH86QUxIe22c/ULUjS253XQ+Sf+Trd8W0jHWmhI/5eE8kWOeq1r9xa
VtYGX05tnVq51VCBN5SDThA4z8VOTD+KO8BYLQowzHQ5uw6HF9DtbTzt+wSgDFAqqh15ghSwTh4K
ZtA3SJjHth6CH9X7BS1zGku8kzQi+rPXYxeya5AQX4wR13nmjkzwOXhDvLeS+X10TafNwQkIhQGn
bG5AFEwhLsi9pQhtHxMed5SI3LRoAcaLQxaWXHaL35lcfdG164U76+8bZE3bg4iys9sERo2jJN6h
LnajnR8TYn9dbGNonE0T7pxX7a95Y6REyiALOtV3YAOolqGRWp0L3fR+EryHT8ReZfHVdLtpQeEM
FT15smZOtBakwfEpgdxMAsJsUVqy11fiZYdFvYIf/6Lmk7wSwRXD/JJ0s808faWdtoVswrn2GVDM
5t7fKRrIsX5zgrzRJCFcPCNhfqbLXJE261YnnaGlks+GtRE1fYpgoXFWtykQKSoEUkdsUWZjuxjt
gebRh68rtHfZsXs7tli8TqwrmgHKu71+cS0FnK76Y4U+dmymdW7umAP8eHMN/OgVwXkN5u/agZaF
5DcvCBKKUjEtJxT23SgZcaobaNlvbj9b1xsKezX4PMxYYAO9+RpajHDNYsn/49UuAQl8knZ8y4xD
y8gHAepaTicXIg678yVp6C/pRL2jEqnS2ezmWz/RNtaPmidrgxDkC3p8hmcgHjB10V5Z/x1w9mh1
VcmLTMIscqJRgvUKC7F0UrmJoVeFg33Ei5NYh28jS5JW8y2LxMU5fcr2iKS/IDT6mV+K9iCnXiyM
1aJpXAaBam+7FF8yNNxbZwEt2PEv1/QAD3EW8wADsaD7dF7fgPtVqBwdFIJHyfat16qaDClugY2b
W300hr9FnNOi9m0x4Xs5E4C7RBRMafplBUSMSPfEUD2eT3PGqRFxVbND8/dJPfsbOs7cwdSJPUhv
BOPavcFe8DLh5+J7g35BFODc4uDbF3wT65ZxKVY+QoMk2647mKsFjO1adMrSv4aqkqslXvj9KQMi
Gfq2qQmi3bBa0msOlAedBCS2gSMBv9P6xG8YhQr77mOeJOugx5K8/+/sQbFR1qergpIVu2Bb/tEi
vU0ccCohZwtqIseJc4vNXi0eoxkW+BEwRr38DHcq0al6Hoe3CZXWuldCkcF+sAGiPZRmgISpIZG3
F7FsZe45UTGTlwtCxu37nHfNBYs0Bciq1dV/BbQdJWj30OTWZVdJwMbUNFyZpHaNj0lps5cnMYRv
AOFMG+1Z6A2lv074w0yiMpx59WpSz1daqyTCdtar8HDBftNRozWPtPRXAIEZfMwa1TVW8KztZ/Dj
V9zePJSvBf+8KGYKM32JlRC5+LuAoNooAoBKVjjKXLAYAMvOjBy4NJqVVCIW/3dQz8wwij5mgNAO
6RtSjC27ye386X73aTvLu7c6kQBFBJzHHWpU+3TmDI5TZ4SSXth9BmpNPRvL7rkiFFQJY3zWRmVv
mhb5R+LJO987tlRtzDLuVAYZEuKwB5bDIhgpJrpjJfH3JBa6MKgIp4+vKB6wmg2LBzEPEYDIvxCL
kpFDak6CNrIbtMlTHcuL4TZ/U2dpwhjBS9hXjqrL342j5Tr5NN8UgCzPCThwLNgtL4Gi208ROVcb
jdH3QmaecVaEpbKZvp09HBp650qJFFqVcBnh6Bq1AdlC776KPXtK5ADNqMz4W4y4eTs6yqhPWIao
YJ90wz78PanqHgoxetAQ8YI7aKrB+/nptlF2UGfmj/SDovru+NXuHtpshPaxbIcKhY3f045o/0TQ
GR704TaNBdPb06Wt6xRf1od2EuSwLIM1s/DZdi+lck60feJCtBpx/5FDG17ocp+eWwPdyyh5pnBX
vfwj2MG8q8arMKJQWQa5v6L4zXeg2ESimKQFuqRBPGDvM3Cw/0LxFaGTaIYkTpieBEu85Ld7+RCP
baN8r6qPeB/R43sjLJA1ZYVsrLXHbQMtcMLrlPQNgH+Pj8oYyIMCq9UMDLE07WW0GJ1e8z2pLppI
BkztDUKxFFC+g5awux7VEZMNH4VI2bMr980wxNZawOuCD3/1sMJI0zwuNUpA5F1NWn7N/vVrIbRp
t0HXYFq0bTmHgrpd90ey/FMFuYGJJxzgnK7CkkEvyufp8qT6pRT9M+7tETyxDC9vF4ZZ2vQLVmOD
aPn2HFPpi335QSOJBPNR4VwjBZA0brxgYPDAlt6WtrMbdpOqVFgllegIS7GlrxS4xCnidl+V27zN
2ZNcVYboEy59oJbAHCwyMrga/9UTJNBoTvyfPV9F+LzvUlMYls06JvuDfl6jxqaT1cMM2HC6m3mt
GeSr1dxVoVJz4ByHiAr+KWOLLbaSXlyhnvExeRaHIn+gh9g+v40Pcrrfol6b8PMLxk/5MvWZl+di
jTbaaTChX47j9HR0rqV1KlhzHmNab5rYqa8Va1Zp7orSTfN7+LWs+OMIN/9seCeLz9rj3rGRjvc0
h9vJmfh75vVp7GoLADR/YhEomFD5ieR2GoZPiD6O2hXVCIPek2+IB1hv/lZIh68/yKHZ5/XIQS8u
mO7PDyVu7zuhWjxzocGYK3VyCwHFPNluEzmKU73ByrYys7QjXGEXvB6Z5q8pWeJQAaRc5BpYeLBs
K7APrzk2fkZNo0cTwKS2C+q7RXkyRVMj0P/0iJroZ1+wm4t0uEKE+bmxCLN7HsUkagAxTjtozKQK
OjKdX5eYeFrFQzEn6UtO0ZF1cqUmFTKwqHhjUze/XuSy1QDYdj4TjWwgquOCjZC9AHVjreu2TLgZ
nViOPAV9EuwHXFu9L4BEj7s70neSRcsteRHP6/lonEt5gnd6owJ5TCvnIotQN63B83ophmKcsOxg
pgzatp6Y9+rowCX4SpC5Qph6Y0ZWwpKkeZXtdy1dnQCmFDM/nFjQOWqpId3+e/4WPwJJnJdIqF/G
Tk+TH17Bcn422FgQDX9z8C2TFtedSaSF+HKyRiFnDD10Skzm1JlCMLFfSFL6KuC7108OaQVQt95j
IJArEKznsc+nd9AyRPHaClHmEKjQTentQGappV81rXOsMhqwbB1j42iqYLwqaf+PlQ1m5XkitrH0
T4lAykgiwCv39YCsXE5jBKiMPKQRSf+JUZC0jquow7EVBq87babMP1ZqgJDEB7/PeY2aeOCC57kb
aLa5nSLvZQWp941TZEVdAn1fSW/B04E7ndlyMPQtnwPJG/XExyQtHZGajA7XwEBc1ZO3wQLKsuty
NoOMKYjhDBuJl0YfS7qHRyF69X8AXSW+F4tUJSob0EzqizpckYT/bUx/LG6weR7smyiR3vwTTvW8
NHxQBYtavOZL/mjEShiz3SCwFJpMSFQqD2x6FDXpOd2K81UBF+6HUFCQR/kmWVN6dXWS/wSpoMfi
JpjmLcr/Y/CTIUkLnSeqW/sj5YyET/0ra7/7Gv9I57cdqbrDcGaDdyo2hyPus+NZrVFDb/gGfmba
I1xjGwOVoK/5xCHA3s4osEfQOKF6WJ4kedf++6zxaETj3+KVlhCuGAc0bFSQ6nzJe/PQ7NM1tpJ9
XDJgHKqOuHK1qf2Roarz1HKig5sjEfNepDeEDm+hhvJ3MEWerci9uKB76L6+cZH/kzjzH7oKp04j
1uJO68cdWqpT35UDd8zd5LrZHPunCQDmnN4P2OhG6D2ofTGrxN2bN/UMQbFkKcDSOnNQGLHq8PpJ
YnsCjMzw0lO7ciu8G1sCHF6Bf0VBVBlsIJankJDcQNhX9t36nS5nRZ2CXLrsIk/VGFgn5NXAamYM
w+v9Tn9DqApM1UWN3f4BVU1n7YpqsEO2JG8wXyJ5avXv/i6a2NDI5tLdQ5k0ajeyJyGHXBH1QkuT
wlZ7SoLIF6yZDXIE0X5PFyzfzR82qEBG3k5j0wVLHJ2F9DSx5JsRPYhzwadowG6EMDSfCgcIW2WN
YjIf8OPgezApQ+vQzzX+uvUSetPzQ1oxpb16T1282cBWz5Y256Xlnjw4BOoMqfsGC0CbDxlzpTd/
C7tayoxmlT7RwLu4cUXrPV8LvTctUhXKaCpgeQp/X5c21HagEuY5jJOXXur4CaTl9NBKNlo3iwGH
advzWggNGHMAghvju7+ItKpRlBlZzSFKuUtnAdbIT646AW7+xnDyWHdahOn0t3cORACoBNWXoOrj
Md39r1JlICWLVQRMoU2HJZZxsmuwREz/klY8d4Nk6zR6/71yYK4NpG6tY/wk8um/lWX7M4I5CNpP
Q/grWBDJ5bHbyb9A+ftj3v4zNNX2FPI+GUTmvyny64FWEKg8XqDCyuZxHXumbPhM5G9+aQhKAInk
Iy//0ByRVMbnN7Hm3CdCt4qzsnMehPs8ulzU8QONhfwVOxsozyGi1Z65QBBK9e5wr52qsUlhDbNF
e64ibSX2FTuLfwWz6lSb7Jl4fF4X+hKpbpY111sqZ5i4jn32ncbxyq0nasA7fsx2wqCYmCl3ht+N
4FxngMEgvBxuOEMiAjeNYpo7r6u9JeerogoF6mtkL0QcDqvE1nD9W356eAoQXkEWqKFucMUnC5h2
WpzoC9t2z45sFe8rkPm38h5ZNcofAvQXiIeg2dmx5H4bZsf1QOduoh0vBwfASFNPB1NNci3r82WP
XzZRtIn6PtT6ESujvTU44qzyffckNfAcEF7zFqOxI4krC9nnf+gfJk7zTvioMxFQSkVePxTwZK7k
Rv+QPzajJFW/jMyanEDqeA15Eyjk670uqedaRu9eNGfpTJQxnb9JI8joNcuD8LUbfTjxygeh793P
IB5KElpPhsnEymbv11Z3oVxWLShYClds/Nnnn5teqI9qr7bPXeqol8zX6UZFIWmFLsAH87OgAloD
rd2J6TwdFqHKpJ/xPNLKFDzkg2nhUi/vDm9Xy3QdZ0ig5m4zwaXDJeRpCftX4FBOL9E/2wJHYccm
i0AEUgNI9GDSd6Aw6f0o0K6ZcXDQZJW41uD0tvefwBXS2Cu3lyDUSH8HrvP7Gv70VRkFwqBBEnwx
Rebs21nQMt4iYnvfPvi+d18w86PAPtK0KOBG4NDKssQGG4Dc6JVqafTOMyF9/xILgb866XJ6Agrn
/RMXhjKjE05IYjD5cRLjsJzHZNfZOx4JD+B6FK4yz5FeuzS0W+4Pv+wMSI4nXYcZ0ZAlQGo6uwcA
oAAnxMXek2Lxy0w/JNtqy56ZAZTQGP8K4MCOHdOlK7B6rQRt36fK+wkec3h/NdYXD0uIBN2Ak5ag
ASiV+agz36WeoJcj19qzfbndxkapEKSnLGkup8Dsr06vCwhicZADRnq8O5TfHgQupESAxLp/DRhC
kW7T4FP85gvC1FePEUr5pBPyku79YyUtPcWqRE/zj6z/fld7nmXClWI+pATdwPxQe1MHPjIQXzYV
S1NBrosn8soMHiJiVIZ4MXgL5NiCtIrlCygfGbj99m5Evs+bQRV9lGnyG3LGfMeaWAp+aoGotAS/
NHkDGwTq3x/sHtwZVyXmrLHb2WgJyYx5Yp8rS6dcub1CLjLTyXdVSiAmy3EIJa6TEZFuTwvrsF1M
E5vRt/HU4buiL1onLlPQICiJbrKOem94idDzRCdmy9znz3KtH0ZNRADG9X+wkr0S7V7bEIci91hs
LntKRlnunWiEu7BJ7RQN6imdCneE3iLqIwLGEi8TVhkBTzj2aCsKHSiMn82xoH3Yis1t72Vbv3Fh
bxGaO790RQ1qEHOyn1fYU40HhSuOIKbfeYHjlvjkzja8TUVpB5G7iYAxvrsDDr9hiHXBK63nhSAx
EnZAG9PS0Ca6d/yIwtO8NV+IS/PVEu25A8w0R7fGJ5a8agsz6cr7JVyN+Vg6v1bxCwDF98BuCDFf
WspPPo/M2sVsuWJWMqbE3EBlmEontTi8mfntAbKGZrEwuctZ763pLNZ7hWMWAhBZvgPbjvV5Ys3L
F85Wdp7XD6dX976sRnSl+gidV4GMiaQ8YT1Q916h7Aj7a94KctAFDD1OkBwDh1QaBEDoNraxJO8I
2Mff5z+59u5PWcoaKcMD3BT0Z2gZJPjWB0sypOGYnQxse99enmiP9n8majqwWfBVRMijhGORwviZ
pcLV/udUjFfvGB64Kbn2gaAzzTyVCmmVpI7GYAWT19zc2zu0YseiozcFQKJ8gk0/DjrPMM4lnUQ+
GyDGFIGx5HalBHxQ5kQzFgQWxsXSOmdRBobtwDx6YTTEb4Txhjuab5j/EGwX2CyxmHyMLClwBn9s
RyGgb7WkczwMvr3/9Nmbo0YTFcnuuhWg2p2VvMqRe3hHulLQZfgZW6LBgAhoMquV+i/id19T1oPh
Zo25way1yMGSqSAVkINm6CYBnA9f8tSPCZInoe9fWoKArxB0VhL1GaQQJk4Q4MCHtBQaGIQhop1e
g0fiikRRDoR3yDT+ZdJdb/wrVBdE/bjJXsM0zaGOYXr6dENZLd07fz7zlHxw4i/uFRdnjYLtFz81
mDx3gOy/qcGQIpwC5fe4La2M5FusfItiW0h4z4grW888/+jpF6nGY7voKNUo+Fbn4qm6AlR97mfA
ohPz9tQLgmgPgXBtiSmTL99+ZM5F2krD/7WW32kbN14lU5Be5f0MQfZ8JHm5RywDl/q2Qzbkioxq
udqHTiWEsuwiWoWls5ygMrzClPCsxQB+dITWLSdh4WW13cuwqq1A2E7c6yaTKyFsCqDr9akNaujZ
PUgSxwDIHsrpBngOe/cMDshN9BGrNwraICwtkNy9U+iY0RFf2E9LPxNPw7T6ALdQNzYbY8cVpFZd
Y7h6SHqZ6C4NvjVqyASbRf6RCWw+gHA19jMF29fJeVAFeKaQ0X07c9VKKFL/fpmwThlyo1DdrzeT
3ULztYumSTyIay901qha0x000c5zWwq2I7xKzL2vFgpuuls8N6RhPsdIM1kH8dI1ZwMJ1kNDukmB
QictMJ5iMRoSsc2Qy8E0pTEsGJcxkbNmZJvSxl5I/IYpMm/Ww191I4GJ+maNGgffKymf262rslxh
1aoaJiO82OwTecO3Lz6bQbgmXLUQkFNA9PkS72nHjgVvgyo7gRB1wjjOtvLujS+yMYMr+CRABgh1
8zxM+HmuNgif6dp15sf33/ksKJG+lsj+N6w0rFcHh9qUuRXFZMSvkfU56h7Q+gAJffYG7Mf9AVdq
/R3e14nNB9ovilddFWDN66iUH7//8xljojhNs6xGiRNQxnhq8F8C3ggK/6KU/7ySZwsfxx0n7/iW
6NxtHeaVjc/t6dtyjopQh7+XegleH0TnLhFX7xUW8fuGCdH0vz8+lzEAB2h6Z3v2Biav1y2B8bWl
ATVvzlSOfTTw8L8Qi9gkRGLg+fI1RXmD7mw0nYelixgFUjHJfQXqhPps2dA5gmpXajYscCF46FUt
zLwwXhuyNp0ZTYkr0vbKor/yJxCN6/Ir2dVNW8aWmWoBPzz0eDbPjq/gCrBtSn44vy3wHwngGBPm
U1M15ZnSiBn0erp+81jVcgKYKkctEjT2o3ZaCwti2BwQN0yaRl5wielnfOlTkBrFhckdfJS+tl61
BIymDF1/T7ZsLmMn57jNcFnTqxW6zxbgpiY2Edjl9x0pRw8dCuY0YyLE3qiRGQmKy3E9aCQcrAMX
f0Pc3GYGyk6wqHkOHfCUaPjfI60EY5odSO5Ul7i9CBea7GIXmKoQsO5EppwTCovnZ7gUryQcPPFk
LbkHV16BfYgabuS3VhHvta3zHLUxZ1TU8RKj5+fbWh6FPFd1jgKmj0VBTTYzJIiIWkSuZ/L+baqx
CJqNjFQDLgMaczVihwNxay9JOLVGMFzduteYXgdZhW5mOUiDjE+x9J0WvxOoJlRkWc0lZJynzwX9
DXrm2lTnPNE4DisYRUr+uERt0TDgyUGjzBjGGeK7MZUQXKj1qq40o2L0kZt/N5S9YRQmkafOubCT
5WD+Ethyg6X+otByXvZ4NSbzdS/0M3bxsbUegOBu6XYodXGLO+aCqZbrFU06cVj/nqNZNOVwi3uD
uOCRbhoI1JUV1+tph1ebWv1PLPYXMcuBv0jgt7eUS7X2gsxCPag4I8awhxIYKjAb0+H5ZZQ8EdcA
N+Hy4BfhMiR0zK/WhhVJ7z6OTpjD1KweCFl5VBVVqoM85ovNK9N8Lmk9Ay4P14JsuNb2YXj90e1V
b4oE8aOTTDZThvLtw7Yyt790lJjSK1tDWE6EIp04nJWJ8FrHneNHpMA0ACCX1nY7CSh7kI1GOzHY
6EzsAMUP1v5YEXBj2gJc0QhdF4f2uE8Zn+BgAvsKgH5swh+szmiNBMBJAau4JWohTv2KcJeh8A+c
yfR98ZYL2p/0we6cmFaMrUpgQlBjHzDpDAjrDUUN+SfNvJi1x4hE2NVTOeEd0l51KPfGQOi53BMn
xIdpHSTosSDlu8TBbDXmlyNy2GzAf4bjkDalVkX82sLdjXEL9o8eGV9SI7t/7iXu9vi62d3EtplY
mI2xMuHeNquxQ3/zbggCKoZRxPQgKWUSbWV+EQ+Niev0lc+Fp4VEGksMi3U/RNawvG8GXiCpv8Un
IoDNFACVSyevrM+I3hijRYKcDiPBXIuvEueWDPChGVTwrCNkjJiFhStMdz9xR07/Y2JwBwt7GRHh
lcqcS4wod1S5l6/pnBkp9KSYi6e9FxDBHl+T0oSNdXWJivSbFfzuByEpt/lKhJNZtAxC8C0oo/Vb
LyDvJ21vrwNkSNwWWUH2J/4OOJv0f126FBjn4BaQlQsc+BaH4bUY92+ieeu+3I71tJFlKh6zk3ra
IqmoXd+w1qeMj20wErNNVgdJmrKuEIN/yZ6H2y86k+3YQW053vRs4clAXcPOpMtUTg4P6Z0zzykj
N5mwKRN2Gn590ZyHF/QBRECyR/oaPJ1QBBPWVLsnkbHmiKmsNC24E2MKTpFiMvrgVFgWJs+/VUaU
DiU5rq+vSdlIQXovccCobOyCox5v4+Qzv62BoVn6eOuhefqwX1wxGZ1amLWpHLGMO01OzLu3txnY
yBzv6ujI6gnCOYNRaP6QkH1N/rGRTRwzae55x2XKDt5p5hbm7QivKDfps+D46L/c5yfP1Tp9wBz3
TrS5288/+XNxrAI2/+QUy4/8JEVFNc7MEASJfttR3wPpaBg53d+B3xlcM9AQIh0y3GhJwkr3uSZi
nDlTM3wl9HjpPs7K+kZuuc5luwa/T2K/5JLnlJVHtO5AqhBLBFrWePSA02n5t/TADUZAp8/3kD+f
BdnQh1zijJ0BtPU/7aa0TJLLtIHF7G1vNYbg8mgTMwDs5EBDxeH1OYSgT7JqOllbyGAnlADje3dn
I8q2JFm2C0tnBFG8/qNjfc3IvbVhPOtJYqSbz3zQMQoDeeIjKNecJI4jZw82lsBAGjpfN5YUziy9
eJyf7x72vwCIUfZ5d66iXK+Ql1/rm3ANC0jzWB1tsk3vIGT0fH3lxprRFvw8AMyKj8aCNvfP8tis
RCmDB0PBF7ghCx3xCEhHPtAbB1cvDmDECFZWbn/7eA6FVQajeGhed3Aiz55A2G0tQChbcrMxda6p
gZaFCQcat03IaSydpiDgN3qLyWgprW9jo6C1Im3d//f5EWGpj2sLYkBS0r1t6tlHqzEtC0UOGEpx
0VU8rHXECF6VC9MbRRh0p5J/n0M5L4jo+adc/VsiNZL/w3DUG2YQYvvl43jdfFq72HRPqkrC/96d
e5RVezNj3M/ObhhZKkSurulkZgqo25CTX85DxpPGpqfbzj0sKJpDvhVfXJx9oWGagR7da09ESOc/
eYWUwuCcuSWqgbjyWcHiQLP+mWXkXSlNRIuYtQDdX6mL/Kl7CJ4UcSICuZceEa2mWlwY9/aF3i/3
lSMocrvct6oUAs2y8YOd4glNyQNy7yLhJIMfK/4fC7wtxKAAoV0HO33x8jGg27KSWbXpE8KRKyp8
NoNFf3ffRda4XXrOpF/lKoxQDIDbpBb8o603TE006MkbAlevhSKf9K157gKGkV8yR9JyeXT7XSNN
UjLb4uZ5z593V051aXSNW73kkwby+WR+SJ2RIdhrYRTRdwwlie0cqXswQLX9Fz+fwU9GY8w3jT8O
3rGV9tY6MayPwF/O0UTqjr+dS0+vel8emid/QvsTsy4HQZhT5Fe3doEahNveM8WmkIQ0GfbCLXJT
CQLUo/jLsC+ZI2H1iwmRjICd5qfnwJxDWtxeCMOzrowwUs4rFOWA6o+wVmVoKuCuupNn60ucTOKL
glOdy7einfqH/ayOmZy4+iWHggrd0tnpPf7dcV83e+UdFWFRax0RGVmHKCKPlyX+onTEI2o5HAh3
9SCtZARx14KhmtEX+So/8AlapDYde2yDGZRQphgA0BkT7GIgDTbQX+DWM5MVf65klSJSA4KJij+t
/ud0SHsCkfQvI0o5O2BAFRLOUNCEKehgJeu2oA1vwoeu4oCwModoMVe0JUs1egjbp8Uu63DxT+P+
fLxS8fWJx5AoZOjHzP/dBGdtB4PY+VJt0omN1cGwc4qwPuQwFux1+gNg0egpt5Nnh5cw5Gb/QeBw
4lTuxBeYWj0/FoZ9aYV0sjn73kvWKuOXYAvV4znt9IpbFeIwTXkprne8tDuxF9Q9vo4LIgnd7g0r
buNzoaNpOY+kGKsQxHnYt3WAICz3+hQxNPYvJZXn1L7a09FSNB8IzDjqozTQ7IBQzbJmOT04nGGi
Wg0N8KY/wP6LO9JWaMijNpF/6Fk0CH7N5Ng+v2zCRp3BZt2HQ6Azzn7pFT5hEx04ZBuxOfN8mgZr
PtcoIGdP0o2gNulRdQYHOaYzKDliWM32miTqaWVAwM5p4Y1YhJI/RHr9FtP+7LZIH0h9ffSLOTRn
y1Wk4HXYHa2uBIuhuY33AZTpejSI2Qu4JADg0F9ueimKlEngOVko/LtiK/Xcypq2+d7gKjMZWkmK
zu7BY4ISnQvYb60IJXuvZ1PtXve79xyHUJYzErpGntWxVZorJ5uDIu/fcrFP78ntqDfOtL5qLa+z
Mh9eBmAGlBrhd5DpE6wbebfhPloXi3N54jHntdLPCw7lfM4s/1QXCk9R+xT9j4ckno9tZ4SjVq9J
Ur7Chp2iXtLkYRFk38wWXxYs0bV1XCO2ebhAKZyL76MabZtQgfIHwzvr0w2pBoaW2fmRTpv6WedH
VgWNmkcZvmujORxm2YU5h1Ai58m936lLhv4p/s+Jv3ACgtqFV5t/lxC2Qnci6pZ8y4db4coYinBU
lRWfof5JR1WqTKgnj66YqgGUN17wS57C3UjgcANXo3rYV+Jn7l21ujoMNCmHUkJFoXBTbAVaebC1
76D0K5wa/ORCPYy7Q6beD6+Mo+qKUUdN9+EAT64Q9JB65d72dnch5rLGIVYkOeY6l92vExI/WO31
1f8u/SKNU2kkfvPGmeXl+Kav9o5Ngq8KlcwvSk12T/eoIbh0mhCYOz0GcLp5hCt4Gk1cfRgMNZbr
6hncJ+SGkskyM2Org9YbL7TAXHBorIDCOlVELYxkVAUo7Ua0m4XLoxVNJ1Vp2UA1tOiUWqhTLc+4
RdZktkVr7lwleC9Akfhv8ekLopJH4A+MgYQNaDc1tMcMKOYciFeLTHku9KjunWqBYYI2TNOxnWSb
tlgTa9pvj1ZzQNLnVXBa1LkMewoUceVxVK0+GRoWJPAJ123fd7sqgBkknNSgNw2VCJn4EwpOD72k
aHm426yHtJAvyTax/enZWr+k5QceTyoaDlR0vPNuThQcRQuYdqbR9UewCFEmwj0PhzzIMkqN8DrO
bGPCC7XcqMj4z0VkPmdtrZye9HoVlMLY9hHpDMGiKPOcVwkZJTEfM7370u9YaWnrhmLf2ICFBH6u
upaXGzwW4x+Vg9JkRbx5kLrwDUa9Dr6PXEKJJ11agsvwsYUIpj7D5lMNBPDGyukSu1EGiDoqdN6V
+y3qQgHJxUcuwgRdqUE3DN+1cKE03Gq8LzBQkW88YXaX4xB6Pa/RnP+sXXbwA502txkfAtvqVk5w
k2j3BwM1v/4nXn7uDIzCmCqfDtCB7ewluA3K8ANn8MJicZ3zclQXaqvGORu3wXVcexBo0H2OG9o3
bruxWppQwHJ7kjgPkWO5BBNBsMJd7hChvEwP0udelAud+JtawNs+HglayrxVQBoh97jhStpd54XI
oaTYS4Nhhn/1kM8fMrZGNC0fReL1CV+aJAGFiOphYzbjIQIiXpqpmc9+404buA6qFN3eKJ1Q7c7X
5KorlkAczrYXImnKIm7yw9ZSd1E99eNDrLavTRDsyAEb1MbWwAfDzwwHp3i6N1zVwQpBPrGcua9C
vN0sb15f99tkKeajynp5HbfknhvwT2qpGbGhmiImutvBzjzP9VHcxr+fUeCPPCnLCEuDYTTWnex1
sYwQMiVnFR+EkOco/5X1Nqg5WIKQDY+QDDIKDFj/ypP+XGfrT80hGtKVw+jEvRnYtKapBlwGgY7t
r6Fq64x1oiliQHhId2srO2Ip6Nh/7B1uEGna1QbpT2uShpNFaF83VFpRhYGx69FvZAEl4pDnWW1Z
3/4qvu82mx8RdclXMLK/rdIeW4q6En/uZq4NVlGxHZZZl5XG5z5D6l9dwsk7rbOcsQV7lhggDAP+
MfwoKOK42fZYVshShwmCSihjysGQLoMKFOx8BpVHWUNfOp4vMqmqNbngicM7ZSiUnYxX8z/FEpAE
80jRcSPocGqeFaJIW4HsMO0e+XEaevYulkrmejIPnTCRnmnfUYsIazdSO3FeVqFkjCcmWFV+Wwfe
ohvnuDXZwyNK65uV8h7nkxONhxzH/HxUGxfiCwMvi59ZILqD97RiSyxuZpIVpOF4O/+xRewAj1dQ
bVSoHm180ZFNAxxXUyMcTRfY+DOT3SdYWIXn4oZj6vjYTTAKu9h5JqPgjBtv8/QPPM/aB3C13P+s
eIjoTTaw48t/6Qi+HMNnjX/sxWEZAwqnPh9Jfmw9M2VMqRt2aqTleUEYhgLM0PQyNuABGa/UzK8S
YbpTBmZ1acxEmP7qkeGC3UCWqtRNyEJ7GalxCsV1nyZYNrVxMiCFjhvqNau/MpFKvX9PGq4blWIz
MxuwssocnqoF1NzXDZzl1uvp2wvnChgQN8P854o/pETZW2Yd2HsI++RiXjWrXe/7ooAhhDrqBOAs
RYfVaiLPPhzsigzBaH1J1t99ERHRJ4DXJ/en/i5+8RG8UybhQdvnyjvojmoj3VVw4zcO44AlYEWP
xnDPi7luxgOkSzZDNNYxq3p5MflBXB1S9ymav7moKTqgAK+B8btPpql/EOyWdmstM/3qXExBl0VQ
nrnc6W4su/Z8bObtL4Vm4Guq4jHzG0RPT57Eta+P8vw9y6RgmMEx2eD8i5f8yDzGp0XYihJe1s7A
0wKklR42ReSh0yVrwtuAhuivJvZC+ETDUHaEQY4RUkwCQHfUishRmeDhw4nqKktJ6am2EKoXN1cb
NerfgVqDN/4spVuzX5JteqXPKMD0csNG0gopViwU0Skf6t5His1EUkO74pUIcgZzJjMoWw1zO/+z
+zzY4sCdn6S8a+YTUFB+iEBJH3pp1oL4Sd2CMysnZXl7zIiib/wLNnp9/bk31ixIgXzCkSRMltAx
pZALPTkBVmBOX9KVs2nxyY3q+YCx7PlEeOBs8HcPUQEnZj7TeyyqbX8cLiKt1RsloF+2A5GS+G1u
6f7+VKu2I/vZHyKL94CTZ5cqi8vaex2nnsH6kddwD62EtXIfBUXtCpeVBg6jfFn+hUslmVz4/FU8
Kbez+N083MARGxE2XzaJEKavGaV7JTTrsBDdH5CoB91uIR8peUutBuU3myH+ITOXnLqgSfzGifYD
bFugzr8wZ4wjUeMgP3eZSe1cfADpPhON5b6YWcXuyHhrlxhKG7sefB1XqO5P29KymVZA2/5BXtKG
Csv2esyu4u+XIbGy5V8rS4i3613szAC6HXLWzT043VtNFLAk/TPUqQXa0SH6VJtrvTXuZOb0PbLs
RbQDRb1ovzQADzwhV3sO4BELs8/05cyAlmvsviBYrv0/hbRC2PqlHEPfXX96gxzl21Q7IREXODOS
ueU3prvAu+J+lZjRa9973pCZ/UGX/MhAu8a3c2kUmRiu70U5uRDPLUhjgjIcVBto22zc3hWW+oSO
jKi0hGUFoDeMDfozaSQfuBt2oNb1jIT4KhxU3A3SDXcknRys+4IQhJPK3cotf620OOZfbt5BIixr
le13zUeId2lD+oMFZWV1NWXz8bneN38GHFJ+I0fAkYqcFoi6Zv/Dz63Vj+7+uwTPeAEFozo7QOHo
2Ybqf8Jc1Xbl90K+wXH6BSHLsxznBpqhiyF1UChbZd1v7FsWeQVyx5to6RgqcO+JEYL4qJXxafk+
kyIpUYcuVniEgKGqkl/Ygzj9kg1xXOiT/Ud95nxcKr8mdFsyA/UhYGgRiOMV1KVX24zbynjHyca0
wdaJPsVxNuiWmKzyBPXJiEz9lel9Tq3+4qG4K2nyryNXKKLpJaBQHhmgaHE871kjOIyjjSlzFXRu
nTV3ucuGCV77/mfwxF5uJMIWbeOQMMOfct2N0bXnFfF4z2gH/gxH3jk3HCqFeHEqz3Xc0B4NB8k0
prKtzWc3CMQl5xctIf50FnkZE8hv9UXAWCDugxOYIOTvQOAoXXgfKwu5AXbjFqwvRU6GI9YqwcjH
dkOQWHO9+clomSzHmduWYvhZDvlCR8t+D0oSWklfhAxiD7duQsTPVju5JIyQ0KuSqpgQm2OV03Fa
NcItIohYk4/yBUbMTT/PW00Bv+GOintRe39+G2b7mU+F2d//jlsgu0lFGKmveZ2aaNbv4Dp9VrZr
o6289b5FyF7PoIj0E1Vc19Z3X9o4cXcvf8woNHt8X3zyQMtbSb1UL4B55snXOn/4hR5W1Yt+GSwM
AX9KXQIrdRErxq67sbjrTm7DTISp6ZyBceubLE1vv3HiMmfr+gyVp3pfDMRRub2hS/AcgbUshGF8
btr+O/4NzxNwNKze2K8q6ZKFaD1xjiWD/m2FIzAYmLIw0YfDPeZqTiBr1kHoM3KCFBjr0Wu+J4VQ
lZ8sTKCHmkw6wpXGKwhioeZLRFSYQRaLhBDNqWMd9yd8giW2+a/BWzHiF7DszQ2OsEtzGzLwV7VW
U2W7fNkmrmLh474HuDY3OOp9oLbKikKrojqytfMXRv2ZlmSgsxzUKtnqauAX8+8xao8BBVKw++3P
va8T9jSXimdHj/2IL+NTAfq+clzvcgSiDHf/LsstxumaBkV3wfw6Ojs18xo2aoGUh4EnQ7wtpmKp
YkOPBzkEIL04yL7ELxZ7snGNhpdBejZKA/3Uu05ZqWA/UKnjo66d6xIV/WwSPCHejkiKea4/g0hW
fGgA+vo75Y83cfEoOLB9hAt29RygchooPJusCWhXphSt2hZZPhSXNQDeKB19a+n38HnO/n1/EUAR
pc4mJ0gpIS97U7yM6vPcdniQE0329mw1Rx2ce19bTbmEbbDqX5pFQlHckfBMAR03riaG68B5WUot
muY0YEx1Kp73un4LRcND4Hk8XKoKaaHF4lY6Gibvf8AnXgR+MJZG715X3ruAP2T1D6fT8BBogG5V
aIx/xsMmy40IytO0c4iZK4tf0Gia8Ju2lHd/Z+9wvjFKXwFXDJeb/+bv5PA3EiKu9XB3jeuiF8fP
uYpFRqNPU5yJtZ2rqaVzqaBde+JdJMNPUCg0+l67AfA86kLaAfDvrC91EgNx80lsTwXEmC56wpfq
yPMnNHouKe4SiaRC02f1KSk4DcMALN7CnWU7LTin2lSz/6jwQK7R2BZB/dAxptA0Tt5ygwCwtTie
LqW2woQTQwtEXL5p9wVjwHus5ZmT+cfgLJ0KDMn6kJK9zlsQg/GNplgWNmUAt3dKViYXxfakKU16
s7yh3ZlTyjMOUvr9eUXclgNz0jUv91s5LP+OmNWh+WCM+HqGXtk4SVCFFLi27aTwfEBW7o0WsEyT
UtxB6hK+8A8dzqXiPviw0W8K1+NjPPPGf0/7jFxJvJv50x8EyU2YhU+J9GcCITjTLAY7yIb9tz78
TLbUXNwIht1+h3lphnFcWGLxo6CEcappU1C3Lcm6oTBPzglqncX8Kt9kMs0MhR9STGu5Ba9SJBRW
adG7TUGYJVTPZZi7NxlucjLYaO/OO3sMhCDBw9lqhiVfPc7U8JA7atcyCGIjJ5UVw43ae37h2yxc
MV+mLC+6zxJHjCrXsknBiHyriAgqOZrK0D/crUXBei6L9iK8UHN+Pac4/LRRAqBrpKYoecZVFo+c
iFfYRQDHwkx72Oi9drVbAZ7jPKqoLY8m5usZXWxV5IbCoSmZuyzmtD8l+RbN+93q066nPRINV/q7
Udxd+zxXgbVauHBTmBnaM+o8iqd3T+x2N6AQxQ5oFjdT+shXLOconuLGWS423R6rtsclM2er4DAg
JhCx20WDt4kcEHtD0g0R3BVdKx9GtgBrXBAOvkaJokH3r6viZnl4yY/zwSMMUcHqWGKvzUtyakXq
rAsKnKKDkrz2yCmTb8gvpYkIhx8srXddykmlL+7f1ChV1wxsSRjZ7HMvomyNcAyJlkjWUP7SJYWZ
jT+iYKalx7e58pFZrF1Ay2B9VYJdMFskc/en5e6lH4Hx/75sCQ+yBX/WIN6Iknv9H9KwCb8j5LKq
r/mSkTKMslgNYbRoU3MoJxAYwEIi/tbx9CjKnZBb43xHi4kuHNV22/TPEp5b7V7USZQEBsMg7BKU
o5Y61OzvIDq2EeOu8xaIpQ8uEbVFKusuATZ92cjbCrtAPNG3bt+zO0lA/Dft/8AZFear+xx5JJqx
b7sdzdAXkCDqErgpPWAcE7nW3UiR3xPYytAlWweiG52yCDlvxyJOfS2TN8r47djwxkiOZA+Wud64
zr4uYUcd1ag0cvqKM8WD+LBd/hNRPcVLIn2h8zXbbGmq99LUCIGNCYBtIWnANOLdkXrKIR8uF2Av
2nz6b7xzWQDweQ4rMWrmKi11EvHCgHtiTgWYo/o6exMMF7WEJ1KG/zwyLuFPHzloMG3cbDjJzu/l
K4rYRFoj9G7UHRDUIVa2M9zFJr7r1NsViqkynHJpWc8OhN0xNtcS0K6bxdBBLTDY5p15ovAkirY0
UW1WODx6LMs6YnrqxTvb1xPEaD4pm9pkMS+ecJ6v5fWsDzrphw1pLkjJYE/QVJkvCHczW16tQTYY
boW1wJSZR50yIFv0/lDmmBztVyZ7Oq+C/xu2u0rNlsKEApZZSmvnqyfM9NDR6MFVKBsNPNHBRBdZ
+ts8DKb1j/avWaDpwXjBwkt3F/TIXM0oHwOB7eDPQzQG3ylm36GQRtRnNEp4Zsqeaiagkja6aJ2m
+g/f2ahoNaFY2Y3GP4jsg/yaIdW2QHHIiMwtTm73HVnR5PUdXfaPrih5NDrdUvSxXFFrLYrzDBI4
ar98ef/FYPHhppHn2hr2/7Kqbglx2uPldoKXeB4DSqGHg1Ot4426j760TAecKuR8cnaY6bRb2Otn
s64Pf4whhxrHThdEuSCIi+mbuzIMiMpueUFTizKW6G+rtPvO24Z3PrhRAkEpx1N07nwYbcnFl+ph
ZiaMgUU2GW4z4FxcHVFUVjsCTggG04phdptghWP03OpDKpvGW6koKeTbw1lXGPgm/wxDklW3vkvO
GIs9raqvVHsbZ0guUlKHePJj/X3YirgyEN6IDonujOBwsLnCF5ZppFZpiWOXnpMXMR0TTkUK3ajU
ugDdslytdPOmrHAInN+NusZDBvJb+nIpEYV49UKVCVEEkRuX/k6Vcc9HoWko+m9jhMbeozxBTlT0
1CeUykJet9ec3XR2d0WQUQ1smeQ0ka93agnSsyTyW3+rL+KCY8iqcvCHywP5e4R05wD/B6wFyWej
3hySf0+jn9fNe3z8etZ//c22ZG+Uj6UskENK9pxbfNgpUu0siC+gsIBAGcXWW6yyK1YsagQhv4m9
Z5go1950BocCPcLarQQRoDaHOngABXG8Qwxg25W5XlqjMp2eVOhs1BqT4x62DSii/bmyyX39Jt8d
S663F8VO/IxQocWAUe2h4BReu6TMqUKe4fJ6Byxtqe9wyT0+0hZUcDIqSvabyu9LCpNeK3+X6bDv
pFnHPxp4HyJQIaTBgm0nokhi66SU/lg+M+Tmz5u1IV5gkVQlscW5dpB6qRUtJ14CvzP7cTFfgFl/
1vm8Xk2KcBlTCIir/MN9c8ClLboTx+nszM/X3gfZG5zK9vBSrtwuvOkVgRdyUtwE10cql0BVipHJ
l7ztQx1ay4WYDOrz+oF17DLGopmJQ00mQm4DWPRPFwqd8NqJTo4oXwqciwAXsfZ3XARBJc5XHe7A
3zQSyC7acAIhnRR16/lDvNoevgXbuWO7GxMyRvbu0hMkPRKoSoOm1bYhGG6OnbrlHZc6l6D72lQD
7RmJ0lCA4k40Aq80fKeZ1ta+mLCttqVtm39nmBvlJ6TV5iEJ5XWPFCKfeA6Y3xlsZaqvcJOodXVU
zj27tt6cnOgAUZv5agQ7DHox5CiNnQGtXFNfVQGu4nH2sXySMaGgYLDYa93zDOIC6ofqxL5CjZ9P
c5QvgWKHw2oSFIgBf8c9H+/h/L4FqASivg9CO28IhTSbYNUmIG1OsVO42SpEqTJmrs3/nLY62OT9
+cfboPHD8rtm+DykyzFuUJHbM0MZMw8bJh/mENjvT3J7DUcp/OUT3ckj+IKFvibFfxgJJt+AnjN7
NFAXjEtOCj7ARs16tlqvVum/kbH701Vuvs/DFyG5zRazZ2DS4KfRfQ5NKy9aWyWp4QkFDWpsaFdU
1Qbg9YPL0yiIVxzFt0SV/7Qcmh63fNL/KfLva+kA5/j0BLRzYC/zhi3MEAXz7bFRAflD8WIMdRc/
Q6MURoC2oKxYzXRyK9O5TIKfeCb/L7gqvrejhx9tmOjM73M18Wq0SUI4sYuT3ygaBvuNO4IoQscq
l73ICsEwPa4Iyw9ykA5s4HqDQ+hG9F6k57g/bLoodCdeQ8dFsPkYE/0kZKKjyGnnq67Szs6zwoBe
0dQkuQ5kuPPArUK4wZQjNDR4mpcyLr25CAmNT/QHEiTJDBhyjlYWk06hSDm/HW17E4lnhSd3OXH3
k+yN40ugjtIOpa7MQb2NDNK+qxGvzJr9R5LCWp1GYaeq85EbyYct5jAa2mOTsrwzawzuh8O42Ha8
/e1R7DURDkRnM2b5f4Gaky5CkwUbjaoEc7A0aHUuv+s+xJKatKTgiEYMmL3U4INphiQdl3eBWaKg
xhF/sR8KJOV8gR5EykG57a2RiGjwHHTYIK1vQdPK461Hj6cNuySfhMpeuAwDgwKl5V7pmICRhgIY
Ex7nwRurWPHTXyzeok92/w81t6qdOMveew5c5a80zCZu7wPFCq6eS2w9305IJrcXuLvyA8WlkbnW
jHdrk9EPBI+cX0O0UyFUDGxKc3hg/ixlow6OfANLCN9B3ohy6RGY6vliEdU/9eAiKteWQ2VbC6Eu
NRZq+ZkDqUjZeRnnX2vBFDSRQlbMR/w8U9j3yjxvUTd0i8Yg46XGGz/A0Bjud7B9axCQFlNgPI0b
/O9DptOfpEiTZ1Xa6VTXqgMPo4ngzGUQT5zYzX7/5BALl+/eN5uErt0xc6erevvK0w4YXiqYiyMj
WUtS/yMUFDkUYwxVyR0vnASrp04q8Jrd/O3UyNku91F69fOjz9qNGHOwtQbMr+c3e5i02HBVS1+S
c1BtGwEkSrml7RUR8IHB9FQXlMLMxvdvKfa1jDwXuIFw8yGLejCwCU8R3d63L++MuhwrN+bHLYO/
tCyuUItn5YuFW6m1sh2bhCsw3mafckAYBaRPBBitUH3zjtvgZUIKp4IFpB69FJZ1kQ3mFqUhHHSO
nbWz3HeXUI12kUDVYJGHeLepFNPrQMi8RJYfYJA4jwUdA8/zgIjDTTsF75rrj22T+/vu7v843zYC
OHqrksAmC/ax8jLpYX9FaHJlrw4G0SMgnM/CZ9ZOKh+QM89eYUPVW8SmBOZDzgY9UshvEpuA5uco
AYSwt9MB1nsfKQL7ngEqdyW1z/v44fTIgVbkBaok1cIRgNeSmhGDep216Sv5l5f+UunLmk/BOzn1
pIsd8bBDOjMYRiBmY/k2R6FLIFGlDqmIt/OYWyVaXCjgBgdZll+qVg3ghYu2dMSPwb7lorv4jt5f
8wdUcfxu/6/oKy1n8RkTOgMK9W9qf7s/pkRR9JqwzueMxlg9inH2Bk4MRZEHuNZ3w7Vb5Qjrew3B
5uuZ00UB8dpnC7BLj7LuzN6Jkj1YBliWryhcfqm8F1JK7slVh4NMJcSgFLHYlF4zl/6qfx9cqkVY
x0W6ddu6+xMzafXmwTF8i1faRNUsmoi8+WdNEgoE4UBmREyJTmNUIRnZR89hHS2ElSO81cTiBcj3
KImv3Ps83oX1jiRJlkfNewDT2tcMF8lieoxJQzzNqmHFb6rImpkPbjw6zv6MCEK9fYwfTqFXs7Km
/JkuH27Wq3hCx855xOMEk9L1K5b8VM8N/zxGmzpeNQtzaSKjiTqizO8oeOwInnUeooq6yrVLwA6L
g2UWY7fA2CYFTGFuyS+3wdCREhJjaDxrNdHk/6HNlhdgIm3n5//B9n6qnSNi/N3B/SQJDoJxlLD8
KV9UxePgzg7pF8rnM3GrfxsyYHgo7no8Lv559pS1MgrhxZFPsZZM/5iYpcE6Jb8yaFMnLKX90KlH
aYosCryeeV2JsKyI1aQn8zEyB1noJ0DyFTAe0Akq7CgVGO8VT24nrUpijGGPfHqGkaAE1DLoGHP2
lHlmbN0iGgJ3tHqhkfsCsPeZZFI28wp36vr8w/+Jk0SvXJH5s5jCTitrcJ+4UFdyC2xyI28XfVHs
IBnGPv+JIqSp3lq4LoYT/zsTilF88xd303iTULu44yyJ1G+gxig7PmsKy2op4Oftfm8HB5Vr4jP7
xm6SNs6RR5zNd0sVIacDl3dVjQUxh/kBhax6wEutJf0h4ekQCgAAazejw5+6aVymcE3HxDnCgeXV
7zh0Kq20TMIcTsZEQcfY8DLgHuMo3/2yc/yf0kjxP0AJHI57M+AOm+nr6lmFFb2VFAZGyQ4PcM4U
mss1+1rDXdv5RDkHWBmjIVfPw+ACB14rsH8J37vvjzOLpxPF0bpVj3msciEX3poJIrBiApzYSdkm
QK6PsRm9jE1vB/6yHGNdOOI/QUuAdKt12nmLom328KhIGynVefqtT2TfgeOEcEXv+wgF9ZRI10UL
CfvmqC6f/Ug/9Tc2ub0qaJ9vhk88UbYJopZhoEKqpo1VhWKuTN5zRvKW6OCf35V9Tabw3YqGptJ4
nDyeWWqg9/471cmoIbdPWhTcqMoyKsu5pCyg1UIuCMK0Fxgf7Gj6yTqTDN2Gbos6lEzmKZRSvcBQ
a4rxvL1ps227CgUJHPQPAxJPt1snBvgab5fUdjkHU3/rVZ5K8uP/lsL91imEcIysJtyi3S1Ym94c
ENP5O13+NulN3eI5vp2XF5PiEXjjag2s+va2tmiVeS28T5VyWQikjd0Xe1jSFRlpYB4elCiV8Nj5
j4eu8fQmZcBY5SOLpHFdr2Owz5roMRzCc3W2AnkfVcbjbD14ubeBxXejjNn7jGCuwBNkgwgycp3f
/inxThwxBkDWFgn0kpOfexgF7BaUI0moLbKaRyfUG06nZSaaVrAgOua+hW5xig2BN8JFEaulsgS6
TpiYqbNxnT6bRF2OJytoakY1Vl11YF5qRWMZaXF0Mz3MLNRXHJwq5Yp5JxSv0OxzzdgWCmNyjkiY
kQfPLRFPKTnVO+o/raMwdQdew1l6lgRE/XK+6Ekg/9uWNn97JS+NSW88D/YqaUhKh4JwV3L57oiQ
0Pu4Ja6XgVPNq8MK/J+drNQXaRZHfApmlRTUFrHjkBYbmyh18PwtUCQfzh8xbD7ywnJWameWUnj/
XvvYyXFiELJ/hEVVlXlwCTvb8OPL87FhG0xIG1AmzQ5Rr9TONv1m8w9NaOKgEqj5bVPX5HO+jM/B
B1bu8ClvqFIv9XqPwwA06L+ReFIDPMuG3dtuQqQXpKr0Wy+DsDN7gI3+EhQllS3Qy1ZNBAhbRp2n
gg46uUUBwtyMccCEpo0Gn9f6Du2bNdj9aPck1fmnGUMYWNyAs6RSgtl5ZR0MH0JJlwKMhwm6D28e
m6YhwNmIh+0NdrFiBtMrJWRWYXPd+Z4l3dgasZkvx8Y3EUvkBGUqGgGlfgo1kc/7am4QaUrsBmpn
zIW8C1n9FmtL/84vSlsDqggfadqD24c9pzD39+WGgg9JDn7lETMz2B6foDiyuddCiOoVJZrLWch2
Tit+pqCqCjlFRQzdpCNpe4T0Bhpgbc1/O2Fs1po//k/U0annnhBP7Weaw+Qc/Ne/JY1J8qcXbSYO
MsIv2GEohaA9EspKC6NKkTOj6z3FPvdMM4AWOqi/cfpz5oG5NE0ggFL/TX1/2+PiO5XMHvnrm1Dv
2Cf7fEICif8Ojr1Zstu8NaxRuDBtO9s2IAaE0qgwvSifiEDVT0Bh2Kgfe2uNCwUYUXT+1PEyl9vr
fkgYpslYrZ95o/2yKDyloBv6/8k1LnE3KGkvkromB0iYW2XEixcHrjGOI6rbfluN/vELHjX7lKM/
0pfaVhF6V+keu1MmqXy0JSSFgnjIL0yBw15h7dZZPLpF9QYrFZzWxiQhIbPa69t170JzehUKqid/
WYGyIXrLAmTBfrMg+Sl84XhObrYjYjIx3Q3WWdfCPih+Y8ktK7wRK8+BzYz2qCSZ3dPqrSHenYLY
4mwvN6wxL1AAdiy3+t6oNK9fdFreVPjzVezgeADB2UkWxakZ0d7XU2Wiqsmt+jdwhkK74O3NEhX/
qYjXmDlIHT4en77jrtMj5xq51ID21BXRQ9AAkFXZrXyd5jHi0+ZxOUEQH6obxkB0iKPd8JeffoWc
C9Xg03c95J9oYJOYdZKnSGMjStMQUjDX3+GiO+lPXJey/nBvDXAieGM53NSEab1uiiZ3cPpHWQTo
9R88HcCJYSjjYO+a+g4t48IpbL7HSaU6NZc//gNd+a7ziq7zLkolagaYJGcEjJ3n41O1/Ax8X6UJ
W1B1NikS/5GUuY/fIl4wUljN0c2OfCFAR1Eg45LtwigHQz07N9H/KC5sDjhX3EXh6Bo1kWY6Trkl
Jv62lskcAAJ9cFCfZXwVyjBOZwlQ1xX8T7OHVL8SX/HddRl+VawEODnkwIjywejM+8olqW6h3wjD
WVxwM+Lnq0npp2ortrKZ7UwI0bn45CO3NWB4asOa0pZ1mnQWauxv9iUkpui8BlCkCSHnN9VkSWsB
Ba/ONM88b7wnXZWhba9yv5yRdZ+oV6v6LMH+GgLbL/Y73f/Yp87QI0nC5Hr+NpEOi/3WzfI6Fhzb
pMmtjmcsZOQqN84K37qnDRVxvrDyQUefjinafi2kUsMU8MwHLP0KSJlphyZNxV1gdaqa0StZkapQ
kZ6BWRNGYNR5Z77WZtsdc62aHUpW7cw4QAHqgFh2yZmx146a6sd3QVq2vd6hheM/P60dqfHnm4ks
5uRqxJMQiB+NB1Adiy/Vm1ZTjqPhLH2dl7wf4YgbFO8pTALN2iWSDVg36Zjr4BFcVnBI97wjkFjj
//YoMPb8FUGNijgxonSFIX/53sqrh5kfy1FdmEA7pAb7+pH+J6RATXw8WQty4NiARYalazXh4M/S
jcx/xWUvONpMxs1LoVEghZrGSTB4Tu1h94Lc2ZSwJf2FGMMsd7ik296VyRRjGQSIyOQs+N53PlVn
gncXqhteNpPxECFbOQFWwzYfLX9Q7E8hnvziE1d+uFVk091tQbAOhOJkQG76FRxkpSeT9Vh/y0/6
BPzaxWgGWMigl1K3CpmVx4fS6r3+xeFhfEFvxy53Qw2vAgKjqtv1989gV0bHf94kydS2o+n4hmy2
u3MlClYBSc2ajjviVnUa3s5Nvdd3jfjh9Q7TQjA/LXdsFKsX9wpUofG03O1TDmNbUbbhhR2igKUN
Xeu0srAfXF1BkTjHasN3frWscDsD7ViW6xjsC3uHwyfWm81NJkwwRdIw+oS2oU8mlt4OZ5sjAfi3
M9ITd1cB4l8ZRQrWjF/skFF+7jcmijmMWd71mNFqfUU2U9I6D+8eYQMRL6k9in9hR47QOB+KlwGx
9lBfv78o/ewFS5oX+W1b1tSgiIkofUSxppmX2bavUvp3H98/FhzL2LinReOMwAGaniLTLtlJq/5l
iBiNKFa31G5onxuqyZZIiChh5ZBtQtwNtgbCwllwAAhiJht3LEddRDcyPd0JURQ/RAMckhCT1Ffq
n9uc4vCbrdWXVsKiCtkCSEBwcXqLnXtugoGNGuyqZNshzm8h/NzsiZ0l9T802j2b/KcfUaH8m/pZ
cQQsJGlh2M9UxMsyHqPusqTZDx3cEypnxpMMowtMipxtbgT5Al6k/F9/ezNa5nu2z+V+Rp6wRham
fuaDeKouy3eHpHw78XO6rhKMvT6Ur/79HSbQUe+ryOlbgqc/q32uRlVcS+rE4U2aWCfZxBuGwRJ6
zG6CZSn1g99qDW2krYcTOMJEJUihomGNf7Nq4k0TG4fBvUQUfa9SrOWtt66W0KvDig7698ENdN1l
Bd9hK2wcXhmS+wjkGDDdej0XZ4Hvi6WvHueGidDbrvDlsZ0KjPtbimG38WAQ9Cd+m1abnAOs63sn
OytEefBSkVUuHlQNk+Jo4INnr1MrpBM+5yb8s48Yjz0pes+B+wlaNBBoaX3hFeV/A6xcnIGnfimH
MRgoUr+36f3UUfwvCIxEyWHXiRMdZwwX4CbQS5YYn2h5sG1oAbrHsoH4BUKr/fzsxYkWOHTdd5Uc
cJBeCfb7Pk9BjYve1JUWhydoWM0c3gJFo9q+XzyINCyyhtSzKU51SKytSNaqSiZbdh0dHz33yUAm
zqztzGErwV6XZPFPUJppd/UR+6olI1RpXkvGxdgvI6BktWuVsVNwT8h7DjCZqWCiyOyZKBPNlFJd
gGROlerTPGXk5flRRRfNzP0y7KucpQc1QpHcNeUp32+voHroEBOfstSw3XpfWXDQBUx4lwqfVKQx
2iNBL+Bu812RXmZN7odvJhU3gOv2kWA3NprDqD0jiWLUiCFZ48HenFGhHebPNtbumhy1rBH2ld0j
CCTrvPfDWCLqoAoFamoZZfpNAbrs478/P3N9NADoNoKz5NQz5tMRT4EEo1JWRDwX9j64NqgA31Ox
q729sti273uLjCjv1J5YVozgE4N88sBgoSdHHtSytxmvPUo5T0TTqeN3iXozL/6Ftk8fenLIdtXP
02Z8f2/ZTqu7kES0d4NEKfAc1TEXQ6PqCuPkTmlxK8N8f3fNo93F1zRraATQnp0Rdsx+TF/Th4rf
C5Q1f8n8h8ZTrR1XyeM+AqbbBp0NYeVZmPU436VGhcDRKErYgF8+Wcr9UpM7DM9k6hYvrWe9Pucv
a5MAc9rYzdvPjuU5FtnSDHfYGxB3ezIHXh9Q5pH+3phmPMU3uADO9RKW5OdwoYqDAoOBXsIL5/Mp
YKbEOU/yHphT1wWQ5J7Mz97WOBoHNemYXFOep3zgobn2cu5VbUulVz/0ExiV1eOVULXW+d0qME6q
0Rys9/RrjbdDcCMhHIjM+kDgcKORM9y3/52613XdY9LRuyInyx+PcJ3AW3pyiyXmOl393rD3b5G1
RsuK/CsqoPko9WPFvMNgCyyI0EBf4tQtTeLysdeGwbq5ht02TTziFN3DL3vj7Yt8lMdnr8Kvqt8k
vMah+lMe0zZO6G+MvruN8nHXmfUe6yYhYhYQRS+ALQHpDRMqWCNcMefoMOrdn2h/lvxg/W8c0p7t
tQq0V75zywH0Q967bb6dC0Zgt5gbCPgenl5ZvjOWVLoFTpf+SBHVJ0sY6O2ezEsiAi9A+sUU+b4o
W+KQPxXGIz9m0w9YkK8cJUCRaoZOsK3lxzvNvst2oxgSdptFCHFLtBS1MXg7U3kGHgFyAOkQuUeA
5wlbexqO/eGrwb5TQxF22rdp559x0RjtCK8qQs+dvm0qH+M55kR4QbSdxIEtTy+shx7kJVMixdRe
kb9dyqE9DzMRQwT9IeoUdX0P03Ygf8slHbyN/Wn/CCXUGiCoTQijpWAU53b13gZsRtK35aRo9CEV
Yb1bMIMmaxW/zS2XR6/i6mMp9AAUMDYzwnjiglBuEARZzllyYybVD+3GyqTnfzpb45y3vz//MK6l
by2JmhNnHPVuimcq6V84SK4f84/3WDXiNgpNjwLRhRm4AftELN8hYGyu+O2aRmb5VqcrYbTQjIa3
crQUNdWaWrenkqVkDUgnOfL4Pm3t1YLvV7P4NoubRxjuQ73bCFmKgcPlanoU5YIjJZl2dkew33wS
QZqOgtJqDpwgtRk1hHvhh4siMs4D4XoexhURk8uBmWL/jnOrVQbGObCAUaIvLRsqOo+ueYX4e6Qd
L+wCQlrxNugv54ro3ioUObd5QZUzuoHOCff4zykQxKFxr3fWA/D1yH+A44fzFcpfQpmbbnlc4/+4
EtalD6HHyx4zRkLOzOra2RsfzPnvFw8zvCaJ3t4OzEv0aYFMiwJeIGuVv/o5B0dCMJ15j9937kB9
cME9+qFER8BrcrbGjCrDOmuQEK/BG8ri2CSUa6eqDEOOWfF/AL1RVA32N51/4VZLF1w8A9kouKsZ
K6ZZUAv4iQbRo+5jqPfvuoqQddeNApdUeMTeQCAO0ezugVNeHxgCoLOSjNnqS08bACVNvl6CVh9r
wvVK4YdG1OSVwhshX+EMYXNyEaG2eUbiPQVUbZDaX4cQC5ST1A33AfxxAp0mcEjYWDTfKHSRgHa5
QZALE7gx4y9e/d/+8zzG6Br8Du1NL10aV12kNc+iIp99Nqn6ZCsJhoMRupX5EvKS78IkE0+xz3/6
MCMbOBuE9wClyXuFfd1/Veui7sRjs4XwCrtKos4yhg9t0V1ECKYbpxmlR05Y3v9xdFaPJBqjjGd4
nDXC3LPGE+s/RQYd6DdYlMW8dnRKijPMq/Pb5DFs46P3pxvTq7dzJUsggcIBhI8aNSwzaB8TDd5t
42hRuKZvPS3E1bXYmorvtIMBP8Qr6paahEsoU7I1zKtgQZXWjyAfadvlEYHfvRHpBOs75VvAOtuj
9uR/tUZS5iuvza3XlmFmANwu4nBdLnepGjSzAs/2jrsEMLy5J/6XzHbNo8dtl9NRzynuDimLRm0D
O+u7JxVdzcb1fn6MVbMytMtgn9oMt42LrKNhR6QKfEiyqvRLDNcclpfMcMWCHc7BLgujKXJ3cPKK
npxDqedDV13mt5RBHB9GvU7jEV8bscHamMoTmt3/NE550ygnvfUGHAS6sJ5UXfm5FjZ6gn2xGkat
8+ki/oVGg6h2TpGbAGjPMjXRdUDIMaOij6oBPoFf5eBqyr1HTVlfMIC6YbGbK1LVzbsFlxeEQlKR
9gylYLRbC/EX/MHMQcPgrCzT6K9tfaffCiGDWkhex9jvIf+6GuPjU/LZvq2+SC6pXTHElFP144Qq
tQ68Z8PCLTltrN/UfoheebqHeJKlvE16+Czq+KAGyL7gjTaCnaRZ906n+AmUilE8sGn7uqP07Z+b
ZMvh9AJPOCw9rCgCtAn6U2gsZ6qlUL78eFCjwfV/nFG3v/98Ubr9LZsGdF//y0Z4QcK1/08q6XJQ
qN84UZZvZEsrm3DcEcfDEwz8IttpD8V+fz765WPIW9PB2DaiB0dP3dYCTVgYTa48K/93JnxWo7g0
2tSfpxBRmZH1W0cg+wVJfOnI97k+72vjrErYqfhojKlp9/As7vcD7qIhcItuwvLq19iGi0kCgBf+
5m+uJi3L1thFED7hbj24AZDxnl0DSjoIMghc5Gp2cVlwFa38XWbTXR3CBH+aIn7+DmunXN1l+eEc
T5xzj/gWvx5nsaXHwzN8iIMx7Gf5W9jfaWNGoVmrXaoLxDnj1tjWVHHePERDnd88rRVpNw5qrJNX
Cz77tuahcwEC0eJ1I8KdAnfWkpG/q0lB5XxAs6bNCpImPf9MASKqlZhxwHigFER6fJO4eeunBU42
OWPlcAJEoEyI+mHcOukTEMBMuMbGMTu9AG2XNX+ksr5WseQFAPlWwgwDEs+JYNUQJGMLSRy3+LNy
oDOCs1HHupsOfWJKUT+HaE4iwK5FSH2AvxdM9R0l6yR9hQVj1+dYjQvwsKo2h9leXpJH/LSwY5yt
Q6QP3XVePBkCrqJ6lv5JYKnHaNLcZsITi1xvJXaYPsApS7ikenLhVIMAuVcbkSi5BTIVEPKgqkzV
HLidpbQOCKmjqYfmVXCjGuRxFMlk5+AjhIq+4VmbVMjMpEmUAM1JJbrmne/KXLRWiVwxHE8OGsMa
oTJPpLZaZp+RqF7Kbfi28v5PSTsIxC5qxubjP29msLdExieTWwGFcTFqEG9RhT49kAcnMxrEguzf
jQXBRyjsEUL5gRphjbhrERyhN/2EbxXxCgx4lXoL/XPm/p6xbcPK31aquFEzmcYRJ6PnjbKbjfTF
8INEW8XLE4lxDFOxoUhk507tc3XRK87KQDIPqED+uo07YSMr0Nv7DsObGLjQTIsT3hyKyp2Iqdom
FtvtCv3ulbgdGp8NTOcUo7BrpaWFKsAN6QzMzSjQBz0pJjBP88ckgT+08WT8rb8BnLvPjM+Fe4FG
wTOAO4Oj7b+pUa7lKsjYUjyO8ELnlwOLS/LRUGKkf6dSp+omafFRKWIZ5wFeMUMCwC9cTvLNJ7hL
cXgoy5TLZocC/Q1CF96huqw+6iGaXLjf/7AmTVwbJ8k/vw7XXhbpGvsQRR7h6XdNkQA5LfhbYrus
UTdxl48sfx/M4c1L3OJ4lOTTgGlBqaCKA2dKCe72XurWW+JMmgZqwJzissNJixkMH7hgycXEDcTy
qK5vn8tDy0+PIyMSY94dzRY/+traAOzOTr2PRIeB7CP5amJYuWvqk/+VLFgLAA1vxHYSu6iVu1nb
EDAf/OuD34uR1ZaIg4ET/kAk+vgsjQ/neUpq6dGXrh7Poj5AQ8p67hkp09VIMZpGjuHy9CbR37ra
abIchN7aH8DZuOVUxrVUD4O0IseJuDE7l1ED+NuF3k1AeKd67IHb99yDW7su+OIIV+mzHaGYlOEV
6HtAmooChu5uG0SCakvsioVc4nY5nSrgw1bmNssh4PAyZSqeC72YWvdhGzSE27XwIQYDs4vtG+7f
6rt1Im+YQ/c51mTWzOgzefzzoXDrWJcc4p9OX05xrER1f0rmSpf0V8hSj1spuicBPrrHGCn73y4H
2VeLH2hl/VBSicftDTTEeIezKwMq6wqijNTCVe0xfHd9ZY5y93MHABUhlB/QuweDp36dlM5znr4s
MeLkxXiqx2/7RculJT7dugtCpfQdIuU+fOEy3+IKaUj0fYkAtSQTQYcxr+wAY+0ryrdhdIo8TOke
Z/jQHX33zo0pxs+H4Pjwa6F8C946UYCTtyGlimlYOU3lnp4x8mpNnCSso8pMLsghkMWnlO0cK1a0
OXQIld9tO2HPei5fS9pZjSd20t4Lj39ideQQff0ju7mIEL06M35MafEUpd59Gvf7FUlbFxvh8TzV
lM8yn+zM8NhUjHunELuNsGjBD/gFVfaPMGbNc//bbHUVRIFHOBNa2H6ro8vefozzhW7xqUyr1529
s36i2A1BljJ1AqERATYQuZASee2pO0NY+rtkY3RRaxz/k90cKb3fTq8Ttlh8mjjanQR+EXhSLmIQ
zXX+eDq3k70qZFSM4oEjP4C1U6cJZmUt6H6uFkHHOlNGb4S2PmwoQUfCawLzaK6PVSL1W2UmEFH6
cBS+8Av2WvNNU3AXMBsQmO2YOqJF+XwP5XeJUPMubqeaPfNb3KEI9ulXKIu/c0fQjVXzSxZCtLyQ
ZDlSHdkwG3dJDsyZ48pgolkbySfhFxLTuBmbOu6j7jsOQN1yaSoutZTwPYS6nTGAPDltOPzVesMl
iUOV0aggwgAClBqaiThsKyKAfmVEeQaggVnYhj0NzBsKWGMlhpFeqahZi8slAaMXnG2G0udiNmQn
Ndoja2QhphWgX0oCALMBzPQYWdADUN/IwH5B1c+kf1AcBd+8B7JulpRIZKcmxRvnXVIOaGBzfVTT
Utb+f0JkmF7V9+sOys5b9kjY9ln7IG4c4axPvxf/uTbpDwuwsZy6Lo0BaYZ04bCj9h3aUaDCfBy7
pKP8BeAzwYSdJFolU9AszaCHJMFLj0Za4Y3RXBCo2pgVqpLpC/pG5BlfT2TrJkm1Wba+fl1D1WX6
YDZKhzUQt9SogibDegEtMZvzF3WiJHREq2+HboRGtwypzd0fDBDcEb1UnfQ9RtPCJZOucrNsK1gv
uj3IhjVi1/uUQKsMJZ951ZK/wQ4imxZdDJp8fGFkirJAE2oV16Eke6Dk81zye2FyI6ryt7SSuxIq
eN7qqZTIdSOSOSEjRH7u7BVLqjlJlvZZbZGoTAze/9niJktsUYir5hcdAfROdpiHg3+jf+lk2Qoz
hqG74YxV3YvN9/PEf4gS2vCyhX5S94Pv+ga4vITkeuhbDsGMGvnCVbGQbCPKYDpkS1VgGy71r9vR
fL/g44EO0CYM86CIkGad8R3IBdjGbrJCKohW2muWZnV7B8UciAbuCKK90HgxBjdc9bUs2NfJR0t5
jd56EVxqGleyR7TxL+0yPTJ7FGJcNeEtLj6pQaH5Y7szgULC4pHGB/fLOvUcpBDLVejeAf6zGRdg
l/f1nhxakZhPAASGDjp7b4FZI9gKMJP/NYeIKhC27iKwjgapZ//zJ8NfUAhQLHipB0k4k6TIv+pn
qJff+q+IoFREOVnZFvVfJPz7d+ge0dh/OURWX2Yaaq9DbkvI58wKBotLkv48pf94/cyhf5DfYMBW
RBn3z/u9f6/RN+GRIKOA+MwbPpsDcQCfx37KVFNOW6pscRP5Qz4sGTOFHtk7ufzXHRssDDWx8UFq
CEQ/tIZXwWIDKmtAW+hNkqecAPI3UqWjmoTGtYK2Hi7bg+sDWtMPkvnoc6FWwyOTc9C1ul9qsOUn
yVT6kHTc8IAT4701Xjze5Z84jxB+xqM9xJrMivfzM4Wp4s2LJhvxIa8uRwaO2OJUK0w4xOmQiYPF
I9RdpDsu3gv3bMxjQbUiOQCrMUrf9HFaFInfx5s3GsYGRaRHmD5Bh8sfZTUb1tzGD7BsiJPClWDn
Q+SpGS+/illVLN2JirFFwFYvmRS3JOytVgI5WBrSwJEoUObGIYk3G6jgXl53vFjQsswtq/NJY9X9
QEcJCltulCqgmUHIkLDBGhZJWJrHWMsLtT7aNgnyw3f5bwV3VmygAd0I2IAF9YhK6TowJCfzsmbG
VjKfO+Vog/y6kDW4/fDXBh90o8IIaZmUajbcUpwElI1snWkPch+YZPfd5n11myGpOg3I+r+ERrX4
7jQqwJWSA5adI2k+rM5QbG5m9r3g8WNxxUx6MDj5G1NoYwnI9wVhx433hMISZnJ+Eu26QPSJrBUu
XDZUYkaUI3YBTPQJeXKTMAyrr+lRmMIDc2oj6/GhizRqKfJVCKLWtnG/satCfg+VrknNemQoRsq2
6812Sw7l1cY5tt2mv2C5Y3cr72DPnpeFoxtG58rUdSetFFuJJa39Jxav35GxfltBG6b75VptFWMC
DW/4mDyhbAHepQBVgX6Gyu4SpU0LERA8spdQGLnUIVIqxu0GwWfLgyk+YNuLE2dbRMErbawyrvHh
XM+bIkbPE5KPAjdOfChnYLCwTUzZhcPeHCH35vsL+865IyEKGlqbg+sPCOOej0oXTnhkIizH8zRW
5pomtDxANGLaUuOLEyOPWzucGYUfAnqIG0UODJ606u/UtDefW5TMPFCruhjgXKddI2SaiNhdjUvz
SzfOfo5GrVkcSNskJywKGn199UoHnMX6A6vStPrhRbqF5nC2vVvvcPnHLXW/NJFkwKPt+0zOb2xV
rbJ/A+ZS2g6f0vI8pn378ugv/N2CcFAdoCQSat0mjLdWdFudutKQCQHX3My1zZoKEkziWtHDICPj
m2lreVUjQ+7llE0IvTdJ5lb6OWLiORWxmeRrfwWKVKefdNMaYUwL2a4P0w7oWuaQReEfF2dBLDFz
POJv9WRXvliFqCsea4n1/DBllPGNQlsfEhezm3tmWsC/0G1LLUUyRDxFlVVnhPsfDE2pYSJnn/HA
kWqGQqWR12veAtky3Wt/je14024y+CtWy79CXV5uq1ivKvPDxg9xv9bJdbT3PZTmASvmbiNFussu
RpBs0piVZARtlz3JHxHegW41T8SNWJBTs0s6amUd2CpTUhVsMmY4cr83Du+GtiTn9PIY4nYQYsqS
VFBaA69Yw8/AGo9j/gGiqoALpRfnhawf0g/V6jbw8fE4KhpOaGmIKwuLVjnluMwf/ukTcwEnTsP9
7BmNGO5pFimgmi9UeTnGYgmFOjV7Zqy41bzxQSpV8BU727cw9r9aG6FzvAaeA6TLohrPMdmsd9oF
wgGynoa+B8k9U7DFWRffjuuiWwqIs+L3bLnM9TmaqOjDbi5Nn6RMZ76ZntUswdg4l4wK2cfrCrDI
jFqesI27tOwZKl87BYh1tcKrV0P0DBwHf7272Mnp8N2jwlKaRynxyqgq/+4bjmlN9WBfS1iGpfWO
AhPgmi50kfyxbjd72NwB/4IanWXF1SnAopVCWKSs83DXxgTBDP/DFz3A3/cc5vUozHrVYKljELey
H7z0qytCvBHtA0N28oko7HSEBXVDxJMuqBJhJb+G6kISt0M0edEqvQuac8Q3zpaLKIe0XGIbHc+q
o+d78SHNHTvB/uE1d4q89jjZ5T27n4CKPBviaMDDn0zxZKxX3fGpAsJF0PLAcBAW1xqu5W26kMK+
ablrW4Aj8+G+qIQXsr0TuIZJvYJhuaDg81cE0mpDD2XLYmhZReOB9nZSGeRJx6eA4XOTTyd8JE/1
nPRwRHpNQP1R6dz7G1DprM1wec+biXXQOv4anUYd8fWGWkTK1qw9BaNDBHU+5KEI78uMFeIasSmC
hLMqhNS0N5QNSvF5YTi2PzQAPxvVc8UD52Hbqy3nfGNhiLizsGvyIlVZvBvgVeXr+SZFbAywfhA1
JYiMAGmK5lfF0bMqqBmT2xiVVOkKcIWENsLtRepZpNGfVR8RqPuxzSgB1hvejGCABUYMyohAs7G4
b7StQhdAp074kPvcW1YkaMx3888BU9v3T8Y0vAqWh/MW3X5SPn+lFTNjH+TI7EA4lMjH6KtcLrzv
33FAJOOh8wIxoWOzeGl0ERjSIHlwywG3V3ehiuM0kl+a5UYFn7FNe+6NY+0XQTIZCOpeeu1BH7G6
G38AVYCmPJ1yXqmJDe5TpicYHC+Lwnx0Qak1i4Gd7PlGVfexI1bVw9t/DaT3K0YtobSaN4RZib97
PB+MNGS0lnsYbs4O4IxbkNjs45t/iUKhpRAZ9dXwFaX3RmPivDUaUNQIdffJmZtBjIhF1t4Ko1Yt
LaYFDB/JsFNgzfA59zHmecmkGWHfv6GfW4oGesarTRw1ASqdRydbM2B/aCSz1mLocInP1At6aL1D
XqEdxmeJ12sRPDPucaz1M64/ziuEvRB5Qn1s59gDzUgA+pOx6ETPYOzxeNH8hgkxMJ2fopdsQPuM
0v3xE74VOamnuhU6D232977De5YTEbbYbQPDfIkSsVS+TwgqBP8uPupvn69VgclwSyU9myKI2y0c
kfUeaKRJzX8T3YVFVmRlFbtJn5SWbms0+rCjzVYsm9bh///dfcXehBVSqIh6V+MXyTH/7dJF0D6h
sn1IVUFma5Wk3O3c3FiiveJ7ET0Pea5eeePkuMQZ2ZOBuOjAGtI00//n8k6zDSnf1gWDKWXxOrXA
vxPT9ZC7l0CMgjN8bzxZnMK/q+XuzmDZr3jveNETKMmxETWmtxZSDaN1pzHFHKWB2W1EldSm22ir
Xnx9XTQm2W9v6mwYrz7NdbYQEZjuIHft60jr5aH8APBwaRQ6dFK2mnbZqq0CXAwov+PI2zY653cF
WjmZelQZ5JVazG2JtMSwEcKVGPgyFfpOuTtwk0jjLw+OAH4FFShzjNpQ06UF5u1/Xl20LdyyH6pO
RhXztJFn2L2eFyErB7MMWpUWhnExyPzoKh3chVseZw2/dBPPJSK/SAgjCp0YQ75baatbiN3QpY4w
npvJyKiNJUgKZejrMNzG+JBF1UVB8X60laxdP6xhezmibZGlm0bvg74qP/+1FZBewW4j00czhHJ9
YRm6XRgO3+fO9pkSKpRHaLfTk9Y6BWm/9GRqqDRr23os3HnEPViBuqIR+0ejtz95NlHrUfBSLwuk
jXTjIi6o0RmS0o1zQc3sH8r9q5JA+Fl6NYFcncWGu43qcUw/SB1ZZCjg+W7BUc6iN7sY389CE2H9
N6B/Uj8WtEGhz0m56JISGFR5UoUh6lAnqYALYDflbvAqM+fvR9gDqftNEYPqXs5wzyEzLG0gLkpG
ta1rwMvbc6FLy/vkxjo6HSoaCyOC4E61V5f5Nu2eCosMkexTlkiwGkewJHVUhFyr6vr50papF0rx
QZcgODj6DFUDfaUOqR7wmweN34NSxbNkq9F+VpKgOJLr0rqlnrO7+iRMQAvbwBtvCY6wdkPdteq8
Nv+zCwIrlcpAfJRBWufboNuzKmVK7jkrCCQzavSyACrr8Y4qRZ3duK9n3cV0Qk5NEIKNrv3gB2++
ri7uFj8vwadr63Ah59tWhrelS9KjMVaxyEcJTeHONg+4uvCHwDe6mWbaoGBJIhfI00h23GKXtV8o
AUVfgS6mwXPY4vU9nMffCF7rMYx0v9X52dV+y7dgK8WxXZWSaaqXDnepdHzG0lq4yaIhqIv2wSmm
e51qt+N3NILb2uiK0HkCeHFvDm0pgd/bquoCGfJVnq2f7iSX63g0/EBwHbrvJuaYBBwHLq9bfD7r
J4qW7kWRvuI7ubgeCYLHKX3ke6TQL1wc7hv9YSBnhR6BFHibbGzejAkSfPcOIiTKnQW/sYQP9aSn
L197OeK8XJvCLja9IslfJGVpJye78CaqReTtLsKtk0USJF/nb0YmCvZF3bCDba5yVrPc27JnkVSc
N3IC2owjSR7x+zsFoK+XPRTmUr/9dS3WS8toYeshupGJnSqwx7Tg991WKmuwm5onK8UESGr2fcNO
DXAdaoF1kUwzKRGVKwyPQwg2q1SHCRhBFL7X31ofmd2ezESHeiFIvmnV+d48to0C3YTxpWykOPA2
vh5AVgObatwhx3ILnKaR2vTzx8E22+SV50oijpZXnpJLkMVW5jtcRLHblmuwSMnb+8kAQ5ct4owN
yh0Y51OGlv3cGD7mmjaAA2WBvEFfiET8KfwrgoHVmtFwfAJUAicGORoZ9W2l2DJsadRTTvsAKfQ3
cRahPhNbTrVaVfTD3+U8rwxS1uPm+9Ddg8tNnz6EbW3DrHTvmVRnm1AiXFdsaXJANXrouWUftw9U
RJLlqRB4i4tJc2u4lnEnYauPr8SjN8VVo1ZCzVe4Axr/Shqe6Eg6zBO7yc+oGVopfW4bBHPRAbPv
PjzWRokhwO39rLjhr+7azfEXGI497NZORvoepp26dGKfH62JDOuuYSxyOZL4a8SSwriu+hsfvs4g
U+ZUVA6iivKsyBDX6Dn215m1Rzse2gJ3iH66RrjKbhpu1ociaIwO307yB52zgSb5AoY2t2CK7Vxt
/5Rm0MMuIiiKpMtx4dey3DRwq/0o16af0YMoNQUpaD3s9ZnU3IVRQG1Qw7BFoLp705UocyIZZroC
+mXr+mjRd3iKWdiwBit7Fa9N3X6MHX0s+aU1+MHPM7//gdqRCPpHalVGJakT+P3kxWaI5U6HB+uS
0lGQumoq1POCXwL9K+EGNtitBS7Ro8OFBU6GzToq4ZqGBBpYns9zs2GuLqDrRR4Ph6XQR27FInXQ
nsSZHXc7vC5qtaQ7x46BOFUJA+4snpBBV8yhUSg60gOSEgU+CdWYwgNWQHQLjTbuIQ1oXBpXuqPd
GghWq9mcTOQBovKU6vs22mAcIK+7Syp1A6FKUMShtxDOp+ljFHdKRiNr+A0mBJsa0ePi46Y6hMCY
2i4zfOpIoxVyYUAYekl9vNC58KeYHcZaZNLOPKnZEP3Hf66y5JGRT+ErvhxvyxUz3DMiNgkF6agA
S3vcvg4M0M8HyWT5eujJWAzMC0BcfiqBkxXteoXrp2UdhL6MvO+ljOWjObQtGlPU7ZjP3OjxXQ8Y
M9N2aPE+KtjO5bOGIDhcSz1pvWBlnPlsw27/x3XmYtE8fkPNeSQZGRA8eQNb4nP4eqmEoGFISaO6
8NkC5+ytiai9a/EEpMIvay29ncO4BiTzsf11dE25p7DJgg2yxDuHpkcIOeJtC8t22D2nW8g5DfnD
9/OLXEoa8sIXGTRIsuPT2/A39Z72XLnq2vXTJtPAKggIisIuuyRv7U61zDyjgM+fU3q2ijeCA0Ek
6TRCFKgf9fCqrQl2B+NrB78glnx86tLdCHE6TB7FcEUdJLUO1HHUFpUjZ3GKW6nz7tdT2bPjRD6g
+XUSHJDS1VuZzI31hCKLlhu0qLDTqbFvyKRGEpQ27M4GPbWn/PGswQEUj48pcNdtTz7qWSQvP3yj
VHCL8ixeepkkJiMxhzO8ucCz6vkiypDYkenGw47L1922GAqwwLh9HwUOYezaaglDuPOibGrQVWr9
JV+l4XhOx2y274Lp8zB/f5LPjVKaVFywmW4nKHXxlmlk8QpA6qqJUOZ3yRyexawSiAOY4wDtbKRw
LaMC1QNfT5pHy1t8PN6xg8iu0MMduFcIKeLdTaQ3/IBaGS/63tJdWPnNE6u4YQsERhP42Uu/tIUK
uOhJTvVGNsN8VSPMZAWpL1FizU7UsG8R07O/y3A3bwhzRe2HUEJQE8+JHnWNxzbShnfmsF3k11I7
djTB53bcM+6QJd1m1NNBWq5k12uxZMnKdSlidND0k/ZGGP+l5d7UoHd3P+WssxR647o97aDiZLqE
HyMMHbvH/Ho1/d9RMMgFt0+wJIwBI1m1uTOcvsGjHPuX7sX21SLCamedyfbKb6Ro56jNUZmEXTVw
09rE6NwR1efGTYHpsDyx0qFI0AKMjy+HhDuxOirOJpqWELnK651VGWDXWDdeGoEWy8u5BUhtopBO
uwSy2VBBxFsLXibPRBypm8K7dN6EVDAxCzkuVx4QRUOVyoUZ9nBCR9qTyzSVPTPbTbYzjp7dniss
rtCfW4kpDkIoVX6lZXMlXJml4JTuv3pifE0/6XbzdW/QhrmxmNyQWAzNDZGejgBxo8RZcYEveHCe
4uS9zE35eGLpJ3sZDKWJjBGuUc+/Nu93oFcTCRRspR5IDVZ7XEc7HVcwharmND/0nfkODHZZKgO4
BtHy3rIiidR28sBC6OmsOM2s/KcJpwWU5HQexPqkqhU3qhBRMgos185BXMHmpkkrqS/g61ESbxXK
wbEVZ5Tf7jS83QNhOLLq0rYWtPxBcGJP7+KN1BgsG2bFffMkxQ9Q17+/OuUE3VpL/6JMO+91xWJa
GS6ULCr1qunQoVf/qC5dIxvbuAtLp2sUxmLCVduoAAw23BBNVJBscvHOiy7wc7YGJLjl9wfrVC1T
72+Xcy/3Zf4Dw7Ou6FUwWLRGftlR47pUpCSwgU0+0CbwdHavjXy1/jS/w4Ytyz6MhcUnUujksK64
Lg4FEcKA6FpEWR++6hx8T9fWacIjfv5aUiBxa9oIMPhr2fX9KeSMwBQy32Rg+NS5KQznH+oE5udU
e9BVanyWHVZ2dxrER1IywSXzNHy1Xlp5PP+Fc/0sY4pS/Jngt8tV8iEpMiXM0OQobXiIn1xhkZDc
DCrNLeuPB5QODQOyOYw6jUH6eUvuTUEdzVDOn41zqRMZSRz3O/inLyCSnC5YqJZKC825TVon2wrZ
FOhzLFmbu/R7tJV7QIQCfqyIQuQNLizau1XmfN6/P+M58k8qE3nrTTOzLwsoY2+DLaxrD7v1V6cv
/eKMQ7LHB01BVuy49Wfr2fQqtoB651ZxB3TgDMLlcc9I5jFtgfxJfmLxeU/uGfKavUPQ4MzmYxVd
lKsnjAWb+uqlj5Wdsjj65XnUZiyKxXxnwH6w7/iQjUw3Wxb+ZSlGlUm1imiz2424m8Z6OfTZ4hFC
2F2R8NOr7C3n/d+fy5o2SRX3L/Jv3/L4oMdIQMVwSoh0B1xyl2RGFU96UWSizRji/oUyuWQPBwPW
ONAgc0JC5fFlsN0fsQeJkRuICoCLQD1decyjRYWrzTV9JQNZMyU2KBLgYyir4A2nRy1yuxwJ9PzP
UqT2dLVRSpbqB81YERcs5hY8y2a8+TQaqGMPNAOZDfiH0u6jJEyPwNezFJAv/QqRNCNl4F7W1rB8
2+4GkY2+qmBUeIZi2a3+E3rJWVnVOZAHfy0sdEipZEUWBP3yc65CM7FLjyv+MkIDl6ksQDgsH0fE
BU3CUzDfmTQIWK3m+xB8wP8DP4x92cVySHFBuPYt1nPIC/JrX2EkvfISnKsqWY6tDp2d60R3vaWR
8AhPsh/WGN5TzTuh7Ii5hFijivZupuo0E+DPILbvHRMgSyAT0RyzdzdxdDtfnM+Ew6E0oPkhuOsk
LRWd//JIrN/azuAAg8AFJ8e8wOdNXT/YMnHeGcd1qfAlePoXSLLuMh2UDJi5CMPWpSx+vZ3FAKGd
afpv3BLkatcfb3ZP3jKLbRJcDWXSBkhUKfaHNlAzGlUDK1T9yXpTjMoRUSAacnqaWU7n4rJI6aCz
wv8d1ZII6NZaElq6ojrevXpOZYJH9yF23cxVdQnpC9wI8CQRhyDJiv6g08AmipDAG/N4ygBLGNXn
o6s9GtTjUcsXc4FNKq6ASLFtFGRgPUs3zbPe8srAxIpvolA44rhGob36YgPXOkFWq7DvzCM5owTN
ltQyINdA4k+/RxXAr8xM4SH6D5qFMcjRP9Qp/yi38xRQPCUCa07aXdsJsyWDQ863nsCx3ml6pzn7
wHdqTlDT2XTA3XPHwLL5OwVPctcD48J5Oen3dL/zUkifT8wpkIJihUAwdy4vef/EFQmlIvfDMMgG
sOpCZs+FaMz17p9fctxv7Bby/KwDqRgkJAWHyktVdcd7PB5XTO9V7n0dP6crd8va8BswAo8WeRLz
xWyxXWahGhcBVTmx6fIVQGUF+VNae0U0KEqn3jKuu3yZeyP0fhC+be3rSuDOe/HOuY7ra2G4mU8k
xbVptXoIc7p67vErvPOBsAOVEu2SPgnk6hPx8Uq/ekBk7vpl8v02QfWHO0Sy2d8Ren9IILyQJAV2
w3j2fx5bAGtREtbgDls61xp8w0nrU3MsFMJRrU2uK7pVda6k1VJ88O02utOKF8SAgB3XKAFUZvcF
xf5Txt8uXowabtnmjql6U14dEXOKZe3lQzjPdNclynQJhJ+/1nE7FcDvNC8B+XqbdbKrS+XeARrF
CimmcG51ravtok7vLtNNdXnVH3uFvRYTiomFI+OmhCM8D8e5bTC9Na6RmpWWTLQk91jUS6XkhbbZ
GS837CUs54DZ/8/e7cxDnoMFfFp2JadxcDbvwM7qx79yVdJDyCOJQCM0ZnKOMmgG0x+Q10n3lrty
yjLnV1X7E9H6vzQw0PnjSk7cfDaUYobPu5h7C1TTGlr9LSQlpyKeoq31DCvcNSHI686yKotegeFH
EXGNendKGDfyqPGJjSfmiScqiG3NWLBK+e9n/247sHkcKqDvd3Ia+B7bYfCmUhWCp4BQ8a1GonQs
uAQZ0KqBkwkAXqbXjInu2SgvvfZW4eMolxGDUOrH8KzHQSb0JcaUGCo3t7kyT6yal72b3UzAJH9f
1YXz5dZZYNWNdLVRYm+IJ7iUZiL8aBx/1uUDGwHjAIeQ+r/6X1qm1UsRP8gRbzhHomMH49fb431G
tvE05CneHning7Lk1w1fLIfvTKBpH7SuwNTCnwCs192WQi/r48HIV4YPYu2hji9zffuZUg8pQ5Lk
dppMX5cVm75CXeA4YoLuGDAKmjGizwRZ6awUBJL+HiB26Vt/WUh+JyGwOVTJrJ1lVPXLKib1vV2V
tP0G91lIjpIc6O8WwvMeuNjiCrLBz8CATazuw8TDFZ+XVNPvlA5fXE3jFb15XYrUApl0rjJFbCLk
NTdEbdsZqicRhpIsAjmyDvwK0ewh6IDl4caylBHNNLwmiZ2WXqvpNVds9DEhjrsOTDvWVuT69pPo
k55k1MzwcjKP+hjEuj9ygEo5fXlrN4lUj7m/bE86fpMO9+5FcNwuqS/MELfXhq/Z3plBhPE2nGJ7
fu6hwYVf4q9888NCyhsPPNk2/jZFoLMdlnDI6xBOmswVry8kwP3LkUZNMr3hMGqdiH1TVxl/d2S1
XgW1p98vp4St6qSYx6ZY5ECIpkPhZsfYYkIsMChvmHbGfJXw+rwCOiGV5xIYNsDyYdHxi6h6OaQj
LNpojJd/XSCISX9ffappUcUydO3IVg08s3SpD3pY3aC7OW5+hyZ7l1wu4U+xZ6Ih+1JI3Kl6yxaj
sa7ruRSEyb5ddNaKuwNnZgZ67jS5EhAZ459mt2fZl+woZ48eIAr6spyQGPqBmEg8uCA/WG+lpA0q
w3/NTer2lr40Ebs2Cv7aijFwJIWhHEQfc2Ou3Nsd2NJLMF8/xUL9OObOtAAGl26blSrGSvqq6mSB
o4VWwmPuG9JxsBWxf9LQ9WL2lrbxweb/pKsXoP65YRZwrrWGz7Bje1zKWFQUYEnV4e4QWxD6kr2M
+Tfz3Dq5YJIQT8hArSgnjSXm0ZVOVMgh4FBvLuFZd8r1puOtrotrSoSjZrxYnMlaPM2pT9nDQxWn
su3ybvpPMEklZ/195g/xlELSkzOopnKqCi7GjbsOFh0ZZa9TCq4FXBgUrCKpZqm6xUsIVLKujzj1
7BpoHlc+jCrYYNMMaeYjMxiaFik4033D8K/agdvtrs6wWf82tb2SULn0ejMQD/uZhPdJG/c8Ierv
L9yIaP8RrqIJgTEQfZc43SryGVCSMN3oj4fRzFXqVmxWQ2BLds4Of7qtbmyyBHnPFVRwdn+ezy78
mRwbXCbaGoVFGcELB7ZTG+ssLzersZAEeILDulVG1f61O6kjAsrDYPnVUYg/X6dTMWXzugytnGj/
b7Qkm/RUD8DOxSe1lNT2f9Mq1Hjnwbmxr2VxIcRTVUmNQCuU+kvxq6cq33o2YlYRr9YFTjXUFsr+
GoCdg+V6SDKEcQAOYeQmN/CurTD8qJ1uEesHQ1LjrvYMvGHgna0tgJsuclA35KP1Z52IJ77zoskM
mhAEBTOVLPk5UF9n4FStZDiXl9zNm717QH+NiWL/WBjWlekE8phgZUu37TbxhaS30U/WjaTl58Pq
/iwPQX3P6A0J37qF7T1UnvtwHRo1XXBkrXaeQ+Amtzy8QuNJC8C+RlH72OJcmmKxk/LNqSUEFZK1
zl+mJ8WOTgdLsex6NM6X9TNYenrAiTIuwk1aY9+/b7c8+cFrBFozIPQcREv1CL9afsfm2lnwtBWR
FAX4Imr4xFB8SjGY0WdpUfCUXEEl9jiKit/QmAX0bgMIfQfMo93WCLPtLxcVvntLW5gSg4MwW5Rf
nbcCDrTHWqG91gQbm2HXaR14cP4UWakGYvJEs37pYaimDMvbVXkrXfslDa3TXGgDRS2OYcwsXq94
Ld/rCc2fccu2CM8RWnkF5mPVHLjFOUc1PswqCO5cVFLsYgt1O1WMj1kbh01qTmPt1uIM9HOOHDTx
2dUJv/9Pg7GjLFR7O9sO1tfkYbY1xQs0Q0KpwfLNn3NIzsS7ckJ03fMUn6FtThMzmd9KstJRRTIN
utWIkp+oy4Pxywf2AaMsRk9cuYS13b2LSrZ4F9DDPL2KcnvvKPm45jSjqkAOPr59JnEuODW9PW33
VNb3SemDoS1AsKpvIQ1rVc+1IgR01q0DR9qhuDh7PpKyjDTx+86fcABO3WP3xEoDMaiGDfxH4mad
MMZ5M76Dyn63RCFXRi+OnMlWyGyIfwr9c8R9mwi/wlZ/HLj/KGXXDXjTO0/Bq2bgUEtbntvZQjeT
v/2hRzR3CtR8c24E39dCHWEkvkp/il0WslorUX3qn6u6JLqGH83kSc8MlEtSqpTPW2rVOE5vSfne
1k8iuP9+TC07oL9VFrF0I4K74OLmBr0yi0/mTS1vlJK3Om+u3/iPY3eWdOS4DFxlWS1jeTGlo72c
zkqZ+xI7qwse/yjmQiBVdYwhTdcqyltgUvfO7N3f1HiHX+QelRtx0CuBIwTlnOmCPaxD5p0bfUVx
08YuHHXBYzNSdB+oqzUWEaRJcSvEoIikl92nNWtv07JEzKvRDbNBYK1QzBVhbcxjw+14ttv6K06E
aWSd6FkLXYBad433eSuDG0A583Fct+i53+Y5uaXecmr0fFb1uQNs8H1KS9g9dp2lEZDBzXw42359
57anlHbBvfzK00mbtAPwcrle9nJzW8lbrENYeWqvAHwOdWVCcICcG0xGTay3GuQPsjJ8UFkUUMhd
R0XE/yWA+KL81gLxT9Mdg7ltx1lgY27BR8F5jidALcg3CUHgOCWC8O3dPzqsyUkgxobudOjBe/qq
VUue9CaUKoGYu3R84cG7gRo8OpuhympWY/YRkMmn6fekGQgj4eMoJ2UT8vFWUZsSlQtmYORse8vs
oYJigrBNe3t1nsmh1V2l1UN73Wh89LnwA4/sh1UPRVWxzQxzG9241/gvhgk6joB4OMKcuI9JtRpF
1xpheAVAA8hlMMRZLskD5+K7XNy2GsdDZGOBNmEdnvqhyCHdbFAzuWXnVET/54yrr4NGFWko3I75
JekF1eze7fW3PMd4ZAn5QWPP3rKyECFG+MliQMSUhzoyCJkFw/offC181/OGO8+9R4XIjJtE2DfZ
Xdcpz6aXvx9PCDAKAViFoxby2dqvMdYOuFCajbiPjRvcRqszC+mnRbdutqNCcYFwnSRotHDFX7uA
PN3c6HCprAnH3tSlQBQeegRA1jcTBTyf0IAtdZLFIKPsh3wmCsSCxJsK0tqrx2xWzv2/8Ob7pulF
OOZGRLOhYwPJaZud6nIwXAGLt1ErXaCje0TEr0ZLxGCXupDUogjaTc1f+jHIy3m7vYAtRb3jXi/s
tRklaDFt78unvBVKTj0KLBVsy+dtGnvx+hMG/rJhDTmn8d4pQle7U2DGzw9Kxym9EtZWpzDLCKaC
Yau1KpRmmGMLfP0ndcVMEMuCy21GY5pHbxxRRJBV5nULa8NdTkGjLYwVj5bHNFN4EXM5FJUPlbLX
fnxA0dEn9VMVaAvO1iqYOCmbt0+JvMPB6+0psYNaK6lzVtFy6VGOcasqtOFDDBznvqGKHs7LAogw
V+ZerLB/DNueqOMJzOYciatGxWlZ8MVW3SMeZG3XkrkK8dzESqYa7WWhnLMzhw4wKvpKiy8ok3a7
PhQqZTgMBkCKNOGb8VJyjy23oIdECnIT/gElh/3JVm7exWaPEId4hg1cL477kymH+KwdaDO95yOk
9EVbE7XdgE45f5VBYYSE+ETEhcBEiLzItyJu2VoFleDskwLnZ0N+8TBM+0fMcAoU6ZVlZ3f/wL+s
cPDgXMYQnz1SwlnMs+EwmXvv2SHvwjxbokKM0lt3jNn7Rk3i0IWO7rq7p9EAdGsRBZnmTdO8vAiK
nWcwW9DpQT0iwpWiA/M5fefQ0pyB0mEM05u7y8KzsbOjIQ7Q7w5NFWYxP5rJF9y9AHQQulitlqVI
5lN85Y/NkobHCcH/npDPoL+Fr4mXUHdSZmC3rTNBsJlwO7nBZPgP1fBuBsRUQntSk8EUU/clsBui
9NLXKE7JnLeGYHPyKmJ+ZZFwPBE6heh11gopQsyCwxmA4J0Jk0xeZ3xGtBnv6om7uwk80NB/R4bo
m8cpbcKZjR6eLwVbizMNaZVk+400Einnm79xZ+U2p+Lj2D3vJgkseJzIqWrBGJsNf/gbtSrJtQxt
7XVcRPjY67nl1+gTHRWwzi5ghuh6p1S3jrsReQ1GPwCQAs+xdvciytAoX5zQQhgDJQ4ZuUq8Za9K
jHgsANNDvxTzVPCRWhK7D4L9kFl8OPa1IrDO9RjPJN/AEnGWLrpwEy2vtMzz+JwepoFPe+FhfZLb
29/4mrxr6z+9ah/XWsyfZBXLFhVCYRXm9PSDv5Z+zbj7HuohdadVr5vtjL0CUhiPuSrs8og430r9
FR0sVWuqHd8imDdF9gZ7OzzwSOdlVJzNU2T07dbuMGUHT2DA9ZmPR92SsgNH+LsMckxjDNba9mLl
ygsx/ExQjQlUb3gyM2rrCTnN7LpiljMxdaNcIu57kCihR1chBX0B2xPPNeLn8XFkexHlzTDkuxq1
EQDBoZTyJebSDvP+TAyd2YvXtmdzSxvZV/rKMbXtxmH6UJynPSZXleyRbxHyUDjUIZAnlf0ModX/
okFz95hNzMiK4LmM697NHP43PjpcrbMaJukplkM3TnKxlbaihOziCymuq8AGR03lUnkAUBguc0IX
GyXDZ4KXkBWw13QiPHbhqISJu2jtQw8TKfEocqWpomsFOyY34AlpdiLOsSiVhMar6x6KAcbsN7W6
HhDnsbjNEdEImRacm9Ah/gjGrFr3Gp7Km4cVdYij0prMybHFUOF1Mgp0nNG9nvaexaSGibo5SVPM
Onwr6CWKBx/zF+3sFqNph8X0HNErIPSS3N0KWKCZHuWpgb1XTo8F89BrToA4xYNY49SLXPnEE+EP
4gZZB/C3AoOWirPD14jDgLs+UheDyFQZaUR32PhM3yDGNo2K9pkVp0GSQ4+wzBG7cWmti5NQuh5V
2e5Zn0AUY6QB13BEHa4RyUNfksNr20bbhcbazK4fCb4cVVM7BhBnyC63AKNosQSTsnuyGwmtMvWI
iG8ijj+/d74KXEA6SLzSKiVfi/T0+s5ObpYTMpuwoc44iRC4MNQrtWq4+31zDSXPnsrp1yJdUnOQ
ex6ZkZYvjt/UorjoHgKxxM8asdTw7uuALe10YrT7tBg3u2IZPLVPhlHUQOugYOk8gZ8BWM8ZEpjd
zPxOBi87iPC6poD5L6+H/O2Qf829XceRxk/JTenQ4PQdFTSC6Ic/J5q0/pjrrFsiK31YaYejCyZe
xDS3XOoQpITJqxPnBIz3Fcz3pFKlrk+4KcSNvc9lFMgB6bnLGOWbyR4wmWIA62nSnbHfQIwPIh26
AL578+CBDoIUC37iStxigdGuRPyL/Mm2ZpuFjhTwi37bT8Hn5yz/RCcRbXcZbiH4hrybZdSXa4y7
LP56KVd4gkykKBEE7l1b280ZKG9TnUBJUqQ3Y1CtchJu8+IQsejTTBQaEYo7jo37KCg53Wkzd0Qo
2MR2yuKiE1ERp/CTKgVQuiA/eVmHpWq5WEw2aoiFDS3nVnD8e2tVM0gVi3lYDbUiTgUA00LERTzR
ahbu+H1TUpnOBnAbeHrjPTCf1ym75nRyDPiAUWkKQxwJrIFxVKd+ejI3HiPiRdGqlg7d7hWzTB4s
GL5xHagSCzSd1HD/Tnz98yk+FzLkSPJ+W3fkjhvjz+yJkeAkdO/2Cps40iyWgiku1yNROxOJVCpS
TOzEf/zbY1Qa+5VO9EIzTagGmaTj/4UT7bvUYe2NJ0ljDWJoTqf4+xF3DSNSxyMXXULoByxHFJ8r
uElT7vmkXL/Jgsbg9dEFt9BWvP/75n/2PQGCfMFJ1TsBEjwcMNRfbn6Xpvzkyu3pLsAHBOALz0uM
X2TD6Vp1BEtufMVjr9O09dpkg4HY1QSSVyIVZEryBD0H5tz/DVbrcXcTMwle5cuULaWtRaisGpzU
kV+ZqPgfB+4/2I0yzxN78BXoIFCfKj3FIMvj6/+Mr/cPZE9ufubEt/cl70sUSQF9krg60dS76OMD
iOepv1cFWku+buNaJFav/tZo/H9FJz/FjFDPEzXqameGWw7IED0zsqRp9vVEPs+30ZEHQ8iltTac
3RYps0hyMyYyqV2z8U7PZlmwoyCoZHq0voQPYryEYPUHUsLsm/1CjbtXyCEmcsnhjYNHONJVADkX
acfrii/T4iFeNhMBvq8vxh3OYujHPjxnwpsuUnx9NTmjkLrT0aFsGzQiLH7lwUsYrzKg339hJiP/
n46eCUSDwK4MjQEOJU1wZgdsg4mukfbXF3yrSx9yIPEgrMPI9kH7qXfQoF/5DyJrRqtA/nurAAPN
P8PyaDcNh1JV4zjT1EzLBBz8yN03njRL7EeNxpdHw+IpE+Rxx3zeRTUTAF+gjgaf2NU8GorhslbI
I8AiaIkOjwKVL1P8UcV7JD05Q2pLQRa9tiQgDmzGyIbkO/dAqReZ1DMIZu7nctWmiCsrcOEhLsPE
IVAR+EZMuXYIcrireMx9UodnCTbu38sqOqyD3RytZ1gSfOGsBrMhuE0lqRXmdMSz6DT95CRTjPuK
A4lP0EhntiDuskraLYZcvPa8UCwKSrJNS45MdI+Te3ChQgZLBf17ZiwtMq+RfvvO2gqsBbD2OkK3
PJCFXFy/LZO8r6DJk2Ki8TzOu4UkL3wvmwCKf3mFxcCVhzFGDK9C4ZJg0rPIleT2IFaQtleG4boo
6K2Wu4WQ4kzSNyGqH1rFIbiQU/7TYJhlhUAKZUdQtL6MeTVPB1HSvPMtjVsHi8vTyHvCXSOofr0h
Kn8tU9t4+mdVgHtpWmbr8DE0BEFNmAMKhai2NSoRRZuKNCqpPxMAUL6ssPODtttY+0WTFXztPQs7
Ewtuv5aduEPwGuV/8UheRT2OrGWzgfmNxLBSM1uNbX75obia2KeYpifVVJrkKMVaPuROY7rVTtod
ewKUuGOqgYCjrSHnr7Gf0+/SOp7KU3r7YTwaCzqz1O5Q9nTcVssxtdrzEjxvvpuaEp6NeJXHhwyv
5m1+o/iyZ/Qdm0j06ez0XxbbiRIs1gC7HMOzbAKrm4s3NFb0wTgobEBHDt2bCDieqOoht05sGONC
UlDArWJMSg5lB5Yg//WEwIDCN2c7qRn5cLfgU0NfINERj9xKytT2UHsTHbHx2fuhA9Bw4BD2Jz3W
PYWPxP9q+CrDF1A/QYkUjVt+gtTocstzihuK9knxiPPe7H6qrvbaUOTSccgzTvt2n1rxEmKXZLsl
aKPdeT4mqUdezbkHcq2bTvK6P+qraUXJF5buEuZRLNVZJdvGGu0Vhrw9+gk8g7Fpx8y53BYAq+c0
n9rZFyB+l0o06bVFdphcYMpiCtDpZb0yUabWfGhO32qoqBJx3kidFrpOFI4MEO/lvg+f9JQABtZr
///n+Km6nKMd9ChfVx7bLz4QzBerp/jhVewNMUxj3fhDSaou5CcR7+ulldakYYkLbZ+wXpKf0KCK
qCDk4ln/pocEAgKiUNX9BpRyVyv50U5hNVDcZOHhjtQOuQblmfiAXZNmT9BRZCGEtQcy+HwpsKYn
BFCFXdataTKFQGaxP0bhZSvDM3yo9Gy6LHhC09Bw9dugUvRGxTwlK/yPdXInwuoQjwZpZEHgICQf
t+KyeVDIQVKc5yW8mbXjUzliPa8XXl9jw3iHMWpuSSRhI8GUvplygwfbbcsz4F2q2Yft0huC2C6H
pItqkIx45zfhRJpQ3Ziq4jXxED85z7kvG8h+kLo1EaiUa3DBtHf0ropOqCw7itiX7HIHc2lRCv7l
sA4jOirsG4d5dh44t8zWEfzLG+D/lP48z68ogIiutbID2CldH8amexf2bp31jowNr/R7htS4a88Q
IjTi1QUYVGhk+4ACPeBwEltjxYhQOKfYUESqFzI9LsalxZ6jwKlR0eqk4yeIobevBdL731fA0qeW
nzQ/jKgLKO2aktFHLnH4437itFcQVfpc/gLDQ0PchyAAkCNtE61KDXaxFarHzzI9A82EaGJeoN85
z8oL21ldivmX1DjEVZ8ctWN2zoZ4vr5+zcq5LMMnf/wOTTdw84asP3CoqOht0tT2OGRI2C2sJw2V
dqFMjNBz2XdUz1x8TzJRPyLV+ENApQh0WonC5+6iJ8Aa3o/YiOGwTh4GmSZgyAx7+S+z5FfN/wmN
uxOJd5QnIsYvs40HzShe8cZpMioglvnrkQpMVLgZZRa9QwgM3VnIZM0jUiU6LhLR99KqK5hyUj1b
KKC0oX4zfttXvQ6fFibSwK+141MZIeXF9YpFsq8qoE08nUY/BfYd3jfHyDQyjgoO+lQXTYoGDsiu
yqNILlXBUbcmToNIxIU8yGnAXg/u/J0ky6BJk9LdiawA1BTEvwrc6q6VWIRUz2sBFB/H4yYxlZLM
FJW4+AeRvMwsgHDUWGleqd/3zESJfvQ6pRTkmoIJpn8wDTwVYzSQblebAJ6xFNUxFk0UF0tuM+/y
8QBtpiWbAgKVGBcRINhom+S+mJGXW7Cffg9CP5BkgYbHnHAgvN0ncjCwFByRPdg1uvQisKgdW8YC
O1gJyJvlWUA9vJOOoELBg9xIlPFY2TR2aKFMJxhf/q+pP05xZ2meFtKWt1IJeW/toAq5BZQQc4Rf
+RDeqc1SvvIu42vegmkGifFAbxzE85CEsDCtiCi+8wfHY0fpgIKLU7zgiMMRbgNIu9rUDINgR/d5
+80ZM6gUvYXBN3Syn1SivSxBUPdatU/FevZ8jI+BCBH1S400sOYb1DFrmi4RZfT4tNIE3Gzrw/fi
0vWcYcptv22nnLvkN5kMAPuDbywkmGc507TBG9/SnZBFfSoIaZxFpp/MrmJaUHiDWjtIresRUxcI
1VvjMsYryIOYajJ0/7K3hd4f/svBD+6P/nm6Ggbo9fE5YRclB1swPlIl+zF6sdIGUxveqzon5Ive
rqIdPPcCzTkTgoHe+fUNJNVzlwB+H65PnEiPICxq/sInWXVrOBZGzexTGnhVqDJr20YhII/c68rF
gJvRvDtYgVFdbl8nFhfyKvUpLC1Hv/DgHLVpXGP+fiZeTDKOpnfK39maUvlrq08fB0bV+IS/9ebb
GLO0Tpi0JEGFhKe1FXjgTgllbABwh7gyXTFT8fbewQf9CB6Lrl6gPCzeWAHLz+lG+VLzAlcPrE+A
WwnIjpS8w3CFsC0x32NyL8errK9m7J1LLML5WEVGqFtjCfR5TJz/y4kMTTT1pAKc55QvCkmnax6X
1ZM71CpQB1LLUoFi4uZIWBVBiUgsICv7Li/OsNtupRQoEeUgX872l/dCZRsm6/qzd9YDbP8xgaQq
YoomqNo9omRqihKKQ2KYR1F8OgOaSxZPMzla6et97jthQJ02xTvvoG3qsp3KSxIs61QEejzX+zU+
B/BOacGI/xULDQqUIcXUFXjHFcCt+Wd4rwvJu65b98PUjbZN7MQVjAKkTw9PqCmku8DzBonNA4PN
b2k4z6FqShZo6At4soWuGkZRh76cuMcmjpq0P4U9CzgaUaoo8miOyH0BM9zQLmLZWT+zd23rd4vK
crOhe+hEByajsDWXBgUm76AiUTURoKcbRImdulQK9Lx1fA3veXa7KZUH++CxcuF/7wZxCCq+ivgJ
yDCCQog8G3E74HbbOQzGbUXtYGZNl65qlv9TEruG14XMm9InfDYz5owp4vayOxHZc1j0kLv4QDTa
IUEainRnCQn1E8pzGAoGcP2s8/0H6zBoUGjucttodDXZUn0jnLv3jD/oSCNYuFB83kQo3vy67lq9
XcWPi66WrfBXK/X7nyX3SavQCAo6ip7LYVMNcILkhNnSkzvzbiBx1K0/hlilMzSZzc06si1Iv+JB
a9GEs41bPIGu8/L/mRxao0TK62w0l8f4SuEVEm1ggcdkRuHpmGhuJ6U9J9GLfk5Jnljw/0jE1AQV
epDqiJka6hVTX6U0OjqfocMHAjMu2/ZMtOaFTQs2uspoGqaCRw9XykokcFWSXEbAztEdI63EKq8B
LcLJrvtCdq0PbucfQHV2X26hzlID2MyYDm7KeI7VJzGv5wWfP/Di2UmXYPT4HmhaVoVJztEadkm9
8DnK46i0DMpNS30fQvaRfBBZst2hKPqrodToZKXIFieEzE0WA9T0GdrTKhv7VxpH33f8JxVncBl4
8mDwD4knHM5/1ablI2ZMxFcAhfD1l2ZA91y0qhS9GeyYa90cteG46zkt0GkgFwoMuWrbsDty3Ssl
CGFgVFaUQlC262vkA2vTyZek559/axCM6veNOcJLWXsmaQx0nF5KuXmwmhzxz/tQAOlyn7tE+l9k
/40Kpl+BJHHjet3TmZWUdVOBgzI1mymO7nhCexMX3mBTjNI2VYgBx+nbpX+IOgUr1RIKshg+RPWt
hb+tVuhg5GxC9qm8s/+4qVrYZ4p4798T479GjcljyfdHRxwnCGePyjoPVYLGMV3L1LI5brYIz0xh
zvoSk2l6DhJoMEndgsHsnrGjXVZvAriMX7laINQOGFLfSeWW0RlHMT0FSWyr1kJViqdbnoLeMYFa
qeCfIVgQerNsH21c3V+ipXaPADOGxypOiK9jD/xbcIkoalLWCZSfMM0y0ub7AQJIDdSbGRLr6i0y
NLNbT1SvsqcpW7Y24XI3kCjUGUk5q8eBwj4NnUUCvXOhuVs8b05T5ErmE5JpIxcxmrxFZas7X0yH
T2HfyLRJ+Lmq5+/mYEf+FlQLRgm0hWSTZjqKtpfSrZMUP57rCEwLFFdb+90SgTvfA6WaBRsfCR7F
ETg5HW/XMyZBVYozDWW6caK7u4grVABM0EuFSVz/rvtX5qyGUJx5s3inCEmsVzJu1jLMyjo2XeYc
ko957mwgvM8FVPeP1vlDEHUmI5w7kR39cFJew3EW+tRTPA/lkLHjlHiqmJ6VE1hoJRdp2yrpXlgs
PhLiZDvPd/z8gWFLeeJ3o63sXclsBAGDxHPbYrvDt5hBhDkXZnUcrK2k2UEWT8ctRShBzsUaJMMw
iILDRMHpltg3StQXTP7HLYG0qdZ74izCKiXBhvGBLNzcuVMykf2M71Uldqe31DMOvWXQuK5hsIqK
ponb3oscdU1pjjd3W9TtF27LHDxISrLmepcJHuQDLo08UJvG1MWqKTn0hd64SuI5UTfaIkQLLKm/
3MMVf/o5rlmpKc+zQll2j3F5OQ9mazAQbbHtdD2sBNsZDUzige6uVesFPL9DpYwa2eForryoq0fV
W3+BEMstSye3FD/qe8gLCimLC57ExLgz50NpAwF7INvum4pzy3uMgQziZjpvbp/YTlEFHnAokkmk
l4jaMCCdcUC9ke431nw+tz2gY2AEBxuUWvFcyZ9N8lxiHB4zykSA5913UGMziV9o2uxI7S3soCdz
yuuP+DzYdTFoGTrlYBcIIPz34GK0vBpbPl5snu0qDy67gF9OIYYwXiz3MKQ8fBO5xsvLq2tCtIsT
EWOhIGMmhTOev/NGGgyjxYKD2+ZZNjbv8XdRhbdrWRWegnydiV0tAh5MDAefgQIsX9n1j39/VNVc
R5KFGJ2MjirdW02xHVfqAMWsluGyYx2FiYw2rE2aQca18bFFntNO084mZdQQs6HOt6wwkMZ9JEow
BxreVFEsElD1x2cQf6mOlkq4zPkb+ItosVG94tllJFcHxjcmt7gSn6VjM4X+FOx4YwP/tys7pmwV
Y6sgU2ADogWwOTo5zN+cqqemZknUtCh7rx9jF61Q9YyL9MO+53bKKq7KufVf/mFGMToEgueynYTc
ejxkyp7pjMCNSsDaleWLwO+RYfTVQWfOVZ1io1GetIEEWr6ARRLV7KCNyrhXdw4xLaoKeKNzZzdj
kIYm0FCOlTEMcULry5O+744tDdMQ5KYOLQDpNLpTgcQ3GvUwmR3clOBpwAOsPz/LWO9Tu8UP0SGR
3wKl05z6NwX7ZvcgeogUJb/9Rpro2A8sHGOSwZD97Fu29/+g9QEBDmdD3GjpmZUGi8TPSFUs71JW
rDyvT/s3rRYDhPc5JFmOTVGnC8LBTljORPB9cWgiwSLOVUFnFkwl/0RQp9+OKcKGzzJ9rasgs0Ox
OVCqry//0WXS6anIK4nrT5wPMPB5ZTah6Cd+kGXoN3XFy8s/HT3HjIUgRcbJSlktVRIJF4ik1w8k
9qjrh8Fbd2lp2/GtLLGmDc/+9lOFtU4sSuo+XgnmgB4XPI7BnAutGI0w9g0H2TLu1kd5RKPWxgVM
8N8t/AEzYT9bsiHx2fvHo9KoVWKq7wa7eevuSLqOVClyazWyaScHnQWPmHSnp7pbq4sGCG4Pedvk
zFg8utq2Ra+yZ6Ea1eENbrXQkXzcwdQsZ0mAOfENAikY3uSAPSP8WowNJaoca7lRmZ7eRPbP2mwC
jCixqOrGTyOajf4/PQr9miPAMLCZNA+/YzRK7zOaT1iadoCb/Uolto5BbuM0NKdizFHrgkBjnztO
fsBZPbRdLs6rVvmsfVclx2+HGVYohViyPsY3DK5Gb7LZsfjDVMd/HV/Pd0p00voh0hzCzI1t8T+j
43MB8hqyJQT0NunO53XWVmfhTf4k7Lyq+PW539ppQf2TOJoO7Vfhdlgzzc89dwmIoVM9iMm3PBP0
JGQ3QSExCGNsSUP74oBl2+L13QSMDeojrZdb9dqBklOtfkxnR7haWwjs7XyiW1AJjrrVswZzJchm
bkNT7mA/Dp1MvJ42DveMoBc4E6oW3AVo7CcY/gIlBZ4vxJ/A9UW6xYKtyhfbqOv0HJKkNpz4p8AA
/b0rt/HZD12osRovLIUooQUtmF0tu3lwVTxikcgKdxCP/y5wLFshk1kgRoaUpuBwgDF/JMRYwlAC
RjjDVfksoxsj/9pHL+o6ZHa1ybxEBgHlpK5tEz5A/n+rSLnxbpxsIsGDZ0G2bgx3+OSJzyOtYSjT
Do2GBEjOncjUJxSXywalbt9MgW9PAX9SkHqB5s3eXkFSZMFMdGBrBGgXb0pJKHcqE+XIGzcZ81l6
Zs6qMrW8gcKtGTIqZFlpyhpjHkQ6npaIIybX+dKPFK7wdNge9i50sIRZZawIiZQjNULdQ4PcTO1s
q5nQavPt+oLD41XeSxJng84KzXHzF1mFe4mlpxkuQjU/KpZhjCffz7tgKs82leF4wrP5h/NR+Fxo
V7NjZ3w0vDcYymZ5UgeCNGxrW7EA4YGrnM7XAaIDspnR1htcXGuJ5/r7ZBntKwJv579VJ9WUkXfu
+kK0qpnUqIoG6Xrzu/Cfg5u85VwxeyOnzODUCzIBsQHSUl6U55iMIRlC/dyP5pq+D0vjXhKNAjTH
ojpAWoz5Ni2woXZNKpHRns47LL9fbbiDM0dC9I496JJ732c8lbHooyytSIyRlH+t9JWokpNA4pIr
VvKmkXb/Y5AiviKOrD7s0HH+iRmqltf5hHGPC8kiup6Ys6a8PXdaYiOcrKC/3h52ihweEUTVE1V0
Xew2ZefFgDxkvqAJizjIde12+YKsQljlsPm93KBxUv4U2QNbQse/NtBdvqX54R+wIP/elbu8zWZp
haXlWLWxITZ8tNlwq1fctQAp89d8/V2uumEFeU5q7h9XrQdDCTMQ7Scnqz9nBBITCc/JpwsnrAm5
Bw5/oQYneLBV6mZ8t59ouNvnBwYTgyItXD7zRIwGfcRUI/G8v07r80YCqQmKeRUciRXxCtxPJZca
4hUmfTL8Vg6JEO5smr/s1Cdi/hPQtKNh0eTY6Gr7KWythRmoFbdQjfosgUiZ8OnHdm+H8Z+Ky+EN
IAVeZTz+Mu5D4qrFohr6cL7Svi/6qdQxqOqiYZWqeYBv4nV8I+ULUcRUkkTJmBstH9tmwZbTh2IU
ZObenhT6KbcvbZNSWARH4LabACwtUvE2a4LPthraLeBwne7dMYy3NPX3EVI/m85PROBHMGgmJ1jf
ItfNcf6iemlc+cIml0q+Blw0TZ/kXUTyJvnyJtZzMkxZ21U3yeyUjT74yjqYMgVkwtzjUskNGZcf
ZIPQWrJfbkk2FhiYuz3a8AYKH6hZFrmHfHizGs4dnmFe7BFT3AapxoPjdL7/G+Akuj3ouNDHZR3d
AWAH8nlPL5RO1fXhfGAzZWwnlRH3LriyDNvevEBtTU2oFnV/kyM7N4eDZC4KzJhumw5zY/1lVxx3
CK6YxmBxGWWSLp/p4xzZdoG7bdO3DJSy1xEOKj4z6Dhm2lLBddw9yze5SNkiF6RDKVf3/M0dKFf9
+yibXAjncgd60O3J4QN6Wjc7hZLS6vO8Z/tLQmCb3kOPzAMj2VpM4KfA06bkHT56GmfPSTpzbX57
+Bpzpi1ya/yLDU94QdlNB4tl1+MrRixKMjW1X8VFESx3LAbfngn0It3o2a1UiBbmPDGrM5kmsfDu
33VeQd1GPmrqZmL+b/HcnNSfgAVGHe4b3mw5nxULXfHbnWBrKYSUU3FGIaNd7m3yjfps47mkOn6d
312GAfyvyUzbg1nBCJc83ycXFqo4/tSzZP6s9ippm/VSIhZPRDsWc4oIyMSk8BCqcrBIJP63cSZ5
1/spifWoTUMRd9gB1AylnRmxRgGdePgFLXd6QoBX+Rkp+kFEwxod/jEKBuWhS6houvCBnkz6Po8z
NrlFNaSG2Im0SR8zl/wXFPSnqSaBU2PbgoeTPWo0UTmhfFR/wslKSdbefKAwdSjXO3sw+KW3DbYU
gXRN0XvKyzUp7CBnDmTdRaAWZxEEplNx+/ykdWFQQys6p4zw0ZPEXuWMzyw/eNWvHJWhn8RJBoUR
iGEz4iDwf1zjxR0SLV7pjdcJm05GB3gYGxCu26nZWeMNuRTfiWcrs9IIxwZ/Kw2jt+Yylzee14pF
JfGk+lpMqZ7ddAZB1M7oUo2hxx+MDsYiPsQiOwxZCReEM4Q5Ts0SXxnSKdJev2ejnuHYRMVuP42s
UCktVx4JrOUAaxxcuBCnDN8x60nmfp174VnxmJM+FyfgFQExN+mLUpPEQ1Flt/D96/sSom4gvJrt
5J07xGb++Xnye8h6NYdScOkLnNjvVJRq1YZ/d+vlLLHdFexKCCJ2dmlmIhffoQGseF/gYB2Gm1YU
/RzPzYnyreeBOknB74HWE00y0vW34hTaPgbJ/Ao6AjbqwDNSlUmqsbRD41qcDYTXe5CoJYUNDaaw
/EeoO+JCwJDmDGnfRfi7Y9qqF1JE3RiIUT5jNxzV5K2dfoanSauUDzwA3WnpA/BTXKqGgZTxE1At
y/69bmBafaCxNV7UJ8fOWQwBJiU3SdolUmMT9sJCATwU1RaC5ylxAz5Era9uNVfhk7xJvxiKzRhA
jKos6qh8mLsgBjw2kfc3jCRkpRjCnLANY626dNH+Rw1jSxGJWEad/w8FNg05F+edHwJC4NyAcuso
UkNvjhQGWnGpWXR6+wldikaBBgBP1UB7Ov9TvnP4T633xtuBiOPCzTUkwpwz6L8Cf3/Q1UOq4q6t
BcVU9xS3+ojt2GwWGZ7VWFJDxb9hGIz23lmiAs6HVsC0/nqgf/VDwtcaAHk8JWFR6hGAdz1UpqxV
qBLmrnfwlfpmquFjThrnJMABca/oTgAFOvAhRi4zmplh2jb6xjoM+/a+pD++Q9OCYorH6/jr+o0Q
bVASgtZd/jWw1t7yPbsmtG+SDWWqQOpuuzvkvGhwh9gLpvNevODTBoHwhDwSBmUsddqrY7fTWmdj
rGxctuq7L99fhFl1d6p/CyRJiZKoq4BTXyEqbrpZ+EGuqHi5eFknbQq7gY1S9GjTIXEo26B6x7Am
Cy3YIUqOwcVVJycEO12UosH/uTlQCdQUjR/ZOQgUJboNgHJTELtQBRTvUxzgMuj3IdMBcrP7UG3z
dVLNdSrtTuPar22d+JguDHbZqruKZIrU1Fwnx5S95vWjAoEJ36+OtJWGm6yg0fqTBTOvR4Mn/IOD
VFUyA5N8Xw9wkqiuw41dL6MuO7V0JnWlWS9MRp+eojWFkrE4PcEv7ktd8AsFFYTxHKDqqZ6yrWMr
Om4+WCYDx8dw16g72tq4jDv6i0GeqtGsfNmow2qUBWrJUl+Cggu5X1okLJSJXafF8FNXJUfB1RZ2
W7HjNR2T1+NOqYFuLVh98/QUguKDN+ueyp4PHlPWdz6rhd+T/paBHasqeLjaGYerVrV2dFRpcOSL
hlOPxiO6xE/RJtosd9SuRP+3+VuDpy7UNJJ5izIYVfZhjyOm/oHsBL56WPYMd8xg+AWNHoZ034VV
NpLmA01RnJU60K4R07I0vXQKXtHDS+NMSZR7ZqSTICRSODL4SntUd0oleSL+/ZdldtLFeq/JG6VL
tOzoZfxDpAWDlJv0EjqOJYLwj3QNTq8hHZTF1MRtdGhsYcfT8blW6IX1PuUbU8MVTldZ400LcXvu
3jML6stdcPWLQ8Wtmi4rm0/ZUxjpaxsFK/i1mQlgc+f0aHIpLEnF/vMd5b5caU0EkpDZM9YDwnfC
e44SCgoLDcTaHnwrU3XhuDaaPWhFIp9ZbTBNdTPMgY26pH9cGkY9ZB6l3se41eY5lWvvZCX9pO/3
XkxgnbyoRZ6wv0NhbhiomGp4TGHqS8J3j38z4xB/p3Z977xaFftUmgXMR7Kjy7MW+jpr62n+S5Ss
mnoSRgrt1oNBXaUz6vZYHHuqBvZ2x7yTEeLLKaxum9Ot6pbdWJVqRNOSVuk628DIW3+G2mP/DGBn
by1OwN4jvxfI+bbD8WGAaSLTb5Y07HQGcnXY/pkWiVLXzz0Ayhfd/di014pvsdPb/6s6rzbPrDFF
C4sndsscsKyJuDmp4804llxrHFzQpIBbpaBWbYGbCws++FGyG7jlXyEzs4ZZe9tLB7YEVvg/UZm8
18FkYroeS50o47YF10BNCmZ/1jMpfWjiwrga5YbSolleE8L1oeNV2KZrGJLQspcQKMTIZx+TNn9/
zlEmwXChNAfD7PSfGC77kKgMUUgWmK3dZh7qC934OIg5WCKEDspmGBMOCij2UgDH9QiumT6XL0DO
zlUf9+nFdsX97kMvRoOyzew0+Kkv6lP8UT34iG/FZZPJGoR/9nxmS5U2/7iafqBzPlrz7xEpOEa1
S/+UER9+4UrD0oNKXls63aebK+HUY5sXE8FhWoKNHCtkTaqgKuEwRxVpNa8quSv3aVPGA0htexn5
TcTXXQ7J70Qj6CeaSnc9/eIrl8SDN0B8hHYu6QOXt1s2vjU/IUdgiSNqY22UT67bg2BoPhkQ2mk0
gk5GCN2U1Akc2TLh52eNdqto2jgOuen3RsyELNlni1B0ZJN+QV94lSEbmJlnFy+y2Pyt7/w9FeQw
0fvQHdChBYo0I2w9OKi82ACkw/Q3X9z3o1NvlmZf9cVkh9Al2IRe26XGk9Km+nw8E1mGOJvAa38m
GG/O1kwjGColn0WUU3Y+bIbGu+yKV9v5OOJ9aH0pBhFjCgsm2YkdJIbYx0t8iKDoedhgU9+XzgEm
MSjPGsfJzpMrCl5tR/E+qSqEcaFCfA586OV8nHY2MU9bX7IIqNaAfQa6VwgJBP1pSsoFTGKUs+U7
F/X/nXPkOMd38itkfLFp8faXC6+t/arq+R5YgVVKHZ3scnEKz64tPjDUnvKcT8Gy50YivV4FCOda
BW3Jw2Tjgmrk53Ho+UdYGUF6ApE04ZGv6mywyjdJ2T1hgO/eKocMAGnQOZq368LRgCBSWpyB4nlu
Xlfw6jG2j9R/h5DD0bD4kTM4St/u2zL07dnA1VcJTiehbxhnxYI2kCLbygnnizGCONllZsYl/Fwi
RLDL2haG60DrQMsov25t+Y4rkFQgFdYBPcF79w6C4pbUkZlW7McRJRc2YJT27ZdHIm1Ae8YI706B
zVc3sS3iFbTgEMAIGxHpli972yd6dl9Phup6xIoLsRrVcs+nvaGaO0BbNcJ56xy3NHUDebjWcIyb
pUb+P5XAVwZwSeZ1tq1suZ6sBQyXwA7/+wtMh9oQkbaIHlAOnZ8yTyY8S4VF9/J3w+0t/oQO6im5
fyUg+NNR2OiuejtyDrGfwqgnT26YbO8F8r9BHtIK7Q3rH0/DozaK7q3rFfClUXmuMJ5kX4lyW7QI
bI6fdQZD0U0myxfQR8ltj1xl7xGkuBJVf2LH9GiQPS8BTKh7hSQjdFWNxiTEoU7C+hMjaxYJgUzt
OAgpoTsWv34Z/bS+cY38O9RbKLawrAAO7TJwgmw3fUMGQckXrM8d7UkCwLQmWtx5tdUYBK7MXeeR
/OjWNE9YazsCigbcSKc2Z71e4pA/HXmfygluXPlKmDd32fppN+DbhyMk7IEFfrRKEr2Q/CDpXiAs
Z8secQuYXrJ75uVTDsz8Ll50fay+M0Qt194A1rECLGl0vlB2xhSNqlCUDvnHKfrfboljS7QWPkQE
ZG4Vgvla+6acvoyw5AWdtum+5fXDoGKb7k8zTD3YEG18JFyJ2pSIIunL6Mm2dB9UGx8IwNlNxNts
fCSio60JaCPYmbWFnqtY3fvbByPHRhAnEgIYnEZNeoMg8PKWr5Na74CO0EOGGE7vVlMWoxKvMdDM
ssh/3/A7fWYg9h6uwVlEDyxMHej8kYVsqGYxeNM3donwXEcqFMKo/gzq3cQ4WU9SgFC2SYPBJux8
uyRItbiomoqgO6boxQMTzq/BPXbVGsp9ZbWR4mBE+0dQiskbD0NEeysEuJm145R2/soB9IHwSdQV
uVSJIfeicubR39vZ/pPFtjTzooFCHUW9EfAr1ZFUTN4RJottt8ardmfXzj5lfOWYzd3RF5jx4JLi
zra7Dk0V7jrHooiZOpTTply9InTJZFfI4MReKQPwdRHnTp//WAVRoc7cVOadcOxnB87zqygMiO1N
Qj9QqbkYt/faD7u5XpaioYH3K29GqAP7SulFDmv+6yB7bUrHgJnds3w/NigkSTodvEhGlWheH+Wg
b+QbJ2XOUi6Xa4JXNLj5y57i9EFTOu2MDZaMFwz9kfqWobnCTKsxlRwQoVO0H7f6anmTGD8pkbeJ
pUPwIkas+6qrXiJ/digGCjx04r8xKPgeVhb+W5/dcJVpWllokfxYHPWkSN8NQsvMFrfRedD4kQH3
dfF17kctBo3XqY2tf31AyMJKnP6E7yD6Enc6udXn1cbmbAudmXZtoI71Q1IArZ6W8LY4wlDlz1Qr
5iHZuFeXMsBylzmtdyaujhCEeLC/gWmz8XTO1+tHjKvOisbPEra6mAOWuSGA8i46shhf9D1NGX6U
7N9MDkCj/Z34sC4+EFwXhMP170go7GCX8mKZbJATwFv9zFvxweH4W4B6XjoFbmacP5xynBd6w6PX
/IGnGj64h1Jchl3yRu25M5anCwLey21p55M3Rbk2Ld51jh7QihOTymv+ztW0M3+Z3gSD2fxoIeAB
ljF/iTu4IDhn685zy4JjWyCaEyy++r/bby/4KlNTCkeETVc6gZS2HTTPQlWGGBWHvTwT+gkHG4EY
TIGnQ4lR7miHfMYFaaHBnGsUG4hZHL4yK161rej716n0sG/+vcSK2u3onZ1oqByag79hwI61TTRG
SDgnMGrFD7X9GcSpDk0UB4P4Xr5XDBVc0lQVhjQ55tI9RmKLVFEBpYOoIqxLRnT8BlLuWrvy77c2
wBeFpGTa+R3riwoVc+y8zs/VTfYnrWgIjbKXMKRkOZ+9WYVWph+Ff4t/OfogYuS/YQtJHlu1A65o
ykyywG+1avtYVvpQKA41waSTX8yosqX3EWLr6x5N8MqpH3rhVH7b8vSfZlhwbC7sjSY/tlMk/Rv1
4g/QN17Jqfzc69y2J+7WZT6dxdf8M1ExVPngCKUmj1ycZMU8oT4TPhxhDE1jlaykNKiiMgaRY5Yi
KXJ4Z41iYCmYkrhd4amjK4rU+hlA/waw/f3LyCtkxeTdVZiWK2qhtxys5RpsB/ifq26vcrOX2GOu
nEWWXBsteTAWqdZ3Qu11w/s2CQrCRXUelWw5R9GVIQHJNHMDnDhZ5p2GKjas45sZZqOnUkKzmrqR
TeCqEBkK+VMJKAI94wratz0y9O7zDj0HfaJKq+hJq0XvJGxzcClY4EBfx+n71MiZLunxqBF92X+M
dOODTC/QYi2XqYZp2Q7AF1OPC1PUIRbyTRgpIgbuymPq6nv0ZB+n7Vt9rCnsqWIc4omcT8h/BUlx
p/f9py4Ey9OOc/nOSZ50W+9RXTTyaBNp4Ho7V77p7QcOSsObWm8vCw4rf59SrelhBQVrg73TWAFo
4e9d9StzyiuXeXfhJILgkXbwRIFiwIyzo7/V4j0zw6fODDgQwkKDar1NGeDLWz0cIiCtNV78Q2Kc
htRKdH8vOtYGDHptjzxUkMeIbV3+hC9fQYKrf1sbui0zHM8pYYlUulsgzwy6Sh0CEthsiqxcoRIa
Xn1gpFgLsPME87BiiphorVdahPXkBL8RdB8b99crLQEXR5VEnooXQ8378MQvKNu8rKkYF9dzXBTd
5lBjKgWFSPgMQs4h7mXmJ1i453g9abG8jTwGSxVYp+0J1lLTKilPChgs5BJsw9wklLQK2zQsJH4z
RsopTJg5BKMU0qsK9N5JaKHxcCXHBTgP1zLog7R5l9UxwyYq4hFOdrkvsPJ3DkQaVYNe8eyXm8DD
2WTcPUxT1QFcq6hBjPcInZyQqaXAWQz+NoCC1qG0Z5xumDx7q3uMyuiPCa0QsoWzaopseFlgwBmW
OUinv+lWCY0VZ8IrXuc7v2k5Y/Ma+cCVvVMPbQakEa8tbnic9/ik+T4fqE/nuHRHdMs+m65deE7v
4aATmI3t9kXS/ATf3zf2mDXuhCDT/5z2eVaD74o/r0AeZLtoZIOnoZPyiu7+gTnpFYvlvmPElKVU
ZHVz3NsFefP3dLyYr/x5DymmIzSiWFKF/bSOYTlf9hQjIIk2aVn+i/44iAPzRdj6eTDYwAtpYH+y
2zUn2b2R6dEFjWN7gaVz4F2HnpczkVnS7v6Q3JuPMOOxZCTUsBMhobJ2DD7q5REyoAQllBoBazFJ
NzeIvRxICBEHThL9GxFILLSPcpBb3Ihd+wS8f0WqTRy2h0gZSUNjcdn7AifZE6z6fX/+KZM4/+T9
tb4yjuT2PZSiUAA7vNaQFX+K+qdo6GLDgZlXmg9O5lHtWkt7zQQ/o3gVIkSkfG8mb2NYBnT/+cJX
Mk0jEY6FeI0E1JgtzTF+GdK2mSYjGjbua4SxrP36LM/bMRNxknkx8K0kwaq/rbUqOB2ZXrZa2AYR
knGS+yyKrghai2mp9yPsJFj3CV2+qhJP6RV+0cI5Ajp7Z+GD8GUsOw/T1gciAJbeLDx400/GE3gi
7nrBetjnxFIjkPnQoT/Hmhj7IArnews5iguGB1ukvONvrWFx+KQqbgqrHmTIsLzwUIi3TKcqyQnR
RHuZRfnOILwFl2nWGC3Tt68+oMvu7aZmPEU7N11US/CZqRYPuw2iWFYExh2/BULChkJURXTsIgqW
4+RHq7Z8dQgTLYyFS0Y1O9Ml/zIgGs2OJjx4hakYq6Vub7BgMMo2668k+MPFDKWZ3fvoj39FOsca
gLdZat2bhx7l19colz8LztXJ7s4PDZpEXo57Hw0g30/Ypg4PtEcvuWGuVbe3DUhHZ/K1K2anI0/n
Xygaew5AvAwxzICeXFoz8mEjKeMcCNn0kyNcv3XXMd82p13s8+cDM/dACUZ69PhjjainAItLaL+6
7r21SWtwnWYp+4zy3hDRnAYvmlU/Zylc2NJZ1oWhVS5R8155hrwgBg4rzNEpxv8oWKUDirieiRys
mWRP+axB9+oyoE4UnCwzHydyxDwOScRRN8bRRIM5vP7DbY7xQYZHtE3Qvit5LHENjHeaxfzrYg0v
z09uO+jCKkOA8uwS9zjuu8q/Fu8NwdoiEfp9DlKBFME7OJNhuwAbCRw08y+F4sbQVU+GGR+1l0b8
DpF6HR7+tOHUb0An0vWXGcbO05q56kGrMuE43qGsQd3Q0I16Bp4ccWbxjerKjclSKDOzh+FqUPBh
khW4THMqhgKTIhfk4IKNbx/ejDsnHbUyG57m1naPVV6HJpAXPqiJ/8qN6M4sSPGklVADM1o0QWj0
igix7w/m3w6GUvVOmmZf5oE/Ncc88sI7OqVcrdp3gL6gsiO9WaRIgd/SILDj6RVKwJtjMQAIffqX
SF8w7IWg3QirrGr+3zmGDpuJpul1do0IuVfVvcXkUOVYH3z4ECHJdQN+ZFeE0nXueME6bQxeGKgO
Pi9IAu230yZChZzRjD+JVk57WfKU1Sfooh3cTu7zQsuuUa4ju2rxperSGw+5zkcD1jAvAuaMuHz7
2x0LpWZRryk5d+lzFy0zZO+UmayenHcPmJBzDHHxaVl2JFK8vtT0DQ2yORCutXfoqvdXT+g9YndB
LjC1tVmLWnlE00LufqG4PbXrZW3Lhstq2vBoJyG5HgQ0i7MXsHauCgmB3N2p5oNw6cqa1OZYFJsS
7awFcSm9LOUyi2nExbCAosbw+FRxwjSryIP8LtDMEGw6rN5icwPyz+4pQHW1EHq9ppLIp5Q7HyUL
/Dgg2vdRV1lMaeGGk5x2vzTfbM1SUK49wzB0lHOKdtFgmSTyM080SvX4zvGEhNPUhdv+QZaRxJR4
0tMINUuqAoL98h90jAS3fbDA4lC5ynXd2yjxD6mY4sfPoQU7pFsvY5ab5Cy6RYbuAaFNEzCND7Br
Y8d/CKNRbu/7pm5QNSPMPePjn2juK5ICp6BO21dnnfiN4Y/yiM+uh7U6R1X+CRKhBXVAcSnvwwKU
BB6DHUplRHs89mjV9kjC52T7aKZiRNQdpdJS2WvQG4tH/4ZuH5B4D8wBUBP6MOD6UPEfp5myo2o2
PqRS8PP7mXTRn+PdMptbTd75CXLbS+pKaCdsMMGa+j0t+cna4EngIcGqB7HQpnTpu3Yu/Lm/eiF/
CuujUAKQwnEn3FHDicknJzAyMwlB4sccLROdjuLvaN4Zm1S6TEdsn36q5lyxGubb7qDg1cZcz9Do
GOCZJGMe/7giaC0v7e3S+e0NN0pboN0jxauzGVSZ3L5VqTac9CQWIiuXjcYiwEzcqnNdN5r/b4IQ
qqRocLAS5PfymfsvpxHQbwexWytwGEyJzzxVQPmoR6oMhYL9kHNtVdt61fg3wnM1vIDklx2fCS9a
orjECQNO9C6va5zD1D77pyMlcdT6azx517a8BDEgP2XIIxQivm8u7Gpl9scx8cHmPfi8oTIXEtHE
8ehuJ9tmG/WPnaXkifuXHV+41BFfK2A1IDnYph5Wn8CD0RjjEYgPhH73hyI1hv5dtmtunA9/RGvQ
r8ROPXi2YAB5hdZ7Q/9lJ2YgbKA8vMtj0GBJkQMQdWQ3J9uRNlakiPKWmKS6wMbQ34E08NuOpRhM
5Z/57eCDns+VGGyCNQOaVosQjFGuwyypIB3KXyB8ODeE8VHKxqxq/ftZ6B1CnEOFGu2X1PehCT2F
HTKR3WSKvpLhloqVCM/r4ti2MYbsp0YhAKvt/3QIH8M6gGzbS29auOJ9Yx/iILKvxXOvVYL3Ny4j
Lm7PVY+a8x+0xulplFJT6k8cM7szI/GpQGhgLiT6NTnY5BFWKmSX+zZwDnKUsDAJzXRCbbjqkM3u
YCyDltwFajkoBKv4abmin1H8MDtII8sfxdQTUouE9nnUWTb0U7ySoLEj11Hfotubv7Z4r61ByNrU
32xzjpTXmhKTOnPp8v39oji+RWWxXLD2EHAEeFssUMd9t2tSPvCWISeAnKbJZvNBIK2maCFeK50c
TGHku8sv87EgKweXiBxAkaN8YnxN241DguMYw1PqlGhTwTfBRLr+iPTttYO4/B64/+o40FGxr/ey
X9kReyqJzAaed4X/Tt/3NyFbI0/doEjzun/H4tdYUGD3zGnkb81qM/TOI+7ag6w1tb4wht5HsBvf
4B1pR/QonCSm3XD8tIThDtAh+BCCCqoiQpKNwtAa9uwo1ZpDmt3y+m6Wj8flOn27j9uwizpCLXx/
iezoq7cFFGAt493NS6LaWBWmrfk8GHCCMsfhGqnjeDASV37WoCfISqpMWl4t9odZodg2ZqNQBxih
zsNNv+HB/aRwR/84jeaje7D8BQqZbEhfjV/xjq+Uw5+nnSOZq5GhAigGBw2S4dqYHJ0wryi+7nkP
dHcXw8L3OwfvnyWIrZsyQJqIp7cuSn7DoQlg4ZKCo4MlOePJ8FdG+Y+bWHsC5Z3n/7sijSi1RUJM
v1DlM6oIgyyF19l8D2cOyE0vQrpIwPWwzht9wCa2eMfT4Lbsoe/g2Rll34HHfWQki2Mg4Ze6W1Z6
H3vw7yTf5mL/9zjhbU0OKAB/zQ4P5zi7cfq1Bh2AwEDAOXrQ5tOUMZYDIHJnsmfhJfYYLBEmO44j
JV121VydVBcr0GaVLUQEBUs8/5MV/Oja2t2DoIOmO6fqFDheFsk/Rek+YBVMnNQ0mYFyBlzB6fvj
0XI+CePdguEUgLMj2nROEmEYPbdz1awrhbAN8nrms+74d+b9SVjuJMkgyhgiR1FWlofKtPr7Fecw
hCVEfdrGm0ZOutK8ROtLhtHuKp5KbyZ2/n9vkjtCsyL9TNDGEnbvHW4njymhCvz9a2Nix7EsiugT
bjMHPagivl67Dc6lLuUkxmMvrs0/B1MJDfCOOy3RcA029bFqrY9h9sHI7U7aiWPLg55FKCk1tz62
3WZ3ZQq0CNsVayf5XAvldid2wmge4isQEsTwhuGknGbrzP9qE5qBrOmKr80w763FjCPUXshNpefp
9FsHk+LaZgkXavUlG3zh7T+Aq4VWaAEdcLY9hkyeBPiDUm/fI6z79tLw/TaZLCyblkI2OUMdEoKz
mCrTGkcBjqHX8W78n8T/tobdVradu7dUyTxe4NJ5tn+IwGTigbtA8+QJlYEPHGNWEmVixDJ7gtCf
dl9qdHl4hXMEZQmLzs2dO1rYYShmSA2G45abVHcWB52srw0F8F84wCZRitfI6L/NsCSF52E6XknT
LBYulzJupYx96b+4U0xnUNhBSbbK4RuoelXXHe2VhjI/CMY7IZScB+7kRNABX5kY6vQafNbIeYRi
9cgsg6FNjwlygNlnrznW9p8T+rh4QUEUUD9xLsJRAXObvaRqt3FTE224r4rYr73y2ZZTU6rQy8c2
gtJLqR9VrzsBIW0zaz1BaJwCK0pTIXZZgo6bgUGUmYQ9zYbLridv0pc9bNon3/xEVf8TD/VNOG76
7Vu2nGDSI7lpHjdOLknMKosTF90ulWYIBfSXWvNPfzlAdMABh81GfCBmPCP4/pGg2zojz29RTXxR
puorEMvSeUTcUcBDPql025jgraI63jFabVFoxyCJe2mBxQdtcZfrMf1ZFOvAIIfCi7ahAkKNUx0P
HN5iv/d7TdhQCKrs1Kg5qwrQwUlAVqdlpxrWqNaRjUhNo2xDW7+IZ4wiOm8QcVGlGvLdVSqAWeNg
Is4PJat69VRCVYLaO1bz3o0MBEQa22UdrLL2PNmbZBHkAUm6SNcU/Gq4jjeK46BewRB+4mlFVEM4
IpKVXqUFeiQh7Nj6HY7wwx4Bdhs0LZgGgS1SPhtFNGXCP5kr7Wa/4+YIdJSDfPWF4hAb4MFqBFh1
UR3Nqrxe8s582zF8suwBib/FSTsGpcBWaJ6ZhwYbW6CajKpYIP/Sp0dBVpAajpAKIoqOjKilbQsX
g9uc3jV7wM8lk3S/8hlzbUw3zQxCEjJY9ShUhehBO8HOvo/oLf1wvi2I5B7Am3V0l34oDT8Eka4b
xFp2dUHrExNLg8uIruO36S0tbIRiDcd1UL+UjpYY1kKt0Oq2OpjKGRbaTCf106JElEjZw+NzbpNG
6hYjnl0fzzMmJ9AMGVwufv3G3ZOJO6kBhBG38Cel2hbLZMq/WifJvJFFdXfUlnJSsMS2z9aXL0Xb
2n+pf0A3ii6wCOYx2HgVYK0NQXLn3Qo8eONB/nTPYD/uOmkw0YUAToFqcLx8BLRJeQ5m4isAjQnb
TMp9mB8nkqLhMJ7v7jYgAHA1t/e+xYoMyR7m6TjODuNatjg8usOF7Fj0WgFKBgpH04Tl2vyFXBr1
6Gy6/s8woCxph/b7eHcu3/WA+GTmhClIpPqL2ac6eLdgXV49zXHPIpmAEIJy8wBotIQurVxy2WhF
09rKtJ2QRhwxgf5gsdfa9FRno73YVbDncNR8kLaVMgchYN4sxWPyRWrM7skEADCzm/xDna8LPkTS
SsesGH/YDWnkNcpxISg8umhjHGOh4BuoTuIeu6vhztf7VXsQhmcGxOZFNe1rZlg2GuQUmI6Vnwcq
jQdwwdscB89hgCzubVyGfcl/62LfxbFdSzqzuEAdIqhxziQtkX6Maacdt6GqgVRf2QZfsxGKjPpS
n5GKq4AEqMu77GzoJ4pG46zaKekhgg3vBk7jc6GFsl7m1kBYnrc4bG1qECBi2W8kWIxZzdJgGUmT
8MiG8D1pHDmrANyRuvxaOIHgOHmZPkAHtzIy1GfOfu2hk+LbkOxXDIWFfNitbQb0V75pIXIPOlKy
QE2+XTQWbMmiEAX3z43foHcN4SIqOy09ku/O+apX3brgTmR8RCRoLvUP9kea0qxd8pEjHQKIc6QI
R3Li/f3c34PfGzdUHDvHzPn62hmtDJrc4ZjbUAM1iRt0HNpR38RdzCO1AP1yIypCFveF1a+c09xD
/3bUjDQqY5+EhymznKf6DeniXh4qTBvjDZN5ZQCq67QduLDzGXxZHOxp/O30a2IKKB9aAc3XPEtE
qyWw30QVix1+/tYSRDLs5/LSz//uwcd4rpeutuKrJ+MJQK+ZuP6y53W01V3v4BYpjxBg1gvk3cEP
p081eMbpFUHCfpCiWtliqvov1GU+ELv3qCa9zE30oviRuM6GycJtlAnsk3ysG2WELpSUPqPni6E+
AxX46DHyGcMh8sUQv93oAM1SsB7lBjgLFU9oig1hthpRXPpcZvrrZKVMFToTjUA5v+r2O35mtKC5
HyWc9SR4bn4x8l+jo7i6wnlbEbAuEspsp+0NlggQG9eSAU6/709PhLSivCfSwIMH8cSWQcrO2MGp
JKHAQRBGv3MRZ4UwgOvcPOhXLahehMBQkIHWr5FTZZJEK8NIrtVvt4vQWDcpqcmm0DNJ3j7WNqOd
zPivG8dV07EFWGDfRJm3T7FFOKw1GWXrs6Y0p9uFk2ZrNvn5WKbWSjF0oy5+p1dAUWK2j+cVB1jz
nHZrBWpMA6sKjOKz5EGIa0E3GyvVgN58UgYjBwxZq3rTCOyaucdtnyRP9SseN1TkIiLzrWx2JxIc
60lMjVTxzFdPt87UMS7uB7pv7FaKlN5dVk4hDUbukCI7AqiXo20osF7q8NnJpq8yJ0vU3LKrT0PU
b3FaIz4Fvh/a9AbAPIOaHzoc+mFCcemd5UhypOIMeGua38xGR+PXdNeQ90dATcNPtuFyb8u6Nc9g
GAyRAH8BaDLesVQkvJCStwoA/GDbynGHeCm2JywXD8WkuqmLEvS8d2Vv6KSwZXsJxqiiff5e6mII
W6KopTcQ70niKViNdePISwReechEZLfpDdDkcR9+phj2Y+XeKM8WdmztAEOQ+7QKXSZt+kEzhGoa
HbGxVhqz2EEW9xFdCSzvDWFbH6lPPBAqQ5/3peYaeBPC/kNR7vW3AoBk1uBIbqk1HLqRN98zHRXx
XG/DHCwhQwXyfEba3b9B1DPihD/hIOhgBgL/wtBYHbsLHV8uCY/AWt8ZEqScxmJwHxtdt6HXMnU9
Dp1FfupOa0jLPmuTDvOT0h9YvG7yXFnq8SN/IJbZGhwBQ0cy+v6KjiJ2MJGnJKU9TcDItZncp/ww
yTl2CQLvOdoblNkfQ1gU1m2WfiL7UP5p9ttZV4w+HfZ1u3PR3I9+Fb6NQemUoAhyT7+F9zqDa68g
VUgbng4uIYxgesBnc+IQ0L7YpYap5wRzDEfaI4DhOT+5xqv/4vcJYESCFS5sguIfW37jpwIdQiPF
FFBXZgasxfs6Iar80wqNAo7O2ePfVvgxjd0AHyRVrE04pKDwq4ReZxgMdZ6gQuTpvVKEq38h4QW3
Hwb0GNaUN/EmjsYpLxa0z0DlwgkS3kLlfw0aJLz4jCJo3fVZSioLEyWYnEB5597CjagY4c2HNATV
+RkdQp7GoOJebsZswcgeL6R/eyjDp3LYEWZ4fl6IlMMMde0I/7uiX6d08wpbGcojJMpEOgVXEltD
N7Gl3Sy4sF/uBuvGMBNfzSyGgledQDNTtKWKYfP3HJkWaUZBC6wXRL6VhUPKL6xM+tIq9wQRjFJL
/Xh2Jd6pZ3HYxJ4+8gBCYyRWXzUXJZcs/ISwRrqrkA0/QVMkg4f5VM0vI0/mBwps8C5e/3tD/q8y
0uxTDKvwiEqODy8xb1zyfXvi4Gonk+lzSyanVwMPKAmQw4PTv00sGLBM0y1GKLypI9Dz3/BAqxFc
T9qEGaz0YRsD6S3m0FUtsmn8F7p0On5C0+VB/3DpUqVCE4iSyyTeE6jvjqRdI8TairDc+rHXjpeG
SPBL9eU1qm0xcDVG/x/0oLbgF/5VZ5iOONglvdJXZGMKunTbolfKutwRkU0KElb5Wn5Ljwy2+fAL
TZvJeJkGuFs7P0ipgVoBrZlEsYV5I/k4KBwyOhZi9r2fVRuM5uWuW4J0M8Q3XHQf6AQ5gbDwyGiS
CnT2FpD/Sz6fg5aiOGJlm9jtXmYQCPWWcPE9Oo+lHnAWcwfH4gVVXm5kvUYgXY1T7GhodpM4YD8F
0DCEtlSicUk3MnE3KxEgzLOwBrAUn77/3lSdJaCDqloFJKV8aO5QRBcxgQaiHFDp9tGog3YcdNN0
ZPBozVs9nCeQ8at31mPQdPK5pE2KY5usL+bZrjM9/fz5hk1ZAx6A83gEitmU4gLx1YbWwu95gVqg
TDhxhUiJJ086MR0C+2FVxIKoV4Kv5lRBTo8rhbOxMGAXntSQRKZGDXfRxlcjjMWeiKCrmeu484Ro
i6UG77HvvpuQDjdZWV7cOPgnIydrJFN2krQHEgh5Ks2oPzyuUvvVX7NxLQ3Co18B/zKeQzba4qC9
adtJ0Ubb30i8PlqSF1120xcY5WnljNP0laiCLLnLdtvCAIZ2pdqv3kgw0GPxooMW9R1iD8Hi3xeC
QAZrPlvWSfZuBhbILWj+GP1LKskTRToCI4rf8NBx5304QYwfWn2o2IkezFjz2VsdfmDf8OKFyooU
GWafrZH6O0xHl6FQ5+FztYH34+K7NWW6n4xG9YjtIKdfnwia59JuTG7Gyjk+ppId7Bjt3KWd/XzL
f5U17YRCMJIS5KuHhIrAgC/scWvHVwO24S3cL07YN4GpYdo1ofMvU4Jg2xGFfefvpOp6EMfrLoZy
ocAw0x9a00zTRpuYo52EDFUCuo01BwUyDXuI27OYW9YuK+DxOg25wb0K2bfeS0bfRC67AuNV5tZd
wK3gIn2OPjNYKxi6VbZcaXu4vFzUPhUuUs2pRwLmSTftTQXLnniskwGRYFRtsrS8axCKxG8rNukz
o8pQGeuWS8WBewy1w975c6LJoZDHZouJwce8YVcHvEX63SaPhHDPxw7aExIXaHUQEWZeJX2H8jrB
Hj98eAP7EKM1MIVJwsIeuyNPCyCHaeeUEwVMLOSSjyVthBr4VESLbmqBIBvpyF4vvC1fXmuc3N7Y
WiAZq+v4p9sUGRM7Ldt9L+EEWVDh1zKrku/3MPmxfmA/dFST6D6fnOffOlcKTysdk+PFoFS5TkKz
Zqlo1tRKoyfTpoL3t978naJd1c7uWWTgf3OUFFT/AkatkC60hqMC5DyX7n82qJyC7Ga7uZfmkWdg
N1KqViSzsnXaJkniwtp1xmKf/w1LWhtthjri38GgI5bBHsa0LDXIYzjTO2p1BCI7HoSx44zBUWYp
QDsTOj/2m9vZVCgs/kCrZJEa8x2WqA7whrn9P2WHlqalBVRp1YTfZuYqVdYWugi7WH17PF7kd8MI
y6r0dxcXCI9mQi7unUdHkKflYSH1BQ6pSHlVrPI1tDvmXg1pjHNxHToob76+P5ufKDW6JuNVxVb2
GiFpZ6E14Vqy90jOXQDR3qTpPjjQBAYV+xbnw13S0Q4Kg96fKtOsrY0212HcRg4Vg3t+chgqO6aF
CLkRURiUyeDXrnn6C1wfF1LcFEEO9OI0uVFct0JD+ffUfmNdgsp8I32S7OnFdEi3S8iY206kWqdX
gOqaojFebRJh+e9yuetBExT4c7G3E+bUtkT92eQIpcUgtZG0EeY3azSYpoKB72/9w062Lzxx37SC
tdGzwfUhKuITbB7Ac6xMgY8BucPCEOySXKVXgLOekWfvss6ukBUKJsttbmVbKmxxqwm+DV1rQb2w
MTkf2j9jZtcUYbpfUWVQBx9oajFBVeo8HODhwbUoXFcc8oZy1xIu6AozoL9I6yzYdQHsnsh3kCpg
VnEvvXqx8zpC/qXPyzyWFJLCu6zhLAQg1+gZJ29vzoKAi1+TCixEadIYyGG/0pDUigMzndcV55Hg
tLTuaHDJ5dLUz8VKQzwsca7TR+Q3iEZYy7T0yCfr7BEZEaaTmUk/l3pOS6wu7QBMec7cZZBDNo1t
xKC2LTXcb3detTiRdJeQmq3OEEe4xUOgblnnkCrdpIA/NYxZKi87PwbbM1FtYaJ6VEKX3K1piTJ8
tW+VaEN0LJgTCx+KOsU8EZJLe17xDZxbwea+Boo1RMvaPRAdg1L0uOpWfxc4XycGXMY7b/TgwDGQ
0VBS3eNzJhuDvyJsOI3m+Ci3YzQ+T5As9yj8xcaeuBxw6JP/7at8r4Vyu49RJGSRltres8SRhivt
l2K3XHbBVt94BffjcqLwtbv2Y5v+nN/h5ZclIMZugCZh41nRsN+7ShL10+DqU55x3WtEVwsXt6PV
KyZooSk4SvhLukA5Nkc2pTCsKc7PJQ//s8RkmzuM/MzWtlZfXLaXeObvrQJIC4g42wT7pidnCLDl
CzHxDIdYHs2IlyrKJTnpNmoS1nQC9yhcrhiP3P5C5Sv4vd2qvpNiExJC0O//0PA9fLWuUNuVrDFZ
RhPjqo5ec3c6gmMBgYV14TNckH7EolcvUPWnH/msQldK7W7pHQ0v+n3ry8308QKzEauI1m7CTFmc
185f0jNtdX9hLIjnwZ9EZTXBSVZ9OrPmNtWNVTp5s0k9vZzzLgx3gAtJZprlp6xpbG7C1Ta6dDZH
MTcoF3gtlJCfdnsNOZxdAiXihtxzIgcxxqMMyJpzwM7S2OiOhoyxZIMBKpP5ktOfIkOTlSlp1TUC
FnwjH22zqZXePGmX0+OaSHo3X4eE/xexewiAknxzd2XAweRdZyt36sNar7Xir9xS+IgaejFf1OoY
peLk0g+/cgsTlrkgeRNQac5A79RK3suoLdtIMgKXpDLJZ8CxATus7nPhyNypOsRqTC76nmmrnm30
MDms3bvtfaoorSj+5nIuxfEWXQcquaKdv3jpc1zD8gYUsrZvRlZY7t4Q+DiuV6sjzqhIQkDvWRRl
z6SoW42JVUq56yf7yuiAgDFuchJWnqfzlQoo1hdbkK2v2TrTjvtKWAGag131+aRkTtnNew7y1pHo
mDKNTp6ncAJ3DCmHKSmpWZDIDlIkc93vvYjdTnZI6MT5gewCFbggRMoe+cn6Zhub+UNoarNCdG1u
mW75A6cvmWBnPiPYwXQowE9sXIB1suaUGDRIDO3DgT0KiCadiBsTE+hwVX5ar7FNBKxU8INFrmoY
wxymTLPODf+tFxaulbq0jUts9fGP2f5giel8Zn2eRoLsWoX0RHCZlEvAvCMDdJ5LHWODooFXCl9t
uPQ8V+PPUN1fiA3Kqvp/VFpCYLm+usj1zk8vma3iPGn3W/KFWyz4Ln6pO7u9K3n9c4yNSmFmxtHl
hlJZ3b/6dL/Wlz6KzJjtqA5ZMpXFjkB1OpEFUdpRfM7C5tG7c4xyKoK6BrjGl3zVjiiBedGxzhTl
QLpxOtDaaKrUxiNFstVyn+VJ2PQYvz2Wcx7y7cE1PH64glqbrCpjeXnQvxxBkc1n9fm2SuwYUCRv
fglSlKvB2mmRDpHbF089ox2ORudhdcy20OZ2tzMnD8Yk/JjIvOLX9pd6kq7EAZEOIu5JZITG2Vs/
0yDSyJhEvY25DAmilqtSfzDF5VnBafzqEQ6cYfkjdGYCrjUlv0RBXXniUrMKJyAVjnGWFQXLT14x
0XqMd2CrCjZKKoOv/viSB1aTFZf9M4q9j9SChlaH6P4tyiFSeEr+XRwHx7BIHo8qDpuh6Dc/OeaQ
RgryxTfytSIL/yC4YUEc/zHqsgOuXDOhlwZCN3Zbx4rb5Bd0RQVhLjUM4+pz9RGoxgGlpXrnZpCk
T7jFK502c5Ua/mPb1NJoSSqvFjrPTpbd+Cocb6Y1lZynAF8Jbprn8OJV6pWjyrtgmwt8pTATRHqw
YKqSazu08XivOQ8ZhN7vnRhEiZmQDWHKV9Sy87IieDY8rHcBxr00ywX/f1dcuUZGpQBRyiVvNUpK
tZ3ZnlKosyDNrW4EjhRv9ANDFO2cy38T9R08BNLX0a56uXst7WpvHkek+O4wyPAMK6pmwu9sPByr
Ils0K+P2wmXAKfOXMFtyxBpCH6PzGMOo9fa8DadSPGWikmRoY0BzzIzZFZOS2WbjkidSxO5ux8R5
aYy0NuIs8PP/8aQuN0PyknLA27EB7dv0qNejHt/IvKk3Fq9nWCh2ZlvTZSnMfxgwr4lZjXVpPvqC
iUiBaVyZGRBXJlbVy1V6ng16j5jFeFdSkcv/+ccYl+tv2VVK549OYTJ+TwPMcyII/4OhBCL672yI
7ZY/f4Q6isBAY4oUguyCMH35HMXrPvYCgseoyGdJqudW8yvurlpKsnrwX1CNb3f68JRiZYw3Lk+6
DzTn7g1ZheeO+yhyy5t1NW3B9B5HlIKNtYSpubEFi+wRNgaDvjJttwDy6GrS/5i8VJ+8mz0fRz+4
VuB48cZP3qv+XRtrV9T0VcYjeXXcdxCQ6ofebnRmu133fBmGrZTGz6m95HxVjvnHiKeKtUknDGi2
PeX3z+sK0jU3xtvrjdHR1LzABK697y+cpG8jOuAF4IU/Myl6AdW0565E/MH+z39rsHz2+lF44/Dt
MQz7tl83cnSfLHVkb1hySOghaAQV++943QjeLJhgjisoKreHIGhtIV54RdLxqVaeqcom1DjS8E8k
2uzRC0ENnwDQ7q+4HyPgjFGL2ry/lBo6TXENmor8uwLkQYFCNTU4QMClBOI9i9q8/luApnyovQ8G
S8U1eSSZk30kPeOydPDxNEbVF0mxtqAqI2gDCao7gw/BYJ/AO3rwDytA5imC/cjJHV90FZqPmLLV
GWSeCT8Z2/CpknMv1AsqzcFrRA8/qLgzN58kNGe+KqzqK1dd/o30b7nLrymRDOqvidqu2pGWuOev
WXIft9VEMf+xGOaOUVamF0rfzqvVchk+fI/xkGBHO4fFny85FCaVZ9GcCdFKt6Oq6ORql1Z1pc2Q
hck3aArsjwCVuelaSUYjTrQlxQ7y1Gjm7zXIcIRx+zNHssWQKwvZTB2QfAxv/LM4De0V4F9FC6sy
BxCp1N1P+CcZ+xpraFzxJ5O7j99LCb1Ugt0qttLSSXGQ4goJYudFuREEr1YXsNGeIwb2pkJYjrev
tmKiTWfe6tE6gGpv4WHAAVR8z1Wms+KVpHfQt1bjMz1MvJ3uXqEaoihBx6EwwWOSqyCf1PAedV+x
FeMTNXy/mBBJtmbEJD/3siSVsNxPa2IN6i9tx8C1/PHcQpTMtFinxDlaP/FOjncgbNl2AodWUaQd
4u+7id6s7nJaiH+JIK5zi5sOoXUM6eL2vL7w4MyoTQKYu666hCL6FK1HJ/ybCLpYQqbzVrJRmDrT
Ffn6SL9tqJoFv69sVkf6AMiDa9JDqCKvs7wCm8lgDPqXsxUUIJKFHY7quNVbEByep1K/lS+elFkO
5vQneJJrOO7Bc6TTkVRX8GIFSTJgY897CMBSbqqPkW9RpLjxJF0EZg1DQYZFROIadcKRB4Vy5B/w
9TRTmOYp+WmVenHeBmqsJ0bWx091gmhZimAbdUkwxyG5BH9NsHkhtwOzx93fvKak/TKPy3XvguG6
LjJc8IBqhU3JAt0Dy2HSYkGtAyyipORx/WLFUvGPU7JsBp6/dI3WVjhhGPlKKM4AFj4X/jG6G4iE
aWtFH4SkTd/UmEV5zGUDF2mUMTRyG6Ua01N5iYLdsOe8/UfzhzZjF2ziv9hUkZveeHRWl2el327F
WZVm0V00lsgnpduR+mr6gN4AZFq4EK94qMM00ryp9ynNGmmtgOSqZhdUneFu32C4xdNQCvlm906B
X0khWZca8IbgUmMcVvza8Y03BCoapT4I1pP/+lFABRFG9ZO3FLmXe0i/5VsYPuKXUWMV/QdvyyG1
RV8qngQbCus92eS7wrvodBgh355lZOuHWUq21OatJgB4MJ2cRQPiBlQDJsDmf53JhT+hafzJ4PD1
ySObSpn3nV/WXDgULyzQdrp6hsHSg8TJqjK2R55CPAqBoNHNG+bBN3QOX9Sm4UkCfdBVsQrnevMD
CCyc3DHNN4M3AUjoaVdQQ8J2TbTNAy7q6ci0pNAUlU6nfxa/qDPKzaYDMyq2nez571cHVhhQ/8RZ
y0YBI1v/RC05knakHx0PPmu8e/GR322KlOCb8buMn5gngvXZlYZYDrXr4duBpGlf3euaKflKuOZX
puNg1/GkYsiaRm8S6EoI789KDG+zmPvUrZjQARGMzqEZT53zDbIgqGG+RdAog+HM38UMty/qNaqy
Ty5GDGnAKQY/6P/G3eMpIaG6z844etCPfyhrQEt51P6tvt13gXOvY3fN3wB9QFQfppe/l64PDMOy
K+D2bWuxplRP9HF9zShyUM9jCUIZeq7xKuaUOUVqGlY8eASEIj2xhjkZ621XKIFG85xRLhhBvsdX
BWcL23hyasUkmnRW5PKbIMJjZvxJx5ove9VIexoKM6dow732ZkvRcAAKFCWWJ2HGVUZjap77xWGA
Ebq40/ktA/SfkEWD5Nx67PTlT+fKTN7+y89cmHbmlEPfmb1mohbikXJz6LgrevEOw6Lb1TZ0a7bg
1pj0LMeeb/elUdmsBQrqkv7jXf4UeMAUml6LAx6iVYsPch/KEpLAPqh9jN0jNd0t9ONDLO9uU8Oe
bQ6t8iW/rftbKl0pmJ93PYCb4BaHSoH2wtDL0DWZVqfEAahdQczNjGz0M12WWqbJINujokK9TCty
/GNJF/+nZVjtDFV0LB8tApgdbYC+P2iNMYl8dEaMO5m4ScnCIn79eb1sn07qF58et3AZomNmcqPV
cjTBWyk0YwstcQdvGxXEgwog0tGyNfDE5JC8M0mFTND6ybR965WvyzZsnPxsYsoXlWbQzWaTphbO
Cryp/bMclRMqzw8jd1g7gGrkdsfGofF1gzEsi1rVmBgw798nWzvWuGV48nBs+gYYvxkCDAyeRwXv
nNJrFun6RZCHD5+c0stkC/SrGAym3POmSRc1r/pRlkOL94oXg/lnP9Rrmzt/36L0k1e1V7QQi7FY
aYp0OMnNRCjLLcoCxj4Z3BRhGHDkAJSSix1w0ElaDm/EVtyAiT5dFjnUYoeTXTYjf6Le8+u+MtL/
yMrUtBNwRffSoHZQaJFVNX1k9vLIG5pcFkvVM1LpRSw1y3PekvtjefL3nKNP9TfihGEGqyDNS+Ia
hG0cjIEeKzibjzvBsEewdZZ7yETyxq9S8rHks8Uht8yCBqE05/dflHRrKPJu0Lw12T9EvogVZI15
hPfcVo8359xHSVuayP5m7zy6VIlc0BIAylOIphMOoEjbLTQjSuiOd3Px+rzmfqL6uJxtP40F7yDF
fEAOJpVWk11/ppnC22jxOUDkNaE0VcradoUOSqnfAOI6OW2tkr/dk6mfbM4EjTIqwSvHH5C2nqhq
MrI6nJzlMeBO+dWDQuZqxxtmXN0rsG1pU6BEkbiJua6EsfCfU/4stCqDk5cGnvB1SBt+9fn+ejPk
6VsmdLPa6XyxS2LzATb/NBl56XJiTPLq3VxW/Zv16OFDji3Q+x7gHEUOYA9W4pwgmEvhgm1N+X+L
oyuf+2EKY+7Dole91M9xGdLii/4WStrAhRqsSuxAdBXA3GdDXAdemzCdBoBsWoFlbF/hvkI2QH+C
fCWnwGXmbWKfuCn1jxczee4QExncghE1Jn5xYvA2SeEle4Ed/8b0uzd8Jgt2JMIh7B/jvEN+/PhU
ElGRxn9WkhrtSMnHxERYSBCSoCV5ZvWhHQLDo+Pgh5X0Mj/HE3s6yhJO30W409e4M6RgWUg6WCqF
VSGnFoI1SoCUCSql5nc6Z3OTuQzGzLIIxNLlhLC6f+2wK3OvGLgRd4daMomUq149sb9Vs7ilfti5
dhL/DYLoJIeXzUxYHReKjmpgN3rdet4oFTI9kfa6fcnMxRRaqOh3nIwWDmuQ74f4JuPrMCRymyHV
+d7rr0MQ6Ka4aPqfFK7JPFAZqe8s9l++ay66gJc793hBVVf1jkry7fYBW6H8q82Nymx1etsOAk6m
slRB/1GmBAvhL2Vrw9OG0WX2IaSo1sVej7T9etPI3Zi4D+TYAEEAEACIswhqd2TiRRLtwYrtcPh5
f6rbA6Daxossutid0seJBlQDOjy0mbnLKG2Ii3AJn+TEUshVrtUNR5sN0quVQdELqVIy6LRkbcyK
BQdUw3I1mJ87y3Uajc85fJ7a8I/Yo8/2KQY8yLoYnK1lAduiGDFT252dwVY01B5cFmuvHttPBhTv
IE+afA9A0qhG/QRFC/wRfVsTNvw6lqJVp3jhqwkt4OyjvLrVhBUrjiHPU7WsXL9b1ctR7W91aUPR
N5UyGBS2odxlNW0djz2I3QUaSVAhTOBv7DLwdhtKaUoXtwMmP/4eqNZcQITXUwezBLTVIGzsaBW7
frVA3uhbxCRwofUmfbjiASdt4ut99wduHZC8LeFWyi1WNh0GftUew3d50RnlyomVi1wUAU67sEC4
8hP1af07w1f0ICfedTSgy3JrYVduoYKEutj6b08m2iLyxR7Ssj30cY8iZknV3oODoKhKZGFO7Lih
d1Ie9+8tdoLeLYqnlNPCk/JYiCotNbcTzcQCkgQudN1rkW8/pBQUklCNpSR4cq6HgKf0ncQHBeUQ
bEnHh3I9Q2IV9tAxoRddOv28FtmHTXFDcRlFy//PghKi7iLDSUrcEdvvubHdR6x4DjPJC68YwT6B
m0MDUd2qRp1vofaRfzizhvLV6enQuVoy8j20fUzEFdSmXA6eBDiPc8EZ+aBua2y6y4BWBqajENtt
HQ5EFSZASGIiVIbcarJi8CHn2poGeTBFuBC9jBe4TookiD1Ag3LwGZnm7W4MUYn+p/JB3s6eCs98
oxeFvSiN2hh0j5qMJIS//YBqosA3KiQK6ruyTZc7hYg6kXmajsDhGO+MroUfjlzJqcowFN2rZqwi
S2Mb/vMy3Rg/2y91QJ3DZUSUtPBTSG0oZ3wXf6QSgyt4aZ3SOrJehOoDDCx0/ZiUnbkfmRRZJs2W
YAoqY39iTTnZh+UHFybZYZ5fpnUy3QC0DCa3mG8iIk/JxCSnhXIqhgsdH2Dna3vGQLGOtx6du+xj
mycPzY19V33gsIkvY6zZfRdMhnEVMk9a/D2phmjT7IbVBseD0kGNLk2o6VDGEXWAykpiPb04MQvO
9oGoCiAmY0bTOT90/P3t6XT+7gFPCdDX4iI9I/XXii1yCoJkWUZYM0v/01vr8idfw8net+oyQOXO
L6U7+Fo2QJ4HqJ6IoI5dI80fKnenLs31iB4NrRL0h5C6Y4CrBqKl+ghM3RNpqPGw/c4HFXykvRNN
AIy43R4FrgmbdNtR6zevMICagcaywymL1CqcTvy7N0NDkBDYL/B1qMnbZQMzUJXMZwWa97binAnB
9VNHnZB41HVvhYh1k3Cy2wogWqm3tCRrByI0+mOSDfXKFdPSgnB++vP9gSbfuEOXKKYXAQkfUbpY
Uel7PZ/DN/M0a3Qt1r6/cmpnmJqH2HB1xhcFl2fJZTRSf7gakK9vBRV9YdLCGRlHwfaDAz60cjxj
yT/Kfisu4Ag7OE2CGlMztINjbepucV9mr8c7TysyfIVE1f0NwG3vTxMntXdyJQzewjvpmM11ZuIS
MLorhpZk2jzRwLNGBDnvnugykE8/01NeLHfGzfaiY4LpLV3u9lh8S6ZlEyclsQ9P2ofjPHlZlcOb
2mn1Zaks1jnA+y7/H/DivYw5NC9iJG67sBqyh4xJzqagiF2D1GE9bU0aHULjc1e23c91a2v2oJrH
7ufR2h+ZrvRQwqBlViRHaWiLJQYhyX/Qe1ib4Fq9kIz2GZlZMzw80xPdExowhmF72y5H85CE66SH
QlMCrM96Gm0TJffjw5fvLZKeXtLBWRea4My7sxJ3LfknwN51MlhtPexoOF7XL/ruYChnlvIgiKsk
R4YaKEmXCf0i1j3oYK4jKOBOaTO8lFLqBKjOppW8aeIBCgCfujX/Vb3lBm4rpzTL8d5qeCKxahqn
AzIAyMw4T7kgItXHtjIs9tNRTSppFRwrOdZb7fyK3p1pms3WrIT+YHsM+wQAJmkl1rmfBGzBXUpv
NtZNmqjHfgihavKtFqegw+bhwcAenkJWHYRczV9N6MpaBntmvWTBLVp5U2JJdssEFg1sULGmArsM
5FxFSAcozt1Hg6QAYNc6Ksbdhuz8kTMO7jsejbPi+K7tlWfHcOeK9sAb1KAOghUxsTBEBvMZf+vL
fP8hhzoh6Tiq3YKz5EKkbQuYrC3QV/FAf/52EGAmslspB854COmAQEVnTGKJ57/0Awj0eNYUpCGk
+RTakWDLk/M/PRGIhjsZx795iqQ/0sTcYmpAkXTp5Klz05zPz5DSXTWgWO/tJJV4ZWyDjkLIF6rR
Odl+nFdlmMVeCryuFihXDiOU/6YZY5eETS+aM6YLgbaJbHExsYXrk6WzjEWw5Whf7m9MJnKFkK6n
NoXcrbQc2QwNDN3rTDKhXdZowxhdpZ7GpNGgS3kBWlP6QQuY60FWm7pkbIxejMzYXCz8U0JS7b4d
Oqsg2THYkZQ1zx5YRIRkpcrJDGejNhLkAN91eL+vgWABGaOmhnxq6kXKkyMMtPjHsIWASjns0Hsg
HdRBUJwpyzUrNzM8L7lqM/U1lgLmnB1SSPHphaZqoLFpSIMWK5TSDRBJT6OYzHEHzYcxwL0yGwFd
Z4wpqADb28e5I3ksC5uuV57Cl4K3Reip+Qb808WlUsGxfnjNfvF+y0RfLAhV1Rr6IJpdGOLhXH7Y
/B4SKuELhcxJjwb7EQg34asbLgaXQmAvUbk79fTRxddqgkiNmIJyEZytoN39/SMm1EfEROLPvWb8
UqaooazyuK5Fl8qiTye/YnjqRl1hmas6tMsiooBryWzrU/xgLJ1Novv4Yr1it9tZkKxmAn+5PD7A
NwF8kV53rK9cCUyHjX000vYOWBSxO3u9ZhzzmbzD5lMx3AkN6BEaKJybRf23P49vybogMPQnauJd
1JWRNAlx1Xb/gTwgVblktrUxaVSEiTRE3K/tuapL98fDm4eNpXgwOlyku9gPfrFIo2+5Va2mdNd8
R5i4msBW9coBKJ8hesZpbyRnSf2wf65VGc6pC54lx2qtyONhOW/cd/E0od3tn48slZS5cD4CT3pS
FZLG9W0V+IaFjc+ubgltXLIqQf14/PkNn7Tsl2574BRq82tXNdnhmCSO3dstu+oUrH1BNZasPckz
EqVNuYmZSNtCBX9ylp9TrE+rSmZt4gg7IeirvQRmxgx9eh8cCchFWHeUPuba523YZ68UG/tDIcNX
hsozOYENU0JUsOcI73GdKTkPUHcLZvNKuv22LPggTjW/l8WIH25lbFm/Dlv9Jaxh7AO+skWAqn7K
Y2p7bYF0yccKsNbnas+pALeHbaEvCdfp4N45gXwxRIFX7Uzh+Gl6nSLjaVPuhohB6gD9LVcdCQv5
XDRLfGJkgmiSj8DyAA8MXFzKbieUwjFrq0HvOetMWocLd+QwbbenA2RMIuN3YHKSzZs48bNp3IaS
DubCfI/6BKyHTC9yItTpDWMBRRZyxeYJN5w+BsKhKJAVynta47reP0P0TKUxhOGewgYouoTHV250
ZjEgiAJQ9pEHJRalp23lwMYOOOFR6PzOewmMcAHO5BBiEXcZ0TsXKBq1Z8LdpXauRSaDq1NmPpJ6
fdMxUkNm5GhbyOaNbsRozho51b+/Qj/xZQ0v9e/HZ4L/xtqm9YFgLKVfA0jVe4I3BkjPoOptwwEm
wf4xYzrw/CuCie9NJQoep+ac/kK+oqavdPaEejCeFe97Hh9wmR91zPe3DakNUzZtNq5o9y0QW0M1
4VwkVZy4hKp92ELrEj8+hCHSPp/c8jkj7Hyu755kzES3/y2LDhxPmVfqm7AIbPkBM/8327QP2qJ7
9SCxL4b66SuiILadHoCWSyH3vga1ho8HohVO9n3kgJkp0SFRHNWfEge8DASskSCmt2u6WO8Jj9nw
ZorBlOGPK8i3WDUzvvNT18PAcjMdp2VIh3FTZtQ2IIj26wih7PIZvLVO1Wq5gphcbw/PChkT0dam
U0VcJ+5eA7TeMsLsAwtWvHQdnBfMFaqs6bYtWQuXYf7SkuNoi8ST1q9i4Buo2U7AnKuPGc2aYh1R
TirLExZTRi1kLYuLkRiodE6CCHEUoaskzwD1lQROBE5+z3fWwEIPZCjz725rlBG7HcsgGKaE2WRJ
yOxaCgl9WkyTYV2fchnByzPSVGsrNLTfewGqtDku3eYyJReOaoqnudtyL3bz0Hnf7eB/bB1mzz6u
j4PA24obgtgZIo3SmVGHfRvFdVDfqwlk2ErmrbjZy9b6ik48QQwHV/bSrFPresJ+KI43fNb3fSYL
XDc0t+uGZRFbVZmhURqPn+pvnu/7xNOjU/o1lzk40N1I6uEYn/IqITb2jO+EkbZGvPMy3SVoIwid
T5ni1qXh6+YzURM8Mc4mLUFrpD5Y/BHx6p0AK9o/jnbYqDA+GtxHsX6Q7eVXzlVFHTuChUlNvvfx
WUu3anGDl+RVoPlwEoA1xgGgR7oBfKy9usWEu1x2vdVK5aHR+daZthUr6cNJWnJ4E50R8AaW05Nr
MOgjWI7WtcDimcvr6f0JaKCoa5EiJaC3F2+d/sz7xiuyxj5nKITHFKHOwma8BBf4XeiXCXg2M53O
AIoUZXVfgi+xF1ej4Kjdep0O7KqiLWPzebn8Oq60CfB71XF22hI7XbaigNR7/Y8Jgnet4RxGFQue
1zpu1pZykdogSxnvY28KnvU/J71/AjVG7pMJIaL7xWbvRovEQwkgp4IvJ/8h4L81GvJ12U+nGzhr
0oqqKhC6/89GYuvE0eRFouYn8oBQts7u7GBPqyuKYZegRdGdgxZjyZSrvhrZj4Nb02L7vv0NCbfo
tASDPlBpVKl1QfXNcjl79iAtEblr6HMurKCDGOXKd815aob/8FbdSUMTMtl//1ucEBXMaoK6qK5y
P1IK8Nh+oUYe6lY6cz81yf9KpVq1u6OR6xfet1VATiI6p6Vj7PIcOeNo1/YsxZsfPPD7aigEHA3h
G0ose174Buz864pKD1aiC2UYSvlZ6qtHSc6iC+M1MkVWBnlXozfkQlFzo/0BGJ/wmqLhi38z5WOF
M1f8gjdXUzUNaSON0VYiWxtscIa9wpzT0TjQ0aj3mVQRyfIrH2sC0t2PtWQSB4LAZR78lzEXDZVZ
/TANK+UqeBhauuK1jSstoWvc8HGmT7W04df5SWl9gzVJpYe91K9+0O27mLQ4MdMaXbgxv18oQCzO
zTdpbQ6uJrkOgPb252NbNtyEjBx/GTrs1x+ilx5Nr/D42QRTMk+8+ARwzbcruix2TnuE7IzvcBwD
peCFqhwaFOeGmZhfRXJ5wBRr549+phcrorfm+JterfU2d0KCJybqIKshqaPyvtYcN8kC82Zc0UKy
GQpH6S4uVULbV5SeU2eWy0Ccf92MeodeXWStLupgqFu7AV34goNA+TRtkLIX1yc0sRxYFI0mUsPY
w7J1ZHGwQJ8hkLMO5tzFRtdQv0QeGhrfW6TEib8TJ24EtsZm6ZGYMZ+SPf6Y4O/m8WssV6FNWu0Z
3bbVxLbw5cIp9m+l3bjSce3WbyL2FmJmLOoxnBRxBfaPMmfUGNnHiAyWE8KSPhwP7OdHzqq6KlBz
VVm0eZ6ILBBb0/LfjBfigIukSTxvaG5GBj8Emero3skWcrdCBD51K32PH8IsWSjHya8SHXv0Xkcp
TFoTBgYEG0rLlFQKwHtmBrh22QItfYUyncZwEUva8crZYx1wpF0WrnyslPfydN35gu3MtkMT6sXb
enfqf/SP+W/oU0P7cJYm6PEoAK3jTC0DbAgZ+iou1rFwRMpnqwkZ7/0S+hp+lddNYPy1mXIhpExy
ea1dXhR5rY3D3LzsjB7cM7Y50aOgvrgkZERA6FPgbboqsDa3+wfmKWgGS7GUK5n+xEen8q6VQPte
qwhAdoxGwmaNRMluONaUl1ppnB+WG6KQajJLXpali2XXBBUm85Nb+a5xNPyBAJGvS4Tr654YKyIw
zUmim2GDoc5rHOsXNn/RyGMe1rgfjZK7ZPzLiEpON8LAngKJ8l22iGW/JpFvXrTESfahfBzd1yMr
6kYZJzwO1ydBFIFO8EJZXbaFI4ls+vwdO6drODYhXbj5vFOv2d4i5qp8xQtWYSjPbHCpUP3Sn41/
2esX+PY+EiHZDR6p4mZ5O3XPxX9FQDAlEg4wVhcVND9bkyNeSjYNa+DsnWFbGwug1RqpvdSjAFB1
Qgo8UT4yV2P+eHB4rq9l8iI7B//gS/1p+Lb9pIwcgrdTWF3f8LSa7OhhWVtZU4m4Ex6bK6TL3H6S
LRi4OV7Rc/JBGlkaPND7zarJsjlzXv0Ii4ri7UywKFADlRDZAAapaRJCb9fxw7o7C3LCuNKiW1QX
7CMnYft/24fnyeCprJh0LqxScHbO47eYnrrJnofknIZ6HCviwKXkkyJMN02jv1iuL5EwKt4IoiKE
5UK/yp4gaFx0xP65/4hzJMI1jiYJn9ryr3NPC04umetrO0TJS+VKWEu6Evg49MkKavfR1HW+jl2X
ZYOeYVrtK/jM640xB2d4ENdCgjkQk7tP2xGCSIdlpqFZy6E90LkhOPA2cBv8XhtunjvBw0kYAW5f
2vV4bFWwvlCkMej+DuMmB9lLgMKas5ia/uPJy3YmNv4uDjnBu6H8yPRDbUtLFC2Q2Y3Oz5Qv5Mmz
3y9SpHfgwsbJ9heMSCQQc8hXTZWBptmSCMTpbW16eoHKmq5aKKYhfNELtPIpOPPJFbK3uzr6p/5t
lFQbXF4hHT+KrmSqyapf4Ok2ME+91/fYkVyzrdYoTswaXXcydF1jzm4KX7VtwNHbk2agsqTQapcb
eqdgT1mr+qZigAeoYEsVnowZDo5p2Dft9n+aihxvfwa8d26qRr4An3YVPGl4IDpqSqshQgMfzm0Q
gNiYeUste9+N91cCJ6isORXu/XVtqB2hDZtLLnwf5We3uIgpV9w2+ss/3ao3xuI25g4olVaxv7HK
T+gsgKZWykvY85IKm90JX8/I0QKMTzB5PHTjZmyejOs6C78TH8s3sCoxM4lnPJ3DTWm/Mvk6bhEs
oKN/Em/90lWSIrj6awYI3wV0AS7qXgjfzP/hYc2MIqJpc3/IMgQJ/LXtvwyxKBi8Lm8tsXv5NAhr
4eKZkOlZK/3zfK7mg2bXSnIHZNtjmQS8yrDikAXvj4FLXLhwhlRSzj/9RzaAV8A1gbfp/Wyf1m+n
mWKnBskiYmb9Q3+dJHs6v+oFAJHR6I2/y3OfgkuNxG2O1MUfEiW91rBrJsDJbVI9oU4rp2Q9fqib
+M1G68gVNN2pXe1vBu0b+MS2o7OShBatOPBQKlPT7Of708B/7Jm9gXbED4u+l3qrWWpeTui/8lAz
QnWj5zTP2BDlMS0pQofMWdiKgKUaExL/OV0hK0ncgQYOPGlpiUsvzCoeJvzwDVUI97CY4baEzHoJ
q3qfiDLWJy2ydRsWHev10FGyVXwpe1jNGglfkXvOPYOwDSyploImc5fRggWfluKwpRbQzv3/fKfJ
pIXjCiOJAP7IPbvFvW5BlwvaJTsI3sheET/3uwGFg72n+sUvTk/IkgZePYOD5PJftqfiYWzszYk6
y3XgtQUgdyTQ3rYVCRMVCGaibOXrL/Fwg3xeNlC7KqG3vna9m4A2CqQ2yZBAgvu6F+LY6tE8OaaR
1VjOkHXRJigRm5mhGSEisPS6jm0HORrdjYc9dciP8yMzea+k4SC86xph5tWS5JIBA8sbhD2N274K
NDWGjq2mJfFDHh32IXOOlB4ktUvsdSL77OVxmb4yL6boONhlKezKIqzM5l2kZXH6unncJ5F8tlg8
MqwoM4vKeeUXGhvKP0Y9e9XOl/ssyRoONZYkMoQbyKxw3E9mjqjlvS4n2Yp+y+64SjYUrx0t3Jb0
MBlRlAhsRFdobCPQvFyaIY8oFlcQicQJuSigM8i7Nnad1HDgb3V/hAK2bEtsG3mkJ/becYcf7G2F
UFBv5Vl02Z419mPDgzJdyqrStipard0fpHL5Gbmq45ocDDTkHMKA1NlTZC6cJjIRAH7Rbym3s2xx
k8HJaj7cHSVtq883OOi068PsJHSjL6HFnLW7Z9ySAKfFCJalTEDQ+UrdtrcS7GSSYmxq5hzqjmKK
PqMlAUcL8/h7gF1JlE/z2wehQ1kq/0tDTUZgo24F56wryEUvZOFW+gGJaMuriur4aICQ/RCGx6Z0
fhxN+6mWr1yKAaQ74WGsTVEHxOJmKHElOqlB2HhWlTqMvzjefu06iwNXAkKYkyl9APsRLS9Yqm5k
fQoHPlUlzdB55KVS6duXt+2qXo2f2iOFviSFQRl3z96e69c+AgaXyYjv8BPYiLhiPQvIOa6+VFmm
0gM7jlW8Z760/7khFreB0lfpXnd/l5n5IUHlBTFZ7Up0g10efuD8KDuz1rNqVYXo8jUglOaS/10e
92C05fMg0V+yeV96fKBL7a8hwnXJGMONR5YonnNz3M9EEzY0qa2w32dCL8b9q97IIxgGgu/hpD+0
I8guswz46Dpm9bCLhfZep9M63s6kHbH5jvex0ZgaGukRBfmVhrQPpwBTRemODrjwo/R5a0eGkIdQ
sdWaEIPmnhERslk0KvVnL31ASc5A/tExyV0ZQJSoM31kZYVfq+K5bMuhqD4WYF7DueD+JfBHCb8g
ZhpgchjYsxBLUCUnS5/tlqU1ovnvOSLtX5x++i+ucr5KaB/NPoL79MZfTu+v5pnnQ7NdfjHp4uzh
fys41mfW0g0xQ5lC5YGhPSSwV6PfudkA2AxwsE9dwgI9Cq7vjgUSoVXc0jSxvHpNejca9gX+G451
JlJS0Xgco2fhnqIAz55gjPLShBbGd/9WVB03bSm7Nq3yPujKXXE2WQwxsYDGUG/flCTOFIoQ1cz6
bpBtbvr2cofdRVlRs0fustHE0qLKmvQVGMoFpm5p8+8NHPK5EMDI+0/IeBtuwRXVcJzoWUGabB4f
dSE57jslPPdZgywH8dRyth+ASKLdlhnAWPsQ7usEevZPFuMYKtcjbqzMOZ6VWDa5eKXJ34sQ2S6m
FTzfyQd3QoUk/38TIwY/jV4aDa3a08zSNym7uAPBTapxW7Wilr2xqzjubq2yx95e4LBPimp6878I
OGxzWhz6gVPz3tM3QcpAd1UD9AWUGsSa5xtfVv6hlM21j0+G8kCEloPZWXZ2Rvqef6QXy4U5gb46
prZO32XSxwKVXydSqZkjYLPYFKmQCJ8OU/9h/8y2bDxohW41CmcNKJfm5NXw0jJHrRwB48QPuhmO
jKpdGcLj98gQwczCzPpafTCR9zdtXRm+KEE8L5k/o2kST+DBKug0S+Kl+LvU5d2FtuEWXOrheiov
+N/g8CgfEdfyOHb9PRM3eAoXGwH7AIP8jw9SKSgJ5WZeb9bVSSZTrfHStEvL9PJp+GJ/Wp9n4zw1
p3YrwaG7hL4PWig3i4+QTucwfMhjyUJPF7GNaH2J+WM9+X51t7yjcXuqmTnlXhCTmxJ1polY/ovn
gYYG5+Poz6PuQQo2/4YMKNMIYLR+HgZBHIKsGHvHTHJ+N3Y6CPcCOIiFan08vBzoJxt1zJ+c7nMZ
aj1VdKAQ6UofmlQiTO5wwXpsmredDJBCeTq2LBUzspEnnuaZ+FW1TaLQkGMtScNh7ky8l390zXjT
scDUpI7eb51FHYc3RyWsNF3tbEhoAb2r096oOvoneFd8K5ot+ngY0saqvgZQjHws22ckuhjE+I/9
LoqUr1j0aWnNPDa6trJcfuk9rSoBhYaDJ3nnUXgzH7fdrRbwklk7zT78b6qfMpmiweLPEAhCIaup
gWW4haqwUpVc3n/iqpBk4/WHm+FOCaA5XOAVVGq4ufOmWlh9OCVZNUf5acldNlZhzugnQSM4NCI0
01DmNKd0m5QqbeyDCIjES3fq5j6784SLvQUy4BWoNQGX9wjtV0zoNhTgae3ShPpfweOlT0i/8qaV
16tLFyaX17nZxGPhI3C1MCj7ZF+02gHyI/owZO23XLqKDNMxks5JPqjh28EOPiuRlB99Bo2TezYJ
c/CUyQxPGiagmMBu4hBqmfsqlXUAmPrhc/4T54+FMVH4otKGiaayIp1rtAX3ueJ4oBpw4JV1c0KF
BvFGIAl4/7aWX0RNHKAw1XFCdOMTrhnc1qty9pWjw0jrg21w8gNmU3Vwb5kXAuWpVpXqYNt/Gtcc
K3ZhxSNvkoGRlmG4PdBxLygZye6KJD0GKDDhcBsnunBsSDlJ2r6Gf/Od7sxTLYOJbjUFlIDRIld+
puudwLXC3o1u+2I0deXQS+7jSDzQIO2VmdnaNJQ2x1f0RP+9y+riRfpO/0FSY50sRupjGVagZoof
9pLfK/tdj9U1ml1i5KGLKrfLak2R9NIEr9fXGV06dkd9m2hzPmnfkHWoYEoWbsNt5wGmIs4Q2yzY
mIHA1Ybd/dl1UkNZy5f1W5bhFCU3ekfS1UaCOF9iqJkacRY+N8IeektLhAi2uTdIpblnWgqXmUG5
I1aeQiZz2IbR/jtA7St2kkQv6yguuDTx+9txipT5MjDKVmboR8Txqkgqk8o88+bH3n183UTd/hFY
/Bm7n6CXBIkfqhKx2oZoYECVylGn1ijvhSB3XWC+55DcWHKrq6kej4Nya7hEbNECEbQ7lcfQ91FB
UG1b8mAHdsjMgfF0GpBNPH+iHsDyRN5kjtV8rntaud0UpBnw+eY75pfNNS93OQ+/J0Kp0Xz/EMtA
Lxnchu9JShAxfxZIeYKNbJB35wP9GAYkb0l73s1tCeYmTOk6cjlyej/o2PFNl2AAVkK6HJXvPUf5
2uHGnrs3dTiJAOnrK3VSAnNZXE8UqmckJz7/C8WrLZ9VnoSeXX+/K/ULdtxWqNTuAc6MuTOTxpcl
5glhvteqXVfmv9yvThunv+aLZu9Jwcau1m+ahmpVBci1AEZwp3rCfkuViZFzn/jdggvdwuT6NIl6
GVtYrmlLHsh7Lhxo/2Fw6h+bS6Nkza/8K/0PElkSnUomNXGAx2hcFqVZDjgccXqp1T2a3HE9vPHn
5n1xuN19BxDuVJuHg52C7me7/3i7vFP8Ew6SldOiWuvpes9MrpQXDstDV4halSoAuTOEpEnV9FOp
2tJAccBuTO6etEKb09lCw3/aYRB1nU3fMBkRxy1mPLMkcWJp8jlR2Wec3V/8S4Nw6Ux0xrqUKis8
ANqcLUT4FI4pZnmCK9ZfXHODZdkT7Ho0/nCcI4kc7t3ZV/8Q9pQmrAt71tpEUCxIFJsrIwwWSjem
x7Cqw4k62wIKILegKo0p7lSnkwJ6MHfhvI6xP+wv8pMQlzLbLpuQ0P0riZPLq14YPdxRmAMEhIbg
FekAgE+AGQLjRQ+3foUtg+G9FXj+0az5k8XNFRw6bwh6Y56jVfW5z42aiY9dGCcZGrabcRWJj8p9
O2oftdssIdKuIOM4pxd3FUece/ASQ9LSdGmbE23yECavNqWq3/kRmwo3wIqU2L9LThy/YhJh++jM
2titYYCn15L+NsGxB0pF1IyrQDhOZWVz+ZDQPlBMfvnTrziKRS826KpCd4dX4iKmn3RPhuY8/Iqt
8ig3aWCaYenWnMGjcGsJ6wAnIVgIQ7jf1aV/RyjcqY/oci4mKxwl7VObs9o8g+jHdULESIlgIGLN
h2Ts4jhEUyS0HfR8rOS1vibS8HfwXYLH68wRmK0kuuCHdq81iNIrYdE5a2nat9I02euyMTFShz8f
FXpO5JJ6Vcm4rdY9ELqnpMOAQnE4Jq4/C/KsIf+MYjEwfILcEkwucpxrVVLTPNBHyBZk9TxZ+8/9
FGWQjVtxy5QRS+KGiWBP9pp/1r0mQAeHQ6xtpWP1kT4PzbC48esVoCU2w/HrIscnS24vlMzSplCc
YJ5HAZFYrHQLLTAV9jFKu6aMUFPrwTbaTUGNcaq4fpJWzs2sf/gxmso5sQ9X9q9/biQkPlQNESOl
Cfxcdn+YqL7f6zQzUDUgRWuDCmjXrIj8o7WeTccTq1lf1yuW7ywh6fOB0MUHir84AEaF76vnLuya
ryRHvKApMJdj5WXF0LnJH5bsQ7Tt/+w9T5t3tKwtqacOgJlycySo3/P0WyV/h5WYP2gOsVQVacdN
J4GmQ/FVBB8/KZFeVOKYvHvedim32+UHAkzwMrxTeMfxBXMKcrvDr10FPKTpPWQaIm/OEMdJnbFu
4uOIQwOOK8WzctNwSm9vCGvlGHF+7cmBKP+xXD27102NwzU+lamfEUlQhd2PJnKGBMdngIHOHBwK
vsNV7nXOVOcFckT69+STsVMR4qasz7M9nAI03p1zUfAIMDVoFMgShhRkJaLWYWUGKd/kYO4Ov1LC
VwmiFZ25zBiFpUWf8tjZoTEUjd7wx2LhBkRg+SzasaXX5oKXDyefiW7Y9L28O/OBj+uW3P5ysFaS
iDkpeYdpw878p8jRMgdarQhDkHfmnyU8Q7q7KPuaa9wssYF44nWE1mgYMD3KPNdwF1Kp/J0H8972
9cO89ynxfYmnOosZwtO6RItqJ1ASZUl4ncuI/201NG5cCY5moGXE5zm9fNGdwJAoaYrVZBgC/IJq
FMNd+qbundXe0U+CAFgEIf1VGhb4Stf0Zh+Gto1gayai+hTpWIZkNEeNYaVa2Q5e2ZxfqieahiKc
rF6/DRWNWfQ1ZMRPwSsVFIYOuP9Xlvx6zhod5eRCWAppTPfrXAlu+Qr6gWBxVMhwhTafDUAd4rgG
oN3fIFRrTgm5cJRM9Vmc11czFOP0jpGJXwbJW6t6p2ffXBXMyqQ/n3JiO5zCwwSOBJ11v9y5xmih
0fWr3S9LUefGKTRo3dFVEtxT7KTKh6/Pj9RwARHjhMG0zx1BTZ5jZF36Tqzop1W2SygtONEHGaU3
4yrr/RYpSTqeySe0cFKU0KUMi/KTkqAv8A1ytnNAUS26SNufKzOw/d1wVcUvSE6qNgu0pDOq4Rm4
p8Cdw627C6Lj/djKgXogHAFb5VBMG9B0cMnrYeHqwPCg3gxoycDmD+YFhSo2vhGdSCVXZAzpNOno
P35G/UeKmOJtKtxg4kX15O2EHuC7sz9smq3X0J1fRg3srhct2ls78jUQ3nwmq+kdTAcGto0oFXZ4
vUlqnZLmog3jnXy44CMYaK6YN2vrrrv7/9tAM3DyWpcdFIgX6Al8AkgwH5Y0N4/HPPnfKp568t/E
GpPtuFF0WsxpQXuAE6ULg+8Y4RaZfzuLI3rHoZllZU4RA+9gwD0qNkCyeG3gQTT236cm3KDoEmtO
2FZdQ0/5fHjYrBMX9gAkFMRUnyQXOyCi3hIvGluKzyT2Jz3y63X7R2I4zCxfMkJLzLu6B+Ip370v
5+EtZBr7V1XVn4P6qs88CfnKW561VzaPy+VGoQUOWz8x/9MTJph2AcjcSoSdCkKHo3IEAg75iMmW
EoXAx+JMaT4bt1fjiF+AcXlwurRK7SbJnVsfptRCdqfc1GVlk8b93g1M52G0/aY9E6TZWN150VRf
MdOR8/QATIcCqqkrAV2+HZeszYwFgpbyBrGpUfp9psODHTJ1hLJJeRGBwHkqCZkMaEdD4Oj9Bh4W
gdK6NK8XKZKOUAoxdymRJmbts/TRMXU1OB9NKrF8ERG5ROWVG4Jr+9Gj9bUu+XfZWEYkrtdeFZmX
wcIIJDaDA6xO5Oc4MlVMENrT7T4DWMhzYsNrK0PSykYirQFeV8WBGDEgc2aWAxDpF1jltNHOGNKJ
I1qznwVT3pAVswpwi7XGnA551s5oYT7aViTd2k9gzq2QnqZrg/Ec+eJrn6Ae8VoJ/A4q5RL/MvdJ
PWIl1YhdHVK2HIo3ALEHMdrS0F8jIJ6/szUmua0D7KLSIHI+Eu9o0JxKTf+oB739XiM0RkpVpJIq
kEq3FNHJVOeYPuHLefHULPlYufBTuDaNamhHy9ggjFXSkQWyeKUssLwFkj2V8D+i8BBH7Hm2rk2K
vnEN6MrZe4tfCj+ecmDv6dgrtpIdLEUVvR29xSZxd4t2WXut/wlOaqZmsCpN4KyhPRooj/oDHCK+
DjJvjQJ4LQsbLT9IrazsF6VHPkAN9Mlq0/p2RGeXC1xF5JskI731aN1jbHQyN6jdesuW/d7jbik/
h+woYGcPhAcpwCUxSyJYRXmcvTc3aNOFcPKycQM7iIKjGWzKvznWAgfE25CsIQe6ALxpLyb37VJy
+06gbdVPiLnDVc9Eb1LRl3gEB8q494VndadEpN+NN0RDeRPXMyovOT3u74dBkLni/s36MgI0rrYc
XoMYRMgUE/nNShYZq5hQ8LndYPsqjuugUsNweLSbBCUOTZXFwa9IvqehrIkeDZ4aWVqdV3ZIay+C
uhW2vZxxSSPOX9Zw2pCCRwZ8oumB4Fl04SlZ3Dvfesita/zkCsze4zmz2xvdsPqYCvitR0rAN/A0
UAklehuG+7lg5gvDYVy8pYYf96pqv9TSxJeh2JNLUAoyIlx5F91zHvc4EsvfUkwS9AExDAO7rLDc
837IpZv0UoUcZ2k5sDbBvnu/JtHu8IGgfvqNaUrZyutogKV+xek29NXtWTIkVzhz3H+AYMR9jPEN
tUXQ4kiycMxQFac5J6dgKnQXHf4EQVc1NkZ3G9mVdf9nqj8P+Hgz73G4MFZvcDOtUbHL0/lwrIH7
D3WVqTJlD+XtMl64MPY6xeDjDQx5dqJy1VH04BsiXTE2vmKDpj4aC+h0C3V6vsEegBAX8jAJG0t/
NNrxnA1nruh2c3Csf0zyDUzDc+fAxnQ0kW5NRBfTD0MF9UOyw/LEycIlQdCnKLvaOasOyFooktaM
cLS8OOhhOiWCHiWO7ZOeoIFwfJWvUcpU5Z8SepzlTU/1V6PmZVbnUbsT9/fIZrUz+adKW+ferk/G
X4DNaS1xHA1QOiKsVHhQ+CrCJFO3pXh3DTyGfcqdhcmH/UW27GXurB+Fp64apq388sy11aNsmQOV
JQZKTlLdio6BC93fhV1av2pGaSxUt60gpKEe0etCx+Efa8qE9HuXCW5rjmgNf0TYcNazbf+4ENH/
MiPbK45jlws081gz23YucpXIxsepTvNtS/IYDj6vSKqv6yn1RBmh2Dz0zy4qBv3OQWnqW0RBAlpd
e3m53yXqAoxDSkk6FPeQGj2V5D/Nv/APJyUXG+CSIC8v+GdWdmpoPoGqvvq2xcebGwkz6u52U/Kp
Ey628sngBz58U/+Ob3uiyxoaErsNR+BGWL5zL03ovl73a/MEARqdr3JsnmmDBeWpU6H9FlBlgmAQ
YkvVDs0tExlZLUAXNOfX7/R+HsyHokCFr3Asf9Gf8SHb4Ol2hOlaZ9NupPtIFRgbIgGH/A1E3jt3
tP1jvLZnohAPFHZh3DyhRxMzZVKCrxpo4RcUcnMCRmSV8PBHiIITvRJFbNs65eMV5SUIHxdUVuhW
oISi78ne3uyChS2bjICXUof4UgYRstwTKeRvEevVXAj//2LHbNHMAVx2e9HhUYNHqAHmlmWGlBHo
F9Dj8LHvyt5AZo9iZAgSTjMob29fQ6yp4/wJhaKpRgizSVBlpupduPLQfiLsFOKReeO7Gpa7TQu0
X/0uAw9aLzo2xw+MgMVB4VpnY5DrBFHqywRoPYdS1mmyWc9sJF3Sekd8dv1lo1i8o8Cwqi3b2PJw
QI3msmRLI+v1UHIGKudLjp/JR//UNidb49ctCjNNR+V+fk5Kk0PseMLLdU2cAMjqOK8w10n9z4UZ
WuIpQbNMGd+eWsXkJju14a69/+1WJYBy7s5I/YvMlnMppo+gC0wIcX0GGz7+FFwEQxzpaUUimZht
Yseh2kUGRbpvzaMnLlF1tdRs/Lqur1TVb85GD4AxAjSg4o7cWSluZsA/C3ae/qbS7ojkIw2GdSfC
y+Ij87FU+s0fm60/tIrX7gSFcG2blWTmksLmzm0xvhsN5KtmfoI4iUrxWmjf8q+dYsg1E0CKuDK8
SR4fvTu1wPKTWrS0g3OMArbRQeBkNuoQhSeS9e6Gz/5XzRMlyj1yRSKbgk/4qqUQqDvKtEeUPbg0
BRS6CzyE9d6MUQ6URjHPx9xnmSuED8AafCAf831KJbka5tbm9cX6too2Czh2jPNP6AymXq9Jxyyd
f7wgP+NO6HcHtR+AbitsUv50ANTRhAmbkXFO5nQj1/XDiD40sJ6a/B9uYr3ykTTwbyhkNVsZBFpE
AGj7DWxk+0P9SDh1Iwazq0n7J4916KMVOB5NDnOxhPhIDnq8QQsEqI58jT2J4p7V24V0HeRkZTHr
D5n1Eo7EP/0GpalZgBS1EARAe8tPqJRv73gBTqp5CAOnrIHBbav2JcHyrhCs8ToCiD0W3a7goj/e
rdHCNZm3Tmjg73PRHtERbd88yzxazRdexTpOHLhKztk+Yq4oBQTAXQoAHVzD3vKZWIkD7YWFvWxp
z8ZaFuf27KYQGqDnRQHYG1x1E7dvHdrzCJqGU0iEiHj18ewpPCVoWndPPZjRnySMwTuwYRGhB4Xa
3xUmsfDHiFjn3reFrhdm6j9CJrFG1nvHNy08TIURrBjOInSWTI3vsg3VoqEvR8rvIO7Sw+8ENq+y
Mike15Nt1E6/SEAuWu6Evqe4cOOqjHRYS7Wnb0w3nJmmUFH0RC8g8Tp+X10r+klPwDo4aWa5PXwE
hyBz/fFfnHBj+Q/cfLTwJe4moz+e2E4dHdj/JIRzH2ANCDwJGVLlLVBvR4mIqLexalkdEvesqt6D
+8de19PVBd9l82TD0b/q93jhkQmzk2nWJLi3BS/0DjvvIuA7QFjp56qiDNBqJYxAcu1YRJeSJ/ap
8pAQQpeG6jePgIWLILdAzW6JUZmowLA/jKrgraayGk+ytdKMmencnJHiuQGTPPEbRA0NYSzjY4Y6
WLg8rW6z6l6I4/KSHaQ4sDOYpu0V/pchMOIDNc5cG31uKN1VxpYL7L7G+jRUypoc+wMDVuUkbH3Q
150LSwdP49XwD2XLAbrTGgaOA24lOMzC9S5rTNQ2jt+lm+nVcBLsuo3vOmZSTJlTSv+Hhi+gq677
2pmKkr/clEVfBbuJnQtbpLQ3VlcAECJT8BYg4eroeq6maBHLQG2FkyHqeQC6DaA2w0vfIZmS8v7U
giOEVgAgH2OjCOb5RGoppRe2UtNpekWUmUhNY+jdExpw3FmJXQiInxi3zKgqDSVPLpEufHEQICIQ
4Mc+yEHCzKeYGIzKM9XhMvqalChzJpdc2oL/4zaDvQALFVFowSjdlHQKgG+fPpKqdWtl1SayOaDH
5GS906N6q4a/qtuwfMBSwo8kQPGtqzaimWegR39vHSyh4vRP8RrdGc/dfcv/BIYD+odXPb1P7FhK
TEjD0jpxSzh4aWjWEbfsu5xlPfnU2E5XYwc4xSu1gCvaE7hv51fffJlK4TcrulPjHQAfBKGn/LAw
llizJ5nuXK50CkNhdJFxAvmdTYKpG3NWXmkwM0WWKiblj1O0ldF7T67YSFKVWoOZuUIzOPvo2WfJ
fRQkyK1oazGYmbGku9TglE9geQpA7Lu5tLe2067yFpzkQbonHacO1mv32b9E2jhvoGmy0je1s8DP
KqnuPnexwczPl4xBh4MJVn3b5I+txsH2tKTaIpiJdKPjNM8D5+n+9DKEqZrAYk/GU1FwEj5RZWD6
6+gQYuPlhguFAIsJNg15/BBzg1COCSC226FOQkku6wcWzLo2sU65K+uzVGWckeh9+YUqT+PT7fIC
4eqYShvSNoPzp29msw9FvUBQfjRjwzJgkABXk15Pn/Yrnuw0AO26FOIYUxksTujQ1bIjxjIAeBaK
rVKVysfJzCnRn1JGuCeNIzUX3CcThJ0ZtO321o5nPabuiorTXDCLjtcJjg8x1BkFtE5ziIL7yi2+
LQ/N8vwsI0uPGKdUUA5tEnpp9NAc1QfArvV+oALYhuE3fvOPt/NFy1/+1zoyyNBK8IhbqvLY27wo
TqMeWGG22iVyNgW0FJ9Vvm0gUItP0LNNjzhrDWnQes8LKjSwB16Hw0gPZUPiCNgf47LMrtwzenOe
BDozo3v3JhrcllTArxDJcGgob2RYn5KptciNQ/RMz7/LZCfdDAEGaZ31maN+0yDs/+V8aytwwiy1
5QYA4pbg2T2oduPxPBLPMojcpIPkzLBJdk5qgZ1RhUSFEe9Wq9bmY8EyoPHZBrsV97pGIhYUlzkD
Aw+N9x5hA5YifFlJs9+iNILrWNgg2YADr2YjTX4h7DvoqCwHPNqCR7EEIXV2Do8L71TPRCx+P38Y
/ZX/EFhG+ITw6mvZVev/Ka+FMWoYUKfs9xFX4S2yuElNeYO740Np5SIStKuUO1bqwaWDtrMPsZe3
TsWUFxfyfrpgfb+dQVkXhvJr/kwsnYVxpwmB8kFvrXNOvlxHff6R1Z1B7BBxixAqgCAqdUdZGPGS
DP7GnRYbS9f0wX3CPfslwUqv8Iku1gHk2kaO0C321yJDMY7ayXOGoIPyBsEbUyLx6M/CM7abMkFl
jG3b8QnKpFHaxynMxHX29HA8ErvqrpXSXn3PK0gWfY//xJDMDpITfZzNGz790Wjlkh7BBgweo/DG
0epwTXw17ZgvkVEeH2RMpp3rtXNRp25T6EEUAccoKroZtV80EpwE1Ww2umMMmowOo0MlXXADAQMM
iolzFbkswchby2mEcJTGUFNpLxhPazV/07X0KRFmWCFcGt4VVLfA43FLJWROXGO5TRaJL1IxzKpk
ghE+E+6V2LQ9LHB9w2dWW+SPdDl+k2phd3kZlNsFtKy352Dl4ivoPrzZcGspC4swJn5xt0whpHif
T5Sg8iJlRwjzVTJcc9P45gODv0vbJd38lRFLUiGXBb4qShr+IJPCOalp4dRbVHRMQIW68MklypjS
q1pNLKDvAoqnNk5U+vfsNEE7B9D83+7G/GSe+0GpKRD9B7OjCVDdCNBlkZ6JbePSa3qKjcPt+rOL
nBZSbt8HIrG2fBEYo3C2nXefTbUlfsx/ThabVO8HoSrb/HZpSiR+OslNss+Wo03Uawm+41OCxMog
k6MAwmIh/9SjWQvUzWjcqy9ptktRJqQD/LDKKPznABKkOqfFXaeBRrm0q8xShma2r8EIjTgwR563
HEiNQxyjJL6PWG2DQgcGGNmRKXPb2NAuFLHUPQBZKtdk6Exx4H4cb8gLtGxGoV6ogGPddL1oT/e5
GFwM7L/CuYcQmqagehzYgXXIFr4/XNfDfGOHuVIeEzkxz0eIW0s3rVtLtjDxdkBMgwqV9NWnYEc6
a4mMfgtSrOlXsYJRQ/hTfUicWluAOOtpFuVDqAxTQVY6EMnp2LakZl5srt2mVsmWmFIUF8z36IUj
IuwN6IAI6I4hyh/NlWT2hQAR9H/jO3vSTg0POz/d70SR1w+IDA3Rzfdj9UZ2Wtj/EoWK58XeNTan
X9m/hMVC9istzQaJPlOrAWdcGE0zZPQcPPQSnlB6IpDBrrIbMcjsk7SEGNTuwzq45tXzPvv+WYjH
ljKnYbEJz7jRznIma+fBjC0xoKc9BHYawVcXmshYwnbx/xyDeztEP3DDwQOXhdKLQXOY8UXruCO/
/qM2LbSUQ5MsqpMP3trg2CGWMphNoIyjBgOAUvTqRD4ZbFOzDC3tjJV1AHqtXeMbcxq64dd+qLQf
E/L1VbzZk6meqjO1mercPn3ITZWuV2mExEimpwUzx5+z/eaU59R+Z/jfU9+qP/FZr4RV6HOTsR+n
Dns34BzQaxW7mf5Ypykcj1VS/Jpmp+7wjjS2hKIE5/rJSjgD8wjpD08QiARKCoSwKgX/iWoqM08n
aTKZ6k9FMDx7ygh7fZ5yi+29bteatUa2MX6rDORoe55FKZFqTOaLnWJ0udnwiUqbn1lqKXpGVQ1V
OB/whJjM2Oe6+xZWyhYvItNOnKxMOh5GigAeGUY1UYsS5bz0OjynRlQcaQ9whBt3yWy6yvpaPX1A
v2gToFQbCK+AREsuiHj5ZNWUDxLdJlB5PfJEA2IvuOfh7oRo+v2USJFpmTYxhJ1BB1y3emqi3taI
j9JZmJC+zhr6lU24gyrbKMeConEnmIkYMgcV8lsC9bdo/S9wR6kWZntY9NpzbPCUyPGX5L3ayAk2
BPU6WI7LYrYCTIP5tiqYuglPM0E1yrkFMZiJqWFVdg51FDsEsNX5IxJoShrRBApocMRsLZJT2L7D
4FKrZf1Qs3tH5/tcinmXJdaWMqf5YBpqF5j386n/NgNAtuFb+s8zWbEZeT5Pf6aOOW7W8s+lb62g
7TVaj0GsGMjUZSE+nfwI0uWNsrWZ5tRH702tW4DewJ1LSNK+UDVYDIZPKQgaiqotD7ir5tpdwVg/
DOGCjKyQeAp8z8ieV0xbweJ0eYdXXHVky4xUxfsGnjZOAnvyp5xI20lY3c9M1lyxT/lz5pxfk6kj
FfXQARnZ+B3MWQTpCH/Ffwq9wLf4M4eAv1URxFH9QrLTg0hYlzqNVk/yvt8drn1OGQnVZuN8H7D3
UQrIwNn2rGg4bTrf58HGN7f4jB4jtdO+ub/s5qQHZM7UouJdMWpSFT3dgrQt8+Ne3SxuRi2M9Gye
D9K7r5psHxrEVazA3KTX6A0LEWxRsoO5EPHBgakH5cXdahiFbr3/Soqc82IxGgxHo2ynSNFVZZTZ
GuEdkM65nV1PZpWD1oJd+JRCO9uRcFAzSWlZgVfX4kIHTv9lp7Sm0Hdlws35Rrq4XtekehZvPwxP
HUIYVuIcri5Hp2T5xoCfE2c9zxS7JFxSL5Si9w/Fd/tdKJZ+tBNi3QGnf9GYxV+yHrBlIa1NQkFT
gq+WrOH2BlszE3XlDW4IiSMOWe9wzCDtPMMZ0MmXDytHmHUN3II8qtC/ThkpGWlPM0RFEfmM81tz
njdkycEeh87T+zraFqW7ZqnktQgFjlcnTB8kyrbN8ivRzxaqJ2gEh7Tc4FDfBFSCHQnHN9xBAQis
nG4RZf9RCj3cHay2fyrv+SeItNxLxs8vHRncjrGs5IBxCAs0BJKmsClqpYiaj8gg4Kx1noSxDx0k
GASnXA2+Awi10ARA4d0FIMK5T5Cz99G2rd2pnyleURF8AKQvtBRldzvlaY8WBoHWAwg7Hr0+lQ6s
NOXjA50K0ExkTrAVGwxlaeJA3LzhPRwEW+tAzHseA9V4cTVA2VBzMMgH6L5DIodKNjhx52CnPUPy
WPkFbPCPmoKR+ctE5GwJ+EtKe1fIZCbOQDN+vBkbEPQjyvAU20KZAL52zrwC5JWd60vBsAqTl5Ga
R809IpEy2POtNDdDpNW7Vx4QPoym+rla1a5z9HA+eTKKMkDB5Xq6CVNY8cpOqaH4rd2Wp6Cfejyd
c+7vg3u+y6zOeCIh0cAOGAcsyaysn8WJabZ73RSxITLKImBg3ZvF2o7tAZ81t2UiGk3dKrZmy0Sj
+Q6+Qhi+FApjXWFl96aEpnMU6PHyC84BTutIN2SQ9TM02Vf/EDdLExqpn+ItS2huYHmJQvI2zmHt
aAW8NgFSgUJh8LRbDNqjBWvVnWqULntnl2AeO2yn/7XLQ4E9aUI89/XkZi0xCoREYkBqpk9esVe8
erBnPKLE7s0AvQLEG480xPOm6+pyAc1Vrona91FMGJMu/wD0o/bKWkj2bMcL/WzzDZJYbI16LnCn
wqOEUrNAPGkdsGCBbWvXjQYp6EE/FGT2TvWcyDeSDp5zjgkoTSr9pXkKppV4p+NjsQSRdwYEa2+F
5Mh027hDG8BlhVc+3T1ycBGs6/clBVSq7uyzMOz3bwkPdznXMhGvDNYPkjrbftx8RsuPpDAV+tFz
N55nJdfh+HFZPZFF3MW6xZP+6+2svIcs2oub9YK/UBUyx8ND9vIpuSM1kgAgYrc4fAJbidZYQE3w
sWFaGxGL7gieMfz+4QT5UYhO5L/5eE8aw1MFE+B7M7shxNYYeiE7+7DxbT92rVYaqH+v6vby9oFl
j0aTK17CXeYTEizQw/A34On1uNHgtyHAefEwibGIZGB4sS7BwnHFQKMo5b4kBvkCce6TqefnWZ9i
/WZWfx9uZpMGLAxh4XMCW+zzLYU79ggrTY38yDBfnB/72SoGll3j5Q8YbUYyhL0/NbfwR1eJvfTy
MEBAAoA7yvTo1kpCvN2ayy4HrG0krCnx++yH42+7W7/9R+qOGkSH9+jpWMoNlw9GZTZ982ipZMQV
SxSooWFiDJPofRK1yD8aX6+BgVWbpLnehQsS29ulOrXGxJny0hfLeatjJpr/gN4NG3cBT70gtd26
9rpZAUfe5WoYoGg34yLFu2gVWTWH3KCFqhVBVR/FOYgFhJYcOnTCaQbxO/TkaosJLo4aQ8ghnj3g
BKk11Pxc6fFku8dZjNegcJsVY4wO/pWYq2us0VRpYjPoQAN3wazTQGafQTHe/Vi7nRWZbAYpMSjo
+Cp2GWVv+cSHL/qX5UZWOan2LTMHHPufrwIt/iLVgZCP7Flq+UPDR1FJWEex81cV+3SDYQKA7Le2
9hFjBywY9zQDzP+MAGwMOaxmn9517d2iPtnMWVRT+h8OnEa+p4bp30fNz/OC/PgKTQP/x+FO5RUm
qCdy60aE/X6A4d0+mA5ETIL8ciGeogMUAr1Tp7eDJ7q1HwwH3ihlFrWv662oP2aELY3oMU7pMt41
PfpeIqTO3dk9GvJY6Vd7/eTxNEWVfn5HUmoEQN6dw0Yr2CWuk6Pkzx7esIVF/+GyavooaZkuDvCm
PwddgUTP2MdSBgVmPdxsgiVZ9d9PrE/0QKM8vzg6jchdBWfFs7OC3oI/1KI+fRJ2m+kMJ1J83Fmo
1oGQNXdeiiBiOpTQHL9U/xMPrCJBoOgeqT+xycuyNqZvpGEkNgRREPNIhu0JHkVjurzpW8W+GPoz
ehsA0hYBaEGl+RPYm9yzUZHCHRY9UwIrQ7/R4VUiFRZ3i2Fwp1XQ6iqBZy/40VtMJRbVN8qU8fVc
RQVhJfLL0FG34tguTzpJOw62SDS9K+kLO07lhMWvQ5bVHE+3ZuxlbLiOwfO/TcTMySSYdLjAxnvb
jVoxG8LPX7Kd83NVXQk9JyE4HDdDmFJxpYWdVLcJnSg6OSxQJAEr4O5eUfueRWKNVg6M/gazip81
mPACdg9I+driWimv8kPjUfBaylVQTqMBO3GOP7JBeY8E3v0FbseCWazkgA3s8O9j25Dy6Hw+dMTj
nckf8Vf5g9V+oD38Lnex5iB/xVz7QlLU90YAgO3fjQsQ1/rPd5GZ/rzFsQbqsh4BoFE9h71vPiJf
DUs7F/YJu0ulGWN/dRzDbr40+l4FAUePb8GwN6lzw7pT/qcKfkq2P6FHu47azuVVRsglgDYDdZ6g
9B5JalgtYvGn/Cvsgaln/j805B5iVWIIeT7O+94ZTw8Y7xPEw7Nm55OJ62wzqxepc7sTuKNYEF1L
aD6cJtnpfI3WE4AJM5G5VIg7znusuGmXjPcYwOH0r6GbmRkP/VWI6IfFEnlnD6LDHlu8jyvOPbWX
N93vt/Wy6bJO51Zm+WzX/LbK4B3fbmdzIso1z0xzB+GvDl8jcjkPzwCihddPF7cr3uMukYNXMWPH
9gjNTkjbVFN6oebIiusE/s1sbOnafmXOcvYSEkbzsqL8YR3lPNL6dQZ0tZ0QJKGOdVwCPhr2DhdM
9FwqKASTLEmMMA/UwmedznP96aMt0uhv1UuKWH2FqAFDqKm6ne/RTBQH39uv4J8V2P3GdT4ISKl7
+fKnx/VNzpxiSJuFS8g539NaCTvXjZBSVWspFhFxqCcifqcMUgCtzRm2VC3L0pgQIrUNlT61hDm8
JdxDFcL0VQrvbMJwFo909MeNEvvof6E1FwMIVIWX5MZWdQP0hgvrQIhwQ0VVQ8jBnk9St0hIG2VT
8zk+zSaR17n8mLfpWZ/tJYOLY6i932kHYGdYPdJly7ZIpUwiMe4gbubyMa5ErnLxPlB9p6bCVJWE
WdtGrbTzFK9/v/4MRz6KrnFrZ4Xqhj4f2LsnVTJHcf4pwlwkC5XW3BMDj6uyJ1FBNvyrdHWMZN73
rXDbtfutcDSORYTkCajnWe9DLVGZu62qNcuo5Be04Y5D/hPrbpzAtaAagtSh66x+UbVZ6tqgjOt1
4NQTgyAFciU59H195AlhMAbuWKybETeQ2/sjc5SeSIKuzhSQ2Wy+6gn8j150msNNxHcVWcp5wqgs
za8QrNgvmfnyhXor24AElO+8+SfYPAfzpRO+iu0is6U8BbR8c0fGB82Gtg9gfzJpNzDJVX4nJyxN
jecQMvySlAKsNrz5P2DwPTegeXs+KB7LF/bm4260wUjSCSMf+OH3wH8pM8vX87YJe0BZ43t4go0s
PDegGIMH1Aad38mYmgjYBCTMqXmr2XkDoxtVl6T3DYFG7ZA1B5UEF7fPhkcip7UlW4KvMfTiRHbV
JiAxUuhYEBqSI+ONByFPIW2WnpGFm7shydzBrfovjbBKCdaj3uMkNh4onXsN6ZpDkWFgQ4KH7rkb
/eNaTC5kHLtjvmzcjVv9HIzQIRxzbK2fRj3FLPK4Gkm1v/Pxcf0qBlWzMwu7zMhTNcVk0Xxe4rQw
/+xmobyqHoirTwhRvnSHOveP4yQa487rrx9unJpvhELbPNasRW++yDxX+p/Ww2mcEHzW0zWN5/fb
0uf0yCcvPr7layuqcCugoCI7fmhLMXGJZUqnKXod+0wDw8PDWgqRfKKQHvIH/3MpLqfv9YdkgdRM
R/OOwtSIgtln4nbYm1oKwMFR25IuYtxzquS9k8rtvXSC8nnF2HL1AfgZHUrMvtInLwf4Yolspr/k
SBojPjGbb5zixAoIUgfEZjBJfN3mBK7cWLSnRymQ3FkpnVA60LfbhbAYoDUzoyJ6vg1ZhJ/FbjLj
ErkX0BTbX+7aMEGU7rNOI574p0xujIyAxWLifgB3j8oNIb7OTbSu7gEKiAn8wVOi21uEpgxtTtMV
EJeTfANI5ynUCx6t8OQP6l6f997NzpBCX3/z2bY0CWzOKLzicL2f3VBa8AlFJtpXMmXKC/G/1Qkr
fkKN5gpb8PCnB9B5inymv2WdQ2L4FAKmsxi6neEN7E3h8Z6h3kX7IvLgqMGFlSMPWr01OvcPywyy
Ul9sdWBYOaYuYHlQKjD+JxVcd6C55IwjzauUi1d6rC/iR5wqf/4K+7bflr4a8+4xxiEUD2Z10q3o
9qVabz6Q0K1/HYrkzr3JJy30QszpSq8UIVpPFT5FTVnzvg0rUSmEpMjDA8moCnDj5OmIV2sr+Rna
+Wa4uWkF5TiMYPVVpmRUnmW57vjI3ocMdMi0g025hsItJ1Qmpy4G6qayUw6ZaEd6E9Ck5v0t7XT/
dGFYWYmLawnrR5L9JcPrvpguE1yNBLh5hO5GjTKlG79HA9VeOPPq0yYxABZ6e9jXcUNlTbzcl3j0
eqq7w4dJy9xqLbzkMFtT7LsW/k5ZFpHCiQRx4+iOhiQx1jmLH8ijbCvH4ANr9viCkles4XvwVZCH
2zNkUfeIS8nuyEzq8/1QyuqueL9yUv6agxPx1vxPGGv3Dm9EV56va76dgwNk9UAz72ordvCJDF89
7WBfTjqfcHo/1LqGTmwjnEfJzoonTrVnUsCn0BlEziv25Ek6xfydiBAhoBrNMJKo4dhyikNoGNGv
AHblKKEI1itsrQCo6XH04iCoFpcJzFNsOe6tjqG7NELLgvOJAABCNKXW/JE/zwX8P44q1jxoNF0p
MITcFzPHMwz1YGsNPa+CbbkPPME2zxH1Zhg8gvGSTj6EJsC1AJXST5rx/7k35ZT9FdqV4qGT+cBm
H6FtsozCBcX/lt0DtE3uqEtFlJz7Ndg4fDsNskE18LYWbDMcIxUbfcKhNSwGMxLF8pJ49AbfJp9f
x9wEEqV31i4B3BkrXXyMtGMmvgsu4KHhJSMAGpvjvr3H87BHFNR02nftT2MolhQVCZOwwv4EUMRs
6mVQpyxcPtQrq4lhIj/Lqvug8sCrENH0zb+N+abXi3dD5swlgh9dnqcEMWvf1krbanYECq5MXOpT
ERFnSRgj1uQY0Y+rWs2jBJTJHCxA/7mXZueqFnCt9ZuDUV0MyK/kQBGihXs/4016j1PvCjrXXGKS
ZWMIWpXqsxQlK9QRhlIX801okgAdnFh5OIzKggdhicV0ix3r68eBf/cdFs4DqFNtBEks1qIYT/AO
pgS/yhX5Q948ZQxu80FjZeG1+C+tjJAI0QWJwa30p0x/CZW6ZmsrUTeu8EDG0aS3ir4Ma2eSKYEl
cRVn4eejiHxVbSi/qaZxj0zYheWDl18DnP7X4seaI+lHpO2XNqMwPYt+T3KNkbUOmgidYNBsAKYL
1PJjnEIsLZnHLO3pQFGT1Z4iH98VjWvhsZClhYVn4/QvybsleG7IbEBO1tTJckOS6uciERITyD4p
BkL/N5LUvi7ZwF1OMPp+JaPWXL6iQaEfT/VFxk09e6xFaeL9VCmRRzAjEfuvP/Y/LujzpM27k/nt
uq8bUjV17SIoK0RUXJvKYOWM8L1sF/CuS2HXJppSn/sy/TjIaUy16eWN+kDel4jxl5wHQYFphY8p
hcmwHxx4Fw3JpQm2KV8n3qekiEOEmic6EzzXGjfKaKtdUckVsuq9xAUr3pnOmX8J9xPvGmP7LZq7
BpV0lISojR00WIOwcwqGIN1smT0fKheGFezWcg6vXngOFGqlvNvkE2mCqYQIiJjUarhatlYMZ4tL
g9rl8jrGBRUhSdW1zAeYvAcwqi99Aap8Tr7yrk1GYWVYpwIlFdR/fGk/PzLOBnKgOuHzgPtYEJd4
aFZAzo4FBb67r/R8NLJAydJY5aJN8fmyzPbMpNRFTff5mQqFsW5tY0EFxtu3+Gv40KSNBjJRTGLi
ZyLB81izt8UfbcJ/kYsM11PbfmGbbJQG5UW2nKq3oh7lLau5AQTT0hTC6KQwPgoH9/IWLV6O3RSr
MrgioJ6OnKsO8+xiKa5GWDKP4wSxFXM3ZtZosBfOQ5DiCygSytlz7f3Yxt2poKlH632sr9FEKctw
kvcQTF8ltdYB7PtbhD9/3a6XavGIxxzRmrKKeB6NFp+OKo75Q5IPY2xCLOlj8UkhISJJs9SkG/QN
zKhb1PtwdB5CnKVBvBOiKr6P3d7jlMxypSRGdWvNVCPKExGkqPKoB+qf1Qtvxw8A4J5MVufnP54/
g+1mqh9tB6Ayl+Co4oJ87NUmz2zKjNnbGhgISt/9hd8jeXGbSGuB5UvHQnKI8BCz8yOvE0dMehmX
ZJGg9CTtFB2CvJ/3Oa7Wwl9T9qeUCr/0hFUSh14kVJoeS1g0Z/FWH+u68Xtk7bjvJLtvvjH8RhPU
F9QIwafhqv2cdreZ4ZmtfTIp44NQWDhCJ0ZFoPGo30/rydUN9d7P2GeSNLy6xAuucboe/Zl7llQT
iULtS61E968nKwMt+CZzBeK3PRW/8WzVakw3N+jdzWbGUS2HLMHV5tty1N+kJeFo+uoSiS8Riexs
v+pJ6L4/zW47DK6BK9NUZyLovl1bZO0+MIZDA0MNZ9SEd8zKOeRfVSLVT43aebo4qeAb+vFNQaQP
sVRaLppX5KaS1vZ2+/34gLVENnKj3QgWhidsoxvni66cuSZziglNhXntBYMC9PxketW2xae7vjCD
YhCMiKaUTxVq7ObS+laS2hvflQg/EsBThxhLUGHt1u4qthOhXB+6Es47jU6g54UYGtZS6Et5GY1Y
+1GsdCm5hprYdmeQDvfXJgJV947IOCUsjQg8pKoWVqiWgPm458vGLq76N4rOFq3L8yzzfprx6TX3
6uxLAEvR6f8YfSBHs7shZcfjaZc/cI8hmhaJvHf+nfDV7u68GSsTDsckVE/G0PM0AwPGEEYAoH4d
iTYrcLPamyIt6yu1ImNJRBnXKxM8zSSYkDo/f94AOjnrTPRrYuH3thbuqxO4LUg9xOetfVNAg0MX
5HyqwZxuEFAJKlno5gi2l0kFChlqp8nj74fbuDO5O+IgxsbJvjOMtcDIYRHIqhN9B0UzXdt7Govq
UnK+k0KeYU6p6D/5u9zWAWv9DXxBRvQQChvX9rY40U3/zlJO5pCBeTnLLGWsnztWRg4HPR1KYpTY
ssrUWZDwD0TPNL4vzdCmd5hkYNlf+vzoxBD9S3HxOyjmsqYQtM6RON2Ko6VlTJfo8IFHHziouN8N
9x+FiTxankk0Qe2sldru6NE0egctaLAl8C5Pv3cxqMNVSfaFNHNhP9xkzWT3zoYJukHnv5doL6Fa
Xa4tUTGYz8peplfQhbhiruM5sStC615n335bp0J6vcImCQvxFxRqBqoeehKCCcsoP+Jcn57N22bw
0rxWWzIO8mFxXfcMxzMJ/rzmVEH8OOlzWNREAjPzaWoWU6PS2Tn+5GDb0Zh03c2XuM4rdawfSmP4
dOB7whh7ZxmdkM77+VrUSCb5mh8jyu39VPaY3R44GhxYYFZEpT9okRIUkIL9xZfzaM2bCh0u8gHt
aB1qUmeVJkyhwGD5QL2xA+bV/Oo5IAwusV30pQ1fey7SNh86nUYlsBUKEhwPM+/q3w1LSHC8nMpq
2t+y6M97CsnGq06aMHyk/dIZ/oiIoM4OX6oEKRPrEBC42mcznwL3yYuNZzhNmr/M04c2bJb2rNRx
ovjAN3jeH5OvFZKcm6oKM+FtWd6Wi8ZmV5LIBSj8WjYswgg6sYjezG++kCLIB/v8fWnD5E1GHIub
M4QGp+FJVFr2PWv1fG5wcfAWTzBP5VoDBwkDvOu4FKQgNZe/qkzderDsxEyR8WA1g2nXsuW+Hp3S
an3PHNnMlKMsN8q26O7wAeIIUd0dmJtdQcr6TLp1KwKPXiKhgWKUEVpLawbBjhA7+ypqqBA7qAjT
TyiqGUU/xnM2sswTs80ZvyLkmuS4IMk538EjJy/ooK9/F2vCAn/vx+LmT0ya9YqroXAV0wJvmEtf
qwTaTlYdHSpu8RgIsvw5iTBb68WUJUJMY4EySF1EfqyS+KKuaWO6ZlsyeX4hE2cxlV7JIELtQLgd
oaGg2JGtHy/k6VEod2qAWqARPFXlpTZcLIjlAAr4ubapytXVBCcB4ZpxBvvU+X00NhqhWUY0dXQW
6vhtn+5C5JGRF5SBaNo/kSaGLfu873KvOhK/4W2CMdQ36leLO7CxUDqpdwMC0xj0jv/szYaocWhS
7py4nELLmrvYa55ajCZuJY32qain4MxJIIo1PbXAGUSTeLhSI58wJi9uqPReiIBcSAVtXQUAKZAq
g9znEveBI74T0mo1B4WkdFqeNjKnVkkyqNByh+ZzWSj8lHjqQKwTM6WK9r306mLpTdHg9X+/Ij4q
YSqCr4WEg0JPTPXTXKeiYdiTSkfH+aBVz7uQ04kmZUV/D8Fw4TQ3HQnvsZjIvKGs2uYNxZNph1Oa
xCUKmMLPMzQ5AseYGQez9AndQx8QQp2kEhhI2vA4Ep8jtQEs/orjNk5dwEx001+9U8f5vzpKsRdD
6k5Vbrb4uGk92+8F2Ivt/pbC4HpHsBxiPzjSKAvrfQoRhigJMNR5sxkAiyBtQW/JZ3FAZtGRi/RH
o/wBJKV8mM229WDvAENZTvRgeD+44LbY6miFE2CmLt7vJD8NTsLg9hxK4lWRXQYr81+tSkmllhKO
Y38HiZ4/WK49UzwKx2j8OQgxM77tPSRKyCyyWVxHgqwa7LwO4laZOGtDOTYiDeZmjU3jobkrnA8z
HY5POJcbDNh7asYOZWBYfTpTol6KcbmfdcWnhS/R2qnvyJ6rZnUG10zDZXhfq/q7qRaZ000s8/SZ
+fZexw+1wOMKcHQG5Q7equIaxQgtFBcfrtzKZOX03UYGwCxXY4rvguM/yXb1D+q28xE5vmRbEI8h
ggiRaDdRTGG+BjM07MgXPehoJKlHkmMX7h5/0tFAR0Tts6GJHmljc6nkjxcWSthm02DwoNSjsFsd
WgBkiXHUpSSvSs9eHGJ3Ip4c/XyLhO4+IoAaG5SZnmG+QKG6RMsBOfTZeH3Uw/0NRlr0r3jGt0By
DtbIG6ujKXaV6CqGJp1seR+52yVgaoeM3kTEPl+9C+FRcMB4P6Pc78BWtoSHp+2v/DSeJ3JpxbvP
4Y9CS8wa770r0gDHn+avgwPB6NxI0vBEBILTBH7RQRSNtkEYXUBcHtm1TmgBxXwFiQoIlAn+lCuj
waoHZgMjutntHaALL/ImNUCQYwIpIQ3U13wXNDj9rQEn2RQvWcgqAMcO2qUoU3i1VMqmfR7d+w45
7zh5lC1kwU59y0fSxjMQzwQGXU8OZYg0aY1dinAo/00h8Li7ChdrHD6B2hwmcFrIJNQ72ViPOknJ
l/uyKgM3FABtZMUTzJazPVuS6zEgpi+/xbUq+XfdMlKIyKLCZ+LIQH8DIfpFsp3WKklodl701xYj
HLZIjRhFthnkIXYWvXV/YEgzFV/hSBVe8xIpeBeEfT86UZX+OR+QiTlrButy8P0VozCA/mEuYZu/
3lYugCQT7gv53IyfxZIXJVl18QyvqrWcmf1Q89bpxiThqR2fhdxwmalXoWtkifiTF1TjCq0GbWiK
giXLxp+aPhOl5Urbsi0TPGFgSKA6gQkoo5xcqz8xhvzj2k+nNZ+ejnrYZU6Wjeg098UpWhgbrRrp
gQOcFwFVuoL6McXpuYF6w7lguHdOvSnjXda0oAa0aoC71TOEoguMW/rPre1Ixewz2a1L9XAD7q1j
5DMWV0PsDbRlHlMZNfOwqcGAMdrbH+jhc9ZUb9Lw7fvi1b9xbiILm4cSEJhZhL0rLSIZ/Y0CmYQe
f+QQK/zpnROyRSaQc258/sburoMPLJGYRTapJDFX5CvDuK1vJ0MHtXD+fJJYlGSAylhgyROo8Iiy
F93X8Bfx3pkKD76qgpDDMgqSlkZsL485ZhkIg62D9y83A91sKdu+DvaGIU564cyBjnyH5Ej6Bk2k
jEw0GUu+KOyy+K++f+BjTODSzr3Pq+4iSlc/smn2ChIuq8DufcAODfNbZBOrX+3AQqIunHYA0Zco
z07C7THXll8xsytmDyRKpdnraINCI91aTnyGH/dHDy2l/paPRUIq/nicEV1DqtsY1N34a+9bcJAY
+5a7ZprxHrOdUKwcHKPaTvuF/WsV+jM2WqTs9cVdBJHv1N/drG6JSqci9SHkkFEXx5dJqXthfTcA
7WjNZXac2uRIkgm5FYICXXb2z2m5M7g8Y6f7SPM7XqHpicfK0OOOGv7x3mhbH5GadXuEVTdhaEWK
PeCkdJW5Ww8EZZ3lascsG0fVKxI75Fxa30PM+YkMbTCjW7AXxrDiaH1MEcE8CQY7922LHpmPdcsf
3tuzjbLqPv0Od9/iK++ehtRB6S+DAOyI8cudkV1jragYHES2kefoDe4p/qHmSa1SWw+Sp9vsWwVI
c6n2r9t+oa5zsOISnMxsOACNMOOF16j+XSoNN8Ga93hrhi4fY3IZpTB2NInA8GX6U18KDLmuWULi
EDSIm000RooZAALrrjRn4vmrWY8RSjpqeNz4OEF7PF356DXLtQMqvT2Q+TlgduHOeBWDIS911STK
hQuGPh9KWJiZAS6OW6X/Oy5CvhGtB0NpPogoEhovTd1eibPMl9qN4vjz+mvmJrUOfZ1afTQgMFt+
xJskzRyHGCDeZPX09SVqq9PN2/wDZKYaXzeX9vdJMCwuvqhSgAX7hoSjQTavBSfD37qkumoiDKCZ
OQei7FiroP7FaCLnO/sLZZJGVWVdby0+SGxECjQfVi3g9otikuuURK0rH3gigOJWAE6SLw8QGhWl
9ZneDqi00ScmYRa8epJRZHYpHYzEoY9EwffPq8WEpmSGwDIuKpUPyvOzciGg3P+bavkT0Bnocexe
bovU6W/7h7RrFg6EQtXysrdFA3tOIRzomm6evaQo3PUArmc1KK1pfS3mNjyywXxPMEWwQPSmkVpY
F8R8puJdsCm+ICODnxuAhrbKC6IQ/9gy9JB2Qq36Q/7AWf32gIRrvTveqSNUXO/MWGA+9T/HQOo7
3tTQcq9vcz+7R5+kYJAzj0RJntlmrmbNJdpa4Kd0n/L7H3TjDPl+C7YUZD3bNs5H1qG27GL7e9CT
a5LnYII66OqvYUCULplqinnxptEr5eMSFNfopkFmVJeYPAkqLb4crw5/nnP9dOlXEMlTQpATbmYe
r90nCfeajvyhuLuZ0UiYmPiuQ9tCjl81i0nXFEuV5DYAOYXQ26mpTWtqgsKIEhVqXFHQ5EOEA6Rl
Zio6a4kJEOo8McH5EiL50HzTeHGTBjcONLtk/NSv5SnK35RbixiQLcIHmakWcZ/bJPyp535n5OKw
EhbiSLt8XUs7NO4uemEF2ckoGLfSbbUJg+GruHIZ2/TycGybeILGnQTHTKvsc+wDEneHRve1Cod7
BV7HdHRGb30quP0GcO6fy8Jk7/+++ByTOiztEmt5DSB7xc58E+P4tfgm2mo0y8ugX6SbDYj0vQIW
7OQTfkhkrelehvaxO1uUcroKGApqVXa6uXgf+wOsmo4rA2DzISRUK5yTLwtgGuK9znepj/yFk2xH
2bUBjnOse72v77q7kbpzqLnJnkNR2G9lxrAOxSJRqLo9qR0YufLP3CXLdjkpTmumaIAIMKo8UIiI
Cp8eLk1nvFslqVT909XKrQ3LTWH3e0w6bVmxPqfZHyP8aGvxLRKaTRz2togkOIfH5vLBYp3DnZKG
lDGJVvGxfjTFLjzDIvSwUMX+Q38Taie7Z4Y9Il7C4v5CXjl/9Juh+srOqBp2P3FEXEavbCRJ6lia
zj6h+LUB/wSlWlMX8vDU1OSM7nP7jag1n19DKyV2WmXM3g0PDJ4YVAWwRd6AGOpUVFvQk3KEtlUL
BkUCmhZbOAf4e94RrPlZvPzwS71WiwTkJvENrkGWW6cTKvflTcUlnMAFE1JK2DrTNZa0QoGeqHvd
oamXNMM5a/xj/mVKFsyvEtBC7Djqb6aBtQC3eLZqkrykHxIqfc4xueLCTHHC16K69HPa945Ap0Ej
Rnu0Uj5oH617Yk7l7zEwrHDQH2ayDGeTuBcw1tu6ZT2ozyyfk67OkvsKWftYO1+xrefR4B9O8W/6
gLQ2LdmzNBFyABofOWQK+YTCBmeO49XSRx94qklloar2Zkh/nMbwLfyZACqDTYnM3xxS90DBO6oi
lvSwuFWgL9TYKiatpIxCe/Jo/cLn8UYYSNVr6i6Vb8SWzjZUdnDDtg3Ssglp0Oc75+1livDD/E0i
5PN2piNLUmYJnMYTsqvXQZffqeSAuN2gB70+mt0bhz0NnJHobB7WKiyqwsH1BymYeZ6RDeYbrJ51
qNsbaEkgxmccn2zUP7bauxrxKidbAKBUznC7cbzzKq5jC2rEMbaH7xS1smkMSxAugx3QkIU7RCTS
z2O1No6msO72d5RpTEuuSOU98e65HKGtaX+zMgAyjRVnXj3BlGynp+uSfL6OyJUtQRG5AmcSE2iy
kI3CHLpqAZLSkSYpLiBzlxghgO1jL+zuRxIOvzKotHuHITDV7JLSY2Ti1Vfubwc0IEmbOe2mD6fP
N1sDjdWwwogb3aavWUWm7ioUbPMlXLjg6FQboi2cKT5Im3oePmOzr6XtpjzFvlhBxayE+EBRbXi1
bka8hnYafJ+WIVSu+bEGdjhlgTQGAHPV18lqLiC4HglFxRk1pdyevcPeDHL38TRDpJphj2sLHB4s
0VeWPWt7MyI6QorYiI5awcyW1fHghS6RPuecvAyUXFymleHTSiawEx9j7aXbio8x0hzRXUYpnkYE
KRDD07oZQ9+Vx9Kj41Z6dzwa2aiuXCL0wO3NeGmr/c+J8uy2OaW3II7qImTYBddcub7qLuONNUnG
SdYV1b9s70pMAbLciQXFCb6tlII73iP3OXv3ppO66c+jTYErI2ksprIBCmVo0mFWinekAet7L4qw
aCfh7Z6ZO0BPgIFaqT5AcoUtCp7Us/+FLW4oQjopvMrwDPNn+2pJ8zOQ0u9GHts/BcK4urJrWYbQ
lbHKPwa7OIH0g7mS7LQ9N2y98Mh3S6hmwwkgY1+W944Z5uDd61HE0JvMQzQ1Uz4iOyj6UK5S0RC/
IkLw3tziU2YRhrjIciNTZdibLJfY/ZJrQ8nzV3dB9MJ+jpGjEHxwov4MThMzf5udIK1/tEVS/Enl
BARLi08aMPJNOLzbD/sUPBYybcuqafQVzzQWGboeWHfSNOa0ykOyaWbGI+emz07oAg9/kvxq18sM
nTGEPFFGJzWIXZINSFxceWqPMEL/R6PeH0lKctfPSOPH1r7LkuXgXyhFFkEeXeBUoLy8xxapl0zF
kMHyDrdCP8jU78WyXS+2GRu2vzbFBflTsUF37Q8k/7h9s6a+Iem6XinN6fbaJ95f5l2Qg3yzcYO4
IzyWrS4z7J6SaeQH9VF9bwc4u/EnsU313n2Wywl5Ku6nkJLe37vbLbDae1pkRfXbCYn5GHQmolpP
4Pkb+QAyGOyOBlyy3VLOQ6/Tda8q7j5CH3kZTI5vQTwcSBLD5g6fRib6dm1N/sw17T4PfR1obNsC
1w57ZSXI9MzgInh6pp3tHONLmLIHIU3AUTaaFXwVZm20PQ/rDRV4UQ29p7fV61nqVdL4mYxuvw7j
dS6UrQ15reNXdkT3SVAOkG8vgX4vBGg0SFJfcQ/YGmTLqmkJKpap/P5//eBnbr5LmwrnNWK/6B3Z
xB7ab7AeJeB60smQlGRBivYGtkvK0A2A+dwmHFqxBIe4mbW8HSNBgGRwhIPlQKt9FKYuR7lT7YfO
tzBk45qMjCuF7mGqCkiB3kSSkzGLldpA3DN4iy1KRnaI63hHUdEwXLIQCLYmAF7oruxG87zMIYq7
zLZjIy35Q1d2b1ATtwwseoK3y8TM+lpJxYHrk5LLbHAChwGNvZEwphdzS3/Zgq4+z9WGnUjz0ZG/
9I0yOrIN7BqJKKn7QZ84ehe7+iAro9ttPOZhFx+Pfhgb5ae8VhNcUz9zEYGHt/iZSe/Yf/qJxyx1
J735h8MhEuzJdO7hSuoc24Ozo3CTeIpQRSzQ2IENExWb9+bHt6fJMP2W3jZMXLOMz6n3OusxD/fA
iWrRKDdPES3QaEg/NbkGatinCJGsJN6qRkA5Tbs6U6iuZyQ2AZwhOx13AuPrp+yEOhJrFyvtssA1
254zi9VHeY/JCVXiWA5+yYegg3sRRgPq4AIRrRMt7ej8Nn9N5k6+TfkzWFgCmxE8CzVsJ/XGhhz6
a7i4K16W6A2bwIAxNqOGaJQgFsYiHJVGSJ6rDGS8UUTtWbvpLhcCqgCtJSWZaCIOY1H4USS0aeX9
AongWFTuSGcwXxTPZa2laRzs1ADtmg2H3Qi27o1uigWanj1+bFct5ReaVw5L4gtqzgw/qMiC8XMw
gTwIiLVObZXJT/kIevEBQ3KTSwBBEz18t5mHyMN3sHUzxBORkIarib0ni1U4ReCDcDCNVmBgbkXA
dWCBhV+14ZvjNHHpPBM18eiNO6tJxFlXqVakC9JCHrjE0t+UXrIcXIxeB/B+gFMguzP4pwbAUC9w
IVW8D910M/IBlq3/NFQ+lwOB70NXiHfGf+NCtVSJiKr05YUy45RMz2QIBH1A2qDgPbzAhn1Eay9A
8BV5G/Pl8Qz3j64LFKR0Q/vc7pZnBz2R+jWQLCuyhI+UOLcR2qHUcum9Omud2vWIxssCOJj8nVP2
w6I9nvJ9D8Z0FOoA3JEdIL/6b2QZ4GwIQXk3YNVgAo9U4eHyxOFaB01aWO/pEBqwCgvArpR5SLZk
81frirSWyYcENfidYk7F2jK8U97jEl628PoR1n/Hib+MM1Wrdddn88IJOdJFAKvRFVcsGtc/KkQB
iliOsqJgG8YMr9+XMo9s68Gg4UtT9TtpPHeDwWF6vT7mWi0ASYc2JpKUW6vnlML1GkWNgidJRNUH
M6FoC799wbmF9A+9DnVPTwwwdpNE5Rv+GnbWCdmJLRn9ffyNaiQ80yThUXZH67SgRgvnsSXSmwry
eJyXpGLq7Q+eWMQDlpAU50LjSP5YxAj2a4e1UX4BDyAsuYIT/4OhvXjMHz30Xake8e7droJy3M0t
ol8UZXswCL6npiD8oP7an197QaPmDFHK1+jOIfnYicss8kWqUKII90xEbubFcKz2AWw3KBZrokW4
Al8f278EJufoFzzu45x1eAVBRLm7i0Xk0HJmqPAjZ91hPviTv8zlJ2ppUiia1Qetr1mAGjqKDWQn
t0+9KkAu5/EkWqwA1eRA/jnvAxDyVHx1o/Ty71WOG6d2URMIoZbNHQ4GvR6Tj2+LUzMGc61llG8E
urRCxn8c06VQXR78JvbGcQkTVKepxA31lxAlm5OSwvVcyGyATJ6T5X3GtYMKEYPhOL1Y7tIzjZDq
X4JNoEdVHhxEPrBfAagDw3+hpDRKW70ZrFv43k8Ch/B72hdiNDFNZSNWAXyToNl3NWy54x3lgyAd
EtDzASUkyZzKdRrnJbLlGUye/PXKss0fYiV6nuGNPtSVpIRQittohxDKh+4K3MfjNmLUvKT/VgnG
CGUnJORtVBTAcueoFWt/NhXZLmFMQWmL+SLb320sGA2xEXRu43RTqwkASl6lWMaLm+7CAOgRRiy9
B35Bkr0DDVMzmCzkBDJkpHF9dLChpP8H9t5DWD/Fj1vwV0IipQ91Q63+8RUiy2KWTgxENnq4FeEi
onT9MRar3Jew90kHAy2BJP9Fqv/DCRwf8EelgMQW/jQtnShEy48Ehmc888Rf6OoB0ouEnu0x0PoG
6NoxRTotIDh5r2cUWrgR3mcCnfjX0rWtgmsJa8CbgOGXDQeq4WAt5acnNzIP90Bn5Q1Dsi90lEYQ
uRSIEqzpa79/MXQAfg1vpNgdBYPsO5IFah6+zhH0NfN4XSvfvOfL1NUVQvpu1zmnMuiODMRtUuaC
WuRb/g0ehRuatUx2c5LqNp6GTPIZ3sUsGAoSAabClyjRTASfU252B7fn89Jq+rFSbpwRAXvxdTQ5
EwHPGJxl6Jqir0fWJQOCbJuJT/vlm3HHQ1XvuOc5l0ps5QyYkyfODPR8gtqo/+uO3Dqe04IxTSl+
ex9K2Xa9cI0F7kICOxsa7OTom3sr1UhYQIK2d9qbWrEVnqX80i9/K9TrAb7rzsKfKbazkP1EuV2w
Jmgqr+etDgb8p0ylQrg5tUpUtmiLQFskHr5DCNpd6EVfcfmk9mOMBn4gDmMmPCq5JIui+l9aAZy8
Tf2lsmnTXXK/POo1IoeHDsvsM6sTxkzDu0wc8pQs6oiVxHaQbt34SyogLmrUfE1VnO80j0ZtsYzl
SqgghXioVo0dIsEsGdeYK+TM+QYvvTUW9/VRxmH8587qHjR7n/NlRCuoHYZ4HtWrISiLTdqMlrOm
PVc0qJH8mDnr0mjJUCPwO3WXyrY8aD5i547DGXJ90Q8Nw2c7uRKTeL1GThYvZB7wrxoUpWObd6Qw
j84QVqHeDyPt+Xju5l3a4npBoAOOTgl3rRtg05gyJKGp2CMpdaB6AgcC6Zis7uEuKccB0RrMS3Eh
tVU+PUsLYeXovhHBgLiO3OVvhUHqViBdb3621E6zdNEE9/s5uVAJnHWQllI4ThLi0YfRCIURQ3F9
9VQOjSRskQa3KHYxv0ujnJgbs4z7hH9NP0qzF9LC+lSxxS/rz7EtT3ityiMcTnGk+yuBP34Ll3eR
5qGFb531jzF8e645IRVpYQHKTkedqhzE/cGxCMNlvtti6evig2IjHSqvJMLsL7csVRiaEJWqRcRw
XTVTmJ9SvK1PfCDdeikBJgE38kAjqX091HrSH3YkeAUecNDaIoGHz7gBgDMrpYxpC1rQK6RcHz3y
TvqzPdl5efssmSsPh98i7Cud5eoWleSmNxk6rZELf+n86OCmy0yvZo4r0/JPzNF+JNLw1omCAf4r
7aerAr2Igy9zouKwF8QVUPGfAuauB3EQNUBzZRfwFrRQhMC+10bJzH0hrtD1DoHtm6mP0fy+5fn+
Lm+iwcRc2wq8OZohSDy7EfnXVP5bnUFkeBwVgC8PbGRckwjwfqMUE0d4qw+t0dV768MBjtQ5PJ5M
gvyCHalM3dVcN1fpQN+5naoRNuyDE43jj+sVDUipKebwMJsGay03lAi1NDgHA/zZHLmJTRQS8kJw
48lrXfn/JOe/kF/6s0DW6yz2mAxtgg0N46tG5eFGkCwwkpJAUCldY4zeZn1LwLDUM4vd7sTZty+h
/EtSC7DKYZRf15LYPjCJJvhWykAFYVAj5ptDu6wE1OtCwKexaVZsdoajoKwG6IoeAsSP0rv+T/FG
o5EX8POtqWaIwnJL5N07viso3aEpOkyhUv2+yNGeuXZVzAx91YzsUrxRNw3oewcf7hhwTozOHKE8
w4JHLm8xx5XBvfGr1kLNdZlLLd5QdNG8VMVWc6wVXW873vIr5jC7jPD13aRyOqqckS7ZG4SDBq+c
Abrzw+A9gzISdVH850U/wj+yyG7A5/07GP5RyOccA638vXDRNmA/1MFuT/Vz3wY2oMOST2vNcQYS
o9dTXvS7oiRwBfFZddKy0coqXX2HxpFIRgeWBrfv3VK++kuFtKOLdVDpA6aa+IVh7G+TLe2jqM+W
qxIBWE8OjBtJMPkVn09Xd7ru7UvXS6pkU41fqzdhMENpMKH+cJ5zgp8QSr2EOSJ10Gmhn2SmxPS/
QACRE4tuUMLBkrc0EqCt1FkPb3yd2zyt0Yk2LtldIx6IEr8elv1J0mjfVKsrT2Z/hk9ca/lsYZ9k
01zF2HlPGlk8vnXDOH0hF/hPwY7rkhAgis29t5w7Vl/4lGNmYLFAdMrO2mtY5Js48iJ8mUK4CJQa
mHeLra+pT1/4CsFhiRuu9KkR7h9CqT3Nj87xUcnw7DVEnBZJ8GbCvlS58TBxe1DYGHCxJ19WF2u8
I7fFJIf6UtCfIry03bpkgnKyDuki55EtaBQIS/Y8GLdzuDWTOygvRJDqOael42Ei5qI4fNYwCSUm
rsEURBnt+F6o2K0/glPSjZd1QoQ7K5dl0QXhZ1T/qyKOxgz5Xwl/W0DAsV1LpJVZ2UG/jEl8v3l6
8vcSmi31VZlFK6Cxa7J2cHi8eVGu94Sb5TpFH4zGl/SQus1ztzGLNIKvzJIFajG9+GxTMBZVpQIA
6DGrrzvViSrK4PhUnS1JNeTeoD6ieOMlUhq3t2unaPk0Te4EtAgDv70nIryDJOYz2Srte3sj8a2N
wZNNovN3NL+yHVpuPgCNJRkvL3vRCNuv7obD1/aeWro+dHCjcwjSgxl3faaYJXFrqHp+qM4szfLf
SEqEiJIm66EMhhC5nsRrq8SS0dfeMK9SwioQR8zOQR1sjNvaqAirnUH4INB1Xf9ZeNHkqhlPMesY
FmCLw64xhK+FxsaqAOKb/w9GSP2wlG1k2Bdrowr6kwButRivWaRiUBgJNHboY8UpsSu3q+r+CFcH
xfDbLAJfHAsFHRdBZPglSc9qfsbHj9TCpE/A9lw1b6h6L8BgIghZooKuKsiX/Q+hgv/37nHbORiR
HMwjIl00CP76Ij4MtRn/BM5mesjCkaDZc2pMt9w3hA6KOFXM7HN8+wv8pHkw41pLn0bJV297ns86
9k+6bu6WkSBSsy4ZefWTj8vYxV58qjyqabXcrn6KNxZl9IQxu2w+rmR2GaZExKVFujV54ZLzz046
jKf0M+Ao8w1y7/+/D/p4eSqxLW+GRLLKXMu8LJS3oaKMbsr8yPHA/gIC2PejgC2HqwH3iv6l26vG
elADdkV6p70Qcq69LVXy4Pxd3Yj+OuHhKLyrwuqaXjbbtjPrkXzweecYQ7LCk3Lj28XgL5u7Pbty
LTbD9awXzv57LnzXZDATBDrHe3z3yTlKBUnns+B+a2iJp3FpD3uftpQD7eNVQwXI87GSRvQWR0pP
EqfAM3WzQ5jB/gNo8qL50aDAtuOtQnRaacQ5F20zpwC1uRxWnVEY20snzmT8T3HEq0wDzqP8sU/Z
w1vpqbLZUw6kkvcL05X6g8LYyxHibMNa5zIZZq/C5taJ824lgMeagGVmtm3cf3HbSKWxorV3geh9
i4LIOQNIb9hPXgUifGMsd2eReu7QeFWAFkhyGWeh8+RdBPs6C5Pus5ksIZAeSq7muPq9U4dp392F
dOZ3pE56XLZloMBuzGZppJtRKR5sdUB8v5Qh1acGbNv2RQPf+vdPrVN0hcTGDxtMKgGJHFYix9R9
ptOuLybj68HXIcqhLy0xtAMsZfcj541e4534wuqfHUcNQ7EWwjs2e5N3FXkZUAswM/qnpxcLxtgg
6JJ8d68dg550E48FD9iOpQKPcuhKn07sspn24PkPG1KLJrC4JgCczi5xemg2APr2aypPYeIMM6Ju
cY8UWdIVIdNTN5FRcljk4q5K8NiACQJGI4nvtLoNj/K9MPshaeawmC1A/laEYR4uat47tTmtdDzV
LQPA6lP1DNj3717w2DDpCXqxIA++mmJoi4ye/9DzmPvPD8xGvdWzeDZJJO8j7UICGGOoULV7TXhM
/qHwXJVwvZQuRucrUaTh/apA2JuymclhgWWMdCzoqmkix/e52ohs+ijpr6BJ+O+mv6d82eSfAeAt
o/PeSwoxhOP9Wmg9w1bZ1BuIADXfiNs4YhO6sgtefOCEp4aIz70/+EYkB8htJ3dmW2A2u2/myDwX
nrpVyVvJukYGZS5rquSw9l5Gf6U2MN2w7YF9OzYFZZLQ5UeGpXrI9VTGMKi/TvpoQpRCTSlR2iKd
7+FVyJfsdV9Ft6R+ananZ0Ep7tlximIpqu78UO5kB9Ka7ecPp6UQYc2ugtYX5UG4FVxJoKQ4PKsy
IfN0Hd6QDoT9Zl94uhIjFAgQUHso3Cbmzh+l8kK+Oaj/YpWzX/x2oDNhVgGn8AX5NTHJrpNOrxNl
n5n1Xz1vncjWbQQ0ZK1ZYh6nLAnfBpjyxFfInuAGt88pFne0P5iLnOHOCaS59PGk53vWAq762tsD
i/jWfc8q6mU+mMtgVLNMBDZYCRQNHyilQgdP4i/avJWRUcTxIQ+kJGUAkPVm8vpkvIxHCJpagWeP
5mbAcGXGxzYi/8SJWonZpDqymptkcdSVn93Zo+htaTj/pR9oWqEJ02V7JMOGfEBZqA5sw310D4an
1Bdw4XLiXJv8hSwSID7+WSslPjhQ7OwZvUjEoP5KCAIdByl6rWUJlDbDpasEFhEkpQkzwVUHPTgi
AgZtE/vwaMKt8bls0Jx7/EflOG7LdLWtnclfBU4gfG5V03pFqbn13JyN4QG+9KZxEfNcWnCVZeoj
Yu7kkd2ZwE7SSxHxR5OrrrUONkWpwKh/ful9NFrXidms5XnQL+VcXxZxt00cE0JsN7XiyszmXXtn
yax59HCLzqgeTkwiEQbcwsGoeUOb3XKjM43enfDfG6qq8sw4tbdxhVThU1CUqdmkyhoA4Rit+Dgj
YexA30Yeriex42ycxQUcui9LlhvOnMyRABIHwhmWQZ1Hmh1IfkY5Ta5zfXeuwLB96xHTO714BfIv
3iNabSChy58vcJXNm5jx2jU206dq4gSBWt5JYPYDuOzaaBVD+BE4V8i4ee/ZBwbji5tiTmHerovu
yXJovNv9O2cSwnA5vzzbVsf1NffzsdwyaizhLz1Blf+o+C+geuDqEoNhXGhBuLemT0y+EC8vsGKZ
X+lqTThLT91LkUzIf5ssk4c6U3E1aaHQJLJGmAfPg8mlPHMQ/hXz4eObozGab0vf/gbz5qb2snUe
GQ8/roEc28lwySvHuvmje1oIJi59xR1EDzSsv5jIUNyFbXvLbMqH0oXDnmsWJAx1kX4ylGnVv16I
DK/UM7cNLnBwxF+84vPMBCs8GOk+ewL53B96ZIfyf4pwvAp6cjK4zB8YRf5bN/buT+qAauBxIzcs
tZaiBjoKrAAtbLZP1Hl1LgoFGrH9DNjbMGtu36XrCdlU1RGHmlgAaivL3JrFvbZV7V00KGsD5toa
knyNRIkRy2+PISkRqJlNIWuXDkf7ku6gAmP9uiViY7viTOk4P6DEvSJFwH6JsXQbXUwpa4MrKZk2
7rBQG28E+TQjNOEsBkUDgSaViRXSX5nxw0O4vri3uI3T9Ju1SZHY7iV1cWw9rRVXv78BTa/McPuu
ieSTA272GNWiAQ8j2DhAgBGwTaVcw4yPBRq5BVl8QyI31V1CrRsQb5AfIpOWbTMBt+P1R0jBW/30
BGhLnCjz+4+926ZOqwqebtFl1fl068od7s7iTkn8ZAWuKzSSePouQKxfhtDr5XWpEuPF0wNJYr2K
7DhROiF4SW8x668fb6LfRuR3c6Du0Z825niHUUlYnRMVZnxWdEViXavUmH5XzfGwtruCUyrSUqvw
nOohQ4B+H344xQopEUR3apt9DsByS2N+Z92mwSM61ZzzbNFlPWOaLQYhpoaGEoLCCx+I5pyEM5sQ
6UhnR3XDyU6oN44ngl8rEIXIUf/yRpCgD5v1Rfhw8TlGjrLQ0nqKrpihN1pPXlwVUYc+tTcG/hXd
lAO75Bib+AcRiGK8lw8Mha0BzeBl47XUaEAjk3MD7of9GshxhtsFOHrp8uQeANtvInZ107Oe3TXc
vBEfmc+1c6K0/PJ2XmRbyRzJahIXvVXe4foQzYXO7tJMRm5s48Z+9ywWva5STY8eHvFAS1zFjZYX
cjj5jMAEvxmA/AhDwV3uarG82txWE5cfrLa+gS9cnijRRKGwK6MkKkv/0/sKOd5N1fuE4H+CCaWC
J2T//AHie59YhYey4qFuWomAgwbfraefFMKso+oG8DxgT3jlqAl6/7HkoUEtfhpc+yTwYMxxNY+i
UxPuSKb8gWn2fWeoQxtGTU9EnUChOyq3OPNqkZMp7MAOPwxlTccDnTqFyCgvZElS478WWfoafxkr
TM+HrZY6+PvnwpUEFtl02cF3ZaDDf0DZrHhzxA0CSp73/LKBAba0OyMoGeKV+7SKIJnMjBFikhIS
HLAbVYp0HVHsYzPDLdxRySLk2m1j1lEAU/Fsu7N85XVrytLsZHmmSf6FXQmibCuigtn5QaUgpLaq
YsQTkU3FCfwfysSYsWoIYbSJ3BPYGXVDZWZDTYV5dbT17C5loFHgy0V2m5WiKZAJwkYUNEJGuo9I
5NMl8baNTSOPor2u5iFbklkdy5TwjV7zSv5LaTgxUvqN2MQPf0AKpWoL+3rvAyIVU/7TxZqwuW/4
tqnbnbpkYC7QFLqBLIsld+ipOgJ0uG4lx0xcPTnomVfZTRZmcVstqLtcPJzuJIKAeHblwl5Pl+cg
g6F+2S35sdHnAJyOXcPBnyHvwMN4CL2NXrGNz3Z1IBlj1RKYxZPkjm/LnEhPsKkSJdKUoBTJmuUC
r68sAJYtyX/hBgveF2siIq/sBcv08RBpTrDg0oeGs9Tcg0hC90p5mPFpLWHEZJwRF1ND34otCit9
Q4hyeLFOhC7JPEQbmH2gyWGU40zitpXYg0NK1oJrIzrrOnLqoIGFx999sScQp9Bvf77Uoxq2SdWv
ffcXFlSLg8wT7tk00LUTLo032CK+PKbUESnJml9HKPoGD9x/KB34FXskks5BFQILT+v8CB/bQwKn
VDxnzaItN8NBMCXfPvWXrvxAFtqXUN2heVj+arIXmOJdDIcfZSLd9s+Atbx0sKanA6+/czclFOZm
dZ9fOl7rV2Tipiwlxd4HSKOYNuKc90MxO9Xw6Apr+6vv8PHiVqPHsBprXqNwXryvJUFnwn4lpYO1
JPV9fJWr6UU/90oG7d+DDi7RBbyPCqxp9OSK51oAfomMXcWONOgcoTYpp8M91bOp8sRbjfO1awgB
V7+71we+4HqPXZFVpyIYnu3q8NFbMnaC+QD4JryKF0ORmkLhKYB0HBmUBENxyiFcaPcit1FBPN5N
LzOzhWz+jG1Jgi4INPACRz35D/JfPNHRkDBmCThnVvMrJyOqxsPiy25Z0PYExkuryXibTtXqH8nO
wiTZMbylk0ezGOcLCvAYszo2nD1x2Ln+zStoK5mPhbgA74kMUyqsbwgfbfdeRXRXLqQANOQbA5o/
dAf5lqsAbH5f0+0H9+b7mmY7LYuOET+Op+XqFpY/9zfM0wh4jfnsPnteVtGDs8/XGRvKoqXgrPBZ
SEIGNFM9RuyB+SKyw/9Cwd6Eq0sYtuR0BAnO5N4PImzBmZbDybhTwcvkrlZTPYNntb9WZ5p82+fl
hiL8mBhwnvej+dkfodNXFp9qhnhfbP/s9d6J0hjELVdJ18J0keTkKqErW6YpaCHufRwC5ESdMphq
NO5eSDu4Mk45Jyoqltoc/4gP5WyYwAq207t7p4ZmWkQsrd3UedZb6AmKX+41uag598+eSksCeMKO
2kNbxLLsj1HJUKmXPd7tevaEywi/ZHW6ZPAfncC9nRBOpbPthrX0KTCbo0HQSE2PIlhK81icocIn
MBnr5PpGglx2GFtwTmlZXA/fwdszbNHObKGkzwRx2r2ALEKOJ4ZhxCC2/5300gU5qhei4ui2Vdpm
j7s72Bf3uVP10WBXYxXUdn12+7Vgyhk9dyM1w5S39aEfvqrds8/yu9ZalErJRCkMhDQoS7DFSEWd
6ftRtREOT4t5aLCdpc78A+UPxHECpusLcBdf+5h6tS5JqdkDpZFBh2d2hffo7KeEU51yCHrloWyb
1yq78FLZk4xeLQPm1Zi33KI780GlStZzXHY7mw48E9AUIjvnFuvk0tKfyvCSrlgjEAVyDVMz14UX
DYffJ7CHLxdAEpHKCUkCfCODsY9WZGRIo8vp0kJxO8k+eUvxp99wudxQ8k3olgi9eVNexr9jwrVz
niStxS0LIJQaAc1g+pbPop7GxzKzzQcpBlRrYmtcJ3XpC3fy0sJiQqh+DW2gN22HkandGd+Q1HMq
EFqi7tQqV+I+ptpsi+T4JWGoyvSFfDRngmnASM4OB7CegZe7cwSPIQa9ihUWRU3L3uL7i578AmFF
xn4oCQdLoKqrvAA95dLSMYbyBCHKanATq6fsAcDUcJS4TirzbI1JFi5+VWqGnRkme1NS9e0UkCrS
CMZTwbE+FCPvAxi/SAB56zXjhMQErlocR37l1ma+TAr1G7n0qqTr+BhULkHJdocAYxE8akQEsXzc
+ZL+59/lSX+DOl0mnyC4KCF7WW+fcLvUdK1qO0QUzkNCHE35T6xXjjVnpbg8rV1TWUtNhaVB7juQ
4agFmHpIJaqNDGgvnYfHHXxWOWij8JJTBSEmaSZs8h4VovfLUD4THYujHYJljrAYjF/aWgpqJuD4
K3zLyYHorG3MikUFJumBEGVldoeoi4jHraUQjkMqg3xBHvk1ge7ZP6LSgj0xpaqCaiEBT+kqioPg
vM+nJ8yId4u0q9ibdT6BQwwg/BJeQ2EW7+4kjuyZpK9D1+H7+Tzf8iVpr+TqBvOq9GNNkaHVUn7Z
EP5UbIh+jk1clGaUNbWsybQnahegT4y/91kO8KzosAysSUU9StWv/bdEeXe0JUoQK0BAqjvrmq+V
+a1R/peuQqO96am+NTBCW5aV7ehCIkAjkSmEjr/jbwC7h8zxKjUtvmg0F4/6MvDUIxTXNTcvp/r8
K1q8WcJygO3LVLRAvn7pikeaVOmBC91o+rZU+AdzSr3EkFQFyHBCo2G3fNyofViGGMLBa+0W4CgR
CjjUyJ9fY/gtQRSucqFunzKhTB6AZ5DZMRBOyNUaOMzo1iEmxxWP/71iG7p/nbJu+JZBFmbv8gMn
cPB4stySof2smuqWX5M8giyyN4RA26dIPg4xpps+RX4RIAoyBKu9OZQNKDo0ZDh3vV1duIlm/VxE
WoeICQoa+TrcIdrB73Ef0L61QGxGaqkfWDtuAFbjuuWSA9U30EvRd1S3fGV0MZwAWkscwnjHyjed
deS/vBwl74zf3MykrHHXJ2L4cNjLVLVi1aQQq1mm3e5Dq5OnFvXMSj6SQkiEbB0u4WoFO0dVcOxZ
qqeHCJX3f56m5OEYTRdgHnPIIKt/wsPDBHyNUVthymK4a6V5aHUTBbwknwNEOI+JK07W8xLKruqP
MXnuukAVbCVEnb1E25CTNfj7BkzgrTO/Ow8YDEGY9CBeiEaFqbPldPtn3j90VuMUKV6DsSQfivEN
o/s1H6fenOJnM7RPW4ous/I4e/BgDxSQE32X24r/NBW4KdTciX+CJngUDDhrAHX32qKXgovautb4
Hb8pKGckCVd/NfN2k1k/bewlIfImrd5fbsWGKs5EWq5VW9i6J6WQ4XrQYbtP8odSrWXXVNwIWDaE
hB/xeeUSFFAhk5NxfpYB9RSiQkYU+47dIOqMIYa48e3gg+xiAIjVlHDs7Uimym8rTWh1Ae/OIW5/
bPLfsCZtGHDgassr74SoApp5+CoPHLuD0M7n62dbPhNar01N0CCPcQVR1x2JEEKpdoQX48x9VGD5
CimXkCjQnLxUkwyY/NQ6kHr7fV10GsoaDkGYYaWb4v00ovYVQ+3wPJycQ7oyBxDig2cOsKBgwTmF
DTcxSAShJABg8AR0A3RuquMoAUNFEqry+4Qx8NHT3Itn5tDf/E/N60Ze6IYF4oksXnAunxs4W/Xy
9hOFnckxr6hTE5zs+dA/mM28E1A1Xz7Z/OhFWGEhNgkimHYnHVftkjOsmz6weD7h6jJ32ksesILE
KF68JplCb4WMNqAhgyZ+bBpfJKgX/CKnV81rKPbB167KVVygLER5QjLhFb6ZUs0LSh3sBBttim2z
P1wV/ujAOggVUjC5hiawUt/h8PCo81NOve2Tv8rTrtzCVVLHfHespt8Rts0Ocgle6NMdHQb7fkEQ
tHbBMvGh0bp5iRjSXcix5lR/n4m9us4+oq5QYq73fqzvTFtQ+runesgINjan1awS7cbcJoTv93St
28VKHJgQ0ek6i3WA8dYcKQXsCwQ64bTXtyPKGCfHXxajqj3HevaEm52iMyV1fYRz1Sfec9yyXKKY
C2M8RwaVkcHUmCE1cV3buYEnJ/ngJiryIqW9i6fDePoesyn4vvFNIxVyJVTcK2YvWMc1u7k2H6SE
rvhusK0fklIpDwmAzVhBI0olTHcYbp5UEVwBX7QwHukO0yZH6JTNiD0HshFi4PBoMofp3ri5Yqyn
UkCCf7PQr2AvbTRV5dBe+zctihqh0SFNooa6mZgrovkIfA/9sPxZvOWCcXJEPh+u9PCvxzkKbaPw
PrdfK0zspnkfnxt0loXJzFSJKk06SZNmm9GHXp/pmoTJQMRhfZGMR3DE9bws20NKMh3WGCCr5Dpk
U/gfUEwKP1qfsjgSaP02EwaXiV2s5RoBpqg964ug6VpQ5shZhNg9VLWViTXivFUQnO8v+cd2SoUl
2vOPTqUEK06v/ik+kwayAHPB8JMi3l4ARpOTjXzFGVW9LHm/N6mgKidJ3T8zqq+ABNNKHOLt+5Fb
v/vE2CSuKaAAIoEkX0Xe6g52MkoPvrp3n0MEL9JDaHdeUi7f5Xo5qZg3QTyvUiUCst8xFoz4Hl/6
Abbls2VoV1sldC3O3omQPRxBsjrJWY3kKHzUDhhDLUrjNzM/ay5J0MzsFetxCoIU4ym/vsVxp8n1
aHW/VvPIYYG/gARkbHssL+z+NiQwmDtIUKpiCE3LtFqB6t6MyUrdiCgqz6Uik4Byt/prkmuEMq9h
uDQ8yDhQtX8eLor0VJAi3yq6zB2k6h43LhGSc1ZSPfdSdoVoIwAZwgw99s/dubmy6oePXhfyJ+nv
YKPOy0UFtSliaplc46UDqgNWnpHzrhvB6BJWuMdqRMnXSSVbrNeTV+9QUeHtBpt1QQ3fXltK8z09
zbiOdaJ4Yx21XSzpX0mN1mQISaFlZs1sYlJOSY9OruFdPNdApt2mos914bTYzTaq6Y4MAzSJNEjm
rmA21UiqPO9P+pN4TzY18b9qCGWIwEREVVlparuQbhydzObwbNb8Sewehc2LOPQ7FbAjm3ZqEsu7
cdKPC62wygKkpzAu+mQQLGwvj6WuLdIC3r+nQgWRJmqdcuyIITetTN/GPAvqRx8VxfBVJVWFjLbT
6FRL8MLNybvLiP6tcTJQFOTuIjaP+K3sNcCIo9uoydqPsLoS2hWSWaLnark+SCLl8m+Ds90PMaUy
w6fJwr5YUiyX1/p0n+l6c7VypooLizvKC1jYwkYbxRbfmQylr7goC8oUAagVNxOI5VrI4PC0NmvR
T3Weoo8uyCzC8MzkTeoQO/ALU7XIisudp1lBJDvyXHaXa7/uu+RZK9Q5axD/CJP2/TxwbnplTao2
nzy+LjOmBY/2sWf4DxoZFR0liVF1g1KGQHxJb6QkgLmnRnzbLTrCM79LuApi2I+bOz7lHdDSA93c
RGLVKG5uQaOw4KlL4+uyIeQeooU8NOTNP8F/bcjCsUFtMe1b3EDFObv1T1G7l61v4B3rNSIGdxKr
nJhtdktc465ETrzcKdQoQqPLT3sNpLmLRc1rz5Qv91Q3BbMju+ddwoE5OofDnvy7tzTkpbm+WAgv
XKW+sbjJXEMer6+CiIfB8/uPPznpq/OdypMnrAfl8UECzFTNarikwsHNXxKJYV0CSSE7FE37ZnsI
GpxAMgl0Fb8Z+xWOHD8vLFThz9VJ0xgw8Kat2P4EYmWjYhaa9eDiti1uGJeeGf4kxJdBrnlfVSxv
GncttLG3E6lCFmFMLNZIi62saPaIPkycP8mGCEwwBfMG4OUilJlj9z0dX3lx5jdWIRuRMnLyWaeW
fk3HLX7G2X7yBGRAhc4Lucnmd7bZXpX3LtJHsnfr6lBVIxWee156k60thdiCS666zDI+O9EsdSbz
igeFK9u3evOnEt7lEdlq87MmwjKg5P0zzKFbJgS1A5rlh0x1tfHgpI7sH1dZQSG2+FO8QioJVTNh
piwqDpLk2y06X5922SwCLyl4vCnaoyVabCBHt1TynWtByt0dH+yNuxqGaACvpa1qldW0xCc+WP/q
z2iNQfZWBGn95Ha0iLk65vxLHwtZ8SIL+6cJvH00a7pGGY3iSpIfFXbgJDbSoujG4LaT3y5AJViG
ZkwAr4tNxEFKP3BRIWm7tM/6RIQVbqkADCiwTQSairAj/kKIvxRdNQN0eYnYjPZqefOIqeE+0odi
fbJTbfrOeWiHN6W0CW/rcaPoX9LfSkRu0jA55F13fWrFsjkVpLkYgSlZZXuqIR5XOQk9yjfayn+H
UzzaDiUCwqJQQA1AN2jdPLH6KcPqBY1tjpNPXgTLtBfWsdiPhoILFR+vfmqk3mdCk6GoUo1+g2b7
CiEcRjH/iE4bSmy3wI0OUY+hbB0+2Kwm2ifEyH3RN7JkQS8cquCsxputUIytkDWEz66iGfWoPkFp
6LiV8uSIliV+/cvR5FABFv00MFtq9K4I+Ap/PcrhAmSjZ5ZKB+YhR/LwZoTZlkQOgoPYLPJ52g0x
z1mYFzNAcw59/YXHGf5tuuEzZr/Vig2Uk0CU8qjLQw4l2DhsAhHqNfXn3RYZpp3M90pm7wpCNmRS
Slxen9F05s4jMWJTUJcxNT0h/NUadpYhP5EheLnIR/rBm0lqZxXtVWMr74uc7wXYdVS09kgAcymP
fkoLSK+O0hDGpXSJDE/U+26nXuezEURxaxgi+XsLKOlYdsdG4O4Wh0fLIM1pgjaGJzT8spQhRkiz
amoDEmc3uFWsxmbtQs3sM2ud0z8C65YyEQDfjM+0SxVY/k3GHXfS8T2otmuht0M0yNfPbiFFsgy0
YiJqEHaCy8XdLb2v6dcqWtRKIJQti4LEaF+J/v6q+Rff5KvisSozo0fmI2mIBgiX9/27XK0aoNyU
z8a1YKRAnfdcbcFlze7l5bqyObJboqwKUYT00nD2LJXKNMioMS1ggUMlAJG5oQPnYnCiPRgqVKdz
+la4vZChVt9pNIFg2rRUiEm7wcAPgU0rvvS/GomO2GseCiuMoXJy/z8DUo7KntnJZ83Mtxh+pP7c
B3+EjGjHUPfZs2vovTmRyQxaJp18bhtfFLX3t+PCKobfdS+k//63yHzIHqvPMrbHdRtA64xo+JBt
dpMufVUX288nXbq3VV4rS1cNcPJKsVP7NQx2Bb1SuUF6pA+6BayqxGq4MZODLzqDvt/2ghl8h3Jf
U1XWosZ/aAydyNuR57UZL+qpUWMYNLg4OOnJQ0JQlwn6Zkejg1C5W7ZKxFTi24A+Z9v1OqItCo/N
a9uZ/lTSz3iN4GX/kPUvXObCLDeSOFClQEryEUpLhqvQH/ujbQNWG6uzHzrnXH8BVF9OQuNsLnKU
s5aCZafznRbNR2PMFLYMNelv0XlW3eUPL0rmupHRRytgwGb7tP8NXus5B551fbX8f9TBlmRPiRYu
rzYNaSFMFRizOZ+LAw/L6sEM31v/DVOO14wG+U/47OGFa80/Rq4ZvsANzG7i95DdGi3wmYC6HBH3
mJIcSsXxwnxUYIcrsXwWgYGmMUZxJwVOffE95EZAYyXnrCuRhPDRYV3+/07G2bg11Tq7VSfmt6q6
ysxAgQvut8t4FGlQtuH5/hUQ++Q5kycpQAb5+UGoqYRgLAPoPNc5NBCduOa+LUD6jjY4hODN/46T
hiWm92DdAoCWYUM8X+7/NaN76gkB1z6gppNm7Su650eOp+pK/Zh3gLmHuLUGcRmZn3daCvZp1bAx
LJ++jD6fzQgkAm+TbDJeANOT7QQvS0M7PY1wx+C7EydiG6Y7+0+ieKSvew2eI4YLy3eDJ2HKWsvq
iTSyYWg9VnuIQsaketg4ivVIi0JbG0MeJraM4cZyQ8n1Q+H+6QQaZ8kftsvVjTsYUcdDtMj6i4+A
In96VzU5rj9CqMC7/5ytJJQc7wPBniqT6h87TRr++B2EcnUtaaIToCbzmXbQpWpQDjpwJndpkD03
nzZ6SiEDAV9A/F6y2rp4szwf5sr+zIQ20nMB9D9B9z3ZUG+s+zuTm6VOPHhqCqxLFbcW3N6AY5O5
COfIr9ePrfIPeKvGwID7FIcKJS/2Fic8Elwzt7+ADobxmdkAP/3Ji0Eon+zLewcLea3G4+mojHtd
thyPMRQ4BrLjO6GyWA/MdXiDV286AhlUK5PjkrrTpq56g9wBEhrcA+vgndljzWYW+r103NASK9MW
ovejw/5swI4lzyIhBbj6FPWma/57SJ/6UkQWXDfzqRoGHyFffovr1hifjHSXjSqB8A4m8YTSE/uj
l4oeZ4XZNAbVxya0S5aLVePchcdr1JavF+sUwLRHkRwfxF9yUxXe3nd+ZTHS0gTUQwiBB6R5XdYn
64op4hJhHAGTDWWcs+8l9n5p9ZiBpDARRgxlO///46CihT2VqYIasyybW0/rY1BEhjH9hEBP0EHT
p66+DNfQ9t1FspboY/32c7cRyYssYQtXARDVyeEq+D63MazmRLAF+5XxvQTeNt2k6CPrKp+g544n
SNosq0ZkNPfXEBPtLqZ7iGVWV40pkugEstnY8cIEsyvYQyL61XqsVkQYXtpyxYeKq6NvTkVDgSwd
DFqiXOMUj0Vl8N7ETipjzMud/n4tdzE9zXBL/Zq79jjBO74+7rh9DpwkfdrGqM+TKS7ANubbDyqV
dWyhvrb0v70iB7DusYDq6BCz6LxJx3FY/M9vKLIaqbm3AtQ8QnV9PGkBeWzkpIPm7S9uUH75sRkZ
A60X49WyrKzDUzHAxAZwMXmiPKbVGnCv1cz3gphmqUN2QlRhfq8PGE40uo1+xoyyVftf4jOcQ5n3
bhO1TFnUU5/wBCqHcykJ1/I7nZ5byDzSCOGJHkk6riV6TdlNrmj43iHus+ipGXHN4zdXJw1HPBC+
1obMW8RI+gnIrrV/K7Q3hzWKSN5GAcAegJoi5eqHCPQdk15zj/5REXDwif7KE9Ehww4EgfyDKZe3
3rqw2wl+Btru++OQwDn4S8V03QjAaJHbgoexO4vV3OuL7W1wzxgfz5LihLxMEApLxJAZOmUc6kab
iBG+CdPzmKSh8IreOdKmH34Xlqc9mZDzgNWsGwDd8s04czGhbkEdJJ3MS2F5kJqIbLFpk9qQkmqz
jX8DMmT+G1mr82M4bdRxrFNA6/bbhdR3n9FhcugRJyvuiHlTV7kFz40Bws0TApHqAw0LPOSdZ1yo
Xw3EJxYr2Vnbmnr3qj5cKYj2N9Yfrq5/59iLdVJc58E1glNRdp0merC8XMjTXLg/2FgRKDiLzLHw
mN466icVpBpF33silbcfD5DbGdGd/Ba1iTnL3oa/anKBBEFTZLt+yS+uOBSL9ql0fslLhnQl8gdt
gm2qKfzcjhQ/9EW0KqfgV9v2eGhMmmOPNz/1bmr5sFx1rhlFD6xlXZ23c8hKCV/I6bK4Bd2q4oAQ
oOC7VTvbQP8F11NYUd4u6sZ+uFUOJeLw8eYn2sGkoeEHJLYIf/4LGJTQkOluDGnr0DpCiXas+yMo
5ge8WTzBHgMn5QQE/4HtaevcFHrBzhpV9hhY0QcM9fvEAVdx6Eqf2xcrJ3CTqCL7zhhUCPssG6YQ
uGfIgKLWN6uy7ljD+aHSZgVT5wj/lCHzQkuOdCEnv80ihknmrFy6faVX6QeNNtNvKqVOZ+ShC/Fs
Vt5i6/No0urpfGUhdF3eO9YNCYMICDDbwozgKj9T/vxSs+z21h7Yaq/UaZ9aJapakIVv/TMDmOYS
JmMnC/n61pTeUVq9qW7US/WvrwBjpZUjfh5SGKF65qtNrLz+QCOGL3aL1D/+nEJQjbroqor4N4a8
40pGMCT022iNoTff8WZdg2UCAvWPBnJihscNGcL/ef31tikAvKI7Mhbo6u2FKT1pZKX9N278uEs0
KmfBNomDs+HqwiCnHDmetaITq7UJyadAbSpMOz1nin3DbDr2okrGL062T4MKPMVkyQSbIyjk74yJ
qVcQ6NINXdAn6E88MDtc2/hdftG5nIOX4Jyb5QqrKQVQwiqV0rJB88iM35ii1ofrarjaIqOVKFIr
zoSDNUh8IciwdFPBQi9fQg7V0d4mUoa1VjZSrGF+jPEaZAUkdTI85PGIncEu+uTlLmo3u4uTyjyL
IW8wmEcPJV5z2RlxL3VMtt2sQK3WIrWP2v+k8E7f5BEGJ9mJD/G959WYvT7hnmIOGscclAzAtSSP
n4eNfVqB4IPPKWpqoHuKlQUMXGssVGjiItc1aHTEuHV8ZDbZpPQIhoMh+//wwwhopAog1/9eM+j5
MW/9oj7uSJMYPiVywmvCK3TK6n6Ka+9TG3qQjUzstJtPdgQxNIR2JhRoi2YDQQgEXDdQQmWGf20K
1IHpmQwfEtmWQ9LvHyyneCwK/oTC1jATiPFMmQyfq5yZ9U0Jmgx7N0gV+bnFZyGEz1//txzN/0gG
ZpmKI6y5dG6Uc1xm8lxZ17R2GYyY6GtOKmWml2EcMX4NZ5RnvEy7ZBDRvbttYaq8K+0I8I1NH/f/
EiGu+zO3sSnVhPGnKnV8+RB+RsvewLIWv5pmRPevl+ZdkI71y8i9PRXX6RXqITNKkkuW+1qjNUNx
C3+IdGlgLlcrRPgwQpiFICdYBA+FW11d2tIgR4Agz42jgEjSGpFRWAcp+iKv2xmuVZauebY9qP0d
IlKoo2l/4C9EIrZOJ4w2K7zPghIuNQs9E+qHLciHp9/WCmSPcs1/elDM6hqlX8um5R2sYDlkwb8D
BxlDh2w+AKCYRO3+Z+GENsr2v05ycyp9/unWm8Pla66BnNNQMbLHEPNIQffZo1wUUccFdwCEPZEk
FamkpKmdaVlf1vaqw9F1DrauNlbC0sqWhf6NN1NHXzH3z++RZJRXyN5gMzmZTQH2L4ec+DfwybXD
SzhKsgZsGpLwGkMPjWV9vzvqkUTEptEVrWEvLgp+Ftb3v/MOSAOns5G5gVqy+qCGY9UKHIWQTZnM
pLnGnWF5+bZ1BpPaWozC3Ok5uW9wL5wrOYe5AE6qVw60Rhtrs72oaH+AvfziT6r0Wc0KTv0Opgo1
RSXa4qzqXAOnn+RMb8iT5iPpYp6wj/9NpO8g0pgHN7gmr45r/+oE23Cr8gT7rGTxL6T60pN22gA0
VgGhZDgm4oLmLM3vEMyPKH0bzgr5KXDA0bTm2vG3LYwdUvQJdBILqQprbP7AGnhF8M4CrXGGmyNe
AdTozablxAMgELLdORwOm9IiFB7C/hA/39BBoL7eGwnZDgB3Ywkor7Jp0Jvs7/g1Tdco/4VrZIQ8
hhKHsp+1kCPrX8R94L+awQakQ3ATuH8GKt0AZeZazc2PG65NM2kxTtUXmrS1UVKRAZNnonnBmDzm
+JQcu2pGp+CLijIE6RRmH2gKAht/EuCLzUf8RA79aH5ErFqkp3WQACcGzYd98T4XZUMStO3IcDhi
gpF46GRw4Ow5k+VzaGB7O1DikXJbSTcEEx0xLHb2KzmV7XgTS3KFrRfKgNDzYRniAZjIkrm13c8K
sLUWltEkv2tMIoHB5fI2fX6X6deicSN1ZQsBbaRkANjgcDF2gJ4LL2W202DKMmtlLhBpqPnt8me7
C+VBeJ3XsLqRYojeX/mUX2A4N5dO3j8eHJtSSFxrQTEG/9VZiITj/DQBI2f1p27QWCAtAVQzoDpE
oRa5d/Z9k7SWuthuBUgXxZ/qd0n0CO+hjIVGL7XUrrH4F2ryRDL3j9qmrV2vpyeCeMKurZv7JP7E
VOyD1+pas1EwVuwnCda5wSRzccsBTyNFXamPpf6A0o+Dkj0+MiivMFXKp/cPDgBkXGkOW/N41WXN
vACKldQMCwt5Q3fXLvq/tVfl242ir700jFQqUCg7BAp8ImHR2WiExuq5iLdESFDyqMTiYI+7c4rO
9ldT+QJofPC4Gz5bBbL3MTHcAyASMvCNRemBEAiPDWHLzXIhK9RSz77kIpsO47AAEFIOaEpGtWkr
5RX2zzWTITkl/V7r1w3V28ZhtffQ1pjpuD9x25p3R1tNHdsIdlJk9hFpj6EP1HHLdSjK9qC5kBHP
vsri78lzh0VXav3H9lDzz1+ypChsNJgLtqux1JQmVX2XiaoF9ukhkbzAvMcRSE/UlHUjF+jiz78E
1Ntu5fMhCvCUBfKktsxBcJM35HaHCk3BV+OP3OaL6d+Ahm8fpnnScKZgdMvaTNEP3y3pPJ6dYZNX
y0JUrJLTtL9/IeqjpcKg+EJMXahiDwb7xN+fBvJNuvqTlK6DShQ7pjSFSeKDhFuhOD9fKU0+bHrC
PomCdJ7gfYFi5zAl9mZu6sE2AEsG1Ifo4Km4zZm2QknDW6SjdZC/TjeZUtNvyeVHElN5/6PrzjlZ
kKI5PiPAk+zjPaisJ1Ql7eIJeiqCN3XF4CNsR/p4tmgKCOKEBddP5Lmpq2urfQz0a1ou+PwXgKZT
lCh8wPja7nAjy8IBKzFbElJ/peULJ6oNwarmE7fty7GGpN+mhjnwjlz7Ab/LWMsGUdRewZypHUGU
2ioMGr0fejuk19zTxC0f+B+WYGgFkqaSznKMN/aDw9DGvmbLmLnOqKEnal/KQiomEpyp1JED9eS6
o7utIbXcrZ/CqhMMx890IERZjFHM/zgPiM7IMMS0mUzAf+KZlxdX6DGFXyMwPS5ecjjUEizqZa89
4yEuJTjFpLIj55kLtGggcDaQIRYAjLi9pVEvfnUTPIaI7ofdNJHmtXnLTf9I0z/gSDB7WLWnI3Uy
li2YjCeLrlx6lZdGm/GzKmyJ0389SAi38/fBAC+9TJjvUZIwtqmgQz3R2Ch8/2rQ8apDr5PYEsUU
h29dDKogm4EStAKeZij5zlleVu8tKwyL+FwIQcEuR0azeZG5INDRNMi3nyj3xhFCPvIH7clYnXJM
OQHXT7ffpeUlVOy8a+dPqHb5IbOh6ADoXVk2gkgHV2ygKUXRuK7NY7T4ymH6WmfEFdH8Vw1MP5Uy
rPAztd5kCyZqDvZYAp6Pr0VBlBIZS1QD6Atug1/aZV851r/dAGaAsc09mNHdbqvfO5n+QEz6HkGs
+CtZIJgBsVWWqJkJRJLxZZ2keRnx09La5g50vSLRyNmeCSrd287NEJ4TqXVOLDmgbHHyX+Z+83GB
blZIgJGWgVjC+rskrLVKf0JLg9cSC3ZBoqqUkENndGARt9szup62k90fTBzof7a75Nk5kpdqAjHh
XTIwbrMAM37mujD5Qa8dqXGDZXtFbrQngvX3Sn+SY27NlCzbfDGVtIsqbD3zu8AzE8vWcN+3pHmp
tdaijrh4kT9Eryp0jAhENIAOPPPYw+/5x/hI+o53W3+byJuDGDxaUWviyyQn16sxMjRZuSXx6Z8Z
gKQKqpH2aM2Tswa6bz1IkWt9ywzguUqcJL5WDsRqn+WS+Hy52JD+g98xb15ovaCVW4KvRVHg1cnX
XiEOpuKvRiq3KF8LXosUIy7eVfM3Nf8+/VOfYQikWI5WnkbTA9L4OVCycTY4qWO4h9GUwzV0XtUo
bmJ5ZTDoH2Hx5c72dFSE0SHMxFnmPwuc2rUldDh0Ifnc1LeuAuPK9TPLNsQWrw8Ta7sz5zwA4711
cZcI2m+f/S0Z7w2re18o8hymquRxXVl1w9L5knyIMyrCWrFRsjtZ7jps170mZNJr1PjheqyJwezB
rYRqPEtmo9Y7M/9ZJh1DbJheiHzqhKUECgYAuIxD+uWPBpaZ46+aY7o08tJeCXL9HcIzMZ2L6+Ik
NkKa5tvJp3taF4H81mbPl680nUVopcb7Az8UnqtEgzDKPgsDgv7BRWdRb3wozpR9GQi9qVWuZ+TT
8D1f+7iGo0mH0YiLe4AbFBCRPVfO2VMX3MbbI07cedwmjyDiaCrygWYclS7ApxLmt0o+0Ryo9sz/
6QEj/tqav48gJ7ZA5sQjY+71hQhMpo4+Z7UtP7qrnvqzXcnZFy4OyOrV7zlnoDGJ+JB7ApfYE2iX
npSwz7kTuL23Lm+csigcAQrI/DlGrESOJ9WifUS2pIM8OKsosweAGXD693aTtCg/F31yQQU6q5Tl
0+bdI2RkQVtdBlKZ17JLG5Jj/w+zNJCaV4dOWygGlNrb4tvQLJuNjhDlWej7AEgVOOHRy+sDIwt3
m+cCzzgTBFhvG2jyRaCtnt8Aa9DjSk5H8Ftvi1lyw0vgvtcEtANgsaAPqQ4GUTmz/b8Q5SxQNIDd
BrJsAK3VHIMWHu8eH2lqZ9CmjphgRBY6B/2MHtz0pAbWus0ZsWKi+lKDpae5pDeplBAZW++23MIf
Ik+dVQ1Gx2d/hTh/WE8xjEcYMCIE1pGoFTpEQX0ZQynQau1ijV2HteyQa0gSX3b0rpChNICT4Y7h
qs60TMC+wRGK3X3habMwNrK6D6Leum1KgKTTWA9a1UWxwaSkTmAK+u7L6JPjm8FFAC0kcuY+Q8Pg
dajGt2fW7bE/1LmSBahU1dhfDbfpj2mYGmeiLiNBTIuYARs66GBS20EjaeUPQL6zXXhDpI4zvqdF
TP3TGpYzjtoVKqPm0r40arN5OD8S3YEj2uVDrHC4vgtSc3hmGPTx2DPzHvZy6p7IEvBGLhzQOyW6
VW3Gi/btL9U+km+BQ4sdhlbW5JTv3S8nxM7MSwKpX+6o5CWTOFSFW+zXtOv2WgVToCVYg8imvEJo
Ef/d6hLXEG1uvsN9NdNhMP+p4P5BJ/AzOV6nDk9zxNMbX18UpEtYlp2AKbVqfnx8K3rUQdtLKjS5
LkiyOP0K8Om9nQO3cMHVJEvgBdP2JjKFgirDth4FLk8QkQueF5u1WHdtGJDlN/vY/sFYz7NHKLWp
bV5Bra4dTJMO29dRLxqg2fpf5ZhHUSBXQaupYcALl/+9J8b2Fx2xYGS3YQ5rAjJgprolAwIQwBmO
axb++WHBSGIdGTmwKKKZGd1kPYBrpQ1Fyj0eqL5ycBaN0p6tzeLEPSM9LqsNwl96V5+0+5o/nsLi
c4aP707713ltJgwD7n9jtlg2yST7jVy2lSXZOdFGQPdm9WrgwfJbWMRmPb+Q1pp6Ud/M0QgJwTq4
v5+BVsnWtrqNOoKkqmeQs3GZC5wi+AmNmGUdRcaEcQxGSjP/PwfWsx/azEzl36wSdm3BxVtWYdbJ
DzuKFblXmmgmn69S5Gj97QuB37+QF3jsVcBytqc7f89X0zvQgNYftkBXp7lZBP+JUsI77bTle/jJ
ZRbPUIU8ks5i19B+LJ4/k1gyd7hEM6vviKqolbBWKc2AxYJ3n8Q3Vq5Oc9YCn/Lb2MDcINvNF7k+
3GIczveUIvCFrfw9LVKM4JCj9MX0aJ+x9NpQ7FsaLSbRhZret9Y7x1RTZy/BxBjdsHgYWENoHErL
PhlaqYgYoaGLhMNNgF4H3oZvp9fj8rPlkZushWz9B7shWC2drGykjX8WO7SX0ElUXErFGqBJMv9D
hMfLVl1Rz1JHbQEJLnWQF7khBYaI+z5mpEGUKB32qmbtlSk4cA6vevZnDdxxkP0rYwq6RKYspcDZ
DZzOn2FSbmgvmpYWw+nIXKmN2mpBIOQEJswv/uYV/ulQUjFBciXoGDcnmiw4slcuL+oPFoR96MHc
VNeaxLd4eULcLjLGmWG7zuYetIW1bqlG9GQ58G6d2IK51qBVTE1tq5d//+gGSeuiN0NjQMTomK+P
/aJVzMIpC8ig1/xwQlrmjBJiNGTdtEPkBTd3gtbSBhVWubE6RYdjJ5Qsu4vI1D6Lh3M8OCyFnkED
NDWRBigimF0JviyON0G/FDPSwY1iWAg4Y/vKdntutiU6Y+xJlJb+bClx8XKJJ7ltY/SIICR+J35B
kf50E7btLLIvyVdgjtuwz4cz72l33CxS/rus38sQzFuvbK98snXrPWfOE4dVRcJ+LM1ENNpG2WS2
wX/BrsDlnRtak5uTV63LxAErBVQd67tBZimiD/bZ/C7ma1OdxkukuEl2oGTF/M/Rnqq+zZTOsQ1B
ByuNHLHE3ILuN4WvHfJvMYHEoRvVfHZONdfIYb9KWZFF4DZF5SPPEhEZUGsCD12GQnqrawsZgsBo
CTL1od9oxwllbKdEUbPVGneqwsbrSZR5YrrRHpRxHR5tQ/bF2VFHR3W8vciuYStadbwN/FefIn8H
G/xDtzO7SKja6HqEq4QFKbgukKkQ90tzMFoBI2wsnnTMePVKPT4wfj3qh7kdeD+huL846t8p7Xcr
9FlmzagwJvrjx5f2JDq2FrBFwDmzrP522g4lJcq01M4Ngxny4G+mh5NKmLriRUzwH+tocH128hS4
+vCrP7wnHsntT9ZDKt4nX4dQVJsOMT1ueBnvLhbgwv2zxA+SQ+B0rwfqCLcFwSw2fsv/++pimdxR
1RG9Qcjx3tkAyr7KI/d7QxiJdLdtgj1IdNLwSuglQFWqfr6BjXIf+2+wVYD2oAAOa6NMwpzJwti7
1e+Unts+96FvTbJGdUpDTi/jZqrcgR12Wf4ke8o/pIhX6bfUjZkcR8XmTM5gweToDZGWKq1q+s5M
1EfA6utLFZ62eLfiu79TfESXBdY68MuPVkNEVaLRlFXdTgANDFrJqpzFXkyaHOt8hZIdGGbK4ufQ
mlFjV3ak0RIHV5Xe6BT3WnJOPmoBSpK3hghQb2EeC4T94mUdZMNYgfJhEgqFinytlCCg9+ZxOM9A
RTOkX9Sy2jtGN/QLo7RXBTMJ2d/aXX/ZAFan0ruriAgaIMIb5sXf1+XTnuhBqW63TnoPkHDrhxeT
oqIr8CWCsv6thcVtKRjkBtv0KgomWkRMDhIUdyBJjoJ+7SZnWT2RCIQkaIkgJXxnwioS2j8eAlVw
dm5idu18PhZCSM0kQImrZrniFOsV3OZbFemroHCuQ93P9ybPnx9WqZwJn2YMauD3wi74zLcd+ruo
tUve7Y87Ej+fyzLbcxAJ4W3GuuLwJiSp429Vik+jv7VZSIloR2DsnkSBtv7HWjfG7cZev1ByOUG2
eyvm9Z2cr6OEs81rz175M8wRPtM4hyieIMLnRJkGYDFVB5nra4Qqc+SeBXZYYpRgt4EArmS6OPh7
RlNEkpP2691Goe7nZWNUf7uKxg17X7DQX+L9/3TlZsjNekw1tl52ucJ1hZN69FsRuTLGnQpElF8p
ewMWsG/1a1pkQ6uNfowlLwcVkW/kiCkjsD01JoUM0YSjAP3tq6NZTb4zZLU8egJh6Qs2TjekiuT5
vEaVbWa1THk+pDiL8Yt2Phj9qNiq1/Odl1i8QHc0Dq9/pbFRMto5KT/lgVdfqEG69Ux5gzBzLGxN
MLJQF/2Rs0xg++ajZJh4VVlWzWjc9HqqAfsuh9ploqx2bU3TEmXKmXpyK3nPkfBQ3phqDX43jpVD
kjLmCGFfwtAhU3sLqfeQ2LyBaWDPx8+XtxMUSxNRtAasDGNQTf4zIlKAbGtTI9mv0vGXbYRfrtI/
ySKHwMK/2Fx03CAuQQwnK2SAoykX5yUppdhnm6MWwvHdbhBGU1d404R6CvPs5OFcuNgbC/dzKguh
PXm5jI1U0OrOFEJDKNHZ2jU17JAIcjlUJsUEaYmK8a2+PyLx36ffIqQQ+GHGAr6MQqK7A4D8VnEV
AmwQI+tabxSXWZvePKdvOeHGeqvUakD7vxiKSS0Rxk+psep99D7VlxojPVxFYDEuQrqeFSVRcrar
lRI5yJENFV4uCetNIkEagA/YXzjUHwrssnlQ1hLAaYFaFweko0GErCPLfSSZTjvKT2EEqFISSKOd
sKlqqlLU2vns070LAaI5qOhZLPgicXEssIxmVvHLtIbjji6PFcq1w+q7EDObJh+OujdY6O2n5ptC
PrrbWsAtpFqx4f5rbi83mPt1sS5IOczeCYgxXtlp8SI6sX9wHdrES+gTavjYqLbpmPo0z7cgVHlp
FJEL9V1AmQ/+hAwqi0GPwWPL6RQinTX81RuiH/k9nOZwfEcZ7njBzpGBMtUJdc/1zSfoRk5Yv0Ob
NCHwh+qBdkWRxnLlxwrutrG7Nor88imRlz0iG8pXmji+myCOh8plsG3QvLDz5y6Ex/0CKGZziKB3
/Klw0Vykxn6Is1iBoRn1LqYPiEAgn4v1hqu2JznqHmFaWLaAP67Fhm4kmANyTnfUrA4ugtFZFS3d
CrcH04+vNvgoD/+cDfR+1wcaLTxREx/J43q5F0si6ZL9yePE+SEbBqqVJzAxBAX9UL0ywMcTJNky
uImrPuhEUsik6RnbJOjBlo/x7AtIWr8f1w6OZoGMTcEDrZ0nwxIKqKPtL7ayQDsYJbmjeu84Y21L
IwFXd+MTyG+U48+3ppYneYkbCnM71q9/ja2IJgiRF56Rn0e9MMsxiRo2wYQu337vChyxMIZ7ASui
uDkeXVilRlvb8jf9UKLBIZxsP+tkRWm5hXneKmS3zT36XmO6/luFEpcumm+SGYBHVMZw+1B31V1x
itRBpXmtMshRVUSOBfJwPF1FSjLamYLLm92ynrxtNxgIJSBMZx2+/P1/mJfGTuqDlUiR/CW/g7fF
73DfzqOEWTW8mqSjFf+x0N2EwpjibDoonXCGLkPQeJyxO6OzFiexdcufiHwI5QzrpUZN94BYaXvH
NlYYpWtHUeNDolH0BryYyWfzdJD4u04Xs87MpVy2l+fgRFDJStY5Vd4ybeQOir8keAkdYgZwMn2A
0+FHRYLZ/F50s+orQh/eQOt6btNmeho58XN5uWS78Ce+fq8rxXfoQ+DtV2GF3Jj5h/qqhi1rH1+t
YbhIscCjVvoZMM2z5U1Ub7p5seQVBT3mrkQzXqnngMXt8uSo6pWNk5+pOs0G4nFYJCpgt14jq9QO
tEYICsO8aLExV8v6xgLk56N1ejle5XRyHv8vCs3nDN+72MQ29gZkTrIzpsLIlRgufg2j87S6dJTg
xwxdK/oEUZkvbUcXw0V+koZe+rZ+HELmyAsQG//R8mmnDToNUK31xkYbY5CBn0NoT90eEIGRp38E
/xLwGcDbSFnuTj9lfJLXZd2cs649Wzw0yVs4ljMBUCJCqrtkuSLlaGms7h/jqy6VEuv3XnulFN/p
5c4doWr/2Wdoomui/8gIVbPXy9ux0gQVRbBG35HCCLv/RQ0ACX1drHZWaVrAhnr26MSk5FxPnmKn
LW1coRxVzmImKuriDptTUzGpy8cZCwsBBVbCF+igyjCW4EjQol7qkcJ7GM5TM/CDG/5r2/qxfDnE
Zb6h7p8iuP4CMhMLDqlti4WfRv9ebmPcs2bnB7DSgXJ/p91sWGW5L+s1YRwNb3LBQq258OTzNLaP
HjRDFCggdXyHKBGILfRwM4/s7ziI/h2mQzmtWyUA16fgr5B+R3v7Wgc+JX/tUHAV9MPvlo9NhaZu
ed0W5+IZFx1CrzFyyP0zHuXs/ImACTA3aPm8v1mgSiHVxc6IYt4CZL+oqO7WcZhJYkdYgqGmOjhB
9numUXYfxyIgFIuytVT/EC3p1RM99QIMcDX7GjoeukStXKrjY3U6gm6ol69fYe4IqGBrm7bnw9Ph
lYM6FwknfWsnKlGNglieJqS+l2mc+Ncb8TIGdqZfjDPatTgPsbeKvOauaHSw8bWjaPAQXH60RhyV
eSEEW4z324DC3MVKZt/Z6n5omL041vCXlACTyTonetZaZK81C8F9w31lq5IS/LqRQR6dz6gJniE9
AY7tf9Rse3ogoKuJCCDt2I706q9uhrNgfTEcsS4spBr5w8QFAb5r3Nbb6gHhk3lLBsfT0uyX2RIK
bRv4ql7G+xE+pAcCpqJVdKgerq7lCGWhcZDc6pZ+2fYeywVVbgkP4bMnovoKn4kq4iFQsLK+Cw/J
CHb+cseMoFzq85PoxS1MIoyP4y6bnRghEBaRjyCGQvivy5QUvhm8S4O3ANCLHrtIvvsFA0VhSqO7
UUvZDPUoeMRsyluSpq92U05ukmuvwGgDxR/TXrQtcRImlai9YlU6LzqEb5W4exfnvjy/O62QFSyO
PeQImeqdvTuGlZxenkxRB/l6eceiNlNPKvblcs9Gv01t8EqdZ2LlTwulgxVzM25W0zJK6wk4RoES
qO5gvlsqCb7qMP+RPNYmtrvVLSbTz0FbmrCQdJ06k8UcUvzr1sGeMZk4IsNJbLAdemzSGt4HoQaY
Z2U0yOVZpzBkD6/mGKkU5SBhVGJ2eHOEmeldlRmQSsaD6co+XMHJf5IUAJIGIRQsshOvY78Q4lFG
Lit9mC3ptRTd8hK7NMyy1GEjkPBCedys2aVWWU/cLvHim0lWWN9KnwjqRxN0fT4uR5M0+AmA7bAB
1Bj3B40KBmJ9tBaS9dN3yV6BdTmQxvh3wwKe+eY/1nSBNOuYIeBzPFNvwmJ6XDA+o/LYRRUS9sxt
70QFCxZDmtU9+jtO/+cAxc+pkmtfGEsiJ//fBjhW0IpuVMftteysiCw9bSVyWCqEgJQOeWUQei06
DMBBDKwQXf8vVdji/YO7eCaBqkOzXL994haTp7ySK23e3mx9Lyp4uQQiXoXND8p82WZz1bUq+Iv6
fYGcEyZSFLS6RRSgrPjFQBERsYoaC/ofMCjmEpbbtw+uiwr7pd9Chwo8MSVwPKLQXpY2DWAXkQs8
UMXIcIt4BwFJS782kyvc51V1RFLUatXxovStVQpzRAGhJBLQUXJY1vm5405bn2lLD9P+HRdMYg3q
Q+dFhq75H5RZH1WLD2lkbszRnb8E+2JGJMpCdzsxkWzuQeYV8xTAuILtlty6JnD7LL49GowzutHJ
KCEfK0ZW46xO4AkmXNNzKgBNqzp6/j/26wor3bv2A79+S8GbUsL1O1i7tdYLTvAiq5r7kIzo3lPw
jHlaoq02xxhBq+5JJRzSghMRV8PR0rMXCBTse4UlfplIoCleaVBOVxrgAWuqtbC7hb3yN4vd9yYn
p3Lz5jpdR8MqkNsQlP8CzYmrksVOz1o9XS0MmfX0pjPL75PB85hu7vQifRdht7DskKfp3nousJ36
CNKpyUec0BlemDpkOMHPZBpJFh9LvPskivK6EOVK61EuGl92RvXS5jEtyhWS4BfevdkZK5KSmvya
GjmfKWFWzJIzFGltlRRhU9xeajDvjJxhmdETMkJRyuWIGIzptY46kSGwFJylct2vnvNvNdgIoN87
J20WklCSlmOSXT4XV2fBkCr0m2URPJ7h6x8DZfLP/U0ay27Lb62ovqctpkxqbAuugCwVeUGfNx5n
nYOp6Qqlybuq6hYGxWlAawUzyPe4diYvHxxMG7OHBt9qs+qjR3MvHqDlxOkf8IOkpDatVw+jFLVE
cqLo7YDB+03hOK6ZZgEzwPFc5EgQTs8gbuPXyMC5BUzWkDQ+Lfeh4qahpqhRyGyyqfCzaaoxNFDO
A1C6rRZY67RjjsVQwtiee+G9bsqFjxid7zUOuj2dFBveejXe75IfparKk94En9FO96kXFOKLY8vl
d/rFQ/stOM1laZApNhEVER8hunzpaiUAKyZZmunLRsnLyt70Rwq0NQNTy8VovIV15mxGE1GXPl41
Bs0NkrV4uNvJEyMLA8dTYNL+LDHbDjzeyCh7E12YHuds/Pk0QGFp9K1fYoUZHRJA+tlrIWLbJyha
eeFVruorMvhZOtF0q5rkYDEK7UWY66S5sN1nk7xY32oltX0SAIu3ZjOoNAQ9fkmLzdrvY7G13Qov
Ib78wxPDUGAy8NwqEqi+3Qp6iGnBpOaF75VzuCwHFkTH3OdKsERaiBSdle4VUGWdVC18S4xaZxb6
eYNrvNeEmN/21hmOdbqfIWDuzYv+TVGEhJ2tPAr7dy+FY+1gOwPaGIBIiwOihbze5e+guaHoKwZL
di+EVbdfZIeCk54IFhP6OH442oN4lITIabZASKuWMVjeVy5drNUFQCPEegEkqCK8lS9HUcbBQWOC
Zo7cmZMVQ+rkSlmtGb3CSVU9Tr9LD4OdzOt5YQ4avP0yuV6m12sbNwDHR3eTvzdkc1jma2+yFfN0
vonbLS4huQavb6kpPz2xi64wp5JhUZiYKEppUb2Hm1kCGf4MYtj3t+e3gyAJ/warvgarJzxI2ySD
lEWSlNhcJaXUQEHTXcxoZJvKugl4PoUEt2uZ9KtbqPTqcZMbYt04Z9cvPJxip44PPoPu5u+OFJ3h
gD/t9KXB5kamnEG49S9wNRnSbg5bqm8v9g8guhcjSYNGpt9SfTWZ5ZQ3WIQLKkRkQvhvo5mv+/T7
8qLLbMDKIhoMi+LN6l26BMccgGPX24T4MsGR98CxSpYZfTW84zZdb3gZPuYq/qrbbR3JpIGPJ1ZK
4jfLMYVD6PK9AyrH41ys/8CyqUrUzRSlALD5dhz5ODtPRyJTXE4ywjIKZF5V25UBRhh693I41tta
YCv4i/bAKKHv61iKf8DnCOkPJolYj//R9vdw7bK3DaCUCP4STyx0XyutPT70O8AERGBCVlwl/rJa
EZggUSAV5nYlc9C8qDAJBOEliKyimLNimo/ukPSKTeAnkfj74wY3C7+MtcSX4g2fzwckM66+PHZL
uPQ3uEx1DbQbeWn64Q4kZwCCmxM3f9cpiDv3v/+z3TGC2PDE/3rponuC61LDr8cEBf67zXlCBI0N
i9vz0Iv1sTpLRF3YEWz8dVh2Vd5XoY9kP/C8xU6SultcYR4l7vX9PRYZWDqWqkErDrobq1nsxTWn
6ShlFJnXxztxMzLvGYIpgSLmFrMbQmgxxXfGK3SPO2EPO0uecnsMUhzHvTKqZXLzUx/9qtGMCICK
08QsWZv9/Id6W71d0+UxMTo5+YhfEqdpnDxr5ceMlAbWGZCB4s923oO06CPmo/DProEeGpXZJLGE
VaU0Z/0kZQ/y838DD7VQt+g833Hl/Sddi1Kx+C0Zp4kvTOvf2AHkf7KYPiKOGgRbB5Hahq96r2tb
Y9xIOc5fKfrLv5OgJklLSAF0uALr2vL4fL8qo6o10arRM5YxY/AOmVAGEDgPEftTZXZwTqt1Rfib
4UG6sHQFpl04FUqIwm6rinnexwW8mW7ezh76RvcGCazO6QL94zF3L2ypa8hjd8opdqL/XaiaTTDu
3p49wkM084O8LRT8esy2MdEgIna/7MRpSLafZTpjkO7vN72z4vDpC7zDZfgSlzhl8nFdXcoE1toF
KXUJgUzCxIa6QzWSKg6xcMNopHujvNNzeNRvGbzuUQNyv5mwJaV1VHypHtmrCgm1PHc6SGGIvujD
Z7+65JqWa+VVKG7ViJBh3/mZDcORL3R/Ehc0K6O0Nd/kxQu27jvh4YLtxuzN6Ld+m1i2ss7P3Oft
hys35VPPQFIphb0UExTZUdWMQVy9hpBQKksgx9AqE1SVnWgBVHENEn6oyO+dXP5lPjbWfl6YXqNN
XxYZasu03RxHxdX3lRK+8dxE+V5spRq8PpQLMpfyb78HECGjWGXZMrpPUQhLQ5rQmCGMVROPm4bH
s5gp48EtaJ4z2W/CmcDZ335K9WaW3PvLW3KJtzcZaZ1zgICcPYmtIjuDcbIbK+EHhuGaGt99OAp6
ZEzM4EJLzu/dRlRiLUalbojMtHXASEF/Moy4NWdtu88ciRSGpSG9oMmVVX8pAIjUkpEXD0AvbsCC
Z0ZhFoloICU2n8osuR6GmTooz6Z4eKIC3xbDnpV31tU3/bz9/pvtnjH2o2hk6kRMygj56JL2NbWg
YBQYNdATQ2rg1IuFC7Uu4gccrf6RVFiEuKF8yniYcbe0prmKQixHKR4VNZBR7h4m/Ha4ZSEN+LWm
4Cz7BN7FLbq6V6MgcPGj48XIA2TtJ9XbmjrAx9vCArpxR6MDAwbjpOneGT2/MYSZwo3xisw4t3RJ
uUQq8r4FX0Z5QU0Wr4SliJXyKizmD2RO/bdx9USKcvRoK2yTXpk8VOO0OYIkhsf4M6aY4A0tZs8+
oPQlsPg9Ta8PJybEZuqSVEXtIHfqu26E6mB8kS+A1379w8rxm4sCrqsGq3gTxkdMih0Nkn5qjm6A
LDJwa+3lcBYnxbkcGmqqLpn2oBAv0qQnwZYOj9SMg5kcJS36av7+7S/BpicBIrsqKD0lCAF3NIG5
gE5L/MsK3AFZETw275tL2LWY2wOxW+q2smgIXGhSJFsyOU+lOCIyTrjirAja787UQpbQCzFUdwGI
HiMhduTHj38tdwGaFZFtuOgE9z7vXmWHOyID0JHbqZKyvD66TBnuNdA0Lz9+hdqvG6tjZqpkRvRW
oEJhCr7Vo4zYu7w7vrxeBzfpq0Q1BLwlOeCjmvmUvkrunb6trJwWh+zolSCn69UBOC39JbzHAiBl
ibSMPYl8xK7BZ8vKyKd1I6YXxYu9ksBvhWAR2EcDfE5tYOGWLZ+GNNBuGQo3XTxuOmktojExokxU
51lbXNR7ITr+6f1rZEkdJKPX7kKpLSZMe4ckJpHIK473ecBECIoxf6KxMrZ971wrGtK3W0pq5M2x
KsUD0z0hgmT2uVrAjpzFwQ9nCFYrAGgYj6cz2cpml4hOAXynaYLcqkImoBBAf07GYJIWTcHdXOds
7p3qZIcHGhndBMov1jSbfWB54DHMuiAqtYr0zqx8y8kcElJL5ZUv7FIONtsQj221l6CYYPU5Ly45
Rs30vxhoI3FotQDzViCKmjzQAU9FOQ2dSEmgmSXcOSbNfbmDt0yuQnS1N0MrjPj7X0z0DPJP4hl3
cW1y++Wbb1NnmDOMFDS4Su6RrOeyg+B4nM/sqHQKnCuL4yZeEilOQRpat9v6GST49o2x3XXiPU3S
QxtqbbG0p4df/kUyBshY5Dk+G/Zb6SwJW63k1ARHqDn2XHP3X366mm5im/bgQD8n3416pwMBFrup
mGU+QYDFimUA7taTDfi+LtbJrn0Xd/VQxfKR0eRqQwLezDA+mghWXkclYeqcrGqDx2frjfyTtIRj
iBqlwa8oscvVBwqLAwjWO77FlkpFutua5ZjzxN9pnor2h5zHXstLrY9w+xOMIyxvOHAaIMbx4+gb
mVhMOvirwboIjSuvbzBRKQY1HR0aYbHZl6QVSoAYEr/3T5vry2gLkcDAkzjnT6PDn8o0dWlD7GJx
KstNM5dAoODsBysbrZSJqNIvTVwjVLUIRKDFuZ6RO4TVsNAbaXYpUD1OkF7gmfLWbgdeiHntlOBS
daF4XRojIRz3z/Cur73ADSGamRHl6afgiZZv3GAnbqeiCtcE/oKT/i6n+A/KILH2GRSFRwYEMBjT
ZIsl6IDo6WuoEAm19WX/AZ8rzYYSLmGXiI52bdwJnj7HWjCKRpzVWU289BZA26YCNpGPDo6KTiwg
JAiYAmA1k5cooHHr2XeDQaRR/L9MM9WXTesb/fAQ+vmJsiVRQCmbn6lXgSGZ2TfjeOiN+Hd+iPqk
sfU5++LX8JU0S0bAU7IR0Yz9tKALgRbu9Ma4A4p8A1WCmczYLd22F4sgRT7bIAT3ZbRpP106Oxrk
6cekif4YjNV6nioIw5SkOmC39t79Z4S4qb72nnTFb74BEx6HEer2WH2tET4Sj8+Xf00Biqqo/96Q
qRIPZ41n0cNT6WcgtKwpfo5GU/YuGXO/HgwkLzuV8a5P4EIUVeoXxlrAWSlAfHweh7TF0oBPzfjF
WxDm1HhpFgD68F1vRIBIs57pluSJW5QRTOWSUyC54MyFX2IjcjRCCWbaCmP5gVpYBqPmeTRN2oxq
fN/jd//ZRWpd1WaH+VdmknEBi9dv7z6RaqcCCpHdvJSnjgxQbKwiAmiATFt3mZRNkmdymnYTQPHL
iC9030P/x1L/MbkTSpDEA0p6NdHqcPF5to2L8oRKQcO53QCuG+DhWSKbfi2+GMr/VWNmvLNVcJ6U
/aw15F7U31rQYlIWrRVvX2aj/S6PvwwOOLPVqLxQ7/a6UyuXEZvElSp5tye4ymh8OJdTztp+BDqN
0NQxiq2mT4dvrSK50vk7DzABsokGQKjG/7lpYzQHIL06orpOpcUyKoYF1lhiIJdqs6gf8HjLqh6o
WAVIgxPS28yglFtThxcbI5/OHvc+p2TOiw2/PjOlbm3sMeRiv9J4dTaugZtzY6/LponIUSaxaq1g
SEH2PQFvlrFDHBq9zEw3mHwf+W8hY2A0b1d6P3B8ZbR0bnhuxXgqcAnPzfL/uCYNgxL7tKVKO8Da
eYY36tPg4KfWbVf2htPB9PKcz6QGd06throZoKeTFKQeRLN5VrsxU8InqzH8DD/zJ5DzHlATVLWf
Kq04NjW66O2a/mSKhbPV2LodmZsV89qHHWlZcmhwS6zNFJWaDlclzRmFi1MlDe+I22dZ2IwACrxb
Lak8xVyZLhhxnrc+SXGbOwy4tZrnf98QXQe48jOSh9L9jkXOuA8FSFCpBnJYW0qvWhTe0sc8oyKt
G79FhXD6U//Eb8hXZODxtAboxsAtjTwqpdZXSa3FUX86fOIBKB1Wt7ydExu8QdQdCSay2leD+bdH
5q9jc7cH5g/bjeB1khXZoXRxOP6U5JU/W+2PKLG5qegoSLEmS4mV7Zg6e7BC2gKad+SClgV8rPci
pA8PbkBAMj0dsJ6JOUZFgWM+zNvUwzCtvltstN0V/lleSuo89E3Tq2uV62FEcPyDn1dikWJkNlRJ
jFYUFm/YAhlVqdEbtXUtrm1/YG9/RoDeA5X/V3jw48ZuSsC9Ygd3IIU1ymF9WNhqgXzQimF9Mu0S
aWIChsjRlew2vx9e9BIrj94Gntq5lE4PKuzPcIjdoYuMqVrR5C1K8k/5BwKBURl5UepK1hAEsiB2
/eFnUfj5NBSmvOC3UooyP75WBM2ZKPQEz+x/VNC58L4f6PLgrx025mYmJiDIMiinZSFfokeJ1fOq
7bRVBIoP3kGo/qnUo6HTGXAVYyrOHsXzLBErItc9Tunqwl8YC7hM+pO69PaDXNVN0PG+a4rY1LE3
C8cpakgg5ZNqD1BP4e/mm1wyxsHQca75K0v5QLFQ9m950O/rXUqBbGV9W/vb2CtdIZ2itNubnjCX
4KEc5Jv9rS+oeutf3RZ/5cdVsFUoaou7Xa9UCzJAw71CpiJoyRIN4cnlR24RUWJ7b8a6ALtrlhhu
3+8pzAVpD7Qlf4eHk+F454EJQMv4j/RIfDau9e6Q7y5Qc7rbZZhP/GLbLCtVr3SFb/d/9v0klR2J
8wWzUX10T4lmvpw7X8drEW7pHxHhG90MYiVFXNjhcnLvYcv2kE61Z7rL3LJASuYOAWP25vbpl5Uc
I3n0TH2EV9feXu604VVdMJ57XFCgNJjU0ksBj6lt1v3ZRGHpOJ1g0BeM4yyVXL3QTivLgo30wqnp
N62Ehhyzh3rYHyA5Qo0BKH7uA5NQd/w1gpk/ppVdPay8zLEB0+f8dN0dmDcvZhakE+G/9/OdBsLR
Q7/Esf0rLJbG7W3ZN9ZeFGCqdyTJHW1A48eOWrLv58W+N8nKjVY2uw+xz2JMcsyGKnjhXiY7FFQE
ZK3VBVRVjZwM9mz7o3sIxCvwAze0irqWdr6N1XeFjbu4nlvPqJpKGQ33WbR/JBJJ7CUJHEM5j5zj
hyJFYJ+Ukgnx+5g6wPa11cTeRRB8mPTMDH0iZ3oLkllEisBo/O7silW0oxQuFnlRiVkdsMr4DyIE
kSnffwBCA8INj8/HlUz5JR4PWVABcHUoe7ihCLfo2sBInRT7IJpDoxQssfe4rl2iLWaWq8b/gNtH
9XKl5L8u7Ir4sBjN0Lfux3XccekW/EDiKalbmiLqMzCoeRSLSwRmyiOlb3L7WGZl87gCCRUrDBqS
5szt4EfFZG7jY61x/FKOCkNkpuV0zHhkUwQsK2FoQ/f+POXHDl5uz0+SQV6WLJfM+VlYp8pp99Pe
zCn/bZfeWxDSzHX/4fmRZYhw65nA9qXGyn7M4dijXB1QNpE5Za+nCcfNwDEF3OLoX2ElSOmmYmLe
rUCdoVr0aQkrf3bqtWkBb3dK097G/DlhUmE9rEDGNFASVl9JDG6mLK2Rl8ApOcIXMvMU6+qxW8wK
Iw4l5TampqyxQskpFlyDkgbOgbeyXOBDzLjn0sd0z/kb7lYyx76fpjAiJ0HbmBV/GOA6DfGmHVNO
hF5lxr58TJgZZnqSlFA1nDvY7r8lWqrtBgdTsi5EZAvXSvMnWW2AeizEASKe5yWJexuQkZAFZJBq
DO/UkpRlIpRdUYVCX0lvLrEcnuQCSJExDRAEBeBhBRNYVyc2z1By9oR4zl5aLf8M8IUA6T1EOwDP
XzWu5hpBsRnQuRiJWv2CaLAR9/FrXe3itQik4HhJu/9rpvQb/SPCZHri8MzdvuMDvYpvd82DsEUa
xs/nUt3Zv96vnta8CM421Haid1QIlKVL39f8xeHRxQWM81R1Dn/F9JynlcvwjEv9UanEzs3e5jRf
5hgIMHFXLeCi2rjT/b9EgsVENASdrOd8liRw20bsLHkMIpsYOh8wwDOTPc9NItWZF/E5xwWljyix
I2Wl/hiUiIKAIzuckQAcqkhsL7hJKMfwG64Urgxz0UqJ8BLfptW5972qP0DNMOluSLLydPba5f9p
WWJRNW988OWbHUlQR+cBO1fEod9WnnQ2NY3eJEkQ0poplfFaf2T3ZLjPUwu0m0DAdQY1NzVvYWJq
IfogUGx1Mgqs+ZwDbNK56We2zuL0zyEryuwI8f+9641amJ0YWRhYvnJRxkvMeqywL7ExEfTLHQ5t
DqfOFxWX2LUVCqUlGr5Jh29T4ppxg0mJi70/dq51Yqw43wryry6wUXftKGh7yuOwJ7d6lEJqWgMF
rBsjd4i/991HWPQeid6r/HCl/frzBWNH4n3KQgWjRWqxJB/YT/ZUU73lxKq+MyZROz7BZmRlqWts
6NnO+NeLDdYZTl3pDLjh3s/8lvx6MxEOQxl+8bXJpA5lZ/s64nvBoQ/6ov99tVrpaQ8X9f1Z5fF8
PkVhSlF56z1Kn6qYTOYaqbfuzsVvIOWjhf77sZkMFCR4yyI3xqGTBiBGTSobxOVEpj53TJCWvcLj
gdzxIL2gGcht6Zw64voESoUHaECnFtEa6Z0+tNLM+6HLGyWSvBnBZTpRCQvm41YMPiFRmYEnE9em
YtqZgBRUNdZDARDzgvP0qId2U0nRXrc1b3bjwu0tBDcBHjxClngCchWa0FJ3YYdbwAKSA7aCIwDp
dij4UEHYU59lX67Q9yh8S9lzw2z+kKJeae2MqrQdZet74KrK90Mknj38GLANKCl9yXH+WhiwgbDh
oPqLwkxTogTpLwGWlQ5ksLhBi47wg4s6OACyiLwMKNN0Ogl//F8UN/bVBpVvH5Z1D4Hg5Tgu8eQO
myH11gW9MQOtus2layduNeD/WI0G/Y04CqAemv4OXK5c6GecZy1LGSyj3qOmV/WIGI7ZzOh6Fe2c
MCn4eAu5Lf6fs/Jq5wuH4SdNDoUuBULyDlY92gqsDTM+wFqetKK58aQ2c19QUJw9zQmvxrDZVo0g
HJc3DHSpZQx1ieWC2oge6PxaUHSQ7toaw6St9U8RVlh7Q5ucv1Ih6URrpP2wBsSWWiE6F2oFv/Ym
wgXQAmtNLBKU9YnOkjX3+kfLbc75dh4HYiC9IATHjEImTysGJEzz7UYmtg+cEaXtE+OLZ/NaLnW6
cAyRsUmjWl9zvxletcedXym8SGmn6yPmEl1v1A/q+xnovXFSe1aXBoMwhGiLmCqOoWTBNKPtkqxK
dyR449kQAoBxkCAlVEXudwZL//qd7N+7J2N3HhGGPXh6nH0ffDejB3S9uhbfKR8L15FTt/8SWHQs
Di1idjypt9bM92EwKICFBMhs3UEBIplYtiQNXBre8gF9V9Tj1w5G2w7JKJf6mVFqb+lPBgf9hbFq
r2J2PQyp+Mf7KHVh7MAcJQW/jCdkeDYVcRstAPf0FV1pAc9c8SWZRwO7KpkLBuUpUcZA15EUFwVq
4b7fP6uIbi8eg/tRbi7aZkTvoJ223vUD80n4BxqXmig9GUxYYicIkEo7rwa6fE7jmn0t/ge6N4+z
MJ+60ZD+WenNxUxF6+gVDgY3cN99qdN70t+iLiSq+Z86x7qvpBRPNrKAoIwQV7mkerv9Exc7maG1
DPaKJPQkEM3M9M1u0RqMOEX+DUwOHVwhkhnMA2Mfh7uWEIPyaCyBwBk2f2hJeXinyWvAID8/TSxN
BpOyga0uXWJdnznDc1ft/FLKxVHCYEvlAnTthcDrV9/T6+bEY0Yi+QuV0Gtv0XY4p1fSqxQCyKfv
iBVGx2aeCSswij0OfSBp8iHjLprcogYTJgY3C9E7VHVbUw5YwCzYpA6HeVUvAP8NgYkQKmi8POF0
gt9wEyBLZpnKE8J+c+IPWqPioaTHLjj186pJCZr9nO4udcdon5CdljFWG7gBv13lm8QtCPloyyQb
tQ+bjrTudKFRpC5A2rR+VMRmBkSNZVG6P6sdDgaAl3bvKLbcXl7MVUvCB7M02L6MejTg8ffe7Wbz
7ZwsXkwsFybTj1m+2SMhwN0CftTAC38OsUMIGlPDVcxb+HyvFZuNpygnZLuT6Yq/M9r7S83njrn1
QOJ3WljETvcIatQ+Wc6PyieMUC7FYBkRjTyhPBZN+IM7zs40aGEw0YNIytoQyfyaBZkl9pWi10j6
eCHLOqvTvgIFB6p+D5bE/MesYFTUNSNAN0HFCO4CQH75D8QzI66da5TdAnTtEKqIuuR0tvDRY9FF
gDTnQicgXZdCB5EVRob4eLuP8LcB9n51plW/4fu8Q0yf5fWgczTkBxoW469+bG1XPPs76XwM7kzf
0eDgilNu2oIcpGrR54LqcoN3p5xR/v0Nzhbux50fmgo34ZstKNEn4sWfez7MOxGBl9Fa5G9FLf4H
hMbsLQji5a6g9ZE/r/ifgQ3Bkp+y7whjBZT6+ggx/af20uPnp4GmxD/Glp9d+SqVPX1XdR2qql3f
AYNeG0VeHiuN3a964AlA5QJXoTKgoveVqafg+lZNzo4yaVukU+BfkSKPryrq1aLz8P5Qw9KbxF2f
ZnZvgj2gzQFcaLg7ERl+hPHRYArbEUJ7wFmWlFJZhit2J0UNF+6TjZcoYaQWqh2RJhsL1OhRkqq2
E30ZBmBlAO83k6wEJHOJETSpyI9GBEv1E49P19pCoonSVIQrlotA4X5ea0F9dhqY0UhFM5gTprf1
XDgh6uoivGd4JP8u/tbSX4jSzCX4Q2kZKp6t7wBzv2McEbECC5GJudyuikEUEY0dvgCy0fAq5Czk
aykKLBZWHz4M3BcSvJcJRCfGQb7hDLr28QkVOkH3NLOq8eWR35HefTWKpGzug8aq4v7f9eyfQGaJ
XacuzXBqWmN0j3OP4qrdbaE5mg6QzybZs1FIH6orjPBza1bG5j0K06e9KPmQGFsammBOt5QoJA2+
iutGG6MeCjSWx0IJKMY3CgpnQCfBVDeN1Tud1iJaaFI6um0NoAKx4wKky4muxC2FifObaCTr7qb+
8LMazULgKkQRWq7K3w4vUrS75daj8WIhFSrLafAv2DDIUaIiVwVIv/yooXTpmEDJb6QcSOCtnTEK
ZCwsO2tl8M9nyiSgAfmK/LMAIdSHepzOoShbmj12RiDfwPW6XFyzWTx+l+nH57fomEqm+sN+T0+D
v9Q5eCP0YwaW7OhDzbPgKNIj9YQ5UMGA8+lDr3Fe34nObvuJbxge/qyiUS4L/JO4SOjyrFfoOG+7
rChVyG7IxHwtRPpGhv9zql/kpPB7rVE1HIpIpASknh1q+SmKT3jAN40+BwUluqZBB1Xtk554Dw8b
ncoMMmIEb6WiQJNO4Lk2LUkroLnO+u4NK0Sg95U9LXmHvOGSE+RqEmxCTBR4VBTtRYhRjehpDSV3
P4NZRpLFbcl3Mi9y7+RJ6qp14Jj2RIOtm3i3wQOmdW1356OKPs7oNLdaBhgL6903Kma6FHYKyYwM
ZTJ+ofk9xfVDC4e7JWo98cRmLsvMSngJK0qBFSWE8N7/WQj1SF40eb0WEZJUoupqEmYDfHfQFRZz
elH92wwlM5Lh0Fs5iRoBCSpwhdOurdDIG5nGSpkRF6G1ZAHmDzP7U7Iu9PGvaB009DzBh2ZtYdQn
FYfNhg3yiv4+dY2kv9TbSDYMxxbwxkJCTFpPg29u0mdJy74PZkes5mdTTggQXtyj8KxkRlj1/3zi
IvxPJI4BYAJ8CpXQQbs8ecNNJWP+gge9zy4F3C6vMJQqZVxv/qh2iiaKfe8/nMUjUcsUrSwFIzqg
JFH9bylPEBeBXlCKFRqGsnBu0IBOK1FBNqbn9o2NEw8wA9HRGL4b8kJODs50deRfJrqhij2r1zfp
1QNcXJbux4fMyHn+VqGK+Z5YlfSISVlwxHQK2EEuVq2k1j6u6Vp8gIPbnYHpv8q1TAxkT5f00uco
be7bgJYnTnq6zfEliguU8sRUUHmXcTUBIO6Get9pMB+qF1kqhbjOUhpAaJ3DUdz0WvLKOpj7kfBd
UY5BZZO3m9Cdn9pfNHxlAQgxd5wHi94w+gFKUg1jrI41sa2Fwj7260ycGWCOlZLXN0aiJ25i2mZs
3is3UC7cAN23W5qB3qIEY4LBdmQB3bS2Z+RhW2hYysZ/SDSydm2wD9X9+e64DcIHMm/6TN9SlqjH
Ek5pxH7F4J1QCkzEnsNNPX9CZwG9uJNU4ms+O5no9YPRHctjbWtxR5tBRLokkz+IAhl6/rywals8
eHYfB3buKzh9R7grNSgjGtV7oMkdZrCKpSnGgxIDPwK3TIcBrETVm3Xs9WtmL4lPpxb7TGae8do+
T+HPa5RMjtR5z6TYcT3FrX9GZEWVpGpz7DVTYsF4j3Fl494H7zrAW5y+i6jXFzGfooFoO+eaIio/
GJsv3Y8P86aCIeaR5S9fgZxGo2ERVWRAFYNXvYuE+t+HAwTe/C+JouI6XkLAyik0dLUED5VhzImO
NzulQFTiIldv1twlFePvUdNSKhUgc4sPd8UL5hv6n2iJNvIj7yI7OYln4V/87fhfsSRjXFw4xI1P
Pv32pzcOH9uW2kHzpg0W12EmnCD3EKqAruHJ6ajHj7Kv9UShRjZCdzpAAg0PtQkw6Ls22trbl94d
GTawKPEAdbDQZ2oSF9lKijJS74/69w7nGXAkQYnJXYcfQg82v6GN/EfRL1KBhohY6Hztnv+f9K0c
A8SO4yZ/DvSGvB33fu4iDV+sg75FviSnFt2BvUsk/JCfKczbNSjp7iNEgVkcGRx8wNAJbtBhe0v6
u3XUwnuCrTqD3cMAWocfAmMuMDDp3JCfnaLMNy+Rl35MGvo39FEmOAV9hGBUUpCpdG/mrZh+Xpyy
JHtBOjEyzHMtoRwj4SzNMdyXW3lmw24OneegT1by50Xm9S/QCrffbpCHYGdzYU/IcnTG5S1QDm64
ZhBoxSwy/ZxJLTGDJAeFJBf579+tz/gelEg5/h7bmtEbIsikk4ZDxtavwgE0JeAaNHUpTb58h072
s/i0hy2T2KA2tmmdVsyw/O8ulf09xSGdWnRuiW4pVgRf042HqLyEsAM1vcoHtmHp8rGRFI7e+UEg
GcWxmAXCYGFJ7eQSIlObeGRlDDW5OMNdCGz/nC3whvjO/ceTVvWnBW/u6Ms9rdGcYippup+vqYaL
p+Q5DZW1AtYn2e5cJk7ejwAQkmX0MXB49bb+FYbMXSo49nPhddwszyaFZUa8UHUQ80blvXTsU5un
dmKPmzWulQoJ1u7pa2zz118Jgf6YVlnEE+BrxpcPlzzXk9Q1d+5rxlL9EcoCuO7B5Fd3Hb0F9gsU
w0DMWPt58TEER28xWyzgGbDmgG+H8cmqqRwdUzjq8GbSCYCA7sPMY448m7HyMTBsr9+GgB895Eiv
g4fL5TS0qlK+YCCnwEqf5806hx4b24aNpTWbjYSomla0khetT5QW5zgwVw41e4MoQYwTzU0WrSGG
XKmx2ipbUFEVEzq/FgnHoQSIsFyinwGU7lnVdlgdT1Q8cmJpHG3UDOZIiiW1iC3Ak6gbyGxZxc9D
IP4dQbZp+qatLqx+EvJ/jsGRs3JjK+HPk3w9kw2cBWKLjcfzgJ4YR++vTG1/hlUupefq/Pprodlm
bAvOQdHewYJ9s4c5I5kiiOPy0VX6cNIAYyiUp6QgvrObAxBGM5FzEjppL71raQ/l6+ngkayBL5D5
P1tjVBBhGn0UU9HrmcegEMfZx9zKnnvRUmIpIuysq2rU+qJUksrgwLiXIWcigCcen3sh2+gL3Oh0
icwTv6mSpsm/9avRjuyVf1FOfBkW3SXKV3sr9eiFdDIfbZWEbu+EvixV5kbgv4WAcOgqv2UhcePN
6lRHzcKuHeozizlBlwR6bUKlGEeroBwUA2VU8o0f7Kpm4u7qKTkPxztouomV1XbsUv0lJ2F4MGMb
HGVhVLl7Gp78PMzTi33s0tEnV0g0zZV9bLn/s94/S2d5hbTTxv7jBHxnNrXRyo8nJXNkMxsxKvhn
zTFgA0sVLQBfb/8p4k+oMs6gSfnwMqqOhmViWmjUMoK6v7xdQdT8HnGbPM9I6lU5V4HUg8QIfNwb
FYsATsl2tfB97a//mghsjARg7J8yhpWcmw7yKcs92VkIkYUlvUXaiu7M3r4WrZ0OK4A6PlWrh0pJ
8lD6wks9pzWYsvEbNKf6xbulgXaTcrpYKSlA4vV6d9wRzj25XMuhG2EPhH/n5y+B3wYCM5lI5eGl
7fqLadO1LS8R8wQt7KcLgB4RgMfMEGNTRZdoDkMYzrxwqp59LwUjdu6nEGS/cc+BU4ZRBD9RFaEN
tAl3nqTG3/JypX8eQxGS6/L+++oNpx+R6BrAfzqg3nsfydMPlj7xVYOI8DZNeaucb5d1TUE+9xJr
eHBkl8K+r6qoNuU25UeUovb8tTcPUF2QYWTRGkv863xtadzBruMmxkMJHBrgWPEzyol30OV526Rm
kGKJtMrK8y6lORsRjxYIPt4iXR2Fwao1ewkCNOpsCFhq9FiUJ2F5kx4yFH7N6SvzdcM37ti16g2h
tK3/opF5hYIA0ThiykSq0iZbKP08jYxCRSdERY5A2pun7akKmQ03QbziXDgEqAuscGFy8DfjHyIX
VmqN17wswKza7Qn2mnXY4bK5z/WntfGLUTO9Y3DHsco00/XQX9VKhnHAvjMuJaU7aKx4/uIYULXD
Qwk+ILHRM8yVhMty+sPAEwZ8X4fOUODFG3VF52ob/EnZ8XjRBM1U/0iBl0bWMpSVOO6iC69tYh6N
pHxnjzsm+lqLrcg8HZP4yjIMg7VS7b0vPwRU3O24l15JKCG0Mo9UCXaoZCwqLo7jl2YXfqGUh5ke
Ao5/05d9ZHpxBF3ZiFXvlcZx4Ez9OwedIbBGRTEz5cvcpbntgBC8qnUNdoFE/3JzHIS4VDIfbA0R
o+ZXFknMRsHA+5EIcu8aPH4l40MU/9rrrIJLsdJJARY/erwNBwSeKm30rBPS75kNyB17j8ZB3Sb/
x1VrVUBflOTUZWu3dIFWLzbvMnCZrEwTwhrsGmHHekQiy+uybp3ezo53UIf5vMPvgyyRn0AtB1Va
41oABqXkZhvLUdDP97lA1V6Y2Er1ZtoTkuHn45lmID/c8os6wk9QofuDjcKW4cTK2OSkwY+pFYGs
JYeFaqkfTe7caYP74LzhY/N1WWbhkCWmBl3eYtwNxqgVYmXQFx63yJUrsKeZgH+8pmgiT8cLnZ65
m6O0itTuyzhG534qvfBH1ucsSIB+SntGq0KpoA/YCMv5PEAqKFs9aYCkPaFTDc+BX7inQLx/6e6R
luyHjtDX1dG2UvoVkWFv0zp4XWZ5ZN81+ncjvGit7GJ8b+sqE/Nna1E9d5shlvCixJaUF7IBJiPj
5SU1n7W3Dc3HS3RliQgHSPwqq1Ntg9k5N2mK874UjQP+4riUVibUYyESjEP155OHqr8VjMQP/nHW
/qTzinPTUkU2lTvTzRkAOH5JghgaxCbr/+ztU+DidS/v81XWIRxQAurd9VUVbtnz4rl+hkHVgjuE
hv0ocgzZ0bu5t5Jv/6FvaC3cHH/jzzqxtrIJETbM4X2dNqwuD9cXMwcwa4BeAfE3xLYF0psnqjgH
sFSJD/at1e6UjJkvfvDv/jTa7Grx78c3rSW12uZAmhA6WhIy9DU20W0gjpCW7FiyLk2MMN48Pp8M
CgSNmwGIa5voNMFt3Pml4UJiAzCbVifrM3Dre8u407icJrrhyDrB4AqpQfWgBsVat3btcN5hKXX1
5YtxaaYTYhfVZqJ2rNekad6rDJLA4/PBE3ulU/kw44cj9VFLgnX61xSSY9NA9VqyI5j6NtKoC6GH
GsxfZwTDmoWN5oEwAGIoOL2VygegBL4P3DYFkg8rvo0YziYCVPKlnx2eX7o9FjPdpOTi/xYx36O3
HJYoEQq6opUdsA0pFzxLhpFhVIAiZfx9psfufeLK3d1RJvslxfK1FC7mX9qG09iPTgFwuPBj4pJ6
BJcYVM7Isqv28Rc4Cbeml9GBZRnb0mbAZ2BdyGmTXsd+Z4elg6K/RegWtosERGd8mgwzV2YDFiWt
dNX5AKko3kTKYK+1g91FN8+g5h41GOr36hNg8lc0eFXBkBaQh9q0oIL4ejBZOkw9M4DUokozksPD
+wcgh6RQvds4QHY13aTWFfZ5Ccluic0b2KOgZVMnJ6ZHuVxDlKlHUPfVV7pEe2DiGMYDWwXrdYqe
3cSrzd5jmnaHdgzMO6OBP8CLV0IbzsxyIDImU2WwDe5tQVdxLYDLo88QGhmabx5DmiVtDrnxyKyd
nYLRyLxeH/mKTwAl/n8Apm4j1U2Q5VERy2kzQGtwHNhgKsOOJ2oufkr8RTjET+QOcI+wy0Gqb79w
zj6o9p9UaJCxBf1lxi1rAOONt7k7DlWORBi0xHf5x6uszi/A63F7ff3JvOsdmVMLImylNgUypE/m
hkqjZecF1neq7+GoVdNTDmv8nlc3fi+hgSMLcbiFTWOb3BvFvG63L6ab2sMlVN/P2qovc+fJJ/gc
OZIa7hilew8bm7f1VRrDLZMAYvtXNr2lQPq723qhwInrRkvyjS81BU6CGft6CVLlBGjN5eDR0e69
ogCvB07Ga6kfFLxINkpsUq1Ik//wm2lbvIo8TkkoYnpXu8QIBVF/LS6yt48nWIaUyjKIuu3FQijE
FP1fcCEbxnvnmaARYYhZG1dAfuMOLJmt0iZ2ny9FtLmtmB91K3gebWing3yZr3SKERX3mWCUfshb
8dmSOYNYIZ9pJyiJVNAsgN26fKl9K+uZ47PYDepGXOFMMnACLqzPu1yXef9xwokuZPAWZo7zzlN6
ct49ym+p9LQzpPtkdJcyhMryDjBrpYkC7X4PzYYiY85dgOAvinUJn8FLlN6IWgqro8ig5+oLPQY1
hy5DqkhJ5t7DqH7VUt1SmMi3ldZAMJMZfY/v4p13yr9lU/r6L8LyrFkp9YBjnQFVBIegEjO/1Bs8
XW1cDxlYgUXANIfdi8WtzQR9ZBZTAbwfmYtuDzisNd4FgnXF9LLTkEiTFi8GuU+ylL8cTaQdWGK0
RKXcr+34d11/WW1sauKAiCmENwD5eHu5jiXBzYaxrnfwBEHJCgY128w36zet4PkfKunw8t5aBCNi
er1x8azwNk8sulrUsreqkqXcyZqoAvkTZ4V2SQq8poNtA625tYIMlVjHOm94V8kyi2jPxkvCSKxD
j8WOco1TzMgBpJMs0nKB90yALEXvMzD/vggnPs6ARuojt11otIdZ7lsPKJZEHQsPQipjzGAxP+Pj
tUShAEyGCru81ZAYQAfpR4ECueYcQbu0YZeinkb0mnKVFZVv0Ly43+PK/NRG+fvqLkC3CJMCA2D/
3N4R5y7lr/33GZ6h1CgLqkDHS6n68vmFOyiHNagDOWwAIXxuxO7I2RgvVWNGnQAexLqUZ1/EiT49
x0DZbN57+37grAm07clR8Asjd2X+MpTau5c8K1JXP69kmIikZOiUs2pvm2M2KUPO99davfSLVzRL
YHZ5i5Z2PM7G7tvjIUNKXT4nyRKP4PREQQIevboiyC9QdcgWCAwHfhS0G6/fPHUmH9xPdx7KiVjO
Q5KHerxFtlpAZrGMxuuzrO2UQKEiy8bsQLkRNLglLyEUhEohNjpIXVVF6/7UQgW/FuVmooq+sNZX
QxC3CB5zALS8CaR6zSxuQnG45bM2MRdojKfX4GHkeOHyz2Be+V+b+TBvJuAFNfVBNnaY+0Q6ZJpY
oQxfToAjkbtfFdTRgg51CDcodCr8wsrGgfHU2FNKFV2SpE+N1h9gv6bIAbl7uq6SFPVzhHtL6QRY
qZNL0Z0PvckHhXhD8JPL+pjHp+Qga+0KrwZTJedI/fKVjZMmUdaL47b71gJBTD1X7E/ek+1VHTR6
x3SES3IoGKT/ecyN8ze6lE8tVmNquWw2Elz6Vwv0QaD4WVXJ94mZ1yzHDF2/zGka3OKTDdzexoYd
FqJkc0kdIcc5gZBoA/AN5PVTBfXaoqgLMfUZqQiOA8iTQ3mjp4yRaP8qtYzC8BRU3mguUtLNZcie
33tIAynmOe8nNlZ3g6Y+Sot/KQc5GMoxeYsJssCu3S+hgRUNo1xHfNuEnCzUluhVfSFEFzQ0N46w
6tU/JHcKRRNTBrXM13dFFeb5xGtUax+aucARHmJkkgDOdz+5sw+f6au1QRjOB8qLbpsw3g9IR+cB
riplhAE1jYS2LPYKBfLgcP0g0BCTLoQdqXi0GuDVi16cd1k9oB5TyHEUJeQgIIDY8ZNrddLHlX7v
o4T/H1HLYcJJlNUVPuMjOPstlo1KK/SzwZ72Vx6maeCbnRYo7yweP8qOMskuiCWxSXM2cspQgM/9
dUiEEzk015GZKq0ev2b5kpYkgBwdD6RpzqTBgKl2id5aV4mmobCYz4zKzCWZf1vujCgJFY6SgdW5
s7VOvEvwiO/tQXjm6QdoIo8QrH0l1tWk0zBxTl+5Qi8yoJOTM7uQRFNdPFcOxlw4POE2nzlibUsD
erXoLOW2Oz0gFfd1v10OUxTUaA1qvMI8EJHWjhUkfO1SfmTE5SJXggiUPusBOEPjqWMMnk478grV
BSh8remKpebFtrjL0dosS/633Q7C6oFubG4STnfPUKOOljsRF70/JDtahvLgRShSO3OJ3nbYW5sq
pAEG9IY5d4Ym9WwTIQI6NJ3BPFeWarMdBYhlvyNY/lesWRUMCiWgRf9E0YE1eA6Nm3KMUH9u8HRO
aT/+BQzBhmEYr41+7DO04zV/hQbYHNX3mxBr9Q0jTtQalv3clut7zJ0K/SSZqLFxAhNdGskG0QUz
aXiLwiXmKqPjfbbJfdkvogkRZxjZATwlKXmE0G3E9jUJFXYYbqNqVH8dArTmysoFDOqNnT13cf+b
/2dn7SmtsgqPH7KM8xGKRYrGoJ/4c67vyeZxmfylqTTheucmKGVJl5FpWDdSGhXpMUQ8b9tU3Q7f
vTltUdibQK2Zj72++egCa+yt4gyvRiFZy+26j+BCEIR7r14DEo0+gdFdhwakH7uL6qwEsPMPhJSZ
ThEFkNFdM7bH0uCNgDQwn5BIamMo4f06NuS0Ltb2F8Zby9ZD+xBU06CIYrkf8y+z/f54EShPOPZH
Kc0Ixm7/9u6m2yLjNGr4476zkqufc13XKjKJ3rJZGb5b3JjtTUc1BpUp5/QQZUVj+eF3cF85aY35
/yVqOqavAUbwmYY/iBnlFnnv8O8G28xm9HULgEni88VR9GebQrMr3dxoa2VJxVNKmoLdkiSJ8EIN
xclMdWAwaqwVmc64PXhikoM1jpmsksmHunMybB9fu6Cm4rVjQdJ6ZMzD/hQwWlEzfacer2PYpYT/
azObBai9d2PuuVepRxTbxBE4uYE494nI455gcg5sHcA4jzLXm59Zc74FYLgF0CiUOHUwqQ7tZ39b
8QK9jrl0uROF9LtglRl5IeVB/l8HuFtf3U4qHs9x1wtdmOrACKty9N/9cCnme1IZLf60lTxsZC5D
/1uPGGuJEezzLKqcy2hmCMFAgI2R7HpPN8G1Ur8gXuzt1qfmI7tZJxll/8lWhH/J5qrlKy8KKjWA
kvIujQyhNxW6jY8AVgEAkyXgwhRZcNODGWpCctfuKJmGn+ojQmBu+H5b/2GGqHQ2qFvnmTgHY7kx
9n9UjnYzuW85q0iJa85PvpKEHQcJnoxDuC25G31GZe6KDF9mvLBRqykaNRvczQ45Nju7oKG6MFov
x/OLavWxGmWSfyfNRmmae964E1UWV6gadp7K0PhXdRCpx0UUGNJK29rCt5rzkmNhEEyCkzSsHIJ0
Cz10EbMBnshzZj75ys/yi/hwgn644SxznBhfZdZ9YsIgA5cJTY9WuGDpYIvAs55RcAs8z3wjUTYQ
MQxrvgkvXAP1oyg5PJ4un9lS/b2Jm+sB8kGIA4q4KykrUML6RJtOHYgDOIIZvw5dup0aMDvC17UR
vG+TwKDEDBm6LQ9rL6lVNbYe7h96tDC9AjYl8laMnjdZGzk2hxSravIN1/tB5FAGfwEhaPgFboQI
aw0VPvJGwg+vioBm/hP4aG/eMKb+bHcxeRsSSB0W3CWUoPVnicGI3+2CQcmMyNizbEllIzFK8fIW
tWbAS01bNb0FRFsbqCGg6qo60O2MoF0YZOHNIABBFDxqxmZvdNcQ40jJnMoRyZ3JGvyl9Y/fwb/E
z1oE8XqCjnj8e3EWvnVEbc1R4bR3Ar9BNzS5RiP8Mkpe0YCsT5okce67HGN0gOCtvn0+NizCjRkB
pxap+YN7FCHLZxQ9gXaWy4SFpZmkxOvVPYu6M010q8HWo0x/vTwSNCS79xlglT/ZyyzjrD4aFOd5
Y5bhynJq8/wryC0jKSyGSLFFnAOcekCsw+q/PQaiNLiC45biN3U2xJJK90mub4bfN4b4BoFBEzwM
qqHfEZHgmrQXA0rltRVJQ2rm6M0HYKj8Zz+CVM4iGddS1tL068+xkSrTT87U4QqZHtd6zPK/6ER6
XrhtHtB9DnXBV7WzyfAmROe8SaBWg3vMm3IYy7nAHB2Wnw8J+gyejbPepvazL+DfE2KnoD3/3fzz
vMQY+2G6T3gHya/Ys/AwfSYhg71zCPjevUoHYm6jESRM3aKEgPv4TLyAaATz8h7UuXvdVYN9nQqm
cLd/bGt3ZqAEE+icjy5CCDHwgZrT9tEzYIuzQsgnU8CeqooQdWzsns2YW2QiHE8+1LsaHUfRZRjR
L2oeXH+/2mFWE7YSrlXtc7IRkNO8YbGlXFV/S8p/FWxFMV5vrzGdIl+5LPygoajKmzNqeVCR9QKx
1adHBLefG7PBH0BP3ZPd1OQhWvvBmmcrsNfZnhmQLOcomcXxYrKcrJmMqXzWHK6gFg1p/53hldrV
gV80k9KmEz0eJITPbsH6R8/PotHZjRQcUMv5E87BTg0w+gJ1vPCIhlYO+rHTe873R6EYxeFBHxa6
mafoz0AYR1D35qpk41chKu2Qb8EM0evqwKnixqbZTf5WPC4n0fTjSDf3sPY0owTajFWmJHDXZF8G
cXD6WMxPP/qbIkiy5r4eXMRmf5CrAaV+SL0RgIStgFeojOumavxSOWQAxaE/2Ig4sfEKP/vdHOnU
gsyq7hKitmpyP//Yuo3WlK7Ss7v4ARfGgYlf61CMj0Qw2r1EE9Ej8NCG8FDyZa4b+gTEgd5zTsOm
DjltHbBaO5BZ5Z1YQ9RZlL6cJPOfSqPc7bw4G9NLBV8ZJvSv6uCi6/tfKZj+CnxRHyfsRbEkwdBn
/Gvz+FT6ZVqMPfsqgt4HEgquMAW9oAXbb7pzVkwg9efhfNUHLzqDtfT5tzUmYIs/r9uunhchWtvC
cmVgqsWr6aXTE2Gwkgj4rsGZZcmou2zQZfbyxGqw4bifvbHIM9MG8ZdRrv1OP8X6mTZ/xhDmIb2Z
j+sgiwMPx03AJwxaeESI4pgM5kC1smMw2oIACpST+pQ8Gk6EG6mfxcjnByzbR+FfNihxXHwXwakD
ohKczteBjtuFXdxSfiS4yZD/KZ0mRooTZ6yWKd/UKp8QR6Bnh4e+Ka/vVha+IWd6XzhFZMGZ/72D
/4Vj9c2OKfHs16a1SnOHbiz4VlqjFpwRYXNvIBSROdxNSYB83dCXYsJvxwZ1XGqwzBk7gupYhsiE
R0oaNGfaFNOonmcU1cCHQpeWo+Qdr0boxVj1Vo9riBkteFAhyN5uJHouPRrw0mvI9EwyR2Iu4i7K
WRr3N3LMoOMQY3Do+9CtbpdakRxqHFxsajLbAnDncuACZEEz3KzOJVnAnHKJw7ZOr7G1c1yesEGy
P+kmZ7BEDZioqqhokeAYNvn98xGbn26HmtDm1T8AUoPnd/vbAdl0yR8JE6B7/p2Hkfu6F7Uq9BUk
1/vcW47qCCsMLUAKVy7OhPHvlRcSgdxreoycjeU6VodgWQhIb/aNuCjDH8VXv5F12E1Tt4sFOE3Q
PgvAEX2lbPp25dHGiWvFWslzpRUQi5utAzE5Rp5m8VbPwF1Nii8EQ1LVJJ3h27Hmf60TqXKHK6J7
VnNj237tm8jIlxhCUzRqGHfb1+DUvx8EaMPUQM8RMBeLKlIVjUQZadNI7NZmiFBr1ztIxMG2nyjJ
BKN/80otWivaLZXzcu2uebIMhLT0+yshKrNA8d++j4LPBszIvc71iT8D2tgY9DwSyyIi0VWtuiRB
JuNkwWTE0BqrAYAj9DWVn11xxgNZS0iKyFYXCamS5V0NrNtU6gvZsHyONfGrm8OlA07leXjltTDd
3Lwlmp2mEvOec0YrRjfOeEwHBmKmEHjixbTsfMaM5OrDKzQ+WqKIA/QFQ1rVidogInIhu/N/V+RM
tQg99FHrEblArmLTXoz3xgEY988NvEBamBoEOIAaF4vEthTveIls5apcI+cLXz2bgR5Wyw08h1KO
+chHmAdd3GolJUMkdjOf8mEAqZ4MlWHuoHApAWn+cIFSEauBhDLhp+VsCwJg3vpxfvPz0rrdjJgt
2MVoYQM6xBmvpclaJxH5FVOMo9upkMbUkhFFCCRMZtiozX8ko+EekXnt1fQ6ZOShaPTT7JbYryU8
T8Ydj2/QW9AvGrpX4fYs8ZmVh3Z526LTr1tUPT/CFnDO7su9RSCWCSd/d5QM7tFaFLUIY9oaJjhn
i8BOuyACZ2x0cQ6j+k5YDUOviWXCVJjCJCYy0afC40s9DaQDNr9yQOaW2xCOsAPr11/hqicuHRd4
cM4/hO9X3KPGvLLnt90Xlynys0rl10LGdVHBccoUn1Ofm407P/6PGESHQqTNaMAkFOZvXH0EVfSG
dxiFUKnWjrSa7tdH2xFslV44LuCicECfH5Whxotw+Up6GR2aKnGUawoLddvviR9UgZ7FGlr9i5zJ
dl9Nj76oM/uN7FQkQbMtObw1Qppyv9O0uH9d8N4t4LRV1NchFmAWnLoHfwtr2jN86uFJQ/j8fwqK
dLDQKxnnLPCzTqjtCzwNQaP3EP5wlT5liT6T8Y+fw2ozMZUtOp4LT5pwHV1WEDRgFDWGAoapLRWT
d6OAX/UJ7zV0num2yFO7yfsuKErCiUquUJygtN0h4t1ajgh0syaV8h/e/PzDvzTiMbef1m/3xPgd
LZdYUdJsweBuCa1G1ceo4GUuGRUgp2Fs6c/qG6V1XZwBsLcQ1+AYGEi2g/NTmbPlxXJ5p5nKJ0cV
f0T+dSALTY2DKutEkJ+PqDeNBK5xprhcOgen+GZZO01uiz4NUj8tH4rQBECUszCzir+b4xBrdMKf
mYK8mYw1e0KNDZjPO/oXM1SwANHnNGmhPI/8oL+a1FppVXizLYq4DSPjyemr/pWPHx51UP4XUSIe
SfVXfaNKHtNoePbQlVBQN0fYI/BFfaMx8KsnExYY5oFgKwJ9PsWyrkjbBZQxSn1Frd7IC1FI2ahL
izR/SBdAh/YckBI1i8YYtO8PGNaM3R4ooZnpUQu4eu4M049iz/I2g3o6TEW/fR8g/1VjmDCNQ58a
Ay2Nu9EEEhJ3kkiqtOdNdAAro3nb0zyf/uLK8mQ5XRaO/OiEGhMsGw1OVZ1t5dpdi6zW0zqBsrFY
uT2GOOSZ24zV4uLZeMaL9K2IDMayTZnAIGylks+kek1NrMqtIUxqRmH7Zt7oLri/n1o534DvhCZg
FOh+p3XntcbHMo5ARvq4HlTrH5EDjfw3LeSYiIrHIdTAfoTEf4Pkx3o/7K2dW1hv2IzHhYar4YTG
E0RsffLCX59HGSGoKd4ERiFr+wrageQfNntmh5weqW8Aos5vxfT4FRWDwTN1V4Jp4rPyA9v98/kI
K9E/BcFeYWfv2Q3811JsyTzNsH/gUSLk7z7s13LW3Y/z4SOpeXaIbqfN/2PiZyUOPB9Kd1gamER8
VCageVmXFJYtuxn/N9CwElrb06N4YetDbbF/o4n7lXZCmx7eY9hzrtiPaPpcqud4WJpViJOWihCD
afbVhDznXima09GplZWSoNOA2iukN3FzNBp1XJOLugO4Os/8J086OA2EXm6wBbyATjg+CwpHNm/q
cuMehgCwAUMw9lfTLyDp6cn4IWfLXw11F2zHybHB89kNlHjNjJzQK3dly5fJLrBESEtvSGiXrQN+
IPNbAakyEy/RnZicthFYBQSx+zbV0+/6CAgsMxtrBHx7pAdWuYeyIVUShdmnzUarlyO0VFcx+qXX
kUh5bMhfmtQTF7QiUS5oxLRn/LSJW6e/GEdssO+FrqVdnMrcw1nlcEeSVDo8/9G84imHIWJ5MrTj
1TTSI6SbajBtavQP1CEzYFKdrA4sAEhDZ6TrwAx/TWtrNk6gHt2bUXpfPf2furGwXC/sePpbv38H
pV2eJJfmUF1w9I5H+k9qss9U2Y86ktJdCH3QNc4iW9cf2R+iGq/bL3HPNq+y6/stuzf3BZFc3Ue0
fnLl3nKOBE9YgWzOzz0DXpShGRZrKUhHfSnNlfZZoapN+f2qvET1Qjdaynl40H9Vsq48KQWgshDZ
OYdUh32bUOmumdIvYqVm7b1X5+vgYcuXgbwzbOUKM9KDZe7TmvmRlVn2qvciN4DYhgehMdDWQZLf
Snp54VeKrHyAKg+z0HhbXGL6NvpieptuQG/c0SD/Fm5Nop3JuVuUbCBb2aaEQV3KtXK3wy4tiS9G
jUyrYP73uNPfV71jJtC5JlYD30rxToCAna4m4MMPRmuStYu2mGVb/sWXontcyjuvrV21ctBRxgki
/qAyflPaDXNgIQC9L5+QZfNZ55hGTw2wTEXm+JkX5uq4yxQNQlEr3V09nGi1zZ4Su9UV92n+36+5
P5BUg/q3BmHeUdXYP5fyjdSmP5r1KmA63Eg84eWUpy2r153NCw8rcxuZOHiESj0GoNjvRTiB1ovh
0cpQ1jAp1ufABZ78xcgzQjsSHWLTwzetraQBVGf+XvkYH124LpMPIu0+dgqXb6LCNH9m0Qk4GUPO
PD4HfNEWxSfJ0mh4orUQ3LiyJ7+3uEiqGIHoHbUxC3+nHgQ0HQMLxEEITDrq9FsSPklbHB5O3n81
C1FDPNCCvyHXE71kEe11Cy7EtNbEMgvwzN4ym7ps4HZ+LKfJzC8tqd6UdTowey1Eq+2s7lkRRxG7
hiY7v+Gcqk253fLdC8cwjOyyvs1E7kY4iKPTSIDPTm1cK52BrxEdB7p2DIMNJp7eFmdrmgtwD5uQ
QGm9kiOijmB0oYVq6UW96U0bXIRyI5n67wK2nRNUuTFPPcLk+t64o2QKDV0+C65A0RWL8uHKhPF5
1LNrKFfXuBoqVDOTp2QS+f9ziIr9xvV9ZGz4GW1PMkZYZKBbnOC89KZw9fEO6BbpPXlOzCP+2igV
bDB4TAwPh802TiPeMqBAcqiU4vpM7Y+ZGqZvWRVR0aWo/PYdUpn8IQIR3y1wL5Rtsu2kg0urDoyI
daAgKzqDMHeaiGTLYwX0Rk2ohiG99sYZCZLJPLvlUC29R3vyGIh40rNcQVP7cKhcYaDNUOgcLKZ+
8G7aVLi4rHnbSbgS9iOQppDFkT4oKaERmXZbJ/IU5S3++vrEVz+JUnrdqhssQf0MVAOC1ecXcaRd
n7hnLa5U99OuUtg4K0RBtYqQlQnF8W7hj41TAOASWQpEURQzSThdSYfxRi9uU/iQ1CfpRpcwCOAr
mQjTeK+zhY8qPF1g+Jh6d11uHfVfqQ30Du3yoNVT1VuIxiRDHBSbGpEeZlHKg2FORil9qQ2YuV8t
OreXEVRSFKTzsX04qe1g20ntDytjPUBpsFNDjeCfYGVCH3spcbsjQQJSE1iXPDZDuLIQVWIVAEpW
XFSFsrtKKP9xKdQhof3Z7/Zi6K2fhS181wmZv+hbDGlEHkJ08qD1S/594yX2bpkkrbmWIoz1hZbn
jEqs9Be02XiCgL108wgQ0JP8n1J6xvq6uUbPc2+xK9MMJcEDilpyqT61Z1YsAvc47N80I9fi2Ihv
6Rvd3r3y38ILq8hNFuULAeXbl9NZCzAwYIGyUKCtVGniU2yO+YmSqk7nX8dYOUF30K4d2bxjfon1
+Jgd3XKi6Vv9LsZPOImcRL/dkuYeWpsLvxlqX/+YjjB32EVF1oRIIPG4z74GofW/dPQk5fTDjXPs
rfo3x1tUpRjN2c7w/FJ/m/4nKzHxSt/OrrJwPFxIfKX859XJTFSKcLS/DsSvVoBGkTHgMwwHh2rV
C7VZk1+1NuZ3iPM0RwezkfPiWJq+bmRrUwtRBpUSJVpDFrV/xO2Qp9bddOrtpQLCHgPhH7bLEDN/
VU35eKnvSvIjWneQmKM7MWxYu3SMdOHp8a67vkxtu1sOAq+idxGUplvC88N/mrJK3TXyKaSk49gu
4YvR5Lr5llOyRDqWAPB7dTT4iUL2/7X1sJ410RwGN+BZStRi4FRHWPt0Jz8Go6NHimm/Sp1+d82D
zvBgkzK8U+iWI1WgsycggX9FiR25uHlsXH5ZBhJcjLDE2y3rAiKGGE/f+MIYceWyly1FdrthBMue
SeDvyYZlrrVob21dZnH+v+lrPgIHrrWSwOC2lr2gvKQuGl11njVb8g5pKQ1oq6fAK9fV1VKYPsjy
hDzsGAjSBksRcAlanseOE9iow2xHXir7bxyagdBNFQnPclb/gYmiJnsJJFaWRIfH35cBWvK9gyDg
ncJRIgoOBvKZAQh0ZgFKWp5i72xA8xtaQ1L6U9FNghqcuQv8eVmGaPTnEicmLVJlFEwMcNSGrXzW
JoY2jNdvR4wW8m2WhTx2d0cqp1p4u3Id8KbibpVhqcK/eEDYQ2IFJa+X1bWLDhhxnjb0elSd0t0c
v3utCb4I0SighVPDIP6BbcOXEZYqNYQcJNjy3Wl/VdCMSfPdVlUffgoHtQM8EZvUyNZq3EYkFuSX
zKDqfWMvRemANRXoixxMi/al4laYZcS/WwZBW9WSK02JbzaC5O28jpzYx+fE5mKoQQUy6rgywxYy
JoHsl9jBBlY614etvABbecSQoSg3nWbO9E04BNIvN1Hj8qlCkrFS2iYOTr7pY6vb+HaQG8QrMd1z
0mAlsrpKepSrXAJX5z+ZD6DfaPNRchl1KnHetDGUciKpmX8a8nDR91yIQCEkNY1TgHPoNq/eW52N
833qbnCVX6UHyjL2Eu6/BxUzMNB6Wnqe8GT6Gdcw4ExMjlejCvvHeHmHR1Lu4T/L4SUcsu/OCrIi
udisvhGPQiwnafI5gmsmvq888VthVhzJ54rZdx8DULaeuupK4rUxRvxiJy+1dGyHqo/WalmB2Avh
BVYFBBnZOE/Tifs6TpgA1lXZOQT/2OR+RnLn3GInBVS1QTmrIJD51FXwrdNuHym8FCnVIHDtUY4/
d0DsuSDcJ/Kh/koy9l4IO49NMKKFzfvpdx70xSM3HcpJYiQtqpZKEMHX/NUVTcS1aQ1HpXcK9mzZ
kPI1NUHqWe8oAqd/48mfMGFQHB9GdvdW06BaCOXHouGiJ144/vQIwk4/oosABJJn0HYUISSVlvLz
bTnvfZsMXPrTJVAfYd/yYXAS9RQsb66hW7m1lpqx15BwdkYDs5T496mLCeJKJUHUtQHiar++mJT9
cwzPMD1rEDceGxH0O6oAocJTUm36HGD15Do3lAMvyrXuQ9nDELvBirFq71Ahf5Wilo70nvnSvqiD
uECvRgYGsIgpOda18ueg68q1Lp7AM8KDzj/tViJvIVD8Akxrox27WM7modKgKmOducC2kJKdzYiR
M3k+KIXOErfbA2bFDQKhAjJ0qDbsfImdUZrqlLKyNc+o74W+YoFwM4V8uU65KghVADtdH4vLNshg
PTrdLlYBqU5KhbU+Z3NyiLfa9DbwNPYM7UvzswOsD3f4xzLitSNRwlRlpNrQCGyJqiEy1MmYur8p
ZgikVJn+a/R9o8Qf3F0awmCqXw1zcmke+07qaRNP/mEflTLp0hPuIW7DEXGAvq++4qOyxv7Un027
bTpRzzdDawL4QfxiCtOvXcG72jGksD4ZRw3lPng1hRmm3UKPRD6QvxbGhFFL3uP5NgpkVJG6CL8D
XAVhXal8xkDtX8wFMmeZUImtzxciuR3xibtxkADeDFXDJLq6cF0XpZGw/SDkPYiEZ3qGDRQrGagA
peGe2spFXkfMK9CqJRp12CbfXu6lgWyaHrp1M/WL3NGlrgfx7CUW+BwelssCCUZ1YYJSNL5COzGH
ACkFsYCXhzlkl4B3opNswn1wqrMuVncUpxQ/ZO61pYCA57FzCWSieDr3qYO8cdBqA5i0u58TXotr
MPZJ2vMXngNYdz5ICXK/s/BrlhhR4plka4FLaMFoAaOGMCQBXuHNQ7X+zUQs0vBRXpHv5XoFKJT0
RtuL7F6MP5Fw46ew3Qm2en0Nt/8YWSMTU+CNbO9YiZaJUEdajW03gEkaRPZs+/YWVzwImOG3qscQ
nBly6yACSIvy+JnkQ4vCUlESWa4zQyebqS2DJ0EySp4nKJfu6AP0FIiRS2u2lP0TdGTWNZgp+fd4
/4ErY/VVsRtpENGGjZDGoOOgEU7Kv0z0x91PGFS23+7QIaHRHPf4I9BcptnXtwc8qYwFiqJhN1hP
i1ztzk7fXqAtc7YU6ji2gAwhRZk4y5BLF68jbtZhoOPC3MKs86gTznnlJPwcdDatDKNv+F5jSN/F
/p4uJOhMn9nZNmNPOkgX0zKDyEyG9spiyu9ObrZqOB/WJOvDUhkxvw380OmeMKruWErPmc4qBVN8
tcn+FKVRDqiQshrt7jHf8GJbjWFHwfd4viu/qVZsD5ABu88Bx76I0hx+ZsI0IpA+eH5Uc7xyO7cO
RJV4acJ9jSZrwi3hHrOkH1ESownI5Kc5RpRUGPuCY1eNZE/WdWleq11RKdeuRixTTJ0xyXmLKW+i
cHa3IQ8N4D/ICmi2CEVDn8Efi8zk718j1+r5p/XQhcr3GpcgcmJLKQcKkuXB3HgEN/JInen6Hod5
0/o+jP/yHtkFcFPB2kugjFSyQ2V8B2np879lsdsn0SQDYBy6/T/2Fb5LKx7ZKWKBObbtcv8sb1Et
UUOHKoBs52rgc3/q5uZ+BPpdGEEBFVq+WUUSplM7WleFA2iOiG89sgHgNRZ0b19jsvALG+H1SVvU
5d0Y5EwGJtMzga6YRB4SqRXBddVst0nMWsGBkm7GBGBzW9qf6s030Pmhq4CO5s0k731YfHYicTxK
YOUPmg9kZ+9sx1PI9HUlDxHzaBHJPt20ktNSLMcLPmWQ0vlLcnYtvZZZEuo/jaQUOLatlQLtnjaG
nXc6iLannNZjq5xzxLBot7Fqp7yz2/nS4oWgOYOiQeYUAPr3sZ+/4sCNgjh+p7xhoo8ZxRYDAlZ8
yxSe+jiGzqYztHT5oDGHzd0vLsSYKhInmSyOKocy905D6R3DyyXOI5HIcG4m4CSmlmH974xFti1h
V8HO+/dc4cTyGq5ktewwErkSRRIdcljujst+1JNchJwvgekMOkrDjRe7o0chNAeFqL0JeRF2Z3ZP
DrzmRlVxP7QwP/xs8Xxy8AIK1KGCZspIG4pDK6eocQ/2Wo0lYd/v/FRfxYSC6vzoVnLViwyrhxgx
drvMebeWeA6//ivykchpdgGhnPxq9BigYAn47WhoVaJ/9xOFMUiTnC886FMBM+JqsBryz/yOSMY1
dekej2Pf1Jw2ncgp+z3PfanuxhXkZr/MEZFo8AG6uAG5en/EYZ3ja/hfXUiCWPnumxq5pNwnK9/q
ik7zK77ZvlFz2NhXrbc6c6sDUv81EJtW8viSbdAmf/vhj8qRSvcjB3QRlt00YM04WqjA3dOhCaad
hwckXZ9WnOFTvMGQV55sLPzbwhi36e68QyO34stUWxtDukj750mU6ualwXWUZ8Gq1DbhCmsAgcMy
6H1sgK55TefLXNJTj2nd6TwNV6crGBPmuQvDA3kANXFt5J6gad7UMO48qKkLF5ZO3bmCh3Nt3RMO
ayGu3TgcY2DxJC4MNnHpuokb8u6o0lu4AhtWLBcfBKddtRkyKGCJezDry2+MpcLANKPbg+dZ3h5N
+XIh9qdM2/Eh0P1x5BGMJbXbh3AgXjdev8Y8DbwHN509sMdGNLHlErNj+O/nJbaWTtrG0fWQpuS+
JxJTzv+sjNBWN2nXZTxly7P7kwLNxyqUO7ccnLkl5XBpm1wJndutbrqFjCCyW361h4mEyFsqfR5I
o1kBalvYShX4FZzd77GJjtVHeVq3Evze2EnV57DfgBduLApe8tggDateK0Yl+B+keC1XbAjyQXeD
M+6+cFwo/majiRlezdpKfx5Lg/ZQUkGgv2bkoKsUC/ZDo9DWK/2R4wGJhRQTjwgdJW5yQpwDE85a
w6JF3CpCI20H2GQBIxXGO+ZbqoBAc04MJq6IoIm9tZH4uZXyuRqp+PsmCLCKh8kMsz6osw4IiP58
IYf/CwKqFdLmpFRb8FUQ6dqal8xi2BHTRBARDRx4RwmjGOKLHpUF52cu3XbpOm5a8o28J8rXuIma
Kx2aK3SZ3lZSAjVh04gYV4A8J6leYyFo7HnhgUoJwXHblnVtOJMcGhWpj7TqNJEYGVzopRM3rmrX
8n546IxSloP9RC4V9mz72WHjwDGhATxwp4F5Ei3w8bBAYmp1/S/BoOoNKwSOUbcdoM/N9fEntE/o
1Un4dnebHFaFqQyb6ZDRgGLKHTR+3xxvGfythrwrMgCvqFbZgQUJv2ZVEjvBZxdf4mjDtJUwQTa0
GH0/wBWWYb46r9tfEUrcwLnGOCxgohTiBvgp9BKVeEgfJRPzi5YeiF6GVQeyUW6ZVW6zIueMN/J6
tI7TxwmAZsAj34jDxGn9MuqJjeNxml9Iz487im42o04vj0cHpi4EUikhEzay2Gzfw1qTRIcpHdzU
oZFX7+vrmQ9XWZQBvoRtenBOrtQTVFgCUq0YFpZyRWGV8/1Yaelr8PtCELK8PkmyPis4Uu7Oqt/b
foEBsFJeCjqKlmFxWTAQQR9+7DfNG+3Ne7t8j6wMdxT7m71mQQvPOPPhV26gVeeCps3yn3H6RTdW
p9b2Br7zf+/IpML325DMk9Lfs8fDt/ss8TZ1syFlxGrLqRKD6vhz5R8qtG99aQZ3BNXTIeIkdp/l
00uW/VgGVo2YIQbJdRjiphqj25rzshVCS3uycqMjt0tUGx1mlQH7z0VCSeL3ts7Fl6ubB12MIyLn
1uTdHEgzpDU2vr3j3nsSBeSJfDmZR3kUD506vJEtuZnNBLpsogvtSfmbesktWVUQCdYi1DotG1sr
5ewAjZEZyJFRFwjCYoBl78fY3rmK18Rnvmb6cYPujxrTSVp88/G9D9JK6eAAvrN9f7x5ZTzlUyFI
EFU45nrQMqsxvgjaGr8KWgUEmL2Y4rHuHT2+9LTOl3Xl6oTSDjrsa5mu/6qxy2kbiOAvotpCU2Yb
2F9NSQ+Z1eL6/ZL08b7GFsNgpdtBGUZJ7na1t1FHEDYiDxlqoUNEpSXEd9WvxhDkvKDPe8Gg0GIJ
cOwXRCiQB7Un5G/mQeVrf8w0P7tct+GTBK9tOZsNguh3PVEUEWNCJPwwdHR/F7DwTIqyrCAqJKUd
EsUdNzC/u0muX57zY9LrygSi71qHhEM/aLdwHY6Cavl//IqIE+jAY5vBHVN8KXXF7ljWOTYGWCgR
+FGkSD1cCp2Qnu9pJH52Lzi0M8Jtq6JhUioDos6rRNP6ja0ze/PjezUjWFtoNg/idUz2htU5vC7g
SmKZZ3c9jMna6E7N/0UHG70PisSGG71MSLO6mYS8Ffpp64lDTKfw1rHVd0k32P1AQtOAlm9Zbimf
8Ap6JygxwQyJ2w5oCoHkQ/zoJHSceO/jJoa1M454wdLGHwRC+I7hcILPTtj4eWF3ieimaW5Vgpg/
y3ngaBqGaoedkdhb0enES2ArvAsvdGiUAbLT2kwxZ19kvrSqo/l87qCFHW5LEPjRlvLdVm/CeVyU
v3JhRgaAV3bRWa4w8P063RXcJZqqmOtbF5NhxjZHc65oMyDNFtRtI2LCMwiW8EdO7VYbcuBCCYgR
fPAYbkJpIcsL6CN270wDnHDZDalIUUdPs6sXTwP4gHVwelyCZicJ7sXSLhsxcZ537VHz6R3bmjlM
iMB8bz7l0MQQ2BU0vPdrhE0iCkeX/bqD/i1QWaQwi0rDadlMNQr5j7sy93Ql4V4TJycr5n33D8OK
ZOSN070bq2adboeGxvmO2yuv1EXxmOTt8p05mZW1h7tudf9tUkQmvV9NxSx5deTJaGDn2yYUUCsJ
NUmAfZBR4ixdHAdRj/4pr8HF7Lexp5FQTTvhkQUiNXPjqSfMFdLp8XaieHUQke9rOHyPO4DJOnkf
pIO6lZ1nYNdLIHje3EBnBj01kB+G5mtFHKFXYF/DWg7XhA/E3vJIzkR3MdVhfmNUxFOa8L0tibWF
IZA9kKav/6iexIMjJqPMuafAe6bblt8RZyRDqhq/hwPDxPNDuWqAiY3uskUWNCMQNZf0lBSHlfuT
rVzpJRx0WxC5FLNclM+97zWCfWPn4ph/9jq6n4fRAIJOw35DGgY+CRccZ6hdxriA05DyIxlsxTS7
pxLm8IHH4rkXqcFA5OeIcW/YoodDUMOoYRvRq8CdjcWmXwQa4yAFLY6g4oQ2JzAstGd/1qZKuiT6
o1b9DTG8wqCsyLwHDPG81Pu13GMx3Up4wgAAe7u0BtfXPTB1Y2MtBtNo24hLDJIgGDJERn/7IYL3
c6GVFxlwTfpa/6CGDbHX3uEnarA6ywb5bPnhf6lleh3NfJ18a/JAsby0x27fO0zN7A9Om5Q66GhO
SFLf1Gsi4U/OHLIAnTcZpQ1ReVEN2YZyuEWiI1v5J88sHGtSYcs162goE99qnTmfCmNx38JfTYMl
vNg3ZgSKsa9KL3EH4yf0UdpTXH8F8B/gn/Xda00iTEZADTRg/bJCLG83j387y4nUoQumHowXoFid
YzoHyBZup69K62Y0iBmX5qWGmDemVic37+LzvbqfuPV8JfPjYqujXw6R7VecZW2ldadOhOA94iT+
zUJ+0UjNp3i0y761HK4W2w80ZvSOgpZmD02HhO63shA7Osk43gyx5d0TF132mj4jBofbf9zV1h2E
LLbU9y8OcAWGI/NiSxDquebNYoehKfibudvTifBeVjUqdZKj+BY1/lwpqtA4LZl5UHGv8slCFnur
nJIIybB2Q9+ip8uXoAHL7SI96On4OymJYFKSay1Q+W13bVow0UstTJNobS0b+RTn0EOUwgWgV0CZ
OzUTvWoEBMZQcbZJYfbMa/JblpXoX+sdW8xnIbTCoo0jnZTobr94EyzYcEKPxKhu0tdV2CXBQb9p
7wR3ejkuNZZoJHzvnA9z5Yb9eBy3bWZrtHbKsvnT1AyOTcQmcZMltNX+p866NrmU0xt9mj5zARi7
twlXkgYeYnGDDUEmiDFLhl6np838oiJ6ZYYg+Bd6xS2mxoEbKyV1idEcS2QAIZeh/ezBbFXzMv8X
sP0seaFhpyWLkGpP8njsOtTalk7hlGi64dU5xBFDlpLt2bCqw81JS+DFn0kBqmBvFT5PmzfaL3UB
/4fL8PDryXGsd+UvBSQi7Y+8VaIL9/0I456bfUG0SUZkbhYnKS+CxXckbjE0IZ1jb2NPw8x3W5iF
VnPnji3s01ZTnSDHfmt2b5Mw/N+OkzWcW3dTmzQiCZ1HGHixVlw0piAbDqryOqUsZQB/hLGGW30k
YaL/rJnmBVAlDkr4T/eJtCpkI0ThJvzhzmCicH+Zz2HrZwOtrgK/tPdHLLdfII0TtHApBRPxcNpJ
UyUlSySDAyxCiiCcLulVVAjVTVuV/m5Rw94hV0lnHqpHnThtL7yTI2GDlSlxiDWuZQ4Sgr8AC1UQ
V35z1qNvZpc2k8Ge6cM8mzxfKyS8RENtdKqCB7mhfmQ+3Lv+GVQTHytq3TSt3y7f4Pis1FgPz9Br
kWOWRBeMGQ/alWkG8IHEztoNKBYFsn0e/VKLJiaZxYe+zMN8S/HwOi+IewK++6F583/MaqTeGxwv
hjX5/bLW51nd8Vmq2X4JG5dMZTHUuii4fgCK6MO2Alwrtwnve1I7ysUvnaoqaTJ7AehYmRffh/yH
4wza6qTK+f7RZup9auYGx4W+U9sK+TYaoUT5lfvNeIaB8PTSLy0LE9eVvcjhFgK/Px2nPrXLh+yH
NJf/n8Zt2vWo97jhe22tHKhUS38yclbApEX8OU7xU3360LpG649N7Fb204Iqshxv/HsL8IdFyPuV
Ros/NE7nz5Vd77dCHt34yN53h169aHnk1f6BBJOyB503ZgT1RnfAveyrA0IPBOlw7D8OJddNwyfS
jbgf2Ae8mL+Mvz5igQ07ajW2NYxY6rj71NloloSrRgEs/Eclfl1Gloo+B4fUa4617yPLWbaMkTPh
ci418eeZ+He1rTT2XKHw22fptpcNl82OnHmiTcogTGOVjXFFlcg5PMgIvO/0a7mK8zG/CkJaP1U2
bKwqhFPHIdAlwVjFlG7I6gnRe1rQ1HOLUwhHD2umUZdWn2jnCuOZ5p0wTlMcj1KppRkvh2MSeBRG
7ODgIK0Y/AQWRJK+Luay6tw3iNT2NpVYVwpS7NAWfaoFANGdCqlJqt3Z2eLdk71e3N9PptVYNMVm
T9bs4sJldSuoD6eM292+rfZk0z0V7mG2OH+pvk43b/kzz3Sb9PdQu8R+PQ/HybWh0RyIQ35FVocP
i/OrHB2C0Wb+C6bVwKDODdNU1DF2C4tp6OU75h1pp1YqpecLVHXsl0hdb3k78E9tk8NyKUl8AN6I
S3Mrvlmb3qymyk5izUe5F7NqZSfndf/w4MyLy9lEA3iEIo0eRar0E360Uf5LhIsnAdcYbhbDH5h7
NfxOQXy3qIUElwpRxG72j8iIiEqFRLYKCWE/9i8N/qsjQuPPoJ/dJa+mKY9YqI7q+jmUg8vMLDl7
LwQ7EQTb9ErDO5bhRaJmQxftmRfXARd4gc+Zy6XGsAiKU+hcFB+Mo6e77ezr0bygfy6wtIS8mhzd
hiQ4WbqIeHxPKF4fzw748tKLrEiD+eg1h5no2SEOTIhDPrKj/L6/b7rzQ8Thn7mofgIukRCsAntw
LfFITWxZWGrrHw93R4nMSr85bpMSEKU6b7fUs6V1KMJ2jtIlK5VaHcCU199L2KxI8j9hqijS5zn6
Y9A1l4N9IxrYWm+aJ9a7YzIYk0lUNk2KtXbXWUB9u5st386KGIKyuU//SR9e/JCHC1I2trHBrvhV
A5fib+IiyWUROQ2dsTXZTb0rH09Bu4sjzCTCSqK76BVK1KVDztOXW25/021FRxH9BBde8se09yun
EguHIvUPD5lHWzd9iUO6QbRKokWyiTdc1bzdsBXFWuUFSs3DQZdLsAFAWgWDkBIOfTgxtpYlMunS
MY0knXXHqktpmpNpCIADmRStrQY+nw5izJdqBBqD1JjGfZWOKAogsoQbwD9YFn5T5/jMoDjnAuhB
q0NvO0bPfbOsgpcD9Tzo7yEki/ni3pzOj3c11vwGHthg1CUX26PSEY8cWgmmQCfyY6O1B1pvu/cJ
lqbGqBOs7JVi4nnQDn0opmA7xifJx8igBwvxIRShbqh7hcu05a3/fvWZ6q9R6WZd2IPgXrhO4ryU
4Ic0IBkhMTLiR7dIwU5huOredkPOo4BNEpWQWGDI7fVM0k7SAIJzDnJlodMMDl00s+W45mCWLA5/
r2hyUv3sIUxvkiqYA3+mSzZkN4gSDJCMmuRFFBiZ2HtDVEJoTEg7BC2z11XAOh/Wgmk2hybnKrcl
NLDaoyUgPqYPEWbyoyKX+NXV3eO3stUePWK98BFmi2Y4Y9hAGb0dcMJE46S6pP/sHy2yiuEvaHYl
vaAniGSlxApwTwhRY842+jOXM7A5bQBMUPNjpp5WPXR0c+Aqw17RbtoOXtWhIEW8AmBZ05HgFTGb
COkPE/MvnjIcsdqSuNxQFFuw0r1wcEksFr/e0canZOdOK4jJ4nuZyYAB7UAF/3rPK77o766W4WFl
FkUsvL5Py/pBOKI3bTLi23i2UzP33RtE3I0KL3wyRnucKQBmSy1LGcBnL/JlLA+liiuZzoF7a+dt
5fQzzReq6Y/7E243E4B2hrVxkprWjFSMRIiNyiJpBKL0SepPhRexlfefNO++yNj5pzLyy0mc6TD5
LY3062Tmcu8stNN/4jX3J1oHGS7lQj5R0PYt5f8B32Fvn6mkODGVwVtwCbHoAf1Z5+ROLPTE7kqy
15GnagMYFtHtd40LLzuMXG6rym3XaYnnnRe5b9oeP4rOArnGbnakV2NLL6+1lOuyrxvdxDCHzSX8
JzqwIcOEJrn6kIquDjnJYvt08utRjBOeL6PxDPJNKsriZL8ykvF1o8zPD5RYVtPqpy1TVqexS/az
if4yVfJDEDtQIuEXGl+B3HqPnOTM56U6dljYpdubDO9VPQk4vsUmbYLHbYR+d75Oz5Ue4+SBPVC0
U9A43rOgtIEo5zay7EMPaendLoO8zRzCS5xUlzfQOLgU1HHmDhtO1g15FgSKDjPIbl9YcrX18eXg
q6e/6fsjW8rEFnDBUeWCcKhD9yhID/RC8KpwdVa/NiMWdBIb2jQg5Pas3OS5eFw5SbBVlTwXc9PJ
9vH7fWXWVMhatrNZcHBL0yxzUMcdRWoSFLpv8WLWo+NAIrybDjq1Xdwla+SHla6rRB8uQHCvNlXA
w807KJ7UjLJHW0npiC2Eil2rf/TzEOmHVLCKiV3nRcHVswjsd3CGH+8WHKv+mxbAsyUhd+Y0rKHi
FzvK3Dh4kjQUDd/pYyrXiNn/5n7KPObMWYgJ06IAiNxJ2AC9dmkHaOVUywYx//hPeouMQwOqfYRC
jZ3ueHoCrqCsJ8/btXOUinJgngq2KrK6jTJU18/ctlypv33NIYCEgLkrKzic4xzdPYUX0ZHRPsfQ
ib61Oky5DzdeR59WmlKOsROvIL3UNsPb7QtinDC0nA5F7AB/9rl2AO/FGKbSZk5WogEKaXIdLvK+
F2HxSqOb+MO3/4svVOnFroAYcEVfiafBp8kx8HgEz4w4b5EY78GetZq9O733eHUJz/hRsSidzh+c
7Ig+0wuHuVUJYArbMs+Ob0FSmgBn4JCuWG5UZGXWvt6tKYY+a9pXj3XFyhv73EsScA1/EmAwdJjz
teTkfNvDNxV3xUkQANePH/3G8VbneWxhi2ysCXLP9or5zNK0pXIWdGRfFEBmCB5+S6BjAZ8mFIbG
PjJoX3XzHDpNlgo1hLbyN546dMrTj/9Xrm9mJwCJr5BJgO2ae5wktVEQmwdMZheeTg3QzxhA3TjQ
q9DawDckUsOAqrH3RwbYglBfDjxTGrxzc97Ca0NnCRu/DA7FzDP+f+jZj6lR6k1bbV7g7HOy4fi+
wd22CpHKVkWoDagevYCNuhEapPAfuB3MQRxUe9s3uJVMsf6Wg5XHI+U561Pr2TqgyMP3ysuFFj15
LR9tXuME63PXoOdS9uHsEDMcxSHPU12hv4SgmnDTVL9zxHbStYjl7A12IUJGe9vUngjRMc5v0VtJ
5NqJWO4m0kTGs9kstPBYE2IRXaykosP2W3zdfgMa8XSw6SlhdmYrC5RJh2pKlUS5R908/2UMT8pv
3/eVOVPiuR6V5OMuhqtbuuWJjqfEge3hEK1StOSgJkfRWcPwsHsD1wPCQ/EehPCyn7nJsNhUPbNd
nI537R/kJftTpBmhIiiRdT/p0SiaXFzuUGLEnUeKTHYwfdAOog4LEuso+VpWy2FqhtUkA+RciRCE
/l0rLWDTOvKsTh7asO2KhNmqD3QxlZA57joTqYel3LmutuCEytSu0nEXXp22PU8RLkTNaXyHiqrg
4MZDVb9fyiwsgjn0WvEvA494i4bigyNmVjZnkhn56FYXmsSAcE/VuWZ8L0P3669/opY31cds2Jre
7vTzMSjSITuRGHMkLJYKRjFHtqeGDXuyoRnK7Z1LUGpqXZh5rBuJ3Fb/CK7p3YhMVhlI8xxKz+lQ
lV1SfhOy6bh6LDPCz27o21VotbgRkbNNTJpAs2qYYulJnbh7uiu0yV6AGDUwrn50IM2drhMwTNZh
4dvAizZyX/fVgiJTv5g1BuUUIrrsLun5C7YneuH3g/FUXT+MbRCyR7NFNDInAY8bIjoedKexTzxC
d5XBAvnpONbcFfz1jC6NwTFZGxcucIz5pcJ2jsaqa0oBgGD1NisA1mQ+++TFZgdPT06ZeG48Nai0
f6Tse03KPCSIV3vujc8jCayGHPJvzVXrluh2NM9ZmmWilaa5j7sbyMFWU3ftiPY/LKzV6qLAsXQz
a8gneBU4TRHtBCJMWIi2JCvFJXH86k1ADTZenqVRtIxdJiZUImMtXZqUhvT/zJ8E0jShR7wqWRlU
P2RHpSb+L3yXJ38tH+FWarhtxZ/09qtHsAE+usgKIVKd2rm4UFU1ht6vUsjIZr6mG2hU/IZIs+YF
6mJArvLE/mhMK6jZ6RBQ0MsRmSGMx/d6RR4TGUDkoTH/S0J/CwNIIAY1Qd5RmnEA/J0qUhP/malL
eQ1uyHSHroa4tfZIP4tgbp3LT3hRuaANZLQtYf7ExBHELHYuVrrQLp4kYd/5gZdvZsImsCpYjYmZ
4f3HHCZ63ChBf41Flrq8H7TOun7+IofxPoMxzYUmF+ibiEXVyLZFiHM2ZK21MWADUAvEm7+Nz5sD
dr8nypgx14l1CESdADIOVhvDR7nCxqV7Vf1KgyswUzlSutQiSkNrySCKg5Ap+T2SFXv2UPUidFGH
/HsmwNOaxvBaUkryyJqPhMC15fF/Q2+DvsfGY61bSp8MZu0kci3xPQS0VUbnUpZn7rHl3wQhFaEn
rqrWycfBEVQ7rCoG65AJL1rw3oX8QNb2rEbdkK3yuWzzOKus5TQVmo598i+JfrmyDBaOYz2B4uhm
kKgmbeBTARFGlEQg8yJXJCivM7vXFkRNbQe1dUiLcCL6rP0LWGaZpqyeUSmoxtll46OrbMIULN0H
/0ekvD53pNJ6bTFnhhCQkkjqtw2MUE05uQVPS97eHPs6yldVTJUq1LTrK7QOhZ6KeHPrf3FnmcLo
HMFMNUkiEpOD0gX8fSR1fn85J8dFwONNhnx6qRnbrxGQeqsIJt0suT6yW86zhE1Fuc1YSz5oyAaR
VNDnj6GiRmMsPB0gfSQ+NNBJnu6/oAPR/LqspZcRREkl1T2DpnooT5SKTbeBP/flA0AqKXwcrRVU
6rATaD6HXfCFTXsAVFx+NuIKAKOpT/4h3sSYYXqlTSfPuM7f0maDyWuiJxPSCk9VywHDhTFfhl9L
yXB5J59zl7lGgzlu8d9XY6ro+s1Lf/uIj+0zYPmIa9OCAsqQAl6KBHPAejnQqYP9UsRnpscUopwB
+jJV4rxOpeHCXarYnGVypC/SoLkwMslTbdQ3mggoUtDI5fLnVGw1ZSZK1cKWBv/5ChCo2jAuI3IT
+eximt0UDgS31XuzlF9sI4IdiZM2epwy5MIA9Cl8JYDp7A6HMUzqrnkBxmUKHpGqLKflCSwmVgd1
cyaFXkhPzJtmm4HdfgyAx4UbDlJKhh76sf/lCL5xYqqEwLmQUgmqsLtodhQphZBKhH3r9Zn17pS9
dXPrR2++XZbk+IvDB6IaAucTzfB4/4f06Lg7gJYO8POc+P+9S/sKCmCaPdCuHlHyvGSPPzGfRKpu
eKvAC7RMyGyG4bYSwZEYDBVpwlR1iCojWuN7S0NYPmpOnyHwmWTnAEVjVzUApNigEbUnp5SE9/iP
Eb5ol84s7Xg7vNuY+IVhERElcHmMEkGe5MyQGwKdxJI4BWSPqdPm+ICufDf14XBKhY2vMg6TAK8t
PwEQj8w8g7AOdrRNJRi9hq6QddAKZKjJCU0d4OPw1jvzORn2bL3/p6eUNXBjPn+kV6viMvtiO5a4
nNsMgoaWLcAbHo5qv/Xcwac3F1RmVJmHqNR2mSFg5l8uVaP7Z/6ZWDfpmyV/HwobteJFwHW66qub
EgWO5MTVe6CH15/8xVZlqdbMrWXj6KgZJNVZ0SbHXP2mjkl/uo3Rbf0VMGqjx1oek7ViUwgzKiEV
/bwUo2oDXGzYSdW10TH84NXEWQ6UzaKNjNx7e/12xfcy8k77wS6/Ac/9LbASrmfXE7myzeGBJvLe
FKDJrXjvpYh4OzR7tzjHpUcgFIIHkaLzUEuCkaTm4zqsN1wc8x+PlbJ5KQQt9YLa4ugCW3uEGAFy
RPtHmkOjCQ5BspCbjbfZbFBsmp3QzuzWY5AEu+4ZGZEAciPXpKpfGv81A0JCc72qCWIo1wtSxgiW
TNQeMM5I58L/jHzeHbTthEqX/yfQOzCQoCdD4H0UZjms86m9LJxqQVKH6ISCScdJln8YurLFaR4u
wd7BZJhGORCpAXqMp6Xqyva5p5y7x1oJ87Qe7IJotkIR0Skc2UBZNDRDtrtkRJbMy+a66xMeYkW5
i0WOjJEy9VasYQw3E6LWA58MAPDPQKQ5wRgBXBfAHJvjINdiDaUZJryOyusO/SF7Anbi6bU+r8nN
3iKikjUG+4TZIevhfdrzbpc8d/u9/uFLi/i6MZAOaO6bAAJB8CNTRnYw0Yngq914AMwyxNoY7j3a
sjfm58ZhUAWhfiCl77mMA0xF8MoB7l3lggcD+urMfAi/x4xjjg1s6LNigwRYfhPX6SL+9j/DdnNL
QWAwheHkx9V7K0LQbAvw7fAhjlygCyW1IyRXN0gGEQjb6+ZzErYFETat2WpP+NI2y9RYiCtCjlGT
OP6FQViDNlOAgcriKr159giqW6yLyV7lkBFASbYbpsQxCquioN6Kehqimzb+u7IG9CBxAsSWqbzX
aosD1hUL2clwc7WBvtZMEXmJdO7rbixyMHUeV5k6F64IM+gxWkPlwX2OAH25nceGs3xGRQHeoLGg
sJgS18QGGSsgvZh2tuT1QofyW7WBB5vYzQ44b31U2w9KKPPQX+xwsHQbxDDdMsZQW+TJwucD0CIS
jxv3EXRk+aclkBu7s1kLIzm5CwV7ACuliWDjIKWdCW7zFYujFarPK8AOyaJ9jD+UdrIOkoYwWsNz
VBXejwtaPWMSqfddyZKExsAJ42AZsamCIVweh5iHceBkq3ckHd7yxZningTT79E5/Cf8nK7F+qNu
RhIZ4icAo/SUXSaCla6jDXEwLfsqfaUhE+klyz8sOQuQGgXchlb/qVJz0JZcYpv05NVOGSx3hHON
gEVfn868r7LV52K7l1VhkIlcxpr6Lxonr7/+A94fGl0f5uwgXEBIzeE0yQpdIBw7Q5oO32xdlqzH
lGMdGYpnSUvE84uYP0DtfbyIizpDJQlfrY8b9ZzZv/GxFzx6tp/z1GIvK0xBmBGTLJR0aynFfmQb
KHLjT1ytgwho/yKX8w6ekfxnYAucKLQg2QbeeISviKuwGvvBIfN15do3txiYyMf1tULt3xoy6goK
NWP+dssrHqqTsKKH3RJpTpaZHoaCt2wsFNGybZBctZHX2Qwub2Zh740MiXnnYp7vMV7JM/b3Rkkf
kGXql8idcu9nD3H+262/kF90jBx9zVMWONfAeQrWqzqF6VkdYGzznv/GnuhdSTv09GuYkPfK6N/Q
4OU7RSqYYRZb659AXNbufoJoKDizvXvyq0WGRq8/uXpwaX5dHxyV/qeNi1J32A6kEm6/FezICdnF
vuP4XXVOUnbalZ+u768ro1K+86xu0awGzBRsCV5u+JZSGgHbSJrR7of9eZfLXlzFdWnmFeta52pP
J7TotR8wJFTtiZ3aMCKmnWKJdiXiBwtojRTTUTsC67bJjOdQUNE8fwQyYTpoypwr7Rch+Fg7Qz2H
LdFv39FDxbnxHhookabpz2VIjZYmEVKgataJcOG0x1inRTMjzcGiyoPMydLUsZp1E8WkhZqJX71E
h9CA1TAjqkHy7LJeLN3ZDBNXhIVq902c8Mlq12Mf8jU2lUSR6iqOlf5TmXD7aff4PJiEOwvwKTxY
dVxpWP4lFEwQ/fQQXrZw5qFoUBWd+KAZuWYnbYe6wJ8DK6RHtx/VULNCRqVuV0PnzRh+tzc8a4Jm
JRhEw3mpPROFQZmaoamw+Ap5cAVB/Fv2bcogFe4Mry/QIpNfpfomyt5ozkLZmzJRUly61aOWJYOY
E9Ws1ggf9fd+cwnYqU740h1hpoNyQUlOVIFuOGGwvUta7E3+VtmuFKVDyXaSbUn8IKSigR9SMiP2
C+jlKtN/4gSfgJNwh3+8rYjNpsM/qXQToVaPfHmRu/o620RdNrC9vNAkNE5zXggbtQIIlMgnGCxa
B1faeZCTJrPdS1X9n0kG3ZwJtbPONbjd51CVWhAajnzb+8GcjFXx7RuPuboNyaxPh5cGXsbTTzfo
8AaptChRGywJH+2GG1J+EP+8eQFJ0uZznXEv04y9HsaYL8h9+RmczaXT4eLYCtRexPm+hGkbLuZO
TzvR9otwi7oUEWNz6i+qQXI+OGyGDR3vNwUjwC2HtlSJP4p5AappQaQI0qhHkpqoo1Yti/ztzd3O
yczcHOgFalvCP23Bk2TAKXoUX29uPQeaUzKjKCY7CGEle8lr2LFaOrIOsQ1ofSG54ffELIrBwsWG
peZWvQeo3fAyAq52/ez8xvY4TaVV1OA1raW3nJF/MATH6GxcdoXicKzFeBw48sXlbRU29CTnGZMm
o58r2YKYMbVWUMktDndwmwIhB5oEQ4k1570+DfXNFsy5NqRjR+j34qMp6ao8dEtvvIv6Ofw3NQGy
SL6riozYT4hOC25BV3sD/lqukomfVwcHmZEmeEQGkdYsOgyM6dqK2cQoAD8cfaeiIP+5mMkdvA5N
WEOt9i6xb9Ivu1m/U2wzK0PM4FoTd5ClD5kdwbWxcC8Z9kvqaj6cXO+u1fN0Jpd243CJgTqco4aK
hn5usTAt4ljgkusa+ThwF7fr6pEtq06/LfKGLEyd7EFoCQ0Or5pHkqecyNExDXkFaoD7tVJ4p+wy
MCSxmfdf0QmBUHeLfXGkBzeRtFKWf9pgh8KOrUL9uHaEuGWYlkktrbn4ouvMg3wCCcnbfmFna6e4
zpfA6iMe4L7LgwoVpdOQiua9dsDk8R9WZRnPRznz3so/GqlxW42CJJY37y1Rytw9gD9UljVZ9sdP
42NDkbDjAmePJQhm3i+AdrKZXntyaSciZy1bbWsZP1S2PtQ9euDjqGXbSipfeX+mMP50UY33Vdq7
Na6FSCDaTcBby7swDaYQoOI/MjJjiE4zveJx/OB/b0Y+bgfj7J4gUADdMf3PkJeg3yxw9SJ+GGUD
FGydY6Jq6qBhPAOXYKdbOwFWy8suVzZytznGFI/tyEnFz/JDGhfUo4MhcRbwPhXiPSfmCFEdvbA6
pgkpzOyCoR2dfPmhxu4z7djdy0abjM73xCXJFndxAhKOMVA+xPo3TNtWJqokNxE/CQIfK+0pt0GU
QHE/cJNAPS0f0sUFJxwVLDaQK1naoJe+2LUVDjxI5ebLUvP/5DDGCUUwKVywIbRLgKuEpQOdG2Bg
DgqvXuIyZ4S9PRE2zGX73K8A/RXqxLx9ciCBP2Oi8KqfWBVM1g2yHV5M8trFDRDnPjuot0XImLNX
VoKBjMtm9ZaMHDlo9n1dM1K+v4VLGoE6OjhTref+nm4Znp0FznnMmUDmWf7jsgLk3yxvsMbKCQsc
CznpYVdJ991VLTWPN4hUvBgKb2BDkziF4on3x18mjkmloY1BxVBlJuebm0TRKidPCgZlD+9J6TWG
Z8RDXcNy12w6W4tjA6hIX4X+uWg20aNlNAj0m6H7JLqefE4C8LBWC2ysK308bO46BpdftTa8xSu7
J5j4847n+kcWEu1OwA21dj11IgEATgtHSlCWaykOHXQ87Lpik4aCxn9DpiF3KiQBL/nI5yIyA8ND
Vy94K/t9MmZsOt1mSwXaEbqPLU4t3te6jtlzN8rqVg0TLdlslPrJ37H9CNAZ4k4rox99ZAxhRnAD
jeTXVJDerV6wyVyaeoMOKephpj3A5+e6m/Sr+KAWArfWRTqEvbm7R3tmYYWAhDjjFSfApZ+uR8dh
fUrI5B59MMMhfHFojpOzoWID6ZT96GHjheEt7QBrBsV/8sgFAF/uT/8i0hvOIBHrC5opJeHph0/P
xJg8axxTSt2XPATW1OyMqICa7kjBNHy+GBeaReYfZXgibRdtbZC6r10JegXzTx++UVDfhOD3cXME
J6bg7wNGaSVgFutctl4lLXg+8kq/w9+OM1mg8sd5r8uIY9BZJkZlESUXr9tcZdTJiF6AXEiGDkGP
qFNamXVtCGmspX8JDYnl6/Cg3ZABmy0Pu45TWdLhixCj2PQum45eXrxn0F6GSMnXA+AwUV0FLtJv
UfMthcS4UIj7Vo+cJtumXjhv+3GKqDxw5ffsQyEsYLpzpIp899BKSU68Utu3qkgDPhaJGVp3cUwA
GPWe1UD6y/c6ILlhI1vMNchJErxAKPZjCm6d//mpGYjUMFV1nyK99OUbIEzE2EogcCI7N+TKiugs
qG7R+HM0sCP5+CpP5mR2Q83UAUtT15SzIhMXTCjHGr1oKrOaZgncipll9LtNU2fewMnNv1VTv+0x
OhUidPY0wiHLBKxjq0VBuue6BPcSsYpHQqCtKQVz5hptbrSMCQqRk+0k2Kki4F8yevX2uQXiMdpN
ChAbJLPYelz5UrKpYNXJf+y5fw7Slyw0qn5RZafpQWDO/bSrBXdvLLOAHQYQEDYvN88WANIyPwJJ
Fugmg6TS3sCvbJAlmaE8Iaqdca2vPnTboKRslkX6NMjmVsbx0Nuh8ltwlB3YWXgP81b5I0Rh0aIH
h0SZYrPwk8xS6GyjGqjbgToOnMJPglg1KKxl+p+bf1RxigdaVkPOGPPFqBGHoB2rwozEWqDK45K7
7GDKcrMh95tIOHQ7v/lh9cJrTRP4hDp7R4MLL7ydf6M25tQIpd7H2BntvAZuDPv6umG+/zEjos+D
3kS11dOJLESLa1fHE8F6eVbZVLQQZSkTtJHLW38qFnhWUOs+1MFNhO+RJFIurV6FpfXIz05hlODR
5GIlEpwuOun18ghCOjheBKCErsx+7WIs8PCCOqF4qcly2jJOIXEpAykot9gOlsD8BFbq2ElBrpEz
TEI/eBdHe+87oRl8p+B+H7c91KVe1Dt7ENHc85qdLxBj1s8Uc4fdsjye0JtUhXJPiXrIdyzjuN80
nHf/+o2QsWFOVesAJpTbMG8dtHVCmV8p7DdyhemYJKbK2Va0rGjEN2VaMRbP95b/8yYgcEvcSKyU
RYBMhYAnTvzcbWGd5HHxRDs2Di2cWbkPdIPTNMlGZSGN3kc4E04ARanssLyauwdyJaXmgTXUzR2c
pEHkV4PtMTwsk/kxgs+c7cZ30mNGu4rPbk/B0LK9j0SJVX2888cOtojtGCEULzsJzCqldC0KcyH7
Yd+6/MkWOqyWthIuph+KIlUjUJ2MJQpElkVHaCGKzI77ZSN5hS0h8eAS3Uj3CV4MtjzZPK9BCYKM
EOyPixh5QDweFfpGe8NiFti01kvJVGqGMF4sqW3wq3+ILZmotr2WIRjB8+gt0LkdJZyFQ7jjplES
tG6732MROhIdJ7Hs66ZUITlhpUrxF2F4zRM+IaW8XqwzEaEoMMYRwJBbnRqcu65LLKrAU/6o5y9E
hH7kpgThfst7f3/Oy9PO7fF6BDDtH6oIeW5C80Rbuzqjud3yTJHw0naFiLf4wXLZi35a/8eN79Pe
G9Ff00gZPUk0g5VwReKqshQ3hM6u7svCeDp/ODmK/qcQkesOIfjROEBcOH/Ar+MAF2dyhgoy21tv
g0sRCdRZ/tdZJR6szXS1jOzvYWHee9+Z2VpTxUaOOc5XbuV1C3uowO099ca82U+dFZ4F5/ZUHh7/
SY2PUUZbm3vE+zNHSE3NU10bakgJCrp1D5nr4XWdHgKyxOCZE/fHvAovrPL95bT+fI3/0ANrt9CR
P2AaP15BXvfk2gUpCZ8aAgIQOEyJMpRCga+NDxQOg54phT71hOuYKONXjpJoeKPDGIr4HPZ1ESF+
m853UNH71Bj3DBhsotdskTVp7YQYXujqUDvbfri8aY8cuaiOrUSUoXZvDYlqWeGp0HcoOocNUSCO
wK1sZbFMCwZn9Mp1YcJymV/vRdMsEN0WmGTXcGvf7Sf9+zXc2uoohIsm4IUMpVa7O6SmTcLYv/bp
187bl4KUl7GeJl4oGGxkJrhUW1CjYgleDBGfBy+PQcbgpNqAtHkIJS8l41biaLvhnVw7ViNbWdL1
5vTe8WC/AocJS6auzP718Xle7Bd9fetCJnuzmWoBrPDEzo2wTDbLl+0t/zjKkQjLygQJcOifGPkP
Q7+uOfVpVOSJ3QxAbwCrQDQMQSNDN7mdlJ8mmN26KcArOKkydN8zkpzAN2L4JMmP8xvSTl7RnCOW
iYeNgPP5FGjoXjbOH4WNz140stj45aXT/IfDTgSwQ2edzNAmK9gAw3hvvZ1gexaMD2VAE0XEG4RD
/HfQ8IKO9rrv1dOBnr7IFAjSVgB759CBYVpnGCq0569fnw7exv+4TOXjk0fuZ/sPAY06Ij8fRl8M
Zybd2r3IfgxbWtguZtwBiqm8Rvvil0xS1o7T2HpJgpfnGpwV4Jh8ptrhD3vBJlAAKP/H9cKLiZwB
61Qf4Q25LuYkQujMTAQ/nOW6HFNsawv+jo/DO4hTgHW8MBvV7/xsDiptxEbIzd7QIrmf9s56+1D6
HDcQ+Aj08XRgpdyhFEelRltZB3d08/HcYHtkouHhAaZXm/V7IfysMtf1Yxo8/pDlzdhe3TQEmPsg
/FGjKIyuFDoMLND94Poy9F59xDhUF4pGoJa4kHZms4HWgB8a59zs72aVPTJVRN7Y0fpttTXPY2Dn
newCxlZeZvMCNwzeGAKtdsQVjHIEIqLaEhAKSvZf/AyjyGgXGkqlfW4/tImxwLAVSxSSFh+PlGTF
kH15jSi/sujYdbImljsOnyFbZpCPGhDTCZXjIv/LMDjUuokC4X7+WWZq528Ks993O1RUfk87L4sA
2kvNnrwjG+KDKTDDulTDt1m9Syc84+fP0aWFQT6YHvfOcVvoiYX48tkpZkZEgLH+nYTFqrAe0X5S
uIJvWqEzmgcIfcFb+UChVlrtJsm0KT6+jdcPLLSeUh5ukP4KLrO1MCOBeis/oM51tcn0THMuBSI2
gP/SBBXS1OvoAI3R9GRJ7UnqzSMmsZ4tmpghVhb0t0MU4Hajq+yhi/neDEn+feES75+3m7ArwwFM
3y2sqNIQ7UMXSPZDU/Xn44tJr5G+PUrNko6Bk6zpiWL+7gWwYRrr6PUK3ZlkEf1o+Hjw50MZ6vY5
Evxh4JL6GB7o2+WaBr3edrohEP3+yVvrnHWYmZPB6l2kRHfPfBlj9HkG+OOf0QlHt2mUt/0VrU9g
KiCBpd1RLZQpEnxUK1WksNpWftKJihQCg4rN8QkWcnm++75/2DSYEfFJ8wa2YUxA95YXkjphbc9h
PStytAU1wxgn1hI2yl4Ee3A38FIQ2Y4E7C6C5DHOr0zAbCM/UIKAE9rznj1P9+vW6sMSNMlEZvnC
v35eDkgxdp8CQeDuZJkKQtjJ9kxK+jVlz3U9OtkRx8CMRARGNcztBmtQgNrqKKHvOWu+BMJ0Ek2w
gKKhntRRws4uwYMRU3rN62Zhfr5L6rsbNP+D7WLu9Fpr26iZ9Qu7SS3tUP94a4U1PZ+FQ+6uROmf
vkIANydvqTYj/p7zAoyoNU0DDCtw4g0QVfPropHc+W0rfSUeOELYE3X3YX1gZ5/3oVukcEjJ+93H
tNTeZzZwrojbFYqIcA0cFBwibcei3ujNOcBtJ7AJXUZgVBaEXZAfEk7tEErilNIIRZhRZnI7cyI7
4fq5e1GnLhQXhE85g1gshvtLj+bqXdkJ2NB25ssXvYt7pjBUH+LTRo3QTXX9VApLySsBAgtrc7wg
j8geec5FsADGRukvhsUgFRVKdKuFrYudv18nmSdwA+7pk5Ubb8XgLerg9qMkzqFiVppS4zCfbbSc
+tmE9lTYFaEf9TjyhC7DZQendnW3ljAG+yULGbii1dqP7gkYPPKVagJWZAWRg7QWNTuaaFGFufl3
wJd2p3MmOt6T2+qRM2ln6aBVEUeSBgjXPpEBxbKtIvR+Hnb1XrQCcBYWol6utTFnDfP12ZXIHiZg
eIdrVQ8R/5oqoH3kLgejujpF5iJooNIbcCPshVdNfsepE241kNwJiqAJ3STVkkpSm06rEsa5EGrK
xpJiZlORqxYatNUWv6DY4ph30g6VOEFlGPltRRfoo/9ZQvq3D+1mZwU5VO1BR3+Nkdoybr8U/Sof
EvMLtjMoiodI/6LWcMEarz+8HBxoqCoIVuSUweUX1CQXEr/oazOqUEDj0xFTuPZqTv7AsNxUp1sQ
YBGPGz0+E8K2zxWLdnrBdkqfCflEQp8ljN5f8W6aLJLwNGqdjYE3WhusSHorMFNeOr63QPRW2BQE
TcgjmLTIGldAjXc8KXDSRgxP2M58WVWYPciyibOAfYJWBKphKgKHa9C0rvIC4vZwVNqXczB/1qQa
UdiddjWbrrt1oGjGEBYdy02+6bl++zSdGQrQ5ZGHQbxisK55whQ38YRWrst35j3moNVrlEdiV4NC
u4xWUfdrFc65+aHcLogQvunrswTPIu8kcgSq64TVnDJq1rzBBczgcKFqvEPBqIC/Y3sdJKvi4Evs
84JGkyfCh1JsubdtWp1f/I5IvzvJM7WvOa0Ws0d/k0cm06WsVHMqLyUHedPsr8oB7AzudAQLZkWe
s/dN5/9IivJMr4LHOp1C7J6zWWfHj7T1MCyuMOUmSG2NVvpN6Tsc+IIXuykpF3IaMZe8xGE7+XDL
DU37od37N0b6SSQIS7uGsBl0O+OEh4mjgVu/bnC5WBK0QAXHcHoewxc+6swhDZQeoF115YZc6itZ
NajaznRQfc88TczKVcNh8SS/i4hrWX/6RCsh/GY7sWPdWv2MhFeT1ZoPYuAWZBWqnNXLStsX98Vy
wdYq7/0jNzST53hJ/xP3LrgEWgRQldu5OmwSOHcRkX6KJvllhXMV754rNzn0Di+LUpmaQ7PzDVkI
WwnsqriJdMZVoGH55EZfdvymRFgHeyHIMBOf4H5jNvXhA3f2q8c9d7fek3ZrHb8SVNkt7xIalzX7
95aFuanKbvHpO3BM3bqnRMOgBQGmZTCMlMezrxtjlAqqJzgCf3S1nOhvQ9gjOCRFMi+fYmkUaUne
541Fd8TV50OpQbeBakpdzDpVO+7arLdSGywMvwaEWtCn1hYTKqAPjOaCtU+DBjCfhncR1qTnMLhd
pi4TPHXWBJ/vqy+MAoymPg1+erjJfZl1P5TWOhnPaVs/SVR/OpCuChFsolYTQDi7JS2f8WAqyI4R
ttEn03cUBtNH/t3p2Rb62qOxeWWCuUK891up2QYYwzI2p5GwtgnimbnQP0my53e9GDt2OK+6fsac
vjBhfXdvnNO0S6OyOmpB3qe4WerHV/oXPJppBKN/4SEQXHl5WzPlQalSemnqdjPAyEDUrvj3Kzs6
XBVZJWU0Ultmu13h7omKKGt4ZFLQUcz0nasZwrQGAMZDmskSXvO1pI3Rrhfx8exW4sUY44BhukDU
eZRvaSwtXYo/Cwl+td7pVW1yB0PsaMO5LZJNgXcrCL6wpXLugU2LIuMuKm+PnP6LU1Yf4Z7dsQNA
Tg7KHy3MJhoNnERKa/LqnbQ6NJJ1LFnBInFLZtpZL6OLgXm9/yQ7qREYl4P9kx8NBbf3lpbzLQjh
0jipm9tkAj9OHo0L1G+w0VdJQIIOAW8el4jF4P80tSmkpJki/KDan+fnMZwRl4ZUQk1yWkLTvV4S
J6DSusbN6jooJOt/eN3NaBZlfEI9h8YrESeX+X9nWLuZmOKtp0XOkaW6bLKiAz+ypWz5whzmTr8b
Y2+Ca3eKBg8CI/M3ejHP1J3oCKT9ea3KWpgEdr4Ifejn1guALJvNxozP3ayPIV9GFTiDSM5F+y0f
3cPs8G0QqsX+AIQ2vdVHfuoVcTKNh5IZ2vHCOZdogBq4CPL4OhycjOSkZwYmChmnoMruEP4Ls6/M
3xAEadP6xx5Kzcj3MLfRFsQ8rYeUXBFh3S7++fFv8LsGYc6rnowRvmxCC3y0KL1JHqrzeqeVGupH
AWIbUz76wpcScBxuAyTmRVVI5PvU/UZHi6RIO7e1xskniL4/Z1e68oTPNVQjWiZaZdU1PYArC/aK
LMpiaT8+B5aSLT//0jhLLIkVgpnNHp8MAMUOzcXz6ymCMR61QAOap++F33bxBF0orHmatBjIXaSB
u3do6VBXdg0qAgANCVlSnEXArzf+1LTEKSv2aQYia2nbDUHzPvSfjQ/uU4Vq5h6wr1F/XkKqAoYY
W4zofbnKzuo1Efg1PGiuBKToGUjxpaYRyJjBFOlN1ivDZGMj43WXdIN3LfL+Rc7OaalRizQ/02NY
uN3xdg78+acXQi9vdO00gMzOt3000rO8JI+DBT1kWlE+5rnAi6PLXuMZAxXYdyKWCVCB00zIVQgF
T1CVh1sLQPTJ2/RKkV6aw6PuXzDV1rQOYN6yffdOEd/a2qYkw89oTpdFL3Td7LKOJIqQXWYLyvju
TkK8WjzegGhAVTj1EdZ61pOCmoCVBdYVjmshKc3gKhQHf2p573cNLum5IztlcykRk1SwSzLWC5LA
7+ZK3BVi6F+pwv2uaWERC6G4u18dJoCuVbqGto4y/CnpbRrlDT/NYR8M0l8Smls6Q7d7uF+NYsyy
MuvZemtmzflPxYvaNPTAYiHRMMyDZd/uzW0muqQxTh+DAJZLf1Feqt3Z5rWcNQV7qvJuaOO7qtQd
C7YLuoszqTZV1DhpdgJ2ZfcaOxDrCrkChc9LZmkJk5ZkJR07uBQHkMFHakT4aso/qbzuuuMe6wNb
liE+sh+8DTo0i01v2eTplGgswwgOlF+NqkqJo5vAlgN9sw9WUrFxr7xHcuJGKoPvUCtbseczVf4O
KTikAwuKOUtoCLt6mdqTPngysnBZj8w7S3+VefEq2JO0ZDZ7gf0EC6d1WLQdzOisuEf17AsIbNTU
rs7xIQt4Vv+MbpvqVUQABbzgGqbeLT7dGre6Sk0gN2kypEkNKcNnLweMtWumhwbaIvevsvtHtUXM
s48MUJF2bXnIZXkyEzVHJZb9/heNW7OM53CO8Nsn5Vsp/M9uh0e/kVNy9W1qNFYYZXxAEaaLg2s8
hOIMXkvMd7GBdLmCn8NyLA4tc7zmMSVvYVmqT+p0l/GniVxs1H2Hpz9hiYEEll9QQL8/gZO4W9fz
8PFfBlIvyuohmdUX6/I1tTAEVuai5O9apPd6GXGB8t1wI5sDuUnhTaWtPNPX5uKB7vZrCZ7hsA5/
Wyq+d36pDzH3NYN6CmPe2/5R1pq8ARai5cH7e7yVTX0hew70r9ogi8Q4S4TPcnBA2fWcslBzXhss
IQh+jx4u7Qtxu/KPM21sZZEb8lqZ1/L5m4cOLicjcG9gx/myouYyA6eS9pq2DOV2COUfnf2qlo3D
92XjWgaVGI0gNAmLfXEntqRU6dnR0pW3V9Z9/CUhUyW158E+5B17uNx6S7EN9P2y5effry6CVj+1
Dn1MXoU6s2+AXHofZCmKgAdyY/7yTTDzuDJLQQzUIh1OSfRLO72Cj/3VORCX5MSMdX7RGMjVXEdF
G8nPwUK4JsQ932PHx57OtBQ+fMe14PWRgp6cx8d43KnIqwTB2mFoHWNbLN04jHvg3ilR+/EzfrZC
iVR6o1aEEBrXfG+kCGMuuwuSWijuWSD0jpZYp8tVc4BgaurWMD4aHBKSCaBMPUjq1CdlpuCX+XrJ
Ss0ZnQIeNv8hnebcPKHvz2Zt+yejhuBfBrBtvlh1fpo8V96KOz9+3z7o/7RzCldazsuvKl0/fn1m
LwbJQKwTvMDxFL60UM4iJGOD2q/PiPg3JOsm8dUz6+fItqvpjmX5Kww4TgQPKHYUE3KS0pBCnFTg
cNSFPUTQv5SYeITelqzkjrbfd+3Ss7ON3fmCKa5keHNd9ImUQxkVF03VnbmD6IPHrG5WGDz+t8bL
2HHMgYqo00kluwL+9iiyojLbSN6eifTsNlJuLYXmhw+QpbYrX5cv5fbjSj6EUBq9jz07vmhpUhMo
ZVzREE8Q/nQaZ6cq/LJS19hJ6K9Ek8xTE8qt5oNde91WcGD2Yq5m1gYxNk48DrbrGBV3NJN9xFjL
qnHEssub2sJBh+dELsDPWoqVwi9zyO7XZJD2JFwTYBFBSrvB0UTYhVgt3Jnfd2Vhp3e80gnVF2Xf
/5H6XEpc4CvThZlbaFbxef2xKrmBGUQhy1COmabYjaLVkyS51oSCQn7tcgwEUy9cj/wX4+figfbJ
H3ecUvq1HmtPEu4Um4FfAs9Yx/a1w436pfCqpX3L7s0+uUzjXJevTanjjXY/46hjJUrL/zgO47Pe
GSDRFfqRPlb3dpRS0OHdLounI2WNJIn/jvAp/8SRigtB5OR9K3VRL0OHEhVyvDMlsj5VEKiWWzAk
0vEg1Zy75lm4mACxxA2yEMlNdAgg8qYZ6x4/fDEQwKVDq01KnWM9Tkvp8bgS6itR6fD4ZidtdfWp
oNPvj3vcon4ZSpBaKFKdiyu6ZrdOyKrb3GtQrPxmzumXKMeyB/+9Kzs75KfLHcFpiiKPBtLTC1gu
ZD2oQlBmfE2hB4R+uNEQoYhrDiA6aCxFFRETOX2Ax0wAZRWUZGHGzcWGyiDKVWM9kbCLJLCoeSAW
ySwyPkwIybwcktQCSGbnq4LIoECn64FSYe6p8gFfn5TQo4lTU5/W7PGb4afikn9nIviwcP/Ye/AM
1suaQJGgnhJSOmK6xilEY7LGwufZV9mGAjNhwzecoZz1mU+uBO8Yf7BOM8rClHzNs/MVRj6gksbb
mGPOsw2xMC3Ln6bxCSfIahDm5ZII8pAuAIkZUO0tG85b83fEMj+jvDTz6XamZi4XJ+THdXOsi9Hc
M04A2O7c41Vp6E43Rv0EnJtt1xgyOsWby/oPLsz1BzemiHlkP777kLsciYYzBguLroBN+uP3JSDJ
PjPDKb9o0Pl3WIqiDe6Ik8A2BCJ5cCrPankpUkb7QoMmc2547ESxtg2I7R4Dz8BkmUuqcfQRU7xI
xv3TNfFuVPXPlJlA8tAI2mdKTSHM2VhgYXOL3bVDyitNXABnymAeIENrsJpYA7L29WSOs6LiLQoa
1l2H+FwJqmAypFYmwtGQ5dTcOD/zfBHoRB5t3tTNcBiObCQz6xsp+lGXOpGe/XntCLBebTfOsQ+K
Q3yi4D3krwIJmVPt72u9kxdH11EZ7gQwjd2A/4o7Rn134kvWCiLt1pP6mWuU4JM5olpVJiPPaMZl
jshKtnetkK9sgCHuLlqslaot4OElj6l2vZUq/6nXsAFGXQIk3TldTsFI2pF2LVN6p8ESEtr/J5QE
Jz8nkPcQVACxyPHWPLBoI+MoME1ZcMxE0/Sz52RWKkvFkbFan1SDczjnjT7D5BFLDWBIYzIloZf4
gq3gi6j9jSMADcKr9yMlo2JLIQzEiYYBdMfPTSROJphT+JphmxnselH5KJpm3/scp1CQVB6Wa42n
fF3U5L+uOnqhZ6xlvVJUv0dug0nZx8zenp833eG7XOnAI9yt5TuO96oOFcXCv1s5rcw424Syivwi
r6aKm5nsJQ7Ub4gYKiXQhF7vUCqULz4lhVa2hCCUPFGf/RcdGTe6tg5dOG34F7d3mkGxDOJ8uYLH
8mE9nAEmBQvmZEdA9yh8MLKqAc3Q0REs1wHnef8fvdqf6IKxumfctSrf94gClpbU8Fl6AG6vdvES
ye3E8mdVJccK+emajOrKV+VZT9leB7J3Bx0oM7rvpS7OxiAWjCIUPkknmt9gMReRUSDg9bQsqSGV
GKB/ajklGL82xCCYvvM0N5n8cYGHSqV6p/PEXhQ6SoUfYMdJflVeg24oFNREF0T9hHxaQTzJQ2wj
6L050czJdsX3jyZdm+HUhTA+p1qdZSzAWvHAWJrVPPRpLQDNRSpDToSxVwPTKu39Vc0k8RUwCTkM
WIV0XY5rh7UlIksH065bKcR9R//3KoGIorMLVevLdd39PoOPs6yRQBCxGwEQX/0crWb2Xm2oRlEB
pruY4RbkJuZuKowox7e3Kd7io0SnMnuw7wVP1qSXGuMQjLhydaBetqaEs3XDzv1EEfDEir0kEthf
8qRAlrHGXi6Dm5NqqynaXgGO4fiVRzRZQ/AWx30rINhIU1ad8AIP/UZ89ZEUVpdXL23v59UN2E0v
gHRuH6lvkGAUQgaT+WYu+H0zyYfqOuICpl1jByX839fxpfVBhhjUND7frM0gOp6oG8vmC6g8ZkR7
S+cU3bKk5nVKseE63Ondu375Dvpgx6mrVd1/8bzvNO+VO91DX/wVTR2RWyp1jJ6XayIbdZz9hiw+
I8RVnlToYtxQKIQkt8MaZBDjzPb39ULGBa2bJLlOiS78azLtQZIuBesSkxazf5O++GSPvywz4f/2
KaGLJ+/lx59QUEZUrbjPQADt4uASoRyI1oBTpBHEteQ6/1RAVBmKMY7ISqnwvX1NTpm2IJII0VtJ
y2ifFFAjYhSRlnxKj7Pp0j/QLz6J9wqrDvfNORacwEr/5xhOYAJllmaTD9mbnc7cSeYLnqI7IHI3
tVORA576SbzzYXT6d8iPYhnfhHypsVHEHqEgE7vikABQg5zRyXZOhOeO/m73grkcvUmU1LniO9wb
XIxDyew7+jTpTWEgcKnsB2p4WazZFVsyq0SN9zyPyrx89rJcBr7GNGwIt3+3BOnwY7qo+fZP+tVX
f3y0jgpGQFlkIr8Wign/jLCxNrUztFyh2vxR4zW4ykf0nDCFIWhRQk4To49xFFEVFFhzS10iPLm9
tONH0bbAsGH45X6XofDStxQzOU4m9t6w8x5/IELtWvzMURoXW95sXK0nLyWIt7IxS02HfZd44F5H
b1h+DCw0B4JQtVy6L390R1SQr00TRLKtsU9UAd5aVSGGeiFBuQKpnesQk3WRSER1liohJ3WwREAL
eD4RliUH0+Aff/BoLICVkIzp+zWHznBX8hLle2hFdWI686mTz3XaHNsHtbjzaOlhiCAAiFOKwRsB
hhNi0bVgPL6ziO1zPP5it7qfvR+S1jt5MzpG3CiB77rp6eXNmCvi9FJk4bX4VU7qrlPDHBixy824
Mv6idPzN7GzKnMXtpL7LtaXQobij27vi1n+OSWSq5jSp8o0eegu1BtBnTuJ0eZ4OaVLqW/IDPCY1
quZQfyk3gxJMTqLRPSLbxeYpTEK4CrQnEE0MTm7mtn9HHQavPlkw9BATZkWKHHEcVhuGdNGZ4Mcy
Sb3eeyRDrqbJ0U876knXBEXAyutWXZalwZCRzk2/LjOvNDxFM5vkL6XB5/vy49m/3auw47jR0GOA
53A4g4qn7llHgfrGUdKbKKBPnqd3+j3zjJ6MEbACAvIDFgyZP3S4d53by1QNTNcawvSclkgNVgr8
OpHuurwQlDTHrAH6WcD3ekAz5QABFQYKOo97T0LAFssUc/JD1Qbn/hv5zLKC15L+FvEoYM/KppMW
IqRef9TAy1rsYzjgbXSoMzNg3hpHTwISI1MhIUoVxtJbnjK8/TLUkk7U8C0KCNCw/QGni/+eDF2g
eMTK/y27/OAwsJmt7YTFrDrT14zYzv8Qr0VfisidWnDiPPLbhshRutZxmVw5DuGeVdN2HSKCyVS6
0FPVjMQ1M0ub3kfIz+cTiYWJjsRQQG2e5k3WpnNTmY44R5hA+wj3McI94g4/XhVaICAhxxU1ZyE2
RouJIOxbvBn9zamblV1hgmEvWlvEnPgIDKhJe0qnvT7PN974Jjtrd8h8oeKv+ukd8yFJ+GtE9zWU
LPOGJ+Bw9GxfheFFMmi7RXK7oK7OnrTaLFHnb95y5Or9E1U2Vhn5KaIj7Y/RokOWWF3XKb5Kz6Ut
Htj5j6Y9x0a0JkQ5HlySHbpPL8ECQ5O01D4wP6zp8urWUIadfvsfoDuYWQ+n7IoQY+OvsIpAWCF0
2P71R0Kz3I9o7B6FoItW1koSt7BA/ujc4hUnTvdTlkl+w2ykxKVHTHIrP8RNhffg4rrCE+3Sobx2
4QmKxYwhpC9RTpRJ3QPpooSuPhI3xIHCuDqellSYlclO4pcwThzunyk7HglTAXZqacsbdgDNxCuN
g7ymgIwY9/LLSoSJwMf9evFtxwAcu3aXOqXLCQhw9C53YVSjRyOxPdN58aY9smHvHmVYHXO5703Q
xSCGG+xl/3aPSd58jdQI4Q4ZQcrAoK5S7Ry4aScEfFtVEMVcTAztOhop2eK8ZCZne7UrLnsmUcKF
CIl/0hDz2eNSLITP/dDQTlfy3/TGE/QJekMZxDGrsla43EmUXyyZBJGLHD6l05o3TO0+q0Pi80C6
3GJDWBdKZGZnWe4R2cJcj9nJ4XZ/HXtVZJSXE6qFVLCyb8EsLKaL0Z7i4rD4B6fYyUhbv70F7zdC
Bu7OPst5bbRTuqd/PToensFfLpwclvG3OpDzkpSHN0B6tldl6vvRTPanHZgkvXa7KWkFX1g65b5V
VMxCDvZy2DmZNbih7XknY26c3lMVmImI6tRRkByoKWPuTXQYO3tOCvBSbPEqyQVhqSPOBB+85IYZ
s21im0uxwrbcKRQbPahR9H/0l3YREUY88RCU2OZFbZueul4tG6KYFzKfTPW6thaIutnUcHmcB4o6
o8w2+Kw678+1vIZlpLi6Cq+Rl8OOZsAXOzL4gIiX52RLGBQ2d5uGuyot8RY6qMIHHj3P81Z0W+Y+
HwIFkpXiHdyOk34Wg5RR6Id7EcV1F4Kve8v9Z51jJpXoL0RVFGYUnBn6un9Srw5OimtnP+ak1f/K
s8uiX4QkYuIO9WrIFiJVk1XJlIsYvdnfw+3TnNYUKSO3EQTo4gC0vessPJoE2TDiBg50F7rRdRcy
aTT75JsZ9SuxKwC3qt1QgFPZNs/81kxxeOxY/hBiL6vfsmH94lsYW+1NRwAdeLUriWa0t2fAy1s/
Af0POgd5qgtOdhX5tlmUSQvoMiOFo4bFJAUANhGI+fknBhHDmdhGcg2dt5hKTtiyX4+uo+k9DVhE
O9udbUZb3Mu0OC0abji65ZbZc3v7hN8AIBwEBzQTUOPrSPSoHoe+mlTCJDl4DNtaYKs4BGolGGxk
u6gDFp7yrtRExeM5jSbjxBrq3oDy22P+haQJyEYF4nSaPsUGzd5bXn7ENdE+gFKlGjF855Vj/mIi
TFijVA01PR1g6YJYfyOjLWgSW+l0jX6lTs+L8X0RP4xFi2GXgkvFEaymU4X8d96mnziz13V85Bse
v0Q2fmR0XOSpdzX1nlzZDKwDAEPLUySFRRWN0kUprsyBhiLH1kVLNVXZYI+KzKPRTA/xm1cg9S7D
JXxBvzRED+XSf1MsdPxm/uw7K5b28elv8FqBkULGaK+wygpMbM8eq6V1vX+69QF9iD2hZKkICOAQ
5C3b0+rjernLb9/ATl6eGHh7F1QKQI9WcTcZ7YZhxTC9YHO6BrWWSbKjcas8IkgWzoW4RcoQQxKG
MUx6XhrmaQJA9NeUhyf0/En4TkcvvoEMRenRcOr45xQtim10s8zq7qk7wzdZmAxSaZTCh3ME81Wb
F1mkixlauAqfO4OEcuQ1aq7C8zM0SSrbcP2XbxpIlsSTf6CM12d9ci+FqxzuwGAAoY03kpyIXJEi
4kyKf7vtlxUhdhTReCCF1fpXIEWNJMbT2Fga050xmQ8fjU/qPdAvOg3Aw6YogmlAy/pDWmlIw3BM
/dYnwlMKOri0ERVjgqkzeb5nPYbxD78sUeHerq288leqIhhOZ2dJMRL+iI5A3iiaW4xddmvLb7Mw
wfVlb3Rd68rfbm0VJj4aMAKPb9+WiI3n1GEa77x+9NkQmPCyyszvyrnLSdDmlvvnIoJPxttffYkt
st4Y3oaGETUk+tG0dFRB95W2YnjCE8Vcm9UMvA41VmZtkHK7KnAvRwR1mMr8qQ38rXAxStPI8tRJ
DnWKh8hkRYQ1NvvxCabMVlRG6miR5ouqZKf65+pO5r2UoRdgmDdilyykeK1zTh30FH9AXakQtz87
6t13Ajlbgrc38cwCb53V2CfqJdM5lqEiNl+tyRhDgPTumMlKufBloLJiWPfUsjUNLqjXVOeXHtC4
hPTT/K8MxwlJyOHPtjvYXbKiVCT6GCTVfxXJOBfo/cEhNzxCEV/shW5xdGVjrgGF015mSNgwVP+Y
KY9Ha75BlFgESXa15WP6XRL08c1FyYRlEn22iYHjlRaU11DXpOLsGcCxuezPVbZ+DrRNuraQewrB
PEYmQWZrtoIG0T0VUdUwZMoFbRiyXVXB6zb+eg26HeCBARPPO0YxOePHweTPXofjz+zbGPke47hA
HfzwchVHMmjSApcb0NMhz7DmXbD9Kpq66MoSqpDKrIcXrZG+WsP3NJRhPCk03ay8Z7NBAozFU+EI
SBOvhWxgMl12LOmvqLtaQONOikKeijAsm+9GrE/MsbV6hZYFHaw+LIp/O3XgIIqVXhFYa7MIyYyO
HifqraMLCgmILh0oZ1mRXWqw7NLO0jQjkBNiBd79R9obsxs2OjUQ5uRg4XUhMwNIwEP/6sIw4oJv
ilUVnsVt1anitM/zGFBJJIPHD5u7tehtjUp1jALuHnuDwbAU0SrCkt02fChTF9mcjnd5NdsfD5uU
b39AccHbjVVn26uj9p4sjbDAO7aduERo0pHZOzKvXG+7lxIiNfPMv2MbUSOhDRO396Zm0WZXFt5a
EWlQIrq7kR1IRUMi+GMuSwH7eAHkTwUDWcKZcfp/8qx2LSyzEtuChe8o4X8LZs+du0ZRjE5GiiVg
i98yHnXaBrfe3thdLkYMyYUI+HpK80U+P1YDzejm0wEPuty6wdXZ+u39d7Gdr/Iz10w1rFVGV7Pi
e98rUAtRDclWQjR/LnbiQmhVljpHIxms/m2UTABqlm7pcypLGIw6/SmUvdh/8yTS5oz44YfCz0EX
GzA5EE6AYgJoCYpnzWnm6cCZZxznXwyilYm614Kk9FXCz6iC08U4pVHyZr0k3K98okDnS9nMsV+q
RMqHAEmMozxXUT6ludHhSuiH1LADxfgFPAwAIIevpucCHE1O9g+9AAp8yXEo17tJWD6rZOJgrknX
OSX+qKhF6r/BEp6goeis4Ruw1xTgBcj0LLelwubXG4MLxVJz8cN3wT0zSBZeMYBJ/Aqmq+4SWOuJ
AOZTsaYtT6IGrMbAdfSpSdYkFvbDh37BZya85wxr3SVl9XCO/KnTkMjKHE0XGZMqqDMxgamT+ydz
k9KtPG2obRlIKl0S5aQXO2xMsQoQCQUixl4gIKK5XsHQP4ozefDs8R7VBmPdKXP2xPOvRxHHP2dI
rgyDpvHy3R55CQqIcxhnqhogz49bzbC+sfTelOF4SSIIIe2BDfPlJ8mcTcDFc7fYHW3uKwYaibuI
JGntDX1W+bXueJhQBtmNhx0Jl/aPyc4h4NlqY+Ubup9zTnwwQvkYK3T9BUju2IrTiC6xB2GUp0Pl
NTlVPL2P2FZUuJPw9tQxDH/XUL96GG3G9OAWckH7jyOqvXqyZLfpTi6fVjwkN9rtdbcmlwsJTRFz
Ucep6V+diug8RrOiDiMQ3NPqbwSu/asR20zqYSlmlyHTjJCIsFRIBv787T8+h2wlJtpiE8wHU8gB
H9jrSKRZI6Pi44dfhFSp18oF4aLYxO8mJHDp5grKDQxyZO4g+7KJhdotTCYdrRu38LNN0z6aORS/
CbYibkq5vaxcIjsuQittD0K66MH+HE9KKS07R/irnVkTw91WGGRuukFci0Dm/V7Dkn2FzA6nWu1X
qztvmltnp4BvXIDvH04sSJV1EqIBU57dUFL2m0lQ4q9rYO5QjSap6AqETJLS8aJoHdRGonsyS6y3
7lWotPStUQdUU+7cSiFYb2lSivU1TU7oCRedBFspuFvrRgSL2Fr8+Rtko77qehhdK6EZNVIs0KB1
bd+zBWnTHLu0AUj8OnreGXVqB9jJJEel1xCjFmWiFG0WBcAIQ6wyE29TKDGVAsMsUGLqpEv5liKH
k6RVlF/Twtu71FRTjU5FUv2rKnmgWMzON0qNkLPZjFFFbx8WjRD9JCaV6t7a1ySXiMvmugNWBI44
N3GOlvIh3dy6hdcMOxTBnFVh81CD7TKkCCE9QLxNeKtR2bfK7tEWomkRpBoR0ELOEszMPLUsJ0qa
bD9JdU3Z84hOi+izzhxaUZPSEEizOA7xkGI/2EHlaY9ktXUs9qkgZ6//zNVIzd/AO7MGo7E57ZX7
sdUxqPDLPwi1blqpLua1qbealad7q7MzowLfQY6LjMkZHJyzN2d5ty8974jB6WwNtVnJ6vNZm8/W
SUWKGQk8iYfBrgm1tKXWCbWx8/n23++Jd1XlXSS/uTPnFs+yDQSmtwFnywbe6JKhFhcj2lJeJ11d
FG+6x70TjWnIo96tarlTVqbBmWLrSsX1md5mci9htQm39w07IEc+6zA20jweqWNzGmvnhqFeaNgc
jQNCAY2EP54qhd1JVUG4pvoDkXQJeFBPVXDNED661Fy7+vhzpmk00cGKgqBOND8wdsfXnTcqbEIU
weIGIDv6b+hlvRQSPQ04UtjXhltGddH6onH2dEdWZGFlwMmd/BxT/ArBVtmg0lrDeJ2bZ4Wt05Mj
ET62A7ZdjYEHqbRGGvspEtu18ksbwhRRCWKOcAb3+BuELoet0AEiB09DjTyvG7KvGeTIZ6hlVPkO
k5jiQ2NOqxWyklAbRcX88s0Y325S6nPGlvAR1pzqqvT04L7OS1YtKEo1b5rYN2/zEce3ywNV/9Gh
eP4mXWaisW67Fu+iPpkPaf3uU2EvbCEESEOyQxGxHMs+g+w16QkkKuUp8qdqDNpvNLfx1BlLwNq1
KbC+HsxaFy5JkOn4rH9n6W8oDc3C/uKFHEwyjWKJot+97X59jNl8Hl4MOE8HUxSEdrdAvk2IZJlK
zFXMFaDTqJ0/XXzXs9HZqJ41SgQqGCeMdBGHcxLcJQGoKZKW0lwYy6Zmm3paLPUGCixmmp4lZWOc
lzXRoi8P64CmsfawzeZLKs98umejCMj3Ukepm+bFMYwdkHAKLDHhBP6XveyGhygoDyePhzPpriLk
5YCqcQhyOKh5IDeWCj4cfaC7mGuMQW7OKv4Zymt2GxwNk75oUs0vYu/pmGsHh1gICuavLfTz3S9T
sJK4Yh3RlZry3wSWwPj3YEt17zZ7J6rgEvAN4OqEmbh5p/5Ftu2PzSC2guExwCxfk9TwSbrkphHd
Iiu6ngBdH+n7wERkxw8Q/oB+I9HcLlUKFdPqSJZtcwAhQxGLPAX0vKb4hurOPicWJ5pvjsK+I5XE
iqsUXxvt0xx/6KFe1kZDIjVu0DJ2gIe564vA4qVHZ/KSkibiLBmaWjAfy1fcMXUBeQREN3g4edOG
N7G3NCqtLKJU1EgJsPUKZze2kyTsE/saI4ms4Af9FoE0caKCTuvjyYBF+sAWmwDxKgBH6z7y09tk
qH+bEa/K6NYZgU6ADsIZ/nmLOA1v+kquebIhyEuLKwclnGwHYZOD3MbFFZ6G361+2qRQQRBXGPDA
0IrtOfiao9Vfc7jycAlkTLyv1O6PTK7TeR/+apDeroTOKmH2MrI0gxVKfyPnbVmdNjVfJOUnZW8n
gS684bIw0UHDLRmRO3CLZxXXN+L6mxLby+Vr44MQeluSm6v711+/MmaXTGalIMgyrlDJP9YR/lwg
fuoQFqwAPOf0Q4wfwdTUcwt3W/ucUHKFck2OwExIOUqOMTkotpHMs1Q0PfnZPh3ZymsUHP2LPUOh
wwIV+kwmRNyBn7e+uSeIWl/XD8DePfF9U22keY5Eq2sZG3eNiloKQS0e0VFk5eykPeu1mIPaI2I4
wXUxjDkv56mgE5I86wuDH5s6Q2R92E0N2B0O/xYYA22csLnq279oyUEFnSsNf/HizIPWE35OvQq0
cIU9es2/eaBKkU7unwqxloAKVpfHDIJ8O9tNVbmHTnDFKvOKtKqBu+WgbV/NQnJMqOk6dLR1GZyN
p/GwNiLGM++3TOw1G2E9u9WmoSCH+snuKPZCE9UyStgRY348uQwin7Wst6mONVdNWWAR3U/QjerI
2sDmRrnVpT875MTZLZ0eKDTlaqgImX5/hhpJz8LPQjYzIcx+IWSAoFE+wJC7uWYuYQ03W6E+oh6I
dpg5t54LKEAtYgZCCEJ0R073wAdwYZfdTDs5xMzBzZwSSAXsj1EjIvIfQeeZ4M+Bvx93kLqPS17R
rv/chlT5OTc+x9zU7F7vp7oo4RFhcmvuRPRsGCVC+5h9rCMmcZErlWpidMgjawXqMh1hyMSoK5uT
gCEGYfmFVlH13cnUVlFENjjPfw8v3+tAW1quaLpjsEUVfzbG1kGAMLV34YjEE8REXUyyOWCZr7Mi
jA57c1b9NJtD3QQ2woddUmQS/hS0bBB1DB3SitF0YfDC74EZzbKUL4umkBifGZcwTw3w6ebhGY9q
OhOdMxN6lvaka3rZTZRdTEhfpAgVFePCNYY4NtkuugLdru8waLHC3zOE9iVhxLpVpER/ePcHYvy7
k+EV8nJX+RYZileOPSCNQrO+Bus/7b3CTdaEdSp+Xql4BBLrZ63ZBfgJlcuML5jCLmEAb7SPUGfd
wR+IRFQwgligN4f1sMONT1uYemQhDQl+PYf5w0T6Zknt5F/zPzQNvxec2PEOhYkGnMJeLEmqbC/G
PAvmizlOKArY9U+0L2GnyEh+8W6n75JGx9jFJHlK6y0tqbpkJq+/w0m0IIWzmO160HwsqfWA+lfx
vURLPpgMzuP2szTwscFYvj2JeHSasVLZu1shHwPjurT4Y6yNKOmAYWR74rYooJGuwSOUXBg5pzXY
olUeVOxABzl4Jni2ODdg0I2QDKD3WgUzxbWETJwOI5AGyqd1TtDXQuz+ogMs4JJNqCZMVIqzCA02
SpusOE4Hbqu69bMC4gntL3+cidTdEcqqOmXZA4pvmziqi4Jsv/nuhIuPGbekfGCksgpoNWC5kE6S
RX7NLSDZ8RegC5W6ZxbfoV/4O+n1V9F0aLB2230Tj1l69WovHsMO6bZourrRjKDeuq8qIcVGySZU
eACwug9wdH626WgB1eOJF0Jw9XbR/XTScAuXBGnnz4Zlow6egVPQL282nSQ4Fg86IaaMXbIhs4Sw
bm48fRtFp4srxyQEP2PB69vCJGAw2JMbx/4/a2E/Mg5MIIdEmdxMkkE3dm0e2Jqn3m97b97WQ27r
TlV+WEPlS1STFqT4iQRSGtSHl+8GXM7U695lTEN1PScyxKmpdIw0MTrtUAmd+Qw3t7/HFEFNN19H
AB7Zh7QICMmaEq6yZ23KWrRW4aytoWQXY+qHorT6NfkKHmUI241gZ5SRerbn7CEQh+lulngLkjpl
zpL0dxCpJRXws3pdPPUzWz6Ocy+jWMqtsow1KD2rUarz9XHMNlWevAiHJgletC7ZQ3kRHuj2Hl+6
/jN7hJq9Q9CgqlMxranLtbLLJEGUfWq9XAb170FnfEaJyGwHjZXOt1rwkhRG+RjWoH46MHvDFgfK
7jA1nlbey06D2zK6QspVCtpL+xOeVQC3LyDW/DUi2gLVD2ZNztQeucar796IXPJckYuL1Wgvfo71
aswVOgavmwZH1C/HovPmNlc0Smwrrk/snGI1RIT1mOvo8XODtferiNwPctlh95O2CPXG7V+88qyt
GKNyXs2NDpzx2ooDjPqBjdrcga95afa7U0fiwpYIXvFTlSlmbD+0YmPifrVfZ4KQHRqgl9uFkRkp
1icx/e2xTLANJqOTcoqWMTQ+NDhSUrcnUdy5tKHc8C1tdkCKeNY4DCQf5lHyESxLZ4Rx6cGtFcZA
H0YIXFLIfPjP843o0pHSka+K4GH4oJh4FsIHAGA5d+gPz22/VCLpqEXdvHHMWahfElpYCzLKlU2i
9bKM1bs10J1zsvRkKSv7bNkQLOgaXDf436FbWpvdOQ236FeNrbaDaoG1IUz9j14jH3DPTPI6xEHy
6yea8hYJ93Ql9jR20A4iwlD4OTJjMx/qMbV/LFzBKZPwlxf7qLyjRpH2O7CmDnb8QTqZ/5so3PHS
N093Pj3OxRHbBp+AY3GbfXcqIWj4N80rlyPcyXzaToLVH/9OiKhQ92aEgfpiBaS0+8i44xG0qVhH
5T3In2mGjpOdrvuM622tLfetAVceCn0K1MWXxupfLaTmQoGeTbBIbgsnnOiV9bZYKZbhUmJkY5hk
Y8C0eTPv7mCCQ0rwyRA22PcwqpSo7a25S5MU0VnP2tLhdcMlUVTqSNVoUsxVr6Q396UGDJFGFmYn
ey17HfLBO1nCmCIfMzCFxW98MCtNYTDaflSx7UNl6gBzo2IiKsT2XZfJIizT1F9VJlsplYKA9t75
eX/a86ji+Q9CizwvfF3Rz+plsfS82BSDq49x8MSAvqtMpRd12ngn+PQ5jy+astabMWTgYugpGxAj
HMNNUikRueBny4TrceRWQoeWDqHWWv1If9p09yX3sjtQvsGMnTc+X1jlGm1MOFsDXm8gAKmvMJLq
jzXRdyDMYQwINPunZh2K9Xdhzc0ScUJrZdKS2z1hmBMweT4Dis7m0MtSlpFwpiI05yC92uVkdVqU
U/YeWexranhROfGoC+wC9STTVYIMMIbcMiUemCa0RzzWrjbQe8YYAdDc1vrBaedRgerz4yOMFzep
7a3lf1zV9SqLofGfVppcJYfpaUT3GtVG07C/zXt0eGiPattyaJdQ3ot6YftniqaMKALXdURey8v1
uV4BgIxpqBYh1J7DSD7CopWHnvPZHFkZ6HAU1jOOfiaRD2EeljH2F8/MKk+tHNjsmAdgcvLcfzRs
MD4xBedeIML3OAIJQL0hURyXZCcd8Wpqg214yKncW62sZY7BySmktp4iLqxoWVLnevgfyuft/USv
P2AzrBpfvmpf3FA30HJZXMCxZTD81YkbYqHIsjS9/l45A18r+HT5Lo/dULCozN8JdcxUINLkn0rt
IasQKPB+K9B6dAJhkSTXml4pxmJO+MOw+g4dJVUnqm8kJTDO2fOPHQU2IS7ET9b3BcIuxOf5FR3N
8opDGnUB14v2YqXuYTv0FnVGkE6q6luYaXjpSbN1jrVtycIqTc5kaQSeMA1OwA5biWB+Z9oCl27/
kS26xrnwHaWmxP9dMs8fySjfc9JfeRtBsyqljaUBfNVwd64nghWdeq3jELHBVa6tO+2zkP/3MBAM
yUoUCNdIlHN3ouFn4yTB68+twWFWYeq08sYb6Cfk9fDfntm1rsb0ExcUpTB5IemNNldzhW0s9QMs
6UG+t+exfMUo/E7s8jr284pBAwSEc320EcSMsmtrgOY3pAghC7bh+qedoFOAJGXwe7ys8D/+AeZ8
ndt5Eni6lkajJ9DAcyri/JVpAHmA2rqC14jbjTEztrzLPz7tDFdQa8tsWXeTwLDMrjh4UfotpqLm
z3RqBMcPmyzO16kyc+TDAScxwQrCzO8P4/dEgFalQcaPJw0Z1y+E+J7/4Ph2r/08DY9uRuFFMPTC
4EwX8zr09s+rxJtBbVO7EyF66dorm9vCQ8YLFkYyKLTuOM3HkYd0GpKpaH3zvtjRm4EWIIs9jNhw
pXt37vbWO/R18g8S3D5K8GFLWynxLNK0S3j2CTK3TrP6PxGnfN2ctkeC7rXU4wEcw7DWqZfcAGO7
2Hrw+AraBSfs9WlUu3JdaTiaei3ym+dzeN6BWul5FcWD6aEnB5LHij80BCennTVFD9IlvrTQ+dUg
+IE5j3Q87kaucfFVH/BRONLpq5Vx6AKWQKfVxK55J2Xp6nVUBckY6J8BA8qQtBwx7Mr+YnoeQrEO
3/zwuuXBEf18wQgZIBcYPlyX1XRFWAJNFl0HpTwWAMMvkyv7UVR2z6JLWcyFfgPazA5BhJ+kCz8x
2LUNnTOZ6nasQd9XT6UvFOa4C9lzmGt802V/2gvZhSDLdbH3nPA1Nt3W2cE0pmabSmLRnx3tIMEx
6zjDiuV4s9F52FY0IusYzKuwfSoLI6+ooF1At7qEqMlZx+jkcLP0PE3hLevPPxBZEjlZW+Ce9NvS
tuA69NOVPuKhgt68zxyNl7woNmLeTbwoYhYBpWTnPRlV3iHAi2Z/esPvFqYF0LNw6Vu2xCOH+gRN
yfssKfAvxOGVMKod6Lq7vRnOxpW0gFXb0pPuFl/QSGVf4wlcokaw1vGXZnNyCxpYtIXpyNADlu6l
l62N+9dt8zE0u7+yOUR6fUegMGkajQlXLy/Q6lE4z4oEkAstPOUuTodo80MsZW9OXSuEyoEYR7Sr
eOFHxbu2dGZUA/NRf+VIi75deNhXGkJcXA9VcW37BMfeV6rWqIOHYtT0NN9aJ986YqFrNlF23yK5
rgWSUjymKwCLKjyTr1nKM7GxCfM7QcTupt7UTA07D50MTmTp7GW18z/PAyMEY50Rybuv8ZzPZwOI
kiJkB+AJk6Uq5Q66lE9TyoZ9ND7zB2m8/CG+nTDDeVdpzTY7H2L6wVGBNqGNUhLh2tBO+d5hKzec
oFbnAePsqmBbBEYRvkpdo5TfL0xn1gseTDSNCv66Ddq8iZwp/OyFO3LRkWlWLYIBC9ZK+26bVTQb
JIaRbkgsF3k8IDJ5IP5tzEcsNSebfNWA0yqWSq9OM4Uwa1MIr0s9fqfXTxxQdT24Cjd11U8OLPvw
bh661RwRk8iDYGSwS71rT6nQ9LfFCgoReI70zAEnTAe4yRd016BJPiW4qs5YOiUp16OYGFRurWEC
uXZ34jIDiUPSo3EQ84t+NAjtWeRdSKr2sRRyCFlAFPi4+ndOTlq2RvWaUZyiypob0BNn1MVXO35H
OGXVyX1Hwh+tSrDM8rYRD4RGdlYn3V3oIld0dwmGY6djxwhQH6U0+YoyB64u5rxmT5dyj4Cxtv+c
ejQ7vnocI2e4+/yvH5+QDeVA3/IYduAA2DTobyjJYJMagNvAbP+18zwDlv64g9FObXQJdxTmkvGl
PrhRUvLVrlwXGm/Nm3T8JvgLrl/D51BNzUOl2ONkQdlAjEj1PaWdhjbzAjaAFNQ4aL6uGXdjfFbx
u4k10Tq8lTsQmwTFlH6qgI6XAR0+kq3+4Ytfkv80OTxR3D+TOaLlpe7sdzyW0Ty0Ye3qzyeCKyu6
SdxT+46lMNK0sPqFtq6jrSPwT1npf/smLN155hjcZ3Zj+s14ZvTpTOA5qe0KO88aia/V2pcTfXGb
dVZlUfF0urVPuUJElXBMx6lzqgyJvpZ7rEJaXLvGNrIo1XC8+JOzxLkqSuJs4jYYxBFnz8kNbz8a
41LHX5Y3lqAX42L/0dHS0Xr0+yAW4SUPdeCPrOlCNAROUdVQW8zDH1QtpRwcjR8YYv6U5k7oJFfP
oZmNKupoTcEiY2g3PP820zuZb3c3oyUs0dsV0JXmEDh6nUeVbPLgya7iTz2J2HtHKeUq0XAG2mOk
uPqZM4mUdWfoDC7vwsr6htc0npKnBQlezDqBWKa6yHAcouP1IXntVQNlXlTUwkidTmDUN0F8RPOH
huttLNpzO+h3fF7qMs9e95rEq9NtDsLNhnm6WRbRE7QNp1au7r5P1hHzESYVGDGzkCXiw27fEnFA
UDKmBk9IJiyZM6hAKQy5eD4pTTBG3C8JmAoCHHfpKINHQzvw0VOlL4NLKw56rn79TS/uuNnouwGk
44K1TDXdjHFqbf3vkpLJQqkiPL8Ihh1HXmIoygXrjpGoLBUX5oGAgfdtldRiCuAg+d47tnd2IVW2
WSscXXFKR8t0Bscs+pirgjXiTQLVBDm950du3AeQjK+ZxkhvLv4BTX65qyOJSxn7Xpxbptst+PHh
zSNCLFTw6am2MhppIHhV2GHXaHEhFz6k33IDnaZ9+us8b0bTF9pD+SjzgWeL1CIrrVSd8fthlFsT
UJqWB7sFdjEBnyYU4yK1RgbP4jj6GIJw+JFokO1oEBsfi1vwnGtLdiS0GXqyBiQuFdxin2HLlbcZ
Dp6boTenLe01eLwBk143nmcx1b6kNRq0+pZckUsLbRdmC6ImZ13W5nynCviDVQK32oe177dSSmPC
ykQcpb8PYWevrLxJiEryRu7IgkX3ZCh61dQ4DDuGlv9CifbgBV+WE7GHnfZpxDIn92PB82CLglcS
gxoIrvivrerGk4b2Q8mneKRHD0f9SzOKJ3tFB2RtedC20aryoXwggnYEP1DyQ5PgAZkMhFQoqNr4
7ZhY7LCm8iNRbDFxED0S7Vc6K2oAX9puOYX4dXFtY/Bky9fMXuBp/OVqpNBzlQaKp/mc2b0UsNXP
SRf6X8baoVU/mSvF51/fa/ImMvh3OWANpPwl763wycF+tGJRaceMR0mr/9UyJQng9I2JrA/CdMYY
EGUiYqTKYq53OROlskGKCtFrMYRtb4/CEJ8MxWXVpPYMPB/Y01lqxccAZw73ATHTPdYnfgF1Y92X
St3z+buxVgEDlQF/bMNvOaJvioak30q8QKvkWwKM5TnrKa+9cIY9wHz6zyG/bk/HDmUrcmw9y7BM
XNUCLGptWt+riWbcequcHaoW4cw/sDBs5bHatrRHjjUDVMdY0aOjCHor7BapLsBkb9Lks19hPHWd
1FuHADiSF44FNSX75+Ty84vMVFhiv3Hc9BnQyKFNq0cfR99Gwbf0kAPXG51Hijbf2B6fZvZpnx6K
s1va/c10sc4w1ObaBnAyD689avenFvhs2mBNIwGaIOVPh8on5gp+DB/NQXv2EYXLVcz+hbV81E91
j9n53DkoQAzqAvzUkmmeBbDkLYtKcSrReZv/LEN9VSN6h7+93EoilupM/jTU5apIWVD+AZLepmk8
1Y0u3M2HKzMdP8fCZ4lLcbmQW57pbH8rLsScp7hLBk2K8RCzafnj8VBFaPYpTSinbZNMLiHAvXez
9dT5Wlrgy/q3xRjd8dVkK6hGGeYmxDGXkdsaqF9zTJDNzuisBIa31izMeIA9d62gR6FYrI9X7yTv
xbXQNidtTcoz2mj2X8sL7LZr6w9TlmkGwuKHG0LbDNf2s0fHpArMoI9OGN0mpNxFUS8+fURcvk0S
iD7xYrBc9bESek8nXK9RQzrBNE3w6e8/7Bi7BY4LMx4DwBJEsmOlgp4lPhK2IYlrmvOZUisyxfBH
cgizRPE8/JCkytjXgy0l+NzUAy/CbiO0PmRK8JIWodBXie1898eBs1jdR/+DqhQSW3ho8d0mWfyK
SiFrXr6eOx/to5TtXhA0eSmkruEsm8AW6aJuyUcJB2bDO8y3trteZLQEWb3wVKL6sS2D+lYXZleW
dEyvJdQc6+qIjlNPLg8U13ccdZ++u+fiNcRJDFD8nIqqHelYL7pwfkYvz4ACIqyUUDvR6iZv7AKW
Kr+nMNBBKMM43tKdYifdAFRmn7WHkNM5V9Dvt++UmGnWChAnEHT9RJWC5cfIlTlo94lw2GOMEtob
ttjzuwdu7riqfzzh3XBhPC+RMCHnGN5In4BdOoH6gWO910CuA7sjQJi2Ohy6v80AK+Cu5WlYPNwJ
EUP3bSpyyeWVSRfQFIpHY6upwHZ4NL/Dmcl3Opf0xXcrsMTaDquHTwb1Fs2leXFskkc31JKGoe8t
pPjQDbo8cl091BBm0uQYfyzrCGaJLMtZ9p7lbabwVUB3Y2HY1KjBQUbed5LQxtQC8YSy6vmMRdPQ
wlfvpbTGBFF2P8iObniso5kVLLeahnNGXklmZCvNXCcv5bUf9P+VmRBj7VduWeWRr+vyBGiQIBX0
aVlLBTXkc4zk7WKC3264E7tT9T2WDXPUUxBxBcI3rO8W8ym/7iJp0O38/iRoNNnJgN4l5sFWk3Eg
zrkCH/6Pxjv2GU5TWUbxlPhCx2iX5MxbDActGPerZKCjzrT48F5pQwfS4GAVQtYpYR85DM/O55L6
IYF9XlNvv8MBqDNV67hnAEvssofeC+e8uzU9e1U83aiu+ob+MdwEZlN2Xzi3JdFzq/X7vm8N+Y8k
ngWolbWrwN1m5Yp8lq4LWx8y1EfC0tXwM/IJOIHIVtvYwYxMYCAsnO79eUvgEdhGNaFUFimHWGLe
LfMn4IwJWzX7j44p384Mr6Ito2mIT6Dx/73/sOky45TmSI/xj7SEN9cjzcbkOJVPqFCwUGgUnGy9
qeyQf3vIcHcZIujR5WRRKmaiyxQ1qsT2r3rfFFRvRwzoJsAuqIJR7SOaLOBtC01IvRKR6Nw2SYRu
GRHTf6ohI9JJ+lsP4laIJNZc5fpX1lpkv26WsqScqP53AksTHyEdHSTM0o6DablsFO06tbBKArB+
c9L5YphnHMwwSNHectKddOli+gAf0Ybx8Pw83Coo9Y7jrh1R3WuxnKJv+JU3Q7hoSitmV61we6no
wyrv6G95fYfh+kEJgjX09fY1Q74cesnIyGTbpU5oOF3A1vWSyoQoKYS9RWeaM+3SsYZqhG5IJbb7
/eoYs6wGGR1npe9oQU7qxU2CnX+dOPsdXhmk304Zxw3i4L7PLXv6/HYRbjfTn6poA0QlhhzNnXob
jA04av63Ou8gkzKBSU3egoFEakm6e9jET4wwNA8ljO+M50xOtBtpQQDExXwfypdHdqv0VS7hAOiP
YOIJ7qyvFoztOIWDknZp4SIYBxm1k/c+XuG9jlwvs6LRubVxk5jx5Nb7A8TnoNsWFVlyHZn0BD3B
HDapFLYDL0fkWAaeFdbnMm0fy7fG+xF8nn2FeXSKaEhFKL7zH6/KhxkU4M3X5dbeXFFTZDji/7ab
T0TFQYxkO5oZPjoh1CN9r7yb3UycAXxfH2Jewq3zYkQYlrNhWyB33t0TW3ZdaVu57wpjeeR9V+2W
Bbm83iX55jauWYvEZH9jw5vWqX6prUyEfFhEvMXMzLsi9He7Bi8laB4WKmW2/M2UsBxwUs9r8dK4
cn5i+rFyhJpHavIW2+qqVNOkbVQ1g/SPWNTLiwb4febTVyeeNzB5dc3t1OaTkVPYW96GfITTbylZ
6kPN4Ysb1kSOGxOgJcavhCc0QRKTKdDc1dmUB8BytkCXS8f8SvIZDOJLP7ZpJXTxcQH9SgvisLWD
40aRaAuWjGl4R64ORcKIiqnR9mDZGeOArXMwhduzH95lSo6N773ptknQS1VZbvioPxi52Lyj6+Rd
UoroMRzQHF0r3mTb7NY+GG2by145m2jXo70GSAp+NFl6rEzsPDzzaqAqBhcRozaeTaep3163MHh2
0ZsQ4V4sI4nO+QKaDH/qW9xlGrepJ2xkrr5FIly2ikU7cJCVp8llB/pnFls4IDFYcLX3UlTsb5vH
6CMDEQuVolnMr6TO51TnQegY+yAg1yK/RWt3BqyfLzxeJ7vxbv/1WdMf8N5Y+Hm5Urhg8dBoXuCB
+c23hLTBW9VE8xU8EisyHEMuXwyMeuM4ASRiKROfjkJWYu/A5laRKIbFOEBvKW9B7i94GJweCe9Z
ud2n1iUomTWwPP9vqmyOsaP/EkF98W9vFv5M9PkCDK3rWX+5ZXolgGMfaia+orarvWUj9+1fvnvB
Qkpd3qtYr/puEu35FHILmKznEur5fmL6bMfFldBxe/SAA7rRxyRo86CTPDCADt3+exQ/7j1ZFH+U
cGENKDQsqQlJfdvK2bskqTw/SIpMAerLzDTdJn+GcrTsQXAInVPXjFH/xyKHMIUGHLbv8ZmItyHu
ydhMBmz6TMhhVI7/eEkMPKzPRIUzc4IxdqN+K1dSw6ErLZ9FzFNc0d18wD7Hl3Wd3ka3kBbtK88w
fzj+F6qh/Imi3J0tP6DUh4OTT/FeMJHw7dsy5CzrVj4eyCOwd6v/PUPRqhixdSAVU1wFTme4P4AD
JK9i3uUUi73PcgTJPk0aQuKQMNxaGTiN9l6Y9F10f48rlXUVfZL+0TziTKcB6G/Y9hNjEk/iZ5dv
cfidEzAGFOAGU5QNZYs8t2spWQkNzBRPICHkXE+trmXU65btMvdtP56D473vQohpPrV4tkRuRM7+
12VVmKmxrjJ6kT/9LV1ZKm+/57zxEpQw9gNJnLo3sfKBsK3InZHLIRnlnaafwKLhAjLPdtIkIKN/
5LFIfO3DM28VOyyWrLLbnpQPvV3wrkA1CJ7TndI8zu5WK5bwA/VtWhGfCGJ8lcuy3sFn8HmSrGmb
boAHn/6+M5uSs1Tti99w8BEXPUh4F3C3zbqZgnsBW1BUjJvjs+l2KSY0aWEnS4ygpLedUFBgMkGp
hyFbK+RN09dkDRvG0oFfHY6EeJegY+rkOU4O+fBPbP3OEUIRAgusLs6otD2AD9iAkAXCgLfEVN/T
30/1elaet25tmAiUeaFWZLKWqPDslo1eWd8eOBWiWowPh1SzcsHzk2R1PkjIjqpgW5MrsF/z/QTE
rlsKAlY2GZNelW/D2QI7afTlMvAmWej8fFUspT0JTWHAmrzqMXidtK69RRVC7NCV18vLD6JSWymT
tu0M9/FgSt5nQNTfXDlhPvjj32+rURO1nhpw4GrWs5czbzmMX3JJ2t0pOLa1+vfJoLQhj3f0JzPw
IYWqNiMsVkm0FKAK+eg/p8NrYppSVKLhopkkGXS7wRmB5DyQt2L8zBzt/SraG1DHT3+shY2vMU2Z
/qeJVJMHpxkaMzpIsoBPj/TvqdWPHc7cJgBpuYsgdTWOM7Q3pYmPdXUwY0o5M4H91ix9LLkDgusa
0kh0QYnO5638PGlvHz3jLHewYbv+e5UB6X9Gt4YDNVBiAGcnErBbqmR+XVPyCzXFKMWqi4eT5Uvq
jiH5iUAlfFYRVSQQwN14Q4FFPGTJ4E8eX0Nps5YlZqhW+1peoTzIaYWw45d/2CIkiT73zEOVZgaz
GKYT7zkzoggmnx/VS/R91KOsLZnLhn81+icUJdj6Kl3JyHvt21CKYkjQMKw3XP1OtqqlSa6JN80q
sO20tMbNrPESEKjV5DNMnW6myJ8KPyr6uoANYfqVrDMq1q22KaW1BhPGoj4P7jFdUwGufZiSf7sq
cGxwUz930CNWQaMFvAV8xYFKNfjHUdnzpniuNHfnBU7ZcYN1C7SM6chXtVqBN4wQXCxFyZPbWVKI
/0BehcaWYfEY3Rxrtp6laP8zX0vHwUKjipUyZ/9+CV87WIGcZk5CQ8zA4zVteXnQ87p8dTx5vST5
7NMJ7LZ3iwU4+Lmns214zHv1rgczMC7ffNeY7oCbAFHLtqNuw4HAttVO2tOR8aKase20HRS5nJsq
LTSNuYuGpj/Hs2Cy0ZYXAqis3mptVJSoI/jtkz99Lss4DexJQgS2TDwoOrPlACQQrqHA7mfMwErk
ow6NLrBgoZC0K4D9d/tmABPmz0XLVdYo3R41RfL6h8C7iEPuO5Ic7Nk0dP6MArbveLhjlvLloKfn
xwnj/cADzHq0EQxKu2Pgawnfm87Ix9Q1pMJvBNkC2gfNIVwAJ4Oov9V/yEX1E8fjt3K6szB0x24T
NQsDQ8QmjOE50etVFofp4YBqH+4cWmcUP/q2ycO/OXGmoGE3Swu1DtHWZ+kU/vsH5HmA9juQPS86
U382scw5OIyCL2sKD+5uSIMFzly5Uz09p6UL3ujaTpiqr2rs0iWkJG+Piwt5tx2IwGyObojtUPzF
7ZfmXxPq3zGFRTWnaVKCO5/LUW5Vny+Mk4DprKM0N9kqiHnWNkG6P0vGwOhRjpuu/L46P+1NCLlH
lSvS8tu1SucSWRqVaWt5EZeUXlWr6Fh+tPMX/DnNfUuGqE14TGB/rVUO4uZrTPO/D229vNcxXnCX
KB5Du3J9sWB5zxZB8q2hMthYDBduxCWy9JXwEPaL5Aol+PtFQnH9yFBwgP5d5fckfnnLxrclb5nR
OtyHkhqyPQ6GFwxW2i68X7bj1MyvwuhvKSfBu9KxfJW/FpWl3rFAP3ZCHePQrZlq6D6j9IlrxPTL
V0JkwvKFgxD7URi1SprNzlfk2UcbedKDVFB4KtlSSxCFfYEn+1s23zwWw1ap35/KbwMQ6galep5V
tWNRPv8Wc63p2krY9iZgcrauQH/39aAIyj9xKD+VMm50Uw4Otl5aqMb+TdsNnOZONcbTl0XBeTJx
c/T+KXNU3zI7ZvdtaJK1y6S/7RZRsOgwbTE6Yzo5zC6PqzOTWjC+zZLKfZyjFNTsUXUkOwgvTiCW
SQ0xdXrAwjrcTr9TlJRnnWziegeteLeenAc7b/GaQQqORLE7zx0elEaF38av2A6W9dWbDdZfM2pb
BH2GvC3fpDYJqHusclHhWoIs9YfwQh3YHdQe66Hyzz5waCG/qeMGT8r3mmMG6Qw7cbBv5gqo5nrI
pQNXWN+B7NNvQKOiZC36xjc+ta2fk6fsbIz+i7dngJPUeSn8VbVzZDLLSsKUrTEKgbm350aZOJuM
OEX0/XxVfFCNdo+IcNSBOXhZy7BHQB/BOk3ImLTUt5Nw6lU7MRUzPbgHsmE25awKh9t1UYA8Yl+u
ZE5sCqiJBZbzGweS2ybmd/dleISwv82ivorvc1F6uLYyK6hD9jOY3KQXhrsR79DVw1LO+rYdgqvY
tvQsbe7rq6ySy/ncOeJytJ/HCohPjcr41/rxOH6OZf/DEsITh3oa71eYaqJPQttpxJgp0biHApqT
kki/pEg0CPaqXmjrzofguvrmakfNj8wLffsKqCsVPFNGlHQGKFlAW0IvjTam6FqnlKGMDj3d0eHk
1jw0T6eR0jaRtGLw2DZtJkpYvsErE1lb1BtVwK5lfxJZ+nJson3jQZDmqstNBQq/8zkLWhnjUtC0
f34J7XycGpKpNEBtbAZdyBFIKzkLFNbCUJmAMgLYEE6pChXhF3avJlCM3PLRyAl5QsHh4N23cygI
+Ufd4MNqJUUYXOAX59JQmbwocGxV1nStLMls/JAPjkUzdY6YBTEcg297f0iWX2+dD+bR9TCzxpGs
LARzkquw+r0gWEwbnkQuJo524qM13asHorTiDDn8+9sEEhs8hCsaOB/ujGfIPgg+LkP+fB83pLKL
TMJh2ApGLU5KYJ3frvJUYfBXFDcqpg8nN64wELIsGN1J4Tw4FEbpwaE+e45S+G+vZqaMKuZviqB9
MeColmhQYE/oVIV/i5zKi6oYK1DSgWvCiTitncZ1rWec28YDi/EOw67wxAC4cKCdINpKRrj5ohew
oFS/czJ5qKoAwrrTMSXveWOQQc/aLJaYLjP9CKtZCPb/taw2KAm/3ejEZ4zvmTui259oJp0ff8GV
sVOsjPNsaUe0wzzO7dFo1VsZLItekVnQHzHA4edkD4r4+5usakM9Wok3l4PnP6wRuk/yCZ8YS+dP
chTcgY2tKcmCVlfwC8ZzbsLXHBGP6jdBa91P5igunDbB/60rEeGK64OYStdh59yFId8HUTJ38+C9
inSKSbNlz84Ggrr9xFS5xLJWGeQB4RpBLuNB3mPKlYG9ooT2tJGXu1I4S3ERpWe9xWcWsC475O5/
V1f+cX/0a4tEGh3pt2mAwgmdvy52o00OcjWs9W7jZdTETL+mhSdQnWLi1sYZ5rkDhIKBN5uXgSiH
hKBiZ1WO28FHcYgqC22iNQpw3TDMf3rpUgUVdSAUQKYrX2lQh9/UoI6hWVK1TMIF72DfGzx8aB2z
QO6efNrhCBlyu//gUNn10FYREEGkp4PIxPmU02fT0OfU17n8al2GFcy9BCaLJuW4BmGOcYA0saDG
xIkTwM24fNpRcoZXdwVLyx29QjUsSbh1HcHl6ggLMaiF/6/AFnNgt0jjJPuFfB4ghAhF24hPGx4k
P74p9xbHDUwWwHiNwWPXLwEZu88W5nVXGUTXidjrh60wRxziODXJllbgEw255DebkIk9TCexgM7+
A3DCyS11UD2gjabXXDRbYYYBsCpJ0Y5riReDYIpb8woLPTVWGNYDHl0+6KwH8ABpw9cDzqGznvPW
qy6Ayjl+Bjtr5fTls0Db/8DtIhL3rFk88vuzoDf5V13XynEkIt4wYZM835v1103JgfCwxyVCQd12
ca6F/fJgLSh2DRP/7yUTDjo1kT3chvTDlOv9i+3/p9IHwSgyBKkKbVa4HAq1Rt6AT/mo1MT6bsqm
gboRlz15TigzTMEa4RdgkB2nKHnhr7BHRbQtX2SpPEtR6clC3saa9/zyUYkBoOhBiALlVnqg291h
FQL0KBMgMneY/JCjoplgh/l6asxs8FJRjUTnrPtm5p8Z67y4s/stSC+E4qnMpvbensqItbLCb+Hd
j5+Kjaoi37o7/Q8SHLfc51JZRN/uPBTfq9dtGblQmiiAho4/J1gkKqCQA8dC3Vlp1DgIwGdGIdTg
fs/AxUaiRNCU5dwu7+/W0drln9m9D0Zgxa+eXjdX8Z458nlZuy2I7Be4ZiL2etdSMnbJ5lHJEwwf
Ga7H14hVOHirVhmQKoe4aLOzaXBQgPZzjtPM4SIBJm0kjpcb/5rpEc29W2yZL1pLoBgs3koiy9iR
KrNYgAdXYGJvyk1Fpm2AL6F4iH5AuHbkP3noa6se3JkKFgDQTth81aIF8/XprHZpdIMlEBEa3Rha
4yfCD78IxpaJM+aKmXfkXwB/gnrf+faDa0oCrzqH/vvJtTCSfA6BqAlAMWJbazEqxMpUJQQwSk5l
BxMrNLo0YNcLGVmUBSslEhO7HmennOpofsvWkLnUJLp6qD1v75Ley0RGRe/RcpGGn6oRJ9mKhXOg
DVOpYQEPtq92oyE0iRSY4W2uLJuXhXiYUNfA+NMRgVfdQxO/a23vfkZlJQRGPQ7wJNukTGuOqR1+
Ur786xkTHDF3f+6Lqp44Rgr0x8yhYapAuyeJE7xhSYe6vJ2Ic4A4whUQW92pd2mppdTZMtF3GBPd
bXUAlp3zGwlAkVb5aV5XSKWciAs4EsMFE/g2ccnG5MRzxcgO2OBs9UhiSA+3uPegn43bbcOCAI5U
GyX93FQhHhUI7PLp8T6VDGb2dqmBeaAhCCQdYUoJEHBcMHN7MibS/rwEeOSDeidXf9oreFVIbxYE
XyjhvXsXhpr+1uX2ugEU69MRVwOeYxgxYBAE35lBQaO+LqtXQKaOthS9MlpvG5KUj3NdlFf8mpkM
098kCfSiXozrFoMwo6DS1R/5NECxV5gb4bWnk2gEzJOWwsrE/J/wFX84L44ewVqIUdC3ye2LA7I4
nZC8DdaE7BALnOaXJmARDl0p5oul2/CEqEgACsrpmnyTzaRLLMwKEHk3kOUZkW2n8QAR/0WNeXU9
+EMgf9I3Fld02DXZ7KemO6LsMUGAA+wjcJu67dQ93O/L+G0y/nhX5mFm3RJMibgZfdXGruKcduw0
oAFHyCEbZdfdqxN3lDjZfNgUtQ0yiPmfuOBEjf3xeY4Zwgin2Dfyq/Q4gYlsp8Hr7N7/sMYyu034
rZzm4mwSYTSLkBXPcqLtYt3abzLWUGA3Cwjq75lEmdeclf8VnL1htcUgFtU00uDGS3CMMAMpdVd7
HtdWi34jv4HgUE9DyF/0+e4NQmAMlNsbQlOdQJM2EPq0y68C5l1mN6i7rgWquRQb7VUFYQXGdx6U
ODqoqIt7CA2N7lISj43JuDu0BUle9imwTQvhkUWsF0HLKJT7YsmC5p3xSiy5n9EQ0y3T27888IKD
7e/nmArT+3n8jYgQWS77cECjuMQtWgHvKh9lxTaJr2FycQKl7bZ7ZYxFnZMOv7iwY+oot4HDRdwY
oe2Jm4wJj++/vLzF3k6xAKE3rQBmyqnI56Nx8GpZa5aKnWcAXKmKjKNcdKZJYzfA5RWpJVmY25b0
TnCo+foC0AYdCNkc/IiMAnnu/5Sv2YDZGiEHrcTdDO9YDBZjKqX5apuE77aulnVVwN3EEY8EVQfn
UpwfNhmXcT8B0ZxrG81P+SZFkbzNQ55JBTT5GaFc68vYFGEC6JzJFsi0vo6JzH9kJ0lkZ9x5COwZ
0eo4XGNaA0054TGuZf3jZT7enOy5zoFG878E19RJFBlJ0TMuPCNCraaPv8YGXYDk/+QbFfl7oauo
RQ6kkctwdY+Df0r+E7vPeIMWglG7AqiXh3fGPXtLu0UPEVoe9xoWHu3zJACC9G6Iv3TvmV4SGV+O
/Y4Rl5Pn4SMh7BCL/Ja8CD9zkm+ohmO7da9GksWXd+bnpOunYFhA8cltJXDa8lTb/PWpNm+JEgcL
oyvT1YA246Ti1iHmQm14EowbMxjp4KNs0e4qVoO0KZegoiBfQLvvVcGrkJRirlyHHE3tHp9JixAR
TNlua5O/lK6nt1vbnwquodeYDr6tU4qHjIS4JpAnvMaEPXXklM4x4TVMHbed6mp1MxRsSt2vHjXG
zRKTUEUty1cu/c+vLucbBCkXdh/58Nt+uC23toF/stHDr2V0VkBQ48HLSLag48+pbW06kbsTd9C8
bIFdKS1Pgez0FO/j78VVHN/3+T1T5gMZb+82Ob15P8bYfeFPR+qjQiKTcnc4qYR3NEy2LeUsZHwR
4IWIZ0Pdnz9EIAgt/mdmXNuocUaawzjnCgeRVWklAF3Leb2ki8+zkYQ7enmQFrYUkIocaewI43kD
ADc9AT+biNXsEMDk0N1UeCjj337gnnrbwJf3NOh9J04sa1GH1t8uqMgClqqbUhvsZH9K5pgySI8d
m5Xn6tvKjjqYCfUE93Clh3M67cfX4WWb0x6l90Y65F+ad5se8tpHSYbH1b5kylQ+PTK26tPOk++5
2YvRoylaA8A6qGG9O61yaUnP3rYQoD3TcXfgucWI0B8QZP7SZ57Mm9OTfNO9V59mjfFSDljuOO+r
gkd/Osl07wpuxanfwaSt8q2tHCKXSVf0lelPn/Q96G39JVFsBiLu4nOLnskepgSo6LXc7w1WzJrx
VZZwJ2wFc5nimNtUOaJO9bcceX3MiKcUHPW/535/xjAUaEbsF7sgJOqnQDH5TzxfzkXR+quII2wE
mA9esvZ+VboY8H7/yJnoVBtqSSX6FNjqkcmOADGougAnQ4hXub+ZoHFt9e0zmtsNYEIKCnLXvQ9q
C+WeVI5U7q+wKlMxgYb+GcHo0YrfbOxnE9Io675XvrKxbF+cZ7hGFHt4ZSCUcDFb57oByQyUivlo
EVLS0u2XNvGr9h/ck3vcCy6fs3Vj9hdxH+svzQAowqUAA3POqy/j5vu4OIJwgUG9cdi3K8D1QZmH
QhCnBLDzisn1eC0X4T2+9BbKz4sr9hLN4iJyOtfTYKWMDwHHHBThoLqYd3KHaS7ilyIxnfayIXKq
JDaEqmLNJdaOyDEZsvvtGiXUn6PYKdxgx8UvfAKmXrGlq3DI+1ZabfsC75sy97Zoii5MUL8uYFwu
BidRE98OhX19RTAB+cOq3jAm7t5RILeSjJzIq3GtJAlorGC6GBhDJXEffnbBn65KtoXVCXQv0LpK
1LDVoY8R0wvk29+PiAu3U8k0BSyYlW736jOGFELlRrSKYOyghyqVuan8pF58o4yHKrQ8l3FfAleF
p2Y8ASGb/REtMX8c5bqNhClBdFMc9l/CyF8stB60wbS3ZiL6EOgmlWJfouYgV5YxZ4c+wX+vqbMi
1UDrC5Gd5Ytke1rec7An55G+hcHduZuJyPZ43p6GWztIjNAqymVLMFIT2jmTVSmIyh7zNS7jmtdA
lT7hbAvbGKIu1N2AG2sUrCEteM2Ye3MQmgEllgIgC3qCcXwhnJC8ST7aveROqn1oSy3GP6Ne6hZZ
Z+QEJNVDN5IV2qQ6pmK1phYI/6DtQzpKGI32xq+IzGieWCRAYu0SixkbqO5+b9NPnrJHF+J/OnzH
h0fDzGYD+DcXPba8pPgqfu8ZSnO4LukxwHghoTJM5KtAJGVRL5TTJ5rUTqq8cbnMSiu2Wp0cbQJ2
u5KrYXaNPrh6jgAuP7RzW52KKHsATKYEa2nHf3g5qO3i6qqLVSj1zBmobN3Qx27YiUYEfy+ZfRSA
RRAHqaF5oblj2bhvL/z+FlhO5H5jWrPKkj1Myk/7zvTU1kXPHfoDnh0Y12OMtDeKPycDpLnrJne9
xNyJdJxlc8q4u1fGhxL6WkbMdHtrw0+p02rACl1vjjuhJgzk8uR2LTGPb40G0MMT6ET1MDYrNdYp
F+vTczNmD7+Egn8gBdxjarVKgcd9Pthi4+4xrS64l1vmTj9fQElC4cx6Kw7oH4BAQLKs0sCmQBAt
RsN/lGnGFHCxXT4YOHpHDCA5p9D0oCJJzdoL+PXah9TcufjkTjC7ywv7ZPYWoT5awrrR9CNpGAnr
cTiM9VwmflH8LHfIpXctPg4gyWU+TglOjC/Tlp2Cq5ofS7g4N80r3A5O4jENAEHGe2/Wz5M19m7T
RORPw9+f7Hcut1Cj55kyGl09au5z8jinu6oLje/6rFp5iqaw7ctPhhTFOvf4I1lZ615XRpM5lpnY
dZPcCJfMFrv33TdjGHOmklwx4aXIBJAEn/ZPdI2U2ZU19ZA6K4lyTqV5CCv9WCXu1lHcsAbCCKxD
AFpygPAYuXbMII5HZIJuxCT35nVfecynr6VfwDd8nV+JsAOUXZ1oBdUoM3Q1sxBOvLKyes1oIso5
9SUBUSEs8jqwbYnTl+LO62I5C8zUcmnaPvZeFW/oo14bPXuDiYcNk/kWHK7ZEEAArcixm+scwh1e
Iz1Zw9hllC8PWGNJ0vC6n8nQjuy+wm0PI22OJhtHAJ8F/u3/ZC9vFxrLrE42ygl+I9xygAdi4eo/
CEOKfuxeq0kbsRmrmA0rKgfOcfMNoHYMNSd/MzdeDlMCnhbjc1bBXefffp/r+tfiFti8B07lx0m7
RPy52gmz+fMUYyTmLrp3HI9hPdWzCsFDt3sqkCkPWNCbVKhHhIwcDIOW4IZ64uaTTACeJUw9988R
TMKE8MXusylP092ahvn39n7VnxZzExzsxL0B0A4uXYWGWV4qrVks/SrkT+Q3tpPIqsU4i/xI4Eos
s3nSHjXGT9IQCQPXy4PMPNET/J+aumDWjmCOXL72W4PLA3Ds3kbBmqccGWubdmCzGUHCQOdh4aV4
+/X2tgwl7Nm6ECIer4RDtpqkh0rCV9fd1vMgBOUWG5LAw4DC6Lk3mulv6UJm/Vm/HBJTocvkoLA5
zRSB3Ef2KA2hvCwLsU44vcwi64tUsY/+3qVPA+/gKRDou/uN9O799Vg60BXSq7Y8AGlmByT1ycJo
yVK/MSihQF7dQ3pFfKzMfYBFzK6W0wKWrya9KN6RDM9JoU3S8fSuuVxIGcIL2KJmZSb/wwvZwWv6
cyLNytc0YursvUfioNha1dvg3kN90Y/FXBVq3LE1BDMovAOVB4Kc34YdS4bL77niZwbqkSbxX3Vz
5VtdBdavhETtVtDqMAa2RfHSOEFRMmJT47uFlc6397/NH4amZPPpBKQcke+xlXyDvzFjeGo0c/sC
XmO2JsQhhMu6na4jQMlpGaSVWcnhkWI5+TnrttYyQ6CoGmDqxVOIYFdc/eBGROHav889uWgI8S4S
Co6oKAIBZm0+G1/JKCxEhUoM/+XQGu6CGBPixHPwOnTZuVaFPrMQ3K/boaaw3UDFDQ0R+I/r6jmh
rVUf9XsQSJeC9GXuYeivATvKU9TNYvkz1RQ2kg7QeAk4i4KsjMRWn05iZ/mo2M4E5LGteFnh60XX
g/1jaSXJGd1xDIrcMMyEsasjWpIwTdmfHbrYy8U+OlUXS3cVLSwKMnIUn0JiGA6pX66bmYU6idEC
TmBe0P9yvXD7tOGvz4qdA3qLjEodioZDAQL/BERz+eJZHqnG9n8DeUa51LK33fcfN3gi86HQAtV+
9OdPnndsDSftVtoDMoOnjNYkn+Tb4iQFlOVETuEL5wpnTVVWN6FDd5tV3wXjRwQdA7Lv6B1RlBlo
mUh02Rn1vKHkCD/JTEalwL3T6whQ/tpNqGOdq8J88TkCKacDMin5QEGCN4pgTPa2nuQ2g1n4i/Td
aeaQM8T6p5FmqiofqK7FRKpyRiRSQm/eprZnOcCq12hG7QRlNR5AfjBEW+wI5z6deJ0XYvVtWzjY
cBbUyeMvrNDzOmZFfcKu3vLcR5ICmhNRn67/x2IsoEIhgprtRr1Hbk5alfw7DOi1u0yqPp7EDMRL
3uFnCQ0rVXsQ3KnIA3e3m074Su7UGHKGGcyrAc/Gs+amDs5hLNtEK9KH8apVT3WBNn/P+B5zF8Lj
DgzB74VYZOnPs+cph19bc7dAZ89eCU5FfEYZl/bnE6jfHHtc36PjmjCFmLS92u/2AaSHowIvruqM
kBgg9EohrU7ct4F7zCJkMMF4sBLM7TBQpeGE0RQHXZlcXgz49dB019uqdGCJUuR5QY6a/6u6RNPS
QMIZdKBPIHaad/VZen+4BXrJ59ovJCGMTR775N+q9qL9gUJMetDgJ6gDGjLdzTIisNa1uQRKqvvx
5MSCqsnQCiE9CKzZZczesrrcV0GG0798FICawZH5kRNfFOvibbChXjyE4eMnjlt2hgLYEAtWUMKa
GiPhUxDbyy+yyVUPKHKJ40nktIoabTjz12Xq2P2rOP4jhGPTfSsRTaC5VKJKdJKdCnpc9S2SppE9
QDPk1LXh46/me3GsoXwBfQDJ8qGO7jvkd6otza/mMHW+/Yzo1cRFeSYzGK1miC8WhcE3oBwwDSth
elVo2ztkXXBOZEekl1uZ92+aM/cgsQMiX1s28TtusD32hVz9MObv/6siLQSxtkIac5CgYlxSSztx
ql/OFIY/oBKGUmPGmpJZqXXggKOep1+E/tRK4zbhyCYHoDpASDMTrjR30cRy1FnYDpQfB5ru1yWj
yVLKC6iKafqJ4myz9NQLCUVcqtqDYYNNFcvF9T26vEbXr4J2g0W22da/XL7WgvbPFQxeAsAbeiUV
mSryUYTzGllnAIdD3277drcCoHVIIE9gJJrMQhwDVSP6ov868ZTo97dm9nvUBqITXthV2eXjSsar
PdryVzUx36wdNCvDdOkvbLgifmAyqfndAqH/gSdC5WpCpu68SBGWTC5Dua3T/pFjuZClvUK4ybdZ
ylTkLSDszs2/7pG+qOAzX+CQATSzsxQaZtjyp3p7xRjkNqd1XqoNFDXxEAX2fefKXNUrNiBJYbb3
X6s7JY5SvJ8ztshDyq+S9xV0k0l3OfTTqd7CrznlcvgxlPR8wb0U44RiHQEHIx2gIXq4uBSPXtdJ
nA3JKWfnmeSXl4BEGVdP5ekLJ6GMUsysIL1CBd4vx7ksMfUTedFzDNvQL2X1lC+ua+eEtVwBu/m4
b8eCVY5E3RmscJtrDIjciD5VUZemm7fXu0SCuKoMxnepJxgGGrbyE3BpxPDCFyNuYL5NOuS4tXaa
XlWSW7sMbyYFfDZueITDdhb/lf++WPRBTdEDi9iSmx07pAqloEoJVs48Mm4obwBZP0FHdCd80MA9
qXfvNQhqdc1x9R9wG2VNKPnqBQOT7BukquO/U/DVWVHPmrd9NHHsjnPOM1MUEUvtv5k3LrG091dr
YvyDIw9CLjhuf/Q7sTefWW855z9T9/0ndn9eeDiLLMUINfLSzjhuKFfva9nBRaBOIqSZVxBn4MAC
OaglKoY4X1VXurpabgw0xHOoDVLNJbYFDifPdQhxiezV2rUQBED/MsopAkY4DE54+UWOI2oxMPRJ
q7sgrBO+OSlkRl2L88Zbf3yxqdGMbkf3xzAmVitZBXFe4nzjpVPA01Okv0N0XdnSyWLLWkIMxWs9
NBuHQqy4ooIEB71jtUKmdRcoz5SPcQ9klUM9xZI4oOIwxVEt4Y4R6gyz5IjPXd3GlIRGi7COhDQh
+DJjDQJZk/tW5nYtdwCtOWxK+7OM46B8NDnRbqckMhIkw1aubd+jEJuYIhzRibh0j3Hz6HrotTaV
cgqK7dvr0kJ9k3PU4aZgCkmyPTh+efGcucS4+xfEQ44sTtGyCeCvIB+aBik9j1I9vye4umx7IMOs
O7OPFliOodwUxv8z33e3eLgOf2gvP24wmdq9t7rt1pWP44iB8BCyWTL1vBnqrlnd+bDYNrAuoTV1
+iyEXqGVvX1OYhLweNmlBOCJu34v8MLH57UvbB63WcPAmPq0EWz7CQ3VZDWUQjd2Qb8DYDy0Mul3
ydjjfASCHoVnVG+5Eok/34HQzRRgMlzn7LndujhcG7Ayg6U5D+cHuOkxyIw5Hq9ZZGkhFkSD40wL
GuDx2BWhHcSMprHQrrZRKwEKYrEX7lQQsKpifwy3mmPEk4V2zAav0gYcPTaMzTNQ+dlvae4rn9dG
uK+bLQjZ78KfxiJ6gkn5fmlpGimOj5JxL2JQQxwbHy5WcVE/oLIso3ha98StgqS2p7uOn5zsXXbL
lr8KlyCqimOBSvGf2+eW7FboRh9aWwii548gZdadhvMc3VYIz33DPlnP6EkTWISso7HH8z5SqxIS
L5QuHohbyGkkHo/ei29sKRJJeeztXw5dhk7s9i2ySIc2vULiex9jIirZn41dGBTst6ICCFJl1l/Z
4B+Q/OQBuCx9AtUAGs050Xi79Hj7s3+22YzemfQU6Bk0WKkBX3XcIeNutUWUY+436Dw8ltb531oM
4EKGHghqxxvgSxG/S+Nc9W8dknu0ZvxzqY1qoW9B4Y5XX5NgMfWqZqU7T/HktByeOSFi4AHeQ8+4
FFIvL3ncsTn/VosA65m4cMGe0pVdceSStcAfygORA9uqimwbKh12X0DWpqiz1z4fHSt7WGaxPpwE
cBXoLJ7Zzp3uO2Tg9IQKgezOewPRgHLUDYuWuOUltk7lq4z0INhmGXkntjLrVGT6JgAF9Q27w2bb
y66oUpUBHG5gVcLh0Qx4L795f6a36kplv3vzKAAwTQil0ZX8b7z8/zUgXh+le7v1hTRtrpl5P2KO
XyFu7VYnLdZtkNNzfRqS4dIyXGoamYb4DYdPjX1pkXiNfW4ULNLjl5roF84863wCzQWLWiCtOTs+
uiRfhgFpEjr4hpc9s8H5dKo1W0qlf3BKCJfMAvgBcgDD4Oopgye5XjtEUUiMa1C1MztANhCGh0fL
eXUgaOX2vsS++dEsfwGfZRfWg1ozDFYnQs/9IqE2Th2atFluIK/rFY7V4mkpFV+aaLWXf8NY8F/E
1p+A7DZDak7NuB1IAT6rjyTFgg3OcK/3C/YeZiKAIKqx/ZW8LyIORwGg0lyOW9qRIGiu8kOCarms
Yj8gTq2ZlKFvOrKERUbLTcaUT6Zosvt1GHWU0aOXtCaB5wJ+6wk2ONxx1LGofIkfwuLd1l5BMoDF
ha9W2imYmz3NjjZxLJbFNSNAzrGK1LDiB7uN6bRDD+EK4jkM17bhgdnVCDYRRCPI5Wr2bBqJInfe
HTKe/hEy9FrB6hhUiqC1wvT6RJKvDHK17KfkmORS/M7g5BK6/ElU7Wk8GSRGwzCLnIC9HsA/6Z8r
A7FSCzyY6PUXMURNQZan6PvSCEj3STYXMTbtTz6gXYOAiQbGg8eIuyVpGKXgdj3abRh2BfHif9Pw
SYn5mCiVjXXo40p9SCS3QHQjFR6FKe9/j0bwdojrZ9MydhGXSPomXno6Hc3aLCnXpEwQr5nBPas+
2oiIds5lDCTtPaGBwuCG68RdyRDc0rtkTPuOq0mttx53FFtQ/THsi4CBm5fFserDWbX3rEuD61l7
Rg5xnZonJHNEB7magoM4EnrBEgSjUdZrR4ji2ay2AxaN6W3IOSTihoutmaQW6IMQxPeOFQr4FVnc
AFHdHrunydqT35UFODmDLtIv/LqmrE8bkkwD5AYWdwVqwjgVRRCP90l1Sk4oay3x6hUzy6k33FbL
yD7JEOojyFltYdfth8TUJSowOkPnTSI5t5HbEZk8yp/1SYPYuMI2jSviIuUmrsi28YsN+0K7IOMg
4gEN33swrjaLLax06nDRcC5o6FuR27dIAqbwV8UCDu1jkbfxgyupWqkQm48zTX7TVOasXFZqnY0b
lYG/jEp39a6d6fKnOEicPpaVTE7h3xq397GF9n09G2H5Ebi8sMIOc9xg1vOFT2/yYIvFMM5A3V3r
jIr6kloludubyqGA2DsJcSbu8VnDfT9X4MTNXYYqqn31m6IZZOIyJAi7hTtM9luKsXK7HfcL8Pew
v8c2tOHjkJAH8RjLgIHMAfwa3rND+4fIqZLWISSnG0t/djfNFawCzqRkJYGocjqwmZkRKmcTg4sB
IF0nlsWkbxlzxdDUhXp+WVjVfNwlyA68rWAS/fFRbHsJJnIuItKXfjZNllI47f02bi8TesjwvyI3
eatSCzNnaapcSUifsvwezTdmoSkcSNDQNpMZtROyfSazFOosp6VY3+Lqjkd+lDqzBZquMcJimyp3
rag4sqo4trn67sL+LrLi//R/Z2sgps7Z4KVgilIu3GRP/qDxod/3wtBAZ/5NmgpqGdNVJSs8JCo9
XDa0cj83c8X1hMy9mViRPJo9KuapIBGJ4Gq4qBfd0NUour9usJAwccf9AnlITe3U9gh00cETY1QZ
hjBI73lc01JvwSOUxCauTzOf7v3zpXkKC99u5/Qqx4cW7DSVM64QGFmh9Y/i3uaIPQDorwnyjYJK
MplP5FJSxSJ0+MRdVrUPHq22aBaqsC9ZekjcPJVYVoDX/CPhBUeAUijngWM1f0ujm2/rcLAJClna
n5o5exDJ6Zf5A8KgTgzFUJYE8JsnqAg7xD8Fme/YvNhEwPmiYw71cIjoxCHrta5bF+fyPjFJP2bL
XqHTNJm8IyEKOLqJxBUd5CiIMxGizmlzBRXiK+AkiZGXONAKDOB1/6qaz6MXUGa55IqxOqN6hna2
prhT6DtfpAkjA5Qu2ixqQyes5Qy+78uBxA1cT4qh8OANU3f8EV9EWU021Tu3Ym84iLOPDfp/pSz3
V3QqsjX/8AqzZWj51Erjj1GoN2eFaSpGhu86yqo7PM6oyDl++qgnMg1x24zKOggHl4bPTG96rWLw
fG4dOM2n6yXM7bFc9QE7aoPLK9ALxPjuw6NPAPxy8jt/c/tHN8D2Coeg2hXVSXrz81FPuLfhv+gd
XOPtdjYPO+I46KfIVS2ZPUK9nEN3i40gtRtE6/fP5bZch89HOlMJr5bl6G/ZGzn+ElH8k9I+NEdU
g1qP72hAV4CHMgqag1F7Y8vrPIbV22BjRW+iRX0J30+aZVqdLcYZ02A2xOsXdgly1cQbTB6eci4q
VwWroPHhXF6inVd1FUPmhpJWq6hl1hWA2UbDttax3c5McGMu0HdntX+iwcjZ+R9x6aN1luuvgGEb
0OovIbHxRzLlfMSG8B8vM0aEvGDC6hTIR3q+lRdZsUgX2VUMCPnj7ldkD4afO5n8XL7ySov5LnSh
0DHvj0UdGcuXdvXUTpD8D0eR7/etEA6liiYI1n1wPpchXHKXn1cM/wBT9hLW9gcstyAd8OAaTFmp
jr6cv+toBZ5y88Jbw9KTa03uaz3lxtENlcoBx9hdi3ak6QUZY99PT1z1NtHciEEZAonFDcR/d74R
Djw2eQ5erEbnhsaET54EJYfh53mXWjxb0EfYWP+2/T74iHceQcPQ1jnWt9YOTd42gZKm9CpoTHZK
iswq1fjwcGy7lq/ni3Ik2ahTze7D7YlD91nhRwjGKSVAZ2KtIaUxR3Og3NO0EPU8MwkPLZGPGOpU
XsoYR27Pfac2MC9uaOqWfd37Fv+qfiB57896SBccUqyPRw49j0pGIzr2DQD/USg7oDGdXAeKWhL3
iPdPhLL05yw8GkoObzv7IROo+z5uZCD9NXosI+Tlv3Wf5mIKQx/dJq5uxf3Ssq17vYTz/21vS11c
Msw3inaZjNMME6aRHpMqWHyXGdsaXEuU5d0lwKnNUnSFcDdMneJQ1/n7MHYBxkBZ4WNBRhUGUBCo
25imcyLAuRyjFkJ0BKSpCSQ1mofp22IBbAJkZML7EYEf1vUO4DV+0E1VvgcVrDkwlybvEIt/1avu
odpbRJY5SFhCuR7Msx3nw3bLWefGq1cMr9MuCv/RJfdND4PfISpGP0IOpvWqeDV466YkPNVKQUmi
C4IS0WLt07m25qBMgHcF2oOCzm3tm/OfW0nxoV4FceJHJGbQVV3aEp8zrExeaXTh92euGFdFCKtB
OfFPInylb50cV7YrTiOG44w9CsRAFJRJKq7SPtUDG8jLAQd3bW3j1bpOy/Ut1C4AgLeY8TF705Ek
ez4VBB3LJnzj1qmszbGDMKfy9IyrK4WmzhDju3IaGro30XKDhi5RdDkMPXwc1NcOWacgCBOc101N
Vdt0zc+l3n5d5pm9VG2ix/mlucsd/xgb2o3DAY+fjIZJytYtrBEZTGysW1CIwKUOeHbKYJfFnL/0
FzDk8KafIbseecfMqphF/UoUdT/mGtWFMQh+/Qzq27vMTK70MzjGRmKa94NWmFRPAG1BETMPLbLU
CE4AG6oC+iInHfrb8nCanWJ/LDCdHS09XBlA8rvOkLmUQPiYBDqxXLuX/zI5EWEyU/oCQZVWj7Lm
TDYXljojZ/6NR32v2fOIYdTrqrx9ErCft420x0jRfApfFMaIfeOH+ephhSirg39i0fbHTAv9nm9Y
dSDkM1RzA9NSnqW9HUNeoXmiSCtggq5Dp09cu0ynwGRQAhUNSd1hcHjtNowwNQEW2/CLOg7FXhYg
hIUHordXaFrGzfFiyJLuPh9zL41Yq9D3gpmZh5x/XCJeArtzLiBDPDUW4vI4jQpZBGCCXfD3MFgo
qz6YEOH0ZOlPlMNbASZlDIzwHDGDdyFzOX7uu3hZgOxp2c7qlMWPT/E+9uELg6b/eTBIl7mb5G5m
MaZqGgwftlu3oAU3uJUlPmNi/504EP0NXY3x0KWaP5nQ+KmmVYH1coc6aAAS19/zJyqqvONca9w1
axeA0mBE6hm9PXTGuVexMUQP0L96NtjQLU9liXxajeW8wRwpHkdZLYVN/S+nT0rA+AHeR7FNZG6o
6W5fRBX2pj9dWX0TJ6YWCBhxDXMrQGchN853xu51q1mSxJseZfdaJ6wOl3/H4AE8b2zUWk+O2rj/
VxWS6g+zUNWgtsWskFuv8f+ZpRoTZDx2c6zaQq21lx1X030GTtzwCiUgc9nmCRJsabNt2gx/HYaA
h4XGE1BpWXtieHcM5E0WmS/i5IycrRBPAAckLcAwu6gwHHOEpVVNlMkFBrKUH5pPgLR8eIcNqMLl
s7A8XygYBta6MrGZZzEY5MJ1hw84GwzqN0lzngoqXR8fCWZIuOJ2XFnxEft7hSkUBReUudrkdxLV
AKI2hpISLiCD87lkJW0VpK5qjqmjXpndX9Vy8QIUIccFK5vlhemdcNl5Bs+gwxYj0UB9UZ2YFWo7
bP9LLCAjgeFa3dH8ow+tGbvFbJxjtZDZwVIrj3we6kXHdkxNKFadXqLvgfc/8z7L3Tq9gzANNSy9
eNrZCHta+lnHZvCpdieEtCh+36VzDIYmwwfYXvuB0dy3zsC/IJT1wQDreSOHPyMLFsToMhOm4z/2
bmOrYt3SGiM9jb+Hc7VHXM/wNQZZfbXC2u3PM/5rnEx5sxkHnCugt7WnOaxnxUE61ybZD8osBtVy
vk3Je76qIRXD647Q37Z8+JuAeaAMorMXgpiegAtme3cJ3XMadleXyVETvLQv42+PDmiPznBHG5op
TmgkAUa94veIus4EGf/xQ7ho3PIWTRFlANW6pa07gl3EWQ6UvlUGta9QXJxTYFvbfeYYb1a3x4g1
6PVd+wrwtfqqycm7V71HTGDPtkUG5V3R7vvgy+TvKSxn5rishNJ9XQ2QGMoVeOzS00G43/rcsG8Z
i9uYNfjIOvRFWZRZ+f6fmKBCataZhXSuVIWJ2Sq88RYdb2fGZ/O/ahKaN5kKdSIHRugGyUl9V9LK
+SgHbOrMSEY+vZrvI8oQm6VG+fitFCMZxP5EzbcucLHaNNyVLCXSXVxtXO4AQdFdPrJe2Wt74Yf2
3Kaoix0y5t+ct21mFuNmRCYdJ6rYvw+z8QTZNlAXfxsakDYsLOSGdTBohZfooE6yRuyAvYnRiego
sa4V0e8eM3rjCBngbWRioPzUrC1UMEcnQpQY0iqXlAwKPIyz4lR4ZPnLbDmOYkd6zpy62jym2p5i
NArwoI1laChrwoWSiHp/8HKESRRCTdG4kVEkiiagJm6FIiAqLQqpBpmG+mVsOGaviEL+WCUEKGUn
PIuwzsaZa/o05fIMOdhilB7bnr5o+YwPRehdANQ2OkBioz3tHV5Hlkwk/SyLsLSeufM1yZfWM27B
1Swbpl5efwJMt6TX5R8EO6VdiKmZ66FsxFLVqwD9AqMRsJrLoJxfCnOd32X9ZzAx43SAFQ6ca42G
MJrt3zi+5D/4o+FrRRrwVp6owQo3CxW/O/lmAoXBiSgq4OjLYs/2ulrjOT+TANBAP6sGd6ENw3vT
9IXPx/C9TlxvGK5Toec1YtYfh6xMq/LDRrQR/Rv9W2i4W4p125NhYoovjw4SsKHkEmd3DL7JKM1N
N8N+AEqLAV46pC/n+VHXBVBW7npLA506HYS2//dosiIW1Wl2nq7JfuFTeXNZy98QmE/wm9cvu9Mm
/Ewo4fvxlZ/aN37Y5fPMnxiVdYMkGn5WS5lOa5d674Wh94NWT8RAyPMh8NLy34TZW4te2yeDQZ5O
anaU9zFmb9e4Ii9I97JLPjCGchJ38+pXwxiZrQHMwDM/kZ76xUd3lEniJoOQ+MoSlgroC7wrNtbP
43iLzejCst2WdAXgFFQPpIHjlVej5LtfB3uwaUqSFZYJ4eOcCDFL08h9TO4M4Und1N+03mLov929
faQM4YW5AEkblzxVSPpqP/kXVALh2jf+U6pN46uvkRlOX0lRw08E5WmrBruejea5h24M055hF1O5
1gKf8V3gf/V9zkxyqYQaiVytttn0OMPIgqujJ4cSZ7bN7ulzZbwUO0dJqJnF2C9ref6OpFV2iKCO
8knlwmzRjRyHUIGf3Zzv5Ar5f2KrN9zWsFXRLL+tuKB2csXpjJTAZWbOSrdKJIabjUf5DdZ5UI1j
HmPxMhjuU/d5SQ/4fGBzpKoQsmLFvXNa7KNv4myu+pklNonlLgibLUepp9vXPmEnnSw3gHzoX2iJ
3wtq327WINuKvbjqCuwUY41vBfqszSxRH3+RLR2zoUfjqg/wdWsKgUMrvfYZWijd+PPXDzM4PjMA
CuyUzvVwniochaPgq5PbtFbKjdhhlOGKK5yREnmI+8NstSy+K2KpOtJyfGDdzbBWpYNizkyAhdMd
6Kz6gekTZh8rM5Lhh56qaGA2OEdUZ0H+QdpZXkFwLSWv4d2ngqZHW08hhZ87T0W3jEK72NGkWSIQ
vza025YaTwf0Bbfby79rcuuq/FyVyrqe/mYsJqztZfpRsu7xRp+lgPH86AGy2L6y8h/s/oVAHe9O
Ph+Vmb6lqV4vYKmM6Djbg8z+d7T94uspOXNl3kw72X1TmN1pabz88Qqt7Gw46REZMFw1bqlco/MC
loKyi0csbBlq+P0nWLQunkKrSc/XGtwyNfHfigvJW3HqXz2xhioNxyRgRAeKC3MwtC1urcTFpBh4
IEVbICJ3Hi1WYHXTN+uGRv4Nsz7lOLujwMJ9IiapvWwGkohS2YCNOF4R6dmpA7PpHq0qG/wMg2bJ
TJ6nXGWVe3g8ta4/U6YdCIYmBy5zGT/6VC/xFD+tO5xvF39ZAFSzU9b4LMpHCFJs05u2Jsjz7RVb
HSZHf7iFo7SCOOegEP9SglVYmP9BD21dbO4VB2QdjGnUiaNk+4//NaiCrMVjC4ayI6XVbbDI82Ce
xbzGRTpc3qInS0P38TQQ+pQw2AqaNvK4dvT9FkbtQ2c4iSgjnVhab8kG0oI7F6DonWhXrZeiXQeB
hb78Z+onDgXcdc9WdeDgP1HfpmHG+FcVMN3VXa7FONW6xcYKs3WYPNUS1XZYCj4cYgs5pLxCNXzo
yI3k+FQe8opm1xvNl+/RxevU2t198c39nMTTsMeDExAgs5NTovA/IFH5ZacZ8IrHqUl0kM16C+VG
fI8c8jKgUGNAoqQ5bZQ6psiehgwK51GtBYgY8aLEtcVt9U7SCNiJMgFa3UjCN3TE7f0lW+n/D9Iy
si5juLNWjAnfxekSNbrKz1pfnBmn7aAGJiKlNmsK5dE3SignZW2Xy3Qq6IXtouEEu4DbGyv0LvPg
QbWhh41SZkYzNSIct1fRymWj7YXSYa2wDe2T4z6ty6ocdH+v8B+P6nFS7dbtPLX30ChDj31qo/S/
rOJa8oBS2YqIJ6XnleUtJV8ywooFbjvzyf3NATw5rC8qMlPC19IfQr1ZjHkjarX8lmN1ohlShd5o
5vDeLI9fOVx8sU8iChZAtvN0xLCfGBl3zYNxtcS+KhADGgcdO/kqmdLVkdGdMBD1/zMEZCE2Cwvq
xxpZis5sncxtLumyUMLexMJbnqZiFA2IgqRefsQs3K7xiJEvEO6hn6I7hdr284dJHAjZ1lfImvKB
QM69uVul0/fhC5SEBCO93QPzjEw8iOe9ItKcZmUD91PWdhsX//pjYUwwJ4MQykx3cy2mXszu3TO/
5hnYyst4/Vh1JfR+EU38H6dB7NQgHSDUgKCh7d6tAlFJXSoxju9GWvtmaKhsiqmRV3A2xLcS/BJg
rJMTJUmFrTSghwYY7J5wTt1BG/V/iPpD5pftpx4RUxJaSOJSIBOAI4F5MRKVKrcOxcwsYebJsopt
glfTIz5VKg5TORyhQyH2IWyqW1xVmMjPZyodQ5LBWPZbM+EsDIw8ajG/fEP5Q9IdgV/TCtUyoKaX
31gZJw326gyfEEcesrdAjZHdZ4eaGVN/1H1TM+jtEtfnjEFb2QkhM6PmjOBvzmwDJLVOQaa6KfVs
CSnQ78Rqhf4nhoM07nQUUYI6tKhFz/BKOK3zljA02NxImlJkRjXY6BXfrKYuzt8jnT3Vp8ZkGDoK
ERDtDjoIiTeC4rQk0TFPs1XMXbvF0J5pL89WnEb/rIsoSoEyOiJiQea8VHEUdquwH/javg3DGiKO
Da1KXKjQehTjiyy4RUlR/+zE46DFIXc1AjHYTsIEQZFnW0UyCYyFUqV5WHoym/Vi3LxzDhDLCNN8
/DUUt0j9aXr+aV4Qo3MkwM4hhjyAr6CeUXuKWK4H+QfldSF03025tyOQaIixyyyRyIsMnAwnzxa2
7F0q4twbC/IFin+DiptpNtXhoac0DD/8f6rhvqN+/xFMjwb6etXB1my5vnfUI+oxTKpq1KvqJLY9
LHhqAE3vnhmUAQ6jvn00Roo66NNK49RUKHHc0AELJbUlfBL43YsNlDCYAjxNhotMhBSr5i+3RmBC
cUYLWOz6WwWZlyJD2wW//a/XBrgRJzg0jS3qqmgq2FK3jzYzsGpXOvKJTUTQIqlQntv5BWJuXdzu
bu0qMxjY6sUvmMz266czACwX9Q3fm67lPTmWrhr4oxAr0uqYdV/m0so0cXFnCKesmf2z60Q2rfZH
gobXzT7S1VwSXbs2oqZu80dwDxF/3i8no7xZf4IeXRCFTH3omrKI/qjTI6GrxUuhOO9xuqGf7kR+
QnfY8ReyoO8Khjmq5t7xqv63cH5cVXxTWkV+MY8D2A3qC25brZ2ITgTzf2b7rd8MVVJRIbSDVo84
iqn3p+RJcN3L+y/SBhV00GA7JJHd7wcOpLXE+NTOleGdcKQHES6xzsoljShs9QJ+1dRUkv4zpYNb
VY8r6MhYVD0mtmFYs5O4PQTiz7ubrnSQF7tjdy3xmWCMWDm6NnNzPKmX+wvHtZTMy6/8LAvCsvPS
p4lwn7enDrck/pnwlCYbnhoqeVEHwvOoi+177azIEnevmKL/0vodT01N+JRUderWgHnntACK2ay0
odG7D0JedJQ0MmW7NTXvniwHPstrZWLU/6w6501bX2uPpTaVTtXkR3aWmoqMmrQssjV9laXMXGT9
zkXYV7D7mxocXRK7AnxLogS8Cru5KugR89twpYJTE0Joiq2XuPqI+oLbFSi8hxYbQz6mncTB3exG
78GHBfVv16CL//TmD+zKJukP+F2opxmtH8HNyzvrSOgKS6ofTESaMFwtLufEuz3+sVrSObS7Q3Lg
rBZGNA2vy37h1sHIcXChIQtTNn9b+xm7NtCthnG6CzdDos+IiAkl9SPuH4vnZfFHkuLu8tIz1mww
gFISRxVTjGMjQd9wc9or1/GxuhmIOcx8jcLUj/3such0hr7P0NFN8S84SRGxSvyTQtiy0gIqpa2A
nupE7SQkeiNpthAMxgQm+s+7CeOQ5r3i03jN0yf0ZBdvf2BUjUFYVatkVl1Wx1MLKLg2Xx2IoKUF
DvnFNwKP1Dj9OpPdMyzXnyFDHTpoDuUt9sZsUzrbA68q8TVZ78Fp9IlBNkw3Uve3HabSJ0jLFo57
3OcXpBOGCpRhIhdF5Q3YOnJeffvVZxGhYIA24u+A9IuSz0wEWO9ZgkMfNHEQRW7g0Q79JboID5uE
CG+Aoim9HhURM28RdzAnuirXEgIB81onsHiXhMjWL+8q+duRIzhsjz+t+y7/BQeZFzKpzMmNtaR2
m4G51s9+GvML+r/xnLX4Kf7eEjhGC9Reevcg6Q/AdOuthno4FvofyTTyCZrkgLVmg2UbG6+iN6ro
xFxSVctTI9V6zvSqBWND9H7WSO95v3Fy6OxfNxlypi4klWEYfd0cWPEMVFHuoM45Jw5L1gZzLEoV
hRtYj0P6f5QvCggxWqpY+y+ZSLbmTvEj2BGoVh4zMRk5YxbhvbXgeW8dcXL9uIhZ0+OIcRgFVv3s
uqv7YbQcJvaAoRxdO49awm7KhZKoYg7hnOLBFaBayJSQm2zqzx/3IzFMrXV2oTpk+83de5ZmegRZ
sosCQnCTyAU1v+fDSM9QI8K4l99SYjh7WlnhrgjLJHzbrfH7aHndvk3RJCoLO9X64i8FIi4W5frR
gkY9GCTGG+2i6qrgjzZJ33nyeLafufxqTHeOLNGoKWYL4TrK/AGblVAvuzChrXaU+7FzYfY0HYPS
JxHz5xbLHJqNUPbwapQ+/qVdPx33/9NC0paOdaAS/M3JLQSDLrOQ0ntbh91JIIWfryQx4hGDsi88
PoSpHDcSZPYsVCuq2FiEUb3tgVXYxgnHYk5Xi8RND2xFhURuG6CeLtZpeHMZw29jNBj0jA+8jxmy
I46R1jKywoeNQNGWLg7trvDqbBei20zaM+KCL7Jm6wXSGS5HGs+WOB491YnEayhHQtfmHmx5xvw6
pSbQ2RzSXBvB58YPC3QcXEzbPVeV90oHuOQvg0MFhD4JM9gcsF4NEKLMiKQnvHCznRjcqxrjYNgF
sO8E+lS5OSCY+nGbXUBLQ4WwXrwziBrt3i1AZkfraEyxTF4ukuhM+r60B50hsxKdlEvBr2cvJheQ
wFIFj4eUBq1iKHgzLOZPR6iYIYi/OHTiGxqRO4g40oUS2wsWRlwLzwG4l4bpI/qz4lyQ+ZW5aLC9
yyu9gAY/omMXBd0p+58XtgKKzLuE8fhuw7/dPKatO5uHcsFuG0ymg4zGvTdvt1Esspf1sqrAY21y
X5runZqVI9q+3rgYJf1nwxq7tfDhlHb91KaClvqqxjVylVvIUvs0M/4qwbEsFytOrUBC8EYx2buU
jcRTdFlXSrtqJBmNdHkIUqprizyLKzO02eJvQQ11W/J/1NU4KZW6Ji10pLqys4FsUP8efaiAGTJ4
Lk2BilBTc103wLSKllSm4CnBEk66mhoqqGRZMNx/sef3Knq2BTJGG306sDotmDYUBRgWoTXaQeFs
QOIqwK+QoYFWwVj8zMfQP6uJQapgIsyVO9WvufVgwU3X817prXkBipJ6usXBr7Vx5xGzOer0buf8
ALqC96lDEbOwnxuM75a4Z0OtOpOpwzcZDC+USNesu3w2VWuH+Eoz4vn6OKe43OQgVPvfOTs7lMy8
DtQ9tZ2JdR3ZW6SkrRJlJY7FmlkDm2zEprOCG3VDdB5PGcoH07EDti2LIr7b3ikzliA95BsGGF7Q
AjRHmbsKmODmDAy9h6h83DZD6ZAhT40zuRSIx/YC5kF+qBDhxR632sRs1KezhGKrVmBjP0Ofi+15
GFHY+aBWcEnTWDjM8jcrF3lJK2qZVhInBUbnf+kDh8CsGoMILTScekZ9CPf1VlnIwimYtjU8GTt2
reISig7DwwDRJRcT97HkZ5N1oklX2OL4rQVSvqUxqwzqGReSoYbF7ix+3c+IiHOt6MznzIfmYAWk
rd1peGOEppdNIH6BC6u9Hlyb3WSM9R3TZ0poDsW5dxIKf3en2E0vV5R9Uadq8b8lrCfBJaoIuGG1
CXbl4sGjPeSqTuQGIP6DzTBQ+YPchrWv60NDIg+RGhJKyrteYcO/StEdag5Z44vfKEBBpAszx/Vx
vY2vQa1cl2lS8BKXrxRwheBVjZ94AlWHVD2ywxOdsvMlcWXZQI5Xj+JmTO2KWpxMQ9NE18yc5xhE
UBW7AOqWP14VraHjHSjB7PkjnUBrA04a03L//cN5mfyDTW0NFEUurMAQST1QMK7ozrRme8ikf5u2
mR5/9l6noBBvP1IDtPpr0yZYsu9qR67TJ8rANYJR/De3Gc409+e79+mCFm3YXAwdfc5rwSwe/nkQ
x2ewjQwQPDnQclFTarEKHX8d0qRglXXBQm3otYaY1Q6eN7gk6rpeiYSAaSTD28XvTpdyscZnK9cS
HrA+pkSrSEd/rPmMg93OjC115HjDZVpGfmfGwoHHgx6TrtAitFPlyfU5llm3GeH6Q6J0dgwsaGAG
RuYEuaA0e6MA75Z+JGRS5sa3yp6CcqIWbywq++UCpYprxXbI7xz7bwpzt9EiQGA+fv3wNxq+OZNS
Fu61b+O+E7mDySvYQMTDYCMiDwECjxYI1aTsNp2bhi2gc/ObH+Dode4x+ENKOZWtXGTL4KTALPcl
35wpWuSeAScK3j0nquEfIR7ucFCqIP2oRXMibtaXrJ5hlhbgjh0iIlu/HHnOTMkNzOlEtgnTCz/L
fpGDTMqWLvIdQk25lQa0T50DbyAyKpSHKPqdoBVHXEQf1FsrUgbOehneIaimNGzIaH4+Iv/Liwua
+igjaONwuRNxMeNlJq9d+IAayOdmEx9FrAs7sr9ktNdTvGi+3ImRMV3woCwyA4+9MtVynEP2dmt0
tgQagqaw/IBg25FDH703pqpNsHEyPOzq1frp3iAvDrJLx9BP5hjWto+r8ziKPo3k6/iNOsf6fyJg
TdrluuK7X5uW7eQ5+Irt6Nd/UdM5TLVSN5bq919H+weBfkDV/7bepGlYuMpzQ94Lx8FJgmB3a5S/
tmo/FWRSuHv+MatYIGah0EC7sHHPzXodCxsN1f6hILZ5anpwp1tbs2VOiGTZAV245Nc4Z3rMipZ8
m4lHh0CQiUqipImd6Yga+Naw4udCHil257EyR4rZ4bgRFFEuX8/sytGQcWrkC8ruiIisqQ8Ib5HA
0nz+OZWghH3BLqUWDTZcKJC3eYVXtNbH5lWSVD8PFaM81PqRLoFdRDUeI4NJNouMTkKn0bFl5Q9+
lfx46g+m+AAqKjwjSZPyPyvUxMKXcmrygcNxs4s4jEQQzePkX84xxdXA3du/RapRaXZpSKXiYXEB
M+MhqfssVUfOXD7JyheT8l5k/jmMHJFyLmLLdZOaYJgo4ju2mxEQcSyPFBEayJ4Rww0Xbex+Ns7Y
JrmCUDAoSwFlYNk4rNdlR+AilbvBung13KnCfavKkYUVE7RqmUK1LaoM/qXl+4hS+zb9LLrqrWFz
cgmmRBUkhXFWHvRklezKyvN0gzQvByobC8vue7teYRPNrQOmJbxhkVsUxD67203pT8lRmef9GOz8
DBNsELnyMMHhEUH8tWr3Y2RbebMbVJsxenweGNFyY7ACtLuSaK6EvJyp4sg9MrMPYKhTtEdj1aHa
0CuNFbpeUWr8c+jXFtQvxQEjeG1wiNnGdmXdN5+2HQ0Dy2DMpg2hm7673Ix/tmKRN+QoZAazlVMH
FHzoBMMUbvIRz7HvXAtXAsFDwmjiYbxolr2wcGZWjkLMiNR6eb6Rr6PysP9z/RYySqq/TIJveVTy
GVr9mBRgsdwEyX3MbTBAHHkyV4OPP4bk0dC4vcQGn0flIUzc//ooz7VwQuL4MQooxHo/WNHeDGcD
1LFG9EQVMXggTAy4DzpgWh4OWecm6wRpWSWF90X5lUMYhOkinBYaMZrbdo9WLTlNb+7zAQUmIeJv
BZldbwMMnfSQUI5zvzTMZNjcrMk0Hz4smgCUoNIITv3y0iWo2FlFMm2t9BNOBILJ1+h02qjq53/u
L8qvCSiOy1n0miC2qxj2FoAr4dHY23anve1skvJx2T2fG2eEMVog9lEaoxtil7K3Sx5v4HLtZ1DI
hKilMVpkOO0BptnMbKtQQ36giaH2u2jR3ao2MdEGnUZWLsumfAYkyd4Lvb10GNXRUy9BZCGCbDhX
XSuCJSvC1scBHwfXPfLXr86HeeRXPdK/YH8ghdxB0TsjECh5iqzAi0DARv+RwvC9oVEIryp+rbO0
iwGXDeYQlRBhI+v1mzqPLpa5GqIbG6WrBitioXPIsVLoJ1LNZjVOkI3GrzqG1wSOvg046pTdPhia
56WVi21yfltY6hdfjPwUMFwP/cYfCBJYKa/lK68fgf2wvFhny3Bt7CCrIOCICCqywq4zlVvYdcDx
LUKHFTpTesruGuDd3Fsj5/b8ADOqZGJ/QFHzwCP7tTZPViq8YK7Dirc1QXCfZCZr6N+Z7+BYXNH7
4NCQweo/Z499jfKK34c5gsslbOPVIdfnxpbfUv0ae+tIKtJXm6kTUhaK9t83Z0TSNZS499q3tVSB
ddNBCi7ilWXwWUtUqfXWPbFI2xwAKS/h9k181kZ5kwBNB8PAGv+0WTJhqJfwrfHxyfHWJC2zqKuU
+e/AK6nMAsKUo05XgYp0hI2LxwWJMqn7FaYEV9gjyOfXTByS82K2N4yKy9WJebPblD3cGZVkvB/d
Q6x0uHT/kRN8ZwYfBde4pDmVzHvZy5KRpDFr8qrCgCYNdBZFOFDLZ0334bzTuZaWvPvCSkrWBL9c
1UNhdnDCtHucTgtviX+I1XHnDRXbkKojXYPsCujsYwqTioRNfEXgqY+VS7khVhg8fuj6FLCPrDfm
hg6yP1hBB0o94Ry5f+PKEcOswop4oY3h7pOkmobuKiPH3kXS584nJjuXUwM5Sp+2CElWFcoKbLaE
qYP1BLm21ju1FzCI4RUJd72hvfnvvVDUUqu0ngDVdbb3w5ysgpKHNrumCcFY/Pm1L8udt1+IYlGf
GnH9wYIC2I3rLWO58coO4YEtMgTFKLi6nl/+Pk5gynw56wmpEOsUV3A6YmHoMKiuYXMfFnny37yQ
sPVHBjq8ZnaURh1gqU0fSSDfdfqfaLDkJLoR59S+gRC7NmkOY9jZvFXwDBFGWa0DnkjcgRuSApVR
CBs4VqufadbWo4ONispJknH5H2uPMFFudqDFqVLErFb7zNkXF4DvxkNFFHVsJu7n8fWhNasdOPJ0
eLeALuBt9b7v2W5Tz3ojUoAQUqruU2cwY2DrN8XZ5mzPaXRzd7ZgUMV2In+Hk6dt7jgSXXdLakBu
J5eKJ87AR3KxF8DH5EsAiTJuoHYDfzQQH7S1ye2kryrlW66RFlgboAy6b4nAgUNoRY9UtsV1ulr2
/K8TW/4aiuQI3ntXu/S01JSvqv/ZJsP5CsQwUpeM3guOTZGFeGRcbxB2x6DXK5Cz0MzNdQuAq5+x
9azsAnHDeB4A+hdDwzGPS9LDaQHGofElnri1AdgWmo7Q31k61l/GFRvp2+pkPkCoG1I8/+a3LP5I
MbMMTCgcJcWJjVexP9dNUZFsgy3P8YrvjzWRiTQK2mSVeCEZF1gqdeTgMRLX9xGYUA/g8RwZq5kG
oWIWPJEOPq4Z4oS3JEnK45BHFXUFoTUWgqPCEq84uGx78Uw36JhDwnpAKr50z/vOx5S89IAj8zGJ
bY6Dx7dFE/7h6NcSambQo7LR15qSsFkzbfICspzZxczawlKd1r/S820r2pGPlkk2N1R4iFfBMTPZ
eT50v2GPYffsa/r+idofNu1G1r5zR242irGyw/BopshJxebV2geCYrLeemK+qO7dTNF7HnTzNiO+
Ic+2EzjRT9orlieFpRX0zZRCoE2D896gbo2BhhwfxBh0UD4b8FGAiqwpsRKWsQupmLCmw5303tX1
7r6mB8iE71xzbC72v1sqMFWqVFo7bB0hjFSLpjW79rFlaC3y6n+aFxAGIvYAU0sU9E2B3snd37Kv
MrMKU1tuMmb76aQma5ocB54y4VWjCnHoyxw/i3zt6UNymXVWF7SXjG1Y3JmumRq1ZaXVHV9wYpF2
No0X1zDaJSAZVLI9K2BP9o8s/jnMyK5j9laFO6o7mpe38Ph3GbgkYdsrSpAFnH04IUuuElwVGXc6
WYaD2DbjcL2XAAXngh7uwK9EIZ0c3/oRxT811iVI542a6Ij57Lp9cnd+fRgtOgmXSLwumTetqQM9
3uvwLm1tY3F3Nk1ridDOUqeRE5JroJLd6shTlAJZyvWlwhoa1XkcoCP6iKvmkwqvLjg4XauEm2Om
hFUOcn08It8zsE1fHSoAENGh0ZfWGTwLqr/7DsB4xa49+UAWvFdGYOg9bwVbJNjb6sTxDOqXZq7U
Kh3hGCoqQfGZP8ufzgICs5ngTyhj5iIh+xt+AEFmxJYEqOGwqbM6wjjG6dtNJUmg9unzhmvZHO1S
H/dV72Y3/I4cdgtvG3nu/M2OcLqhiOAP3N2UV+EYCBsUO7ZciysEUgmuP5ZLsqSa/6Ny1D9TOvs/
PoDjqFxhzgJ6LkrRhzTRNNVpcnlwLBn7RjggWgZ/CaBO7BAqMiMDPpqpyJc0Q1kjglacHPYkMpjb
AtWiuuXsszh9jFVPIo18yhFyRC4NAi0BXGek3flxdNdOregK539QC4BtHvk8EFnpwExzAeTot6dQ
57rGbzNMvutBcWMcb7UZ+aaxT2/Z/4B33Q0Hu2ecKewQrBCXcbvv6R7cKuMk9zAVkFMgQp5eBy1M
HkE/jNEXNdcVBmVO/iNFxphzSWObDW5dO1jvFwXRbHVMlgRK+4YXo9nM/XWtjBrsTi6WM0g8Gl0h
H/+l5GwueqPUGmNBxZ9FS1Tn2OMHNhuzhRWhwehxKeK1ZgRoA0kfwMkYN25nddMPoeruDJW24VDO
8J9dPH1VesDJABdJuWA6G8NvVx/FfRd/vRxalPFwe18JoVKp8Lj6Mwqry+5PLomXiv9W6SGNCwVR
9am7cxKR2jpCJ7R2lobxGFA7T63frx/hSPrTkREGBZHDfPO53IrDAWovHfD6T3CB/k7YAi2oFSOS
s/3R5kzUzwuwy4TM4Py3AJMrsjN0Yvly3ptrlHZMsS6thO20zvzofFzouiOeaTPHvP7i9EhPZ5/0
bY3AOH1P9vBIBAEzaUi25j8Nf5JrJNTlgnJecST8Yce5jEs63kMwiU7j011ugH8lfvkc6l7vxXa6
ATSdtCVK2WNK2a4ex2Upt0C8ptigVQaN2Tr+hhDJfPbYLpUsUAJru6EL/CpFHY98oVeHSPEGE0T8
udeXLlyZqObvu/5VshGKJ72AGrAol9hNQWtaC7STjS4uslRVQw2XbZ/FVQyXO4LyxvWl2dTwCd6x
VnQ5rnPWMqcEU6Elj1O6M4KK2tHe9j/5cixNrZJh7ww+MO4PwAZde+1Nj2C0XkctmSRtx+lomOrE
QhJmO8fUD75F0ZE83mrTOiJ3whQCWzRzvo28sOvVO1beikpHtGqbbC/cifFaHs6eQcks+r1VEnLE
LdSA7KFQpKHL/3GkX9c+nd4uVMy0IE4Toicejj22x4nhd0+vjMw1TpWS4wMifeWqDOl3Dq3ofzb5
UQSDqjQlxtc9fqOLXSkx6AqGOw78qmMP95IoTSrCkIMJOKJ+UKkh/fYp+BXSzsi9JIjvUy3IKlfx
SzYRk5yt5TY7I29y+h+pT0EpRFL59TrjqRgmCynPsnRow9sXeSueLHJVk/S+Z0UR/w8XoTYJq59d
BshtYzbS56Q7vQNxWfOCGBUQGCR3gJ7k+P6TEb9KYi4guWbZy/27xLTPd5CxLKywxidpH1gTE9nV
q329BzrDkeDip3PPy6Qerf6JooO5vj+i++qh2O/sngZkdTVe6Ck8Zw+vy9fUcBW/iVBKwVT0domw
+EStcEoY1LOrLQM7m0yOW5mjgG5v7KYtcGU+esJ6pvegXCD8DC4qMWvMAZc5+bHuZYdB3y8mnowY
I6I0yR5rHn6LkldSROOvlTLUbtRPCXaSPVbFPLCXecnFTAr0XSTvHcyeJo62ZbZFD+DCZCODBgOZ
Sqvkiu9cG2EzMxIZdepZ1je07nbawag0s1S2c0YLzEJIEoufJTjQN14vmwCh7n7h2MyUqKZK2S0T
Acrd7lKQmjq3dk9xEEwO4YlRV46/p/ax+zTP0ggi6ekG3S0ybYcbSMuw3q3zYl91xs9RiQ0XUXJJ
1OwD6aOoalooIQqTxSwzOD7a0EQ4o6n5QeY+wfaYFYWlCg9Rj3Gb+UXEKGlp7GSmQ50+vLfnRk1D
UGl6SPlSDLBSw7oandzE/HYXU117op/m7is8Wwx4YawdzOx94W2rLfgyRXwzvldrQTO046Ly0AgV
vUX50q0Bo1XAY/mE+r53Ohfq3F1RfPdKhwtxKwnD28gvncDjm3WMGnyHEA7JeGuZI+NcEKaeGcKH
5ljwubQuuM7kNNqgemgC9Op8ZTwdfyBmYk3u5jGIg6pnI+QRj/oQF8fsbKUhRVH+HfMUxo6JDrcO
e2KV2XNmN5V0/r4POxsaTiQLZmLJ1/p5/Q2op9+vNV21HytOduHd1WKQYkRqDN6FKL9L4pf4o6r+
49zPalQ/xTiptAO/87MZWAOrHhXPLe7NryHVaU8XIURvw4Cl4G9E5mF8/wlVE10y5Hx3KsMQkZvs
AHE5PdPiakoXQkD6T6kGrVsdo4raXqeETtro+HqBIa7gKLEZZKN+YGnNSI35RFdIGvYjcHixpkRP
5IbmEAjISZsvF7x+4rhTKP2MA4FSztBsBGTbfwQaytUvVQqgslPoJOV6JFwFbYs7ChUdz1leCgar
NZ+CfjypT3gHMed1yeODxxkOuCqDwjNN6/d84iW0Ubpcv6Ynlot0PB4aw7Uxgxp0MIfcX8oPLrBc
QesyjCkv7VYytQDkY4pqdgybUu/pKpyiDOdVcQOULPUpp7KTf0TwpOqftTakHg6vZzViRx9PTa5Q
5zJ41Zeb0X62OVh9Buhy5lFhGpaC3P1qkadN6w2u+JtS5IPmtoNoH2q6AtkXHdBnBGTDVJ6PdiDp
uaahgf2CqvNGZjKCHoQvVtsZuyyu8Z1/z4Y4xmsdULZ17sR4fMs+1ZORDAGWHfUXxYmtZQyzLUpA
o5kAwPjTSDLv4wpy6QDbR3knIMyjD/A8u7aU1Hcc/CQkuiJMgW0JctR86oHWD9oYQHcdDSwlegQT
M069vnNUVHaSYqpPgG/doNA0HxFG1tBvm7ZQSs2hj4AtGsZobml9y750GLvb3ki4bmRymtMBTlB0
1op8rPqiANQYp/n3FtfdmskGISOxd2+eA4GEIGSAtH2bprbZ8+onHhwz+h1gU2U0G+BwLQ/4lNLC
xzvmsVMknLBLC/6wGC96i0Z1TLX3Z2ZGiViJq7rJxFo4M5huguv2yK2WhXjwYfB5A/wOjnjIC2lv
frArDLDOcesHc24bhxbDdmiT8mrESCoUXsWlWQkbfKxy1sjT/Ygk+4Lryd+/NS1Q6lHrzkXDXBpj
XluKEY1ZGO+0z383lflwS3bO2cSisZtWk+JM1eCjT56NqLjyLZUhDvJrjyJfRSADtwHQwp0bFqoG
Bd7LmBpiH7wLV42Q5zM1wo6dZZSld7pgmvshSwdlOPlMw8HQmRYD6/ivwZ22Edwc+1pfQdOAp00Z
AcuNfKowctqYjqZsPFzW8vep2vfkpIr2RbGoy9hnf6NdhqHR9U99H8bGrjRLPyY9L3IAwmpnkrRC
vHvLTooYRWikI3nOf4gLUtWU4zrzUbIibF+XvfQQDtGJ+2/RS0fzVsVhRZ+4tXk4wCZkMjvNRaJH
F4BNkPL3DHaIiISJyqIvrYOLHhlLoaLdZUlbYNLcW18ycQ6IibL0sizknFu3NN7RrfHlnYJUwOdj
BLY37WfUt36SDiWVT3+9XJuEIxz0nhDSEGqpiDAC0ruKrNkdqzRGaQAQvuDo9thAjGRZawN1DGja
BJ9FSiT3ggWFfBpEQqGrKsE6DDjCQVLJIV3PMhBXntUZJMoXnfMpAKI6McODfaWElNJY2hT6ETHS
/Dfu0iKEq33UIJPUvB8s0h2W6U0UjJLTTtLRBC8CDg30Kwmo9fPF06mrCgP6kJrdlwNxW6Ju0Dcd
o/dyVenZZsp64Yj531rYUY5hqFk4uwlXC6gfMfmP0Uuxd5uP16S2mJNNx1+wz4unweShAvk6JqBT
lU9hF5S/nvG2rjmVDg+/hoa5OjfdVCJvh7dSYrCw/LgeTaJg9Qk3xYvLltjAHLIt28v5SfbaClqy
KkSUuZLYQpvhsiRHkX+mIMmjbpKFrJZUX3yyTq/Qzzpy3uMf7Najx7Oh74G+U1ArNCXDH5f8rjOS
G0k5CZ8mUtnzFe4mm0yjqGJE/j2eu0pnqlrzWG+hXWbnpzT4nGNqHewJKIJG2ucBJYTCrQEZP8i/
yIPEjavTRfpZTGBRNbIIdahSsfkR6sFoiBK+BcBeTRi5zW+sdDMSCwDpadbAkxCp38b4hRTzILUm
a2klZNqtVoN2LjZmmKM8+3Zn3ctGgiez6TtuMVUJgVphc6Y9MeI2mkSOW3dh1xmpr+TSW3twdqL+
zcdpFWbxNh/nYCoVoUuf7gwxFWIMGnyquGFKq18CiMTYshvPn+ulMeKeR3DPKtFfFYXEh0nJiGqx
dhb8ti90TxhkMJfTWD56BiZkTrOMrisyzlLBMUtG2QJIKCIk7reMt/0kdq4xJgCv8tUjAh+KOo5h
/9Lrsc88IfOB18ryt3BxNq0NSo2hqsdYA6kp4S95NQYBfu2eJbO8ETAFs5m29hu98V+Fpqus/YjR
fVAYmJDRfth7jXBBb0rvwkaLGc3wV3VObJd3gDNQ/c+nWaoUH3DB7i9ipHeBiqil5QAL87PbgZaU
3TQoYKSyrzsPJggL4/2gO2EhCKp9LTbgAdrQZBo8PkrayvOvbqYdSHY7owpkphNVm1Ec1eNvHpzG
INaUmmNNeBFUiS/LfX1AT/vQXkVL1IYmx8bt8T+pLyx+F9QuV768tDbtEJGZcK1DJuZxQLbHoY6x
9zGydZ4Ro6sg5bKBnQJ55/J1+gg7xEOPtuDRh2iJ3zUGmeRJ/j38H34d2IMfy/xQ1fxAj4U2L9XS
VnU5Hr5NUDBe7Skgc/vGKnQQFMCV0zbCM4Y50beTSvWPNblBaX3hKlDMefsPt7siR/Hk1V6jL7jk
dhVphzGBeZQR0RDrp7WTNGomglgRaw9CdCYUeD0NyTAz8xhjTj6VvNpCLKumje3mbiKhRTEYUpNK
+xYuSBT1VwH/GB/Zv6C2J1i8KSC5nzEtFlEsC/QsOaRZP6VUpzp0dDvjpgZZPbss37md6UrCcx/X
gNe/nUk+t19TYSQLNrTfHnjC7mZPGdFxl++8jQ0V5n5epfw03hglG65kI9YqS+TLbSq0+hj86LqX
hQtpYIm73e06zd45OsiFl7/XHJ4miFlSJWiA9kFp+e5ULbAXBpBQC1vJ0uGLg/X6Ao3Y08cvk/K9
y8+yWMEpsT+yyCMQMS5c1YKzaE/LZZhiPKcva9SlTzNuXfhBFntwPfO2IbgSc/bw43w0DU1i9ey1
qvC94+RCetdVvCZ0FoVSFse6ERBHTummIAgYQGVuBG+AwgXlN/4hhcA9KLFetbZpi+ejGVW3R1kM
0bC7M92OT2zk7NHU1NDf2Yrdq9xtIFEwTtRxeI23Td/hWFJfksOP8YPjY7KeaQRbGkRXBJvI2xYN
jCoi3QiPFmfFlttZCDhGdUAzFwnTunpUNfRoyvPwj7lonT6MMpxHob0nFmF3PUy5Lb7QGNrQsUbK
Ods09Z6eVuB8tn4qov0EDggktxBo4hxzYC6G3xHaF2+ZrH3i+Ai4P6HhwVFTSIWVSQYigp1gMnBt
oh+NF9UOc1Yim8jb2NyFRbb2dBS/NaxIDDnBK/QO4PW6DgULBZKArVWDeMwx/jEE6LMXWlSU3NLW
4CXyb/V+Wq+XTzvUCyu3Ma6qdwKlxViqygcSyW2WGFa9GgqK2qVMpYvbzADXLFFmNMJqZ9aEMtk7
WW55URpE5r6+sJuN9nigoBc5HwffWoQzFJy45S22EO/j0BexvAwnxCni19msVd/PsFmhyiCW2mqz
vDHbgGPwC+1jqWDYJYtsGxFHU+IAp8AlB8LowbX+6mYQGkwRlbgggXEJmnf9Qn3OIWHhTUkTq/xN
Gawmy64katApLE4trW3LBXFbeQ4bODK4sXINNi5yS1gNchrXJPdzJh/fsdftZWzSrbvVtXxLCoMj
/zUD1GeWmxO/t1VRPCoNJComf+oyyhzaKEBXJFUPv7BwVGu3ytGoJ/s/DDaTiTQ0S7MEaPBW1Hy8
cT6SWbuk0cp3tgRPAtAzUcFDSgaCuql72Dd74U1d9IKzSvLV+ApeIPECWjiB/4Qj+oE/1oJq2y91
2RH9fUr2vw7Arr6Bc2+vBcJOgY/4Y1+5vshm+s8xTAIo/5jdoLQFlic/9UeaYsPXQDnsVdtBvLqS
TP7YWZbt/HRZ/4d7e1kMHSswy09rJV3y8zhFFqD0H77J9+ko/sq2f1V2+lrrl0MpLiDqmsrjJidH
o1N6hHOUJeKLOtolslOCWogol8TFc0wO635LXLKgjfAux3n8/cNM0/TCPq3LLTrTWxDrmC7Ph/oX
RnuaPa8HsrFZxgVdexoAnmWPvs3aqGlNuDaau0dw+Q3GhEiEgvyPngfqxm+2VH/vf2gmVYpkSDjz
YukSR/wiKs/Zgd8j9ZzpLxPFpiYuPsIzUVANDpp25xTgzDvzIYlJH8kHsbwi0KcTSybOCw3p43cj
SmOPPsWBKf/lmuUjoh8Dm91LxesxAQ9NZm/fPxRBI/iuls1lTSu7h+z0R8z9UH1xmPLnxReKbqkI
oOReJOVh5N7so7DC/6pNePB3jZ+b0x/qfzkvhOuMW/aQI+uKg2sIA5CX6USSYl34fmC3xa+ceQxA
ZXxDaH0IJlZ8mz+pVyXnUmv0W1dHXZ3M15NP0Mk97cBGf8POCptnWD6LN7i8+BQLQob5EMvEl5Fa
sp++2QjzHWtQ5htwRJaC6NTuJJoAcGJdjl899ocdqxIf10cD7jVmctg+6VgJqi4r82H1euS5YttB
a46K0o0R9naXJCf3+L55YantJDsSKV09qb8ohBBul5lQCU644iwk66U2K4hwQ4XToniCe6VEuBDc
W1DCDTQM8uw71qJ07OVj4mV8Hvn/5hG3O9w9jrAmKDaGE6SN4nZiGgyRHpZdwIMLH6daRWR1LRC1
Y6Kw2B9RwglGval903qeGZwVu/OAxUJOZUHXNrD5dx2kDPOpIxldOJ2mZBX4v/Eki5wDtrVr7UDp
ZGHdzl3b1q93cl9EcC/FWvY6teWPd2ZexNTjYMrLIfox6rTA5W7a0Oy0on5T9pjxyYzhfTjhTfU+
qEqnBvCnBnwVjqnM9nEjQ8ii5MZhdjhb0md+Y+NRumyOPPYHJ92pseP9zDSARFzDoD6tvQR6Lg/0
IMnVe8Xlm7WbLClwmaVv8czRyguWKgwCmuuEYdGtpIMEyjc1wdem/9rV75zz+NdN8+bCZhMAABju
9Ly/I68E8YiB3x3r7C+xo/fcQj575xSiFtrsoL0Hvj3W6GdICRa4knqBW8IKUl0NVc7gPfDwhIPr
6gb6HzfxmN22fV+T/wpIioUpaLB0Lbl/UJ1/GPa7i80VBKINtvoxrxwPaiRmpCe+/PUg9rahcxYw
SwGXHM7ZoT5bHHY01xaPAKyyDNnPyYIFamjxwcsBaMxyKiV1XbZwmgEK8dcMKofTZQsVFI+YJFB9
I5m8TpZaUXaf6hJ82Hcsyln8iIm4M7Rc5AtQ6j6t5kukdRJtw9tMrkNDUWNePISI651j+Lkfr+WQ
45lcCUarKMfJ7rmGoA5RLu3AKbOpfX/LSioFfTebN5lB++1VIR82brE0g080E9z17mV/Y5p3Ekz0
ugeXTh/EiV06mgL0fdu7mpX1fHc5moSjBBbc2x6c1H9mlBX0fLitlwIx9YAFZw9AJGjkSkuBTeOJ
doLqnUVcYiBUzLWvO3hidx6b1D+FpQ5z1nS6CSUlWd4XKXo5pDjcuIfuoHl6mhjE6ieF09QClCHi
qz9bX05rMDwD8/Tx4zTQdX/GIDZdLMZ3Vt+TLM3AQ190VyQ3yDNNDQ6TUNq1XBP8gPcK6FcHgOda
iuwd0Ws4og27nwXLt3LnevVx15Ey1eMTEEdSiV8MC80c2EAWxVthHMuBUBW5Va7sUR2BqQfkgk8b
kdV37Mj71O2jS/cKBLm/yxKzBxcbH81c1/4adzLhHV0YXmB5dJDJbtX/2nLNsinCnbVtPYjAEKwJ
XgHJkzwhQuHvlQ/30R1/Gx9t1ewmw4+BJH5kneK6yOqjcU/RpyNQc5rr7nPf4NGhZVRsDQ7FjfwF
OWHFNSH4uWp8zX9/5+Y33qAMUz1QdQ0+vwC2+kZRZEKn0bMJyz4V/TsMBfdIhIbAZDiTf3EloJmH
LRnU/IlYbNkK7Y8DkZ+RRQURqZZkfAwj83p4zTk9V91Xl/xKbFHeN2XcHETf3+9ZfEr0Ly9vgzvf
2XlA4N+UuW0kfpHMabiwpJ3ihSYDoXsO1wImLcwnYNFDpRVhfxv/Rsd23vZJQ+KV8KWux/YmAsgv
OPvEuPxNdh7ZprXoyRYwiwmH7Bp1+iz2OLFPO2c8YXGaD3TE87GQt1dra+5P/9ejVXdCs1OeZuoT
w+MSjrxBjpANXpNNOH7Oti0SmM0LzTUqrTxphP30KTMzCX5zJ1hLpY5Om7ZtM3WO6Ml6x6F1sJA7
5EvCol4rDZ/ENf8jfVJFnBcdJuP/4j/vNgC7bZIfOORex/iIOktmR+00NE6l9D4btwPG1A7Crk0G
9igMLdkTExe/2YpBOvjzqjJHceVrBOg3mIAnmCkroiSia8ZnSD7G6bSvAI0NNQk61/FvDL+jCF0A
j4VUNk5RI1P4+viOQCAeWZAQoYFBvciMqU1NzKWAJ9LgxgHtezBNACzWiZp7VEqnq+4h/j5hntv6
EoLKrAtxtch3/6U1XFrH34ZSEhaqoZvDkTVPj2QDl+SGPLZJkDtWgp/Kl06Eye6t5ssoMmmHdKHj
2WZwPkyN1RDFkjnv+upjOo+L6lpbJ3P3s7KLQDwT8qgAhzKvUJPNqcfFd7tCVK0nGBuddi8pmlzg
crMRAIS2nQFXemd9friKkPtyUjIHe1IUxuvRxKv9RdmMUNCwdlu1BlVx2Mm+4W+jyXS+dDjwU1L8
y88QLP+UN9wIYHBbRJRRoiZp91S6c63fBjSAGIdsqzsLtZxJrU8BD/3epg1KvmSG2XDnKpTquyIz
u4Z4QN8OcUKtI7coUrngnzOgm79LOVW1mEcGlHjSld/e2aIRzC+TQwsaw7hhEG2oVHp8V2WB/3xb
EmXRIrC1nJ5jmJ6ZnyV815je1P5gqwSCQ5vF/YpFNW5vkE1q59uRLUT5of5lfMRQtwiq3i2KWi9P
MGnv7b2rCRWOuCMAM2wcyzoFyEv/JiQqJSIWjd3J1SZ1Bnh2vbjtlhIpO7Abx6wg68D+/UtBKiWZ
mOeiC1dV54rOTmHMZh5QqKBOOL1BUu52t0lgWb1G6teC9SjhTiYlsL8TKs77aIRO606kpANanCBj
fNIU/89RC+SKMC0tN+HsNYaBSNeuyCU4E/+A1hblZolp4nDvEqWc7tezcO3wIh9md2OohOwfrncL
HNJ4qoPLN4gGnFVCDm1mLbUv6e5pQ58aumimPhmeJmVeNJH/eGxB5xxuXnVflaNcZ7uqouWh1DTT
7xLlB7jR6fCFkRHJ4kJEmXW/V2xO9zdscBA1l8RW5DZljyGrjtlQAJ3oGb7ng0/HrAzBiCMQjZhb
pNzvG2dwUzq7KZz5aJfs/eIY49C09N94JIORs7jeRsxLUJw1fz7hNJqUuTIyHy2X9wZCV1E9ACRF
p6jXkinnX8sSoQJlKFPYer/YMdnq33G63Vc9iYkAwfkARUxxlaoa7Z1tFTAzz5Wg1Wmy05/NEite
x4R+jRPEkvUS50U1Rlp/iLAQnFMoy+OWdp+yu8tUsArsUOXFJf8U9qp+QcACHi3HlQLFcyF9b+7k
xxHateDpfcSYsV8OpafshIoIfQOrsN43jupJj6p10lqvH7A4F2saUFFw9ToZmbgTa+Tx1NFeW11/
j8efaBhwmAtT5ggNACAbubCIm1q8qWYrjZMxCslGrU0PExAJ1pHXwk10U+Q9tpUyCCPu1Vi8rCHM
qtqwEALjesCFhFiVNW0T07/rSkSQ/ydUfKGnWt+tWnU8PrM5BpABKjPfZtUIuAeDnG3ELfEWwB2L
iAPtpuMHVP6Cg8UIQKMUvdLkFd6JNo5eM1cOAotq06dDs/iyGGobf4d9Vl2nIjZo5X1py85oWHvW
40KmB0yiyy8XJ3oZMAcSvpPtzvRXoSEXX3G+WCbs/rIbQV9f2Mgi/4zwCpsIOIjjTt7n4KQnWzbM
5rf10Ea500yEGCRgkpC1F0j0L6Z5AIt1oFCEW3C23MFMGZf0sm1l4sBEfbppladPJUaESWvzvXZO
XMPQ3BZNoQtANjAB6VUs59Qd/KpneEicCoxU9JnuUegV5M8FpD2+8rKHM+cvoEEe0Lh4BbD4K9eX
Lj5QKGc7q1N287A2UfpZTXhVcZpdY2poIboyZAyXVrjBEuwsz42pQdf381hERS5pqp5vxGe+IAIZ
QUBsrrz6AFAkT2+o1eDnWlaToCZlHPiZ1BhEfXE/dUP8VzO4jiFqZEuvQcGFVD0cF5jy6VyfzLRK
iqsjEVDlvDECy5nPPCBOqZZafuQVhi/Xwyp/eg4cW7+7s1mK2JomHjIO6O+wc5+1sLYe4LkC5TV8
pjhJ/otKvY7WWIP5J8FDD/r2ckLAzUGUEZtgpWuVC5v5nOksj5jUcr+iOMFjr3Xx9hWEmQaJFs5x
aG0IFjMFEQarzNXnB8WWdefhwu+BK7Bosge6KRHNWBloRdyNFKmGjG/s3dxcWUGIEVOXJAQjceMU
F3iw9st5zmBtlTF9wjd7UsJB22FA0pkYONiurgbiS3s7L/FKZ6OIKyJx5Q4Ce7xbYX9ENLmo0rsk
fZhnhoNDhZ5EuvliFo2Syy9BceO6vcrAwXcy3XzpBYFZbf/x1sQzqSaEvdnbujI8Um7uItGihW3C
eHLQImhoOFfD2OiGk+I3W147Mm9YWgOlF/y2auvfRNJYA1xdmZBVpeBGWeCTs3hgj7TPypPfUO5+
qwJ+k6hseR+STA9mJ+yVMs+T0F2HS9mmE62GJNj99egpY1WbGR/cRS5vvA0qJXZpTn/njEYfhnTq
xnAj+24THBJKOXCQDpf7Q86f27Q7aWdKfeC0M+iGre20kuK145cbI4PvkMh1QbpUV+owZksB1Qm+
UKZtKb8SazSaqNAzDr3/VO2g5cHFmQ9pE/Q6BFyP844DifOJUmF6UE4gZpeTQiPbBPPUbkg47LNJ
CigyFmTswbsAKDzB+f5NzXaJJ2EcNInjfkReA2zdGLt3XIl4s/C5o7/KLPxAKfqMdnpDG5HAApeI
7IkjBPJfKwjxCAjnR4awWrkZ9usRivzfLT3/UM/4MQHb0wXZAMkM8dcM8Dy6WjuTJlb4Iod8PQfc
Wxuwv79v7I6gw5IEjt4WXwcLLkbFojE7P7ftPdFid0ZucCCY/nD9Ax5TrRo2mk2x7L8WIrMOXjN1
ARoCHECZQ9k4OvZWtZXU/AiePkQhlkRc6P4z2TCthYBKPeZgBAWogMa6ztGsckTQ0xFAI0cyGsCu
3SRjzQ8XVvNMTXKS3ZdSSc4p8dBCxIdDJ4YsrxJ9A/JbKjH0hrWou48uJwgcM+hq2vyRvGEzw0al
PDqWfrENigU2xLeYObRUhVFkL3VQuXx5S0GJ+/4SuZo4AtBOJ+lSGzSX3DAspnDxBjYLwxvKxcrs
kUt6U3SgqVPoqFfMX2BrNEMpNIQ6UV4Zhok7EoiuiodwAe9lL30NaSXCp7tDBOjqhNfGs7cPQmVi
RZ6IAfw3KHATGiWk+fT7AhxqUqASUXC3tNgsJvnMJQdzCrdNFDbehcQd/y03iYRwDO6TzlVArPzw
Zfp6GwSiyBSJmdhgt7MaTzMdd7bEVjhqxKlWPOnze+S06ylEkxatvFnSZEH3C6dBrAZOU2fkZ1jz
wD6+DzJPW3Vhdgu1d+6IInv2hoOVTDg/AnGSZb5LFrhnW+MiQTl6RVAMrXzcbSJ8R41EUknDXEOt
zTzWNyWiz1JUlPxnemsWWrI6TVQwem/nbToxui53qCgn3XuZIZX6ievImHqxe7NXwXSOqQFgAH9K
Ht0QUGipd2P+auEGjh2oEo9NTwDqMhKKoooeqBSxxRT1sKfFeTzyvZ6TBbWdFRUbam2Ozvv0R0Uo
z03Kqec7qT5o+MIJ9oTNE5O4nA2vlI87fz6K/NG3+A4JxNiTtRc1JzBVzkA8MIn88fBDN/67DaVH
4fsIp4rj+zj9bkSTSLmGYQ1Z6rN0a3AOwqomyFRiff0Bulg/EzHe1FXnt6arr+WyqLrFgw4A41vA
E4OlVNJU46dpHkJkG4KMgjGsNwnwzwX07/3TJ/l3/WBhOy8AYaTrfSPIcK0itNapd2CHF0BkpwK0
sPr71NxU0BdWFltDH4EDDy5VKEly4MEtRNDgSBXasmP3kqQUzb7HXLkL+IW/0dvHO1Cjg21ucqMn
YYYEMhTrxO1TG34TeXX5cYn9ork6E95CT1YKQnwJQcTAcTq/mw6Kgxx4DfFyxLkD4QrPetKqPpAd
ECfZevV8/fHfCHx8QLBLbIbzsfNvDyIOX7eldVVJAJRxd6Gz2jszOe16Es2gnzYbI+jUG7FYIYzV
uei09Cv3ub+dt5p8lVWq8JO0EKAsGAmflVdRFNnApMU69RFF1k1VoEI3gRPmitwT4l/KcWK569e1
KWJ3qSv9+ZLLNdOFCdozrvy1sSOSodYHM+7WbmMmTF7Bq2o8LeNmyegKvAq/gEgYiRwl/D3/7jgM
MtIgrzlXRFCruj+I9aYjAu2QrSMho8MA4yLrJV/MWE216CbD4rDiGOlP7KoKgSbUtG/Gavmmftcp
YIe62uhLPRwhVOfanDiqijmxlsNbUZgFUjGmwEQWHLUxBHVzfzJsfScJxXWnmNrzlOfzKdh9agm7
rWIzD8kBrRzQBl/w2Pqf2ONEDMCxlqudfYHd5JLmwGSWawS+WlwgL1zBTtScN3ITmsJG13j161pC
6Hneu3lZLgEAte+bhQteVMG8PRYk7EpEzDnSN1iSFRQ1c9+VVp4WjsfzP4IzTsWAUdZncvGkpKWS
deexIpR++7ZbTwqwpdo8yuABuujBnyEK/25NxKOCZ+D2Vfx0RlBg1DZhWvdH5/cdCWBQ1hUcgobd
A6dzMmtsztmOJpmgemKP0eaLHJ0/EO2zsm/ag2ZKW8lz9YxxAXVIgAI1O/8o42kipuEUDihu82RQ
jUDfhg6ldEQn2ctjp7gCdV6VUNcK9/pomap3P3Rh9t14vTFN3c3nyUvoZTcoo4uLRsn8kNciNWB1
lAXZmK/RXdHqeIeTiCfd6UsbCiHgsyZYDskJa0y9/cKvtzh//osBPRL5rLSWV1sj90gRihxCvCZr
ABfnw82G/h2g5WFFb7skJgWMS5y5wukpRSB7aloa23z0dpbVL8cAGDSl3Qc7Ph20TBkN3ddgwUx5
ZO5Ed3GDYDJc7FsOXAOW1VAWBysy7IgddmC39qYFvq5qD30GB8vJL7kBH6NuQFPAKUz4mmIAr3kY
pfoAGId/ype8FLLlA9ByDF8p+dF/nGSpGQ3YkgkvL+VURArFcB4g0PY9l2/tOALKmEhCK1Tw/5V3
61g5wN81tHGAEqvNlqawKgL33WjEjFsic8e2T9Ach6gBb0tJGab9g4fpN2cO+aYZ1BjZQDngxkfA
bu7h+jRHwkzimEPwKttXB8wTLPv3SoJKA6XSGk2nOlVMXD9+odna32ij1q1STkbsHswqILE+fs9V
7luT8Mxf3JhFePswgWHdlIoHAvKia0Dd1ZBo1kRjeLvOeMtpJQyrHKpj0mOofFn17cJI+bWRiByS
rdUbWVlw0oGuw0oHv7zfvnqfl0UqHkryMj7v81HoFsbG44i5mhehccDvOuVaXBvSJ+S3jcLn6Bqp
1DrQlXbQPeUpvOc9ezruEGi8987Tyw9jVjLMX65WfG+BZfowU38q301uJWnHXB7kZJuyKk1YERj6
w8odpRRLHxRufsxE4QorC8KpARazQXB3Z3WfA1qYqg7Q8lcgaNSLr13o1TXRoJWMlOCAx49E/v+Z
lsfXFBa0tcP5kMB2ghCGgehaJyFueQvXvy2lciBu2cCRkXBqeiBt8/HSXOGADvCLx2gybOX2iSg1
7RkxaWuTfZwgyo8WBkHbSoTyb3tTkQTvI4kHAFpr+1jT7yKH8i0SloDMoA1e17ksqINIx+RFiyI+
hDOVxxtrx3/cJ24D2aC03QVqLfc5QFpvfxOztabg1hV/QuOSVYdjco6J5H+qAP3gCANUiEuQk24B
abDuICUge5yF+XyB4FILI1jDBajXXdR3B05cTXt5bkSK0ojCwQN0azp0/isIDRmtmO3W+3/CRY8X
4ROTGfaCQ+RLpMGCgPu4fu6eNzqTa1HFc70HCbHrAAwBYrLhkK7T1L3gn4xs5sE5tLWxEldJ+v6B
eeZ3yUStf23dwrYg73zR0EotoHEjGptQQ1AQeZhJQoIgJbsEWTLOL5ZvEO/dbnc48UA6lKiRRM3x
XLoXNNzn6bC6Z7/GzZXykXU6FALVB/nn0UvmIkAkcNQLfaOvDCKlYAbdvQ3jptu4iEd2u3LX0z01
3UHLMToEfCETd918aGRnVZR7ZQlm0jimIBFxS3PzoxbGHWFYPhOe6LOfAsJPlt7pL49QCnCPGxmv
JOs8MWkzgtMZ5+JBv/U71b+CXtMrm2iDPX7gHOwMWLJpis4pNpUj9hpO8ULZa3+Wwp0drgY9qeSq
k7p4y6I/KS9UoOLHStFSx2+RK2S7bv82J+ryhMkmrOYPzjQXtZ9GzjkFLJWqG3LYCIDWlqcoZuh7
HchEhMh6KSG/wncVbFMh3AADMFM2ZP8+FlrVjO9s6d7EVIlseUggQaCZp+/Mvq3Oo4Q9+6mokKV6
Y7fyyCKCFcP8LDeQpQL0HGXAHnWSrwItnkNd+2eeJ8XE59Tfwe3AIprWLuDaeM/N6v9wG1mcvexe
1w+qH0pT0JKw+euFJVcT4Nxn1WDPU5VsZpceC3yS6+X0aa1lLiHf6kSw4jk3tQrLbONWed/cdsmn
Qg+pmxd1jFy5AwkcGGymBXEsvULL1wFbj+Kh86zoErfS0YURL8nexciTF3fcFQHV2IbD6DY5LfLA
+d7yo/6H+fC8lp2h3/Kr3mPO8bGGUTsPE/CtSAt2PAmTbgb1hLDmw4g/e3gO/SwyPCn7lPQY7WiE
j1TM9dZdmcZdZ8OdU70Pt5Oa+Y5wviBVkUqb+gbtvxi2gf4lTP6Sk31cVOCCkUSno4/V1Y5niOKs
nPO465ces1Jg8mId68/B4xlFJ7QOTR7pwd9ETblR4NAsAcFd4O9CQFcaTKwPC3mTR1J/pgWokNSV
Jacgb3zYDYfDXucDjRi74pBEtY71ziaJMWNxxAqttBf+teyoYxM2feEtND6jhNLYosC7Iqgon6LE
JKysgc30+1CZasJQqpJ1BsFgQrlK9oymenJk2wSse9eEqjSFU6wMbbLyrUoSk/w5KQhRS432T09W
YVFalOlvj85Sss7aiulWxhbIxht0GHCjdHrsSO8AcVJ7Lmwn70HUla2+o0TVU6wSF/TEOmxwNWKm
YT6RphqleGtkEZDcQsjDodGeN/Uzj8V3ccKgtJRVEtGZ8/dcUYQ31tAR5ScBxx1p88DrsGOHPauE
o2AD3txnfHansU+NT0of8jC1n4Hmaf+zFXXk1UdWN8ydUNQAg3mVFLKHwMw0+tKsgLngEHrvH/T7
3i9zesqEc/QZnktfGaq5yZwHDwEhIbMi+YFK08AZEl9GIMPxxocnOQwOw8/DQgfd4QEagu1Z0awq
jFpZFOdJAUVnjlpeo7D2o4q1C8L235HNxUDrfbZJqFPN5/zKkwQbOt/yhSzUtCCwzx6h9/Q7bslv
E3NW2a5kt6CiBooj/3ZXrAZhUj4TnUtAX7Ls2xw3msMPLb71OVZaBb6/Fhv1etzf1FLXGsjr7kJP
jxnNpPylCtq1oLJFz22qQUxW7Qhpx6st2H8A8zIUbRifZgwBEWvSZbRH8DsHGiQmNcr+ZQwzWei7
evVXre5x94Ew0W3A009z/aRu5DxUDH1m1UjDhMhcEGinhVxxQuqRbfSITt6h/ia9llAgXPYoTFhr
Ezil3e2+nRtCYl01lrH6HHJ0/Gsxd5Sx4VVMiPSMI1/UPIchIJTcXioVQRwXmk+ia1Wd3dIQiZ3U
OrSfHAgUsUSUEA/3MCdjB2WiiRpAZRmAf+DXbnVuhvg14mIjrSBTCVN/tg42a0hD//DHO46B5DnI
M5CszVoNZyuK47OoQ1W1V++TRsFLhzHGKeTsK/86g0plsp2JVjFdYslSu2Ja+3/0SaAmpveVtgYi
nfJ/8XKa0oZ02cOASgyoldkP0aDnh9clrvLc1R0WzZUHWOXKR0KHMMqdyp/hvKN9jNk7TOB4dR+T
gYNdLdg7YsTUmCNUD8+ZdHyRU+Aq0aPP4FAS21RpFW8HPe5vD2PE7V8jkHdko7eC8GFYmOg3NwGR
I5YgzIoifaPXCn/SuF69wElJDF2BvQ9du5NsM5mOF/57EE5lp393tZrcFjPZQpWOMT2CFXS6+cyG
Qygxyh37/Bx/+mk7ouWaJdoYwUK31kDpgSUDYRlt5naNNKshntG9FC2t/hOmarPaIn9XE1lZNdic
K3pZtHYDlYMbUPMvgrFe0XI/uP90JjshQrBIYr7CpV0MRvfRiSql3wBc9TDmbJA7ql54Xp4L2Q4F
Cah04zbn1Co9dmbNJLahate547M5f0S+nHmThzn19UgXvahPYWtkTfwryLBlE0Lwd4aIq18LTU/k
zETwrF5E0eUpWS9TPllGA6wGyUm1nOOE0kzPQKMG9uOgvAY/54cpOsSFVP+oDXLGgSmrKmVMJ6vn
bGQjk3Pnr2EjGRhnn5k89BgEnwUP5vekr3FKMcCkqwHf2L+IvZdNfsZ49ZapmGUOiL6Ajlkg9n+t
40uDDFgO1EQXx0mJfpQOFuB4a4INUVpmkc8Jgbm18rpykR9ZSUU2nmoyVwm1PGjZtNw5rQK+iuyu
nvyWnuF3s5zrK/OSew2aOzhfLVv84YqP+mL1CSiDt3iIDsUbMRufuIvvCLXp6lrVY8QeQF/4HiSn
ZXa/z2sbFpv80rFckrhykQKJlAjkDGcYEpbrjemVLJvb3pty59ohVm22WkoCH1g7clsPJxf3xIm2
RwZc5DfG0w2ZwLxBp+0hwxcXBvVjvJL3Sgktjw5kiOxhnpHhcL/bZo5xqa1AUuVBp+QsbnUaXcDQ
UY69Tt18EgVcEQ4LkeHOhP0aZCt2ZhAP/+cOSOAlfIGb9qm3EDIJf8CLRVlKNWkN+QiRismCTNvz
c2tpbXmXmovGgNSNXy5nwKA1N1ZTzx/BUvJGnGk4Mi/khnu8iT9ZOUweet8e2eumciM/B7xt4yYN
HLC5Hfqv7WfLwpOvRx2n2Isiv23N1q0Se48c1Jf0Yz8mvKnI4QnoIxBns5ZVukYRhbRsZCmK859z
c5X3prS6YUSrvJE1PPCwYV3o9bvk8uSvSPzsiW6ifBAK8UT5M+GaUo17t84vtwVOlROkj7ij0Zv3
E/PvyQtAwYu07udrwym8Bb3mWk/9vQ617ROpgoaTPSjLlwPPswFfJdFj9LsGHtsv7Mh+q4A06nSk
Qblh7L+cE6iaMw9g2L6XaoQaDmS3Bly/aCgMqaRAv2MDVbOd+RKL9Eo/p4NaiZ3tNlnFR/Becc66
ffp9k005PGYP1M3keQlZXWD9MLn07agCCg4SFgf47NoW5eckYLOCnQo457cZb696JhaS8Oiijz+J
SzZs26dILJgxxFRK+tVuOlKn3Ct6BGdukwGyhbTwLCC0xSlaRCF0FhmCytmEFQFzLcn6/FsKQIE1
T1Dk9TQBNtyhsPII303a2ZFN39xvFlauhXQRYD+tce2lcZ9CMik49/9vLZ6TNSY9tVFea1bWoQ2g
K+qE3SbcUrhxVhewYwpovJkRTadTEaFMUpxFJFnNlZZPN+D+XDwKxSs1rTPiMO+ONfFd6NEcij/j
f/GYopADLuWGNXwjafHBHgt8sfJpRiLIQTK55LATbekaqNEVrydeSJ6KUOlEibN7Xe/bxxcDoZbv
Cac/wTbnitMEfgakEsUdWu/FvxRR63OPh/CEpG/9I9Wo0YSJH4kx+kg5pTLVQZqFLvHaW+tnWtub
UY6jyJ6wYwu0/lKW/9BE3h+i+C5jPvzEu1Sx90V/VMCLF1+AdIxyFnIJG/kg6xnZ04JGi3YAfji2
7dwAMPX73ABDkFpK+BOkDE8MkfN5t9lmBOwTjyAbh7O/JXf4HWWfm2ONrt4znxPXJAaR4OW4eT+Z
DXB9XBx5lQ3mpNBj6/eQUWMIzyo8KgXvBrnV8VkV5ym2A/Kt8IN+jFsB708b9Vgx5rJMmgXAXqHp
1Q36+VyCdR/c1zhZA3t2FRItKANgFVaje4S2e4h0toLo3sdNVkxVrxR8babke7yJ0dhLfNVE0OYT
2Mts23XInmzzsZcLtBCFGBn+qqepkDaixWnDEbROQ5INnZcIxCBnxI9eA7lMy13bLY2B0SDY1xQD
rFaC2BrE2Mrbi925qqqdnYL5R6odqdL4Q7vFpESQcOaozmdT+TcXpv1A1+LQvSE0O7eGHVppEihz
3fzSamM6l0D75nIfsL/UnlyHUR3S2zBOTMYyjAGDIc8a5aIvhPLlrCP5DgSpnUqd0vcK46X3qAW2
v7HQhhv1C/XnWIy9MLwgGQV2Qd8pXz6Ou9MrcGQpR53HdSXPscyB8LpJ4nuZ9ozS/koMMkgogAhT
2SqlS2a9ymLszc1anhFx4fQKQWRckXo9NKcn1lL5Qby+00MAntrOnwWsDQcM9guIzep2E6RNyCGx
+9BdZASUxxVrk9zRGPrj9UOFhqDd2/3QuSLi5SFezwJefUChQR4HGdxihGuYV6aghOyFlOLkiTne
ShLQeKkGzb4p5kuFw3fSVckdPsIejEXL4e/MTom7WhJJOC9UXAM6e79laHmuqry4aN0qh+Xw9HPm
BcrSPx72nZO92nM+aj1EemDHRf2cDAs87ZgCXdbet2msNwy64QDWrLfb6v6PN1tx/BxHMbvScSlG
T7Wg2zOEXo2ODIq3wcM/3TuZm9dPRJBzh+ra91Zk3iaOslL6ttfD6ZjPRqblziTQZ5Ogo10wOmbi
1EDlcgO3KuXmwtw9M7yI2StVuQyC+sNfYURhKGbnXN/mOnX032AQImV8waBH9DLGR+XKXxvSoxhJ
VuIBEVvTUqRVQflNbKitBRh6bOVc+GqmbxLrydxJQei2cftzb7L72oqITOUYcL3w5Rm0U+saMV9S
zecU7P+POjTtOR6HsqVBiqE9gmgPdy3qDu8EwmncBtvmXAm0IJn+4NOrSu3nhPHXyqxGsM+/HU4e
g2b4UEra5Jjo/2IbKFqnfCXpY91zQUQrFnUpj3Ry7eXGCR5WGo/E5js3i/zchcs20I27LthHc+8H
yIkGcT1LbJxLtUapkCo7KTSS2LUm1eDa/VZqzDRUXN2EuM1Cm0FH2y5kUh2P0rc7tGOloWrLFjCu
VCossP4YEPQx68SaLPBYnLNPEq/WqHcRLTGbP+TAoCw0VRp4xw3VWJ1Vy5M2LCSTCwhygyLzAUOl
RXC1xg7/hHpZvHPCS4XcuHj0FD7gqKaVSyzxFxgpCu4VYzOwUbz+24HAImqS6GuB2jzjUEAsLUZB
49Ar4uUTDcoOiYy4VBYcc+Oydzqe5G4DXByQyaGxljpoWTaYANjt2aJCWPPedQIX5rgL1C1EFS7o
2okNmZF8+w20pgIcTjgs1OdFmRanrYpVV16poVcpZRnYW4bfdsNn2l1jlHY8f9uw4BuDYgRjsiIB
tXG1UhHTFKsTiT5E00Lom39qT2Y8t1AmZgZSjuLXCoqbqx3xmTS3t3gxl3T6/9YpJh6+mSQxf0DZ
OEQMRxFDu5KM8p4X4Ml8hjFsGDNHbI+wTOp3DNtv90wbdRnHP2qz5uV2wYUAZfKmUelQFl93I19B
S+epbAMxggpqAj9kXSzMEpzKvg9jCncGn4SQFbOmhUr0PsIgZwEuxB8HOwOe4zNMEVeGtDO0OtWj
TkfRzB3BU8Vg7fZl7aIE5ol5plW1O/Zf+8VDcIAjS4XPxu0ZytPXc68cVFU9/ZVhWOrmHHtsYRdZ
uGv77+jeA4hZOd34qoXLFjjMMjJSq5ppqBf8g+W2p8yCGfxJnBRmgotD5jIAj2g8JFzJATH6kb6L
jv6B/3QnszYrlWZ7U4XlokqUNKndbBzyIGReKA5bDJ59/9nmnH5/HQJiWnxXU4MLC29ZnIBUb5Ev
G/fcxXX6zYbUf8LibE8Xxc18Qg1mKy2xNdMQoGO9yA0LKuSCwlnBq9lrXCOSqXlt+o/11ApWq3YQ
D6w+iDeaa00kdAOS72jwiofx6C7ix5H/62T85S1V8o+aNld5LGQenqgzxYDrKiz+6nYVvYAUQ9t7
c/8brXElo+0htsEkfX+lazLl7X0qcNTDJb3GKrYTb+uVGmFAKAcWEgUlVKUwwaJfD83vToF8ectJ
DV1+cgURnC/pGgBeaAoxz6rR+gkUKrCQgw01w1z5Jk7vtyvPkptWrD9FM6Mf6z1s61iwqXQpfwXq
djBCpP7lO9gwLXOXoRJx+feDml2FmQF2btvGI6dvW4e13G0yOcTuEzVHjPdAsbLqI4Kge2jDegea
zu2dQncqb/IJOhMMKkuOztOcEjwqDw3iEJG+Vyy8WyIYHdpTQV9bljEMPY/tx4+7lcLYkPmLuJKX
Nck3W8VU5CUSLBnUJaykuCNofwQ9tt1jPQ6jHAEyhAmR1AdQHFYvq6wE0bRQtQRAyLTLa3E9vg6N
pyYiKORE+hjzaxHzZeYBs7N33w80/ni8nAG7+7rhTSMu56WiEG8UrUHu03WgftgjGtwUrrHiOhMW
UZidWEcL2kHEKYqJ1f3SCn6mIQnuTdkuTG0rUDjLWiBSKjNCX/N2AMQA4DlcYYfosh8euzrr7zru
bo6O1F5eQH/Ll244alCI3S3iRkS9qRXmApIydRHcfBrTbVA0Ee4Cc21UwdhviJthXWEWpOD8b8pX
Spgc12tnv0n39Us0gs7Pm+Gn0D69lsASF071UuLL51FMoFB5rD7kCYQyBhwnAuSmpVo2vQprQFHP
KcHrttNwn2U2DufLbzH8fJ0v1EQQXXrICk7zlUsOg9zkxtxICnvyKA08aSW9V0XSdYHhLMtBDgyf
/LR30Zvpvl/t5jM4CGE+bIV+A4HwJOv23Wls9w7kFHwgbZorwDHdwjzBfP+h6nWcijaLkcTWIBDr
TVpf6TlXOIqxrzTTUjTp5qA/bAeK/Pp6zVkxsbKptB5ws1cdVulBOIedIGsZiVgknQxokDHhGMaw
taweCMsCABNux1cPBB06hHdfDvfoUahZIEDVHKPa5s7A0Sgmpx/NbIA96loq/euHfkW90wfkUSA3
yNKJRSrfwZcL8GhC7NdqwQkKKaK7y9sqeAdVsXPkR+Q+h4w5SQvCFly5mjdrURvYKPTZji1CtA06
ZVcsKGvH36nQjv9iLCVvKkgDh6FIzSkSMIkzrHgAP1bFQAddZgfK+hoK7pVxOHFcNTywbBS1qUOo
tovYh5sCBoYVBfy+Ocy3NzTIlpWTMYOWYihU3pNY7AuIk14+HjyNo6FEmPSyu4NJBcMQrUVN5qcH
O5bqyJg5PTUwv2DlXVBexqKUSwfFmq7NSUuRX6FnHdXBONz5fcOkJ3J6wFNyPHAcnnFFY+dE0Cqx
+IbryLmKr0FdFlt3F43GKtM0JsQUX99Fj8GKyiZTfL7z+fF+I6Je8+kCylyH+icKf5e8T0UB6wfx
9mmcvVUqk/D2Zh4RaZrgqYc0dAg4KHB80abP6FbsI+acCZ+X+TUWAGEJs1QCEt3NTq72e81FuQyl
aGK/qf2ucRADblSyUzH42xzdaAPITWPV713AfqGRtEdkf04eN6YCCdyU1vrdZko84L9xlmiQmBfu
YNvmZlP5faH2N6A9Aev3LMpoY3s4yO4OwehTEzYU+34iviS7Qggz4cnraRH5fegKaeB98NW7xsFk
GCh0WPKgO8XLCkoq0sD3YPKmGJKeXbhVqCKzfoDmZrlkVvujlXpTQDDxV5ow1ovFTophKKugt62N
BSJEt69WRfyVw1GCe/0sPzXk3K5P86wuJXKUQv+LCWOslEin9ZD2NwoarlyyeqGdinGDVqaK4Z7F
Ca5Q60R6n8p30HrPZLJ+clOJf4EatLKP2DX1YnpvQ5zGTXJXvsTuoXFYFuwK43qC6+WFkzJ3NKGE
EnbzDVH7Z+nRi6ay+wJzktZoTQ/OEi2Mj9KZEXeV2jQvbdqRjy8lI0vEMFzccYIC/5HWg8bTj/9l
PXQGT3Sag2eUcnNGkEIYOtY9c0+9JSA+cSHt4CYRQ+X2IQY5rm+ryZDn+EePyGbUp73etV+jMnJ3
U/o7dmWTmYV420md7j1G7dufxLSB+hHVBVDa5iJlU206K3IPz0byGXcJfUt7SdpoJ+uk6wN7We9J
0koo2vH2tG7Cb3fJHEJp/XeeQ6MQjQTQfppluST41+SV0vzbWk5RF1TYjQyVGy0OhwkLKe0uJbNc
FqMuqS+JDSm+j1aUjTC35+tviF/gt2Tab/HhLSxfUCyvLKVSnEh+TomXK/EdqMqB6eBxQIzYZe07
sDdgkYf2PXkA10JL1aYTSyW2YrjjjyTi0/BOYiMTIMSOQDCYlBGvPnzkPHZiYlV0NjjVROcfF5UO
gA9Uh2qn4yKG5uNdlEicHBEpETl12jTd7HdUOUi+omLV2us92REM8DY3xpx2/02owZul9NjEcQm0
V7qu7Tnwq3Tp0UYmNTBZD27dJLT3SB9fOFEEecWbf9GSV8esQwZZ+rgZCrOXLGps6xnTco4HBj1J
XiDFdvq2zzGHlfXgCEilVEs4phLGUB+F/FPxGtlpxd66nBUhWY3WzyZB1REVNfUnvmdaHWzoDrrZ
5lrZK14BBhT3h/QjWfExPJr5FpB4Xn+MqVIrpKrc2fuEwnlC1cGrxx3MD7IgUlwv0I2zcWIdzzYN
SBrQHCSDNCOgWvk/URwfL3U2cshu0P1Pi0tvPbLQnz939LBzi0fOkQ79L49LOgSXmrhriD81my47
saDkk106pbTjdtfG1qCdixZfuVljQPjprTlDgWYsy495xhYRUdoUVpcBFYF4hThi0RvCy/Ry2lvk
hp1T8BNEYgLegge2w0jgTi7TJwqD9CTzL4cdhQxP8U6pE4MN4pUBDcXnMhqfheLh22AvRQvEH95Y
8nVzaIapHsKym6SECoT0mAdrtmhwJRfVbTo30dYcxpobE2ZcAPd86MxQd/xKrbbWxvbLwFApU3o0
ReuM/Vy4S7tym/CW3lZkw9bfUoLFlacrucITil+EsuA1zat4So+mTNp8Imc9jhhU9BJzbzQ2I7GB
zOepROxf2rbSkSCdTV/gVOahjE35aAGDfiDKt5KOuzvWKGEloaGj7eNzWrrOwhHQ4yfcXNgU7iK3
1laOkz3oHXd4O4oDnue5QqjNPDmLm+Dr04d1VbhKzirkCeW2Uf2LYtSPJQvgTX4qYOiKts6EZmoz
b7alHv6zehSGaq3jgAAid6sdOVAaJGpfiflBWapfuyAaU3MsJiGhs6ij2inKtUpEjDVsn4V/nojE
eB900PqYSGGZ7NR37DEvVrDVfdpZ9ONGysZLK46nYLqFsO5FQ/n5vw+3UitYwCzPytLb1VS0sXhE
913A065LE0fqJt4ASPyabXWQDBSOhQdZxr81Y/ljUdgACo6V7Izwck09Fhqq7W3oEyQCy534m7Dc
L+rSNPvkxKl/V+ZLtXEgA4Dg4IUoEXjMmQBg4sINeBycJAfEUJMY0sP8sAj27EKUZ7QNg77mCl8T
iasntHQIc6P8/wWZZr+wZWfpVuxlpfJ2vFHIGA1nktP5wEp+oGICvlDdTtsG5ce+BVbxDYKoTtUd
5yPh+uJXt4Xm5sEtF0iXvY08vhwGpUNuuVnwxMfsPvEFbH5WJ+WGEUkoJUo/cYZA73erT/vhZBdM
IkWixrtNGLF/KupolFhoiXKcOLXWHRk6sNAKGrAXLnmf2DIw4eO0oQEXiSYMPU4hpuntO3ksgcmS
iUzzH6U0rNhJHC0d6cW5tRbeBjeo7EICA4xcMToVT7H0wM8IUb/LL/Hz/wrR9ApzroL/2amUmNDj
xXxItRBa19OGX+V1trtjX+6b8+stUFI+J9MS+KB4HIH57r6m2CTDTA8XzYmuPdz2x6PCxjGYivdX
4cAUUFMGu2X3UCuQ83Pc/VI/CQLrL1JYyuXCqcEHh/5NhY/zj7hpiQel4HF9EHYxvLMYPUCBGmQ0
SEXYNMsaWI/SI7AtyeDYt4CKeNj369qynyGfdHlKy6OQjR8sWIA8oHqXBhZV1DKATfq/7o96YT6R
CqDfAOwyuZkiMCZOrPfQym58XDV+fJKsfaEfT/TAriyTSkO6qg9hc4vQVXDsEbkDIADDkUHMwXeP
UZhGasJZm5NfMqYQ/xBlQHqTLIaWqHh1Bq2DBGG7WYrXRqPYh3qoUhI+cY3yI8Eo/9wfBkznQSfN
sL2EaFaWs5YwDsuKlpR5N8lMTYxZ83CczM5b+KPCssn5gRH/Ur0sHF35HHvqZXGedmB04EARRQju
DiQOExfmLPDyfuKxrB0Gzb1lYV55+oMWnalRq2edxZYasrWjKvqyezlvtm4QZx8wfEPlPlB4gYGT
ceAab+Wg14vZdwzQ0EtoHPykQHy9HwzZ7P0cvI7WJNIdDh8I153gygDsZWcB+2Da6KnZKpqWRe3k
Bvet7hMtVSeLEd8G76xz9//DBtRDPDxx78kg6U8UCErPjcOhvtCd72/N/DTfLI6z2Wa9VfjQosxX
GCjFHDLVFi1O4W0fpc7Nq0D24BpkzjkXwBLH2yUbwH5E6ACPKQ2obHBvUvNDUqh53mBeHqJCK+kA
bxrs9/HQ4msU97OFhnZI+ymo+ut69Rf63j2bdv+BePKjXq4HhxL2c64fYI4E8M445nddN+u4/bO6
MhdHyzoVDDDvKe1q/OOPERswMTJhB83tq7u10WP0Gh78Q6xsftCaIqg0hF7uvgWS1YScTh3RRXpZ
pwiXKhT/NhyP28natr+vwHdnoss6mUm/bUjIkU/74pMph7c7V+dqRVafVCori7ViA85LamHJvXbT
hE3nh1yvP4V+zVBciSwsqcui9ZRYyTNmUXoVlvjZioX2TslbNMA77A4SS3G1q5/LLgT8TGYh4bko
AZhgeZw/S1Kc8Dtom8pNL+eIriZ6K6dI2hIuJqziIP5GWoWP8qHgkCtTDKrIbZ8yZqCU1g+jWq18
zrEbJ+Xg6c4dwCYkvW7wB8ABSW0di0eHM12Ed1pHWeABDcgbG8zJbyt/nOL/UeUJqCBJXvPsmIvQ
+Q3+VTUt+eKEovtB9FFADIu1Lkylmm+fiqB5SUDG0wcTQ/17CGibAbdBT2NjHStcJsfFlFnPV6H0
PvoCs4ywLGqnXuME/hV9PSa8Mk3+I6qecORrMsi/KuKdPtWPPPzyRtA1zKXWafYIFfXgJOIL5iVL
wlsml3abgEDy9S5OGMG2Lt3PaKv+ck4ROAEtPan/BP9FFAoY+FjrTKVqlPIpN4rjJjOtnc1hTguw
tmFBw8URqzrPO9lgADlEvPEBpjwnkP8iWWcWWRyEGwaz8aeND79GT14o5m+MKDpmlOi7FEfc3Kqg
j/mP8xJELkcY+DMdHhYFrkmNdWVxWYuFyGgmimRt8YX1UewHWKOABMc/F986XRQKkhAujZsKFhDJ
/nXF8PP4fyHOrP/ZDxc/1afmhBQVZ4fOvtw2MThfBhObZ0AFFU23KnWP8bCE+YXko+NVqL40Vzts
SHUb3N9npUCTsLBeSyOtYAQ8rnMnaFDq7cx8eARW/qEonAAoH3TMTrikixhsp7BT70ikKrUTl1Ga
0j2H6QZUVQfAG9kJUrZwt70rF2QEZ5ZEAGulzWRcxv8vDXa1rCj39VBb3pRav928RJvvsgAjKbKf
t6Xi/ghC61Al/3ZEhjP+LQb5yQ3sP2tq4cEhAJ790jFPm8uc3C8d+MbRLyTb7AqvyxrXPEZBEEBb
hrsLycPuE0jkC82rP7+udZ8JXvtKDEaFhmap/KEvOWdOU9SRjvdskyzmKGqBVq3vSFo2rkfkG3VD
2MXHP6s3s490iT6A2YkfUArhdJWLTJbYfzupjlAGhJrHvHlzsfgxnWqAtlI5JIfI6OS0G8dPCSvs
DNbo6qEbhLgoy5CJLez6A4okD93k4RBWWiooGSaEpR8tSgdsIQKY0nX4N2MzNSPkATGi7wwlMffv
eThnfxpY8baMmL28iSIMrF0T/tTYYn7avaMV0vNQomibvPXgz6AjimaI1210ChQtIHA/NVE1ds/D
fvHgg0epvqbANfznMD957nm2XJ4zJxKbBNtdqvH5NZYGBJj3Amv1Uk3wuBHFrP/uBeC/wXWoEOCM
jhb2pkfZzqQWvRBNzM33oBuL0tHhTsa7S3wPagWJRXvTCBCfuAcHr2yXQh2wILGDuVTcH8vTLdSt
JADJB3okq2k4yeZBr8cM9MAwhUwgxlnuXEJYdz8liS+ko1uIJJMRta0j+42mHptZ5sT2iTnAdw/I
10C71enJ8cO7ntZRP6B1g3zbT+Vk/X3E6TjV3CDDnhps0EoZIhrDON54Fzqqbb4YH6xIOIcEU8LR
83wDasPUryWJmTznUR092r6cf6m+uky237S9ts5k4OFWEGpKHCooLQk5br06Zt/aJCGYAjWqt+uQ
/mq9SgbYNlsbmS0UebLyqpAP6NyZuUUgvQBN9ktI2XVXnWJktHFFT22i9BbfTPb0h1gP5qrrjPLV
kQrqPpM04M1fW8m98qBBOPaMk0dnyBE4SWZF798NvJvDYca9RqK718mz6tXUKfs9muWQfSYdOCl8
EahElZ5yI9o4PUUxq2KU5Q4F3liRFHOTMn5kSBuL+lpoOzHcNamLnfEI9zXqkdCqDOOW77X3rn1L
KV7V+vMELjF4PdPrCq81KqOXbpl+EYmWc/TVO4fy9Yz2brVZ/yX3QO2fhSqsqQtQzYLlcNm7VQyf
28LctNgepcqGBV/lbMphIVqQKPJ3tdQOtnzDxtqaCTgvDpnRp3rrGnbrTxJyinpJA11Lwgr1CVOM
mnNZ2ufitK+QywOykpwO7tUWm7vPvcfxbClHQETeN713j9ttY7sy9h5a7dPjJ25Eh0kRuRY/+TrT
swvu9UN/1RJR8U95E1Y24xeDgXXIBicU/ed6IqAOEbdVbg9h+WBkTtACk87wgbFSgArHPYBczvZH
iEOypYdKprz4hqO8ao7HxVt2eiatQMc271EFxqauI2kH7t2YZMzUJiVJxoz5rCMnWyB7tUTbGtJe
kPdmv2S7dZOycnPhXe+JeFj0WCIGxhmyOUHm1vWTK7H4+Inqx7PpO+1URUj7iGVRxS2Go6fX2IIp
N1jalQxw4dPpdYaDFMfNUqjJuDUndlaJeFI4N4iEkLI9lSeQ/SYbeOhHgbtA/HknC1whOYVRbOja
R+9mEGN6ONsi9xxmtRNDcPzYeI/tV/ABdCEUaN4jhtltDWPuunHoy8eLEU72qHFm27E0yPG0pbH9
R/S2zL0KW9fZNkJaY4Uz0bDQRMoaXw00vD/4rlFGDKSpUh3G//lVXaaNMHtXsk9JbsKY8ZgfT01o
kcLKHNQEggB4oLp6I6xA2I2kLzma7SUJUvkOHyxcHk0O7hts0/k37v8gxbXkylyBWRoO6OQ3K/Ry
BOQfV/nP6YZrMi98f2F2JtJUvjRnflBfEbZNvX/LmKCAizQ2+LwdjgjkK+ByDHc73/qXnvXZpuGK
42Qg0G/Hn3k2nTw51xcrYRHugJ+32ymroo5MDV16ftCbS/9YS/MTWmM/WAoxwdLsueVD2dqitV5V
TQyB43GHsZ+J9MtZ5MCVn4GOvOe555ebv4hjFcRtwKAqUuJCPDjqAJXtBDiKiZOQpIWvGFyFfZa5
VuqVgFFq77rIXUBeBilFVHUntZywAwSbEd0yULUzDQafEPywDlfiSDPc7W5HAZA3Kom4mnDtnvZf
BIim1SbghZpWAdt4E//1oPuHBXwoiICIPwpiLK0/sKb9eJ1L50gKBpoOeLYsHDGrJmfnvkcgO0d2
okH7UktcnmRLXgNYNrwitsO6DvarCmEkCKRDSlKg+rIfS82TaOUqpXk8JTRYiiAq0ToNsXNhoJmG
80KM6zeRekzkGEqB9pwif4IiP9nG1DUHIsR3M2aBEgk8dxRZ2lmga+TjcY0hXM+4vKyy3gmK/Jxp
2gv/xDGV7Hb/MpB8drdJX4xVaBK7L9tUXMGL1jS1EXkrSBoe8V3aNADefZEu7IafQ/p3oA8G8zMX
F0UMayrajVcj+jtupRmlGZU0ItgAbcz+LQJkAhXJUVxeM61J5LdWFeMvyhv24RYJDvhJ3a5G9JJM
Q9yVAT0cZx/hjmhurRxZWEpTnY7d3iyPANSCbqRbCRnHe8KfgEWnLnAVgTah8UF7OmK82hVObdjK
97YLYlmOfmtd0WT681pffzKZxQmO/CHWLrTOGB5R0cgwC045RX1GwQFUCvHLRHp6CVAHdUoGhBY5
VrCaSDMZcZKZDvvyZssQNUOcirS5h0LItwwDlZY1tpgzJxoAIfDTaAIsAyZZMYaDcGKxDRQfcfUY
s+axWLmP/l6YvvuXSm9NiwS03pwjkg6DhEVk2j5wsRzqPCPts/SJrpztGQQGQGkgtQDOjCR//dvF
yxU/+LCQrXGttNf681FfftKZEG3ncD18BaFFYhFs5Oy57uqLl8i3hh36CVO0Rjec8Ax0ZuSa51eV
mNptaxlB9qbQkP9RTpUwD+nMf3xTW9OCdwIOMD4DBhjDyAT8bESDv4TFHhRTUM9oASHm0OgJL4wg
lv91oSyaN2bOKj32Y6kxq2OOdV2TY8sLHx1hgXVT4FYCeZd0Z2EPE3BpRMNwFBofZeLaNd3YE2/g
SdEA0gvJmjc0ZUXquQBjLaXUqWDQ1yXzccqgUKiDCfROVOunI9qv5H16IfWJhgXpulzPqdOLeFu1
eWSAA2lHbQA1QVoDZDz5oaUN0rdu/9/66e2hmKx0sVWc2SHaFB8Ecq8a+Dp15GsWF+nsCOPGehVQ
mQ0CWfc6YdOw/mCiA5cnLGgMEWQqE98zNyYnXp69lIblskjkEpMfgiXOToXD5rOZkGKL8z1QezsR
iqGWiegqH47Co25KRqA3WzWLKeg5PEDyYp20Bxd/2JYECfZOYpW6sBSOtAuEqqUfHHAC0CtzkLxP
s/ojatHWouiv2X0MT0nL4kGMWHQ43z0+qHr2FiCmTAGqcRu62MRfSGSzBl7wlhgkG3ZWa3FW5rSN
d5ICCl+amA8U20n8q1TMzBPNzNG9UlhxNOR6MrpGOFNCNrPV8tf4+ypYRxvGWhVaieb/kOgvikdZ
3yYyqUg5x55/UHnvDxwyuGkmdYXUli0O2D899v7A3cxfR8mXB6kUQlYFNXUs9ibpnvlh8AmjnejL
oZDMHyOcGrfQHdexNztf3L/coGR2lZQeM3vSfcW0kpAyqSrfcfHhuks7Q2Y/bSq4tA5knXNmdPM6
qJwGu6VKrp/FbdBnDOMNTVFJzb5EeugzSJfOc458vwT7OA5+QmYwSasrCFfxrAH0lDFRtzSt99Fd
oJ1K+hai+aRYMozw+Au6uKnZSU6HU+rFommhiZndqoXubT5vK0QYKr70fq4Gg5qIT8XtFtt4xo+Y
FhUtpZqn8uiF2wYJb1ErzhmbF2ejtKHPy+UFXmGQga7oJ6POeRoQg+JBJr+WxzQljSboGXhsgTMD
3rncIoMA40zgzDkK6I0CSz5eTmXIGyd/MfpCZFTMViR/TYZFsh75TUZnnko6fIrALiGvdq8x2Zz8
2ZFxf/ihnjvJUB6abeer/WUEyTFpPJwt/39MAVfPvzbm/zSEGBkwL86QZwg2PoZ+ZcOnOnD2dTQx
75Z9cNYB0IlS3FAprkIL+VdZh35rMojwmcwN0CUnvmUnFiN789n/uUynDrVzedqSpxaThfmhPHK6
f5uHfkwDIJX0XEpg2nVv7EnFXbj8ug2KmL8UjpY9LsAYr2Utcw24CD20/LKrfbS1DFmILSnwqgqV
Ao7qNYAsfwn1W6Q+XHbfg0ytpY8FL9MqUs8W99a5VPw9gkGXAOkKU94ihLHSPWEpge+O9bTiR3Df
1zT6PpQGJl/ZLd13VsuwfZjaogCVtAW1zDU9JxgrDIfTPVX6N5jrXnhSWvBHlUA+V9XzcZP7kz76
FqnjztaPorlixMklAVVfQUOeUiOGBNplN9G2+6+ndMbLRZx/AOO/55TcoPdhTU5o7scpFJ1d+mqj
zqlLTb40f+bWNHWqbPgatYUS5tJTYIxjjqdDRRK+GJOVObYo63b3XHm8u8bz37RIhr+somXA8hYR
jDpR548aaCc7IS2jwKPIH8eHPSUkejQFDiKgSPNzDDer/snn9jH452dicZQiz4gDqfKYbyr21isI
Y5OzkLlTD29huObpPXmikKBdIgcl8VFXZruIP38y0aKUGVk+5Y8LloLzdBpxdlYQmaeY1aXqVw2I
N2cXBs+NxznT9tEF+ckr8sRP/KctAIBdjcZ6ggTSO2arpJEUANne/QZyKzxs/221MMdJFUOYzY+3
A2GHWInhZIrY6S0LvHSElEAyFjmvmzxbRjRAa6zK4ch9bVdcxAiOK+ZzOmutc4rBw42FhRGZrWd4
t5XOa+9tG+DqHNE2XLBEyY4qN7EE4fhPSQ2SXwmaj3V144/r7RqIOzFnsFiMrhdXnL2So4t/166l
wFpM3xtlT/kyqFxhSVg/tN+hoSksO3DqcOwKUh7JxcH5HXlqRyYYR/Pvu9yiOrsPrr6+cMZRbcea
IHP+88LcGc+biZ8uNh1UTKhbnfL22fP4RdQBO9ONr0FwMQRThQpd/DPXN6fM4Ew4BpjtorqPGv0D
mh0cPdoJEQpPJlgLtcz2LagfIGxs04sFOJcDAByGX0zL4kI28N/Q2vAomwA7ElN9oYq+Tgtn1wRt
4sUeQJ9vVXJA45t+ZQmXKh3anvG/8dEN9YuTSMerq5FLFKSK11Uqjiu806svUEJQM9StuAYn9zBt
N+oGCABmJFTwgEld/8doRmHzPGw2NW15/tfeCLv5+wNm8vT4KIiKOqQVqAhvyrNwJReDyeglH/kd
uJlQfazngGBxEJ8Mxww6279vVzjYnOXua7plIEHmzltN7ATByGyimZ2nFTAiIP3tiluUkbX2fk32
cbZ+aAy/UdRKvCRtcuS7LAXP+R5a2Oc48eNYn3JINRbKWsQ6IDXt3HvjLs9c0GvlwS4JPkt3/VcN
5MunlbjXaQPTE5uGDtxXH1yR/NMFbg0XohgjQPPIXumkFvWrQLIdjKL6REqeUPSA0rgR/eH0Bw1q
J/ESkm3ZOL2HDzdtplo8HykK1YQ+MI7SD4HGHl//HEmbbgYB5vr5efMQCVmS7ExKQVai4aHZFDYa
EXZQUlJJv0M0/e5C89Tp43tExIl6hTsVCFxF6dZ/F9BwVxY6/jq9xQ/69Ibm45j0BYoL8cW9L9VN
mHj0WLv71qmlmfvfNsKWpD8GvR8rDBM4yDAz/uV/b9EVGyu4qB4a5qA39X9lGhjgc/UrDNy0XUI4
qQG7duSr0nikSnSPsQQBBvu81e3JdRL0XIAbnUWBQCL7Yv3ASi4IQpyqzCNUUBnscMTuNZwF/07S
NN6SIJLecMbpM4EuQp3YQkuJewNcQcYBDnS7JFxAEOdtGjF9cAADZb0tYItc7pd+O5JODbefCtGI
l002j14AAcKZykor3EhAj9RNGTHOVlM4fHlfAF6sBVyoGgXrLr4EZlFUqPL7y9y8NXZJYCF9zUiL
AvxGTxCphaLTVQ2D8e/TPZw3gn1d/y9G46Y86BmxN0VBczY+iGBN8lk9lOm3jCmV2hF4vCWh/cGy
ZKEVXm6YLhvnYWNf/RUWqKOPGfRvY7HA9jny7fo8VtlNsASPjGQpLXAfKY6/hQg9E+4UdnjjczuO
2DWNvfo/cG/jNl2egzbZQT7pM8ndl7Q/6iFAR3Em+yu8rSzJw5XZITRlA3Mzb9/kmkw1VvDl7GgI
8szJWisXvp/QHxLnETd+oMjYlg9HmzXbttcqvon+M0rEZ49+8NEx75QKbDrJHTcirll996UmEjMc
bMIp1tgi8qQWuESdiEOO7V4jzoMMPHQiKtqYaTm044uucngalE6rZ5QyVjeooUl5Xz6H/6vPB+2t
OwfRfXpKWsSmyRUVzwcmocIAJocHKCTVPdcMVnWXgG2qMADP8MCpWZykOSdtrLcJthwYwS3RxyKd
1SrujWxvqLdhqMBDN4AUZwttsYaDITwiEPpyU1X8jHpckHuRPcYpDrp5w0mfZ4Kj1BA6lOwhpqKh
V3ObuZyv4k83jMR11J6EKMWhZA1lq2BN3FeIR2qPZ6nQEHq3Q2b0mHX1zg0SZc50+v9wXYpaZO2t
pL/AcjxOaKWS54iwjL/xXmJBDkvze2lb8wS4Pe6ed4pkDKjz+TnuQaNUgAIe9EIgr8mMCi41u5Ml
eslTDqbUB6bwbsHrlnxjbgQPIGbHGj9jzkob2rohAKhUol9nCusvhQwwWtj+R3ayGq7VDH3WYSYL
ERFuzRB+3OvklA29LSp/aVmYV7k//xpHeoA2Tebznr/cuTHkMnH2x040FlT+zEdx7xqw0qcZWYqM
WKF4Fs6NzEzPgaSLAk26NuUuP3v9rhKvpTnx22mAHWqB/dy9b4GvbBCWdNn1NBvGkIdHBPb8R/pM
kTQouhtfuEcFgIQcY4YSr8fOASE987xkzBywY5ClU6xfGETjGUDdohQKoRQv3Ojc7NGJTJHAF6j9
sS5kTo39FOjb1OWj4WKwiwmpdBGSU9YH5kJq7B5nkhNE10eyeeEfYoyB9GVX9hd4zbn7oq5/qgfB
FtmZpdoWMooAsSmQxhnGmp/n4kOX7njHnvPVek837B1bFN8u48Q4cy1erhR6WT3RAsUSN453yDcg
uzcrxetP86gOykSIOmhZ7OOGfMWRCNy50GjiOcimvFp/+LAt0nucgjtfs09U68LqYEDRJuuSJ7sQ
ikqCOOk9qdEMGGOVeK5poJyFCDLV2LO7TokdTSw4IexiZsnT6CQjKduxxlYt9YBj7caK1/Ynw14N
UC+peybL+1K6zzR2pZTtCOp4Hu21whO+yMBXI2eyACs7BkQmkdZJ6zL6fJsMe9mcaqNjQJYXm6+a
RHNdDG9UqFjYlFFL7gbBkCk6+YU1Lwj0yUApsySYcm7zRMqLVuASk36Cw97IEkMh7uz/mdkeKxPX
uTnwQTnb4EIw6Jw9VRK1D8fW3qJSeGuq3zWrDSTprtHbLUTl8Z/i4sql1E+EejyVuG8MXXsM9san
lE49zhV64IoxUXGoN4bOPQq2RpnLoWL3MbpwUFk2Gck87p6rVgMehYPfkjZk6dGZAma6dqRBf3tW
IcgCOei8fbvBq7zt+FMJZZJHIU533K1ZgHjB+wrUYwe4JfwTTXEO17nJ7woJAm6vjWs0ubm+wHZA
lahDzTDYpww/dkpR9wKDlUcnhfaZaqYlDL2gl7xgTVmY5Fe8T3GbL7Tu3IUq3F5CGLCA7QwmwqXP
93elhcS9Y4XgOWv/Xp3mhCXXZ8wUdcddmDfE5FfN8518nnhU+iPrelBGhUMYp9WA7oOgjcsPrWO0
iNQ/h8cppKtfBXCariIJlbZso5+Z8h8CtxVfA/r09R7Dcu3/o9546jXMQ3Jf7sb6YUI48UeahQKz
6y4TjZm8pteS4vhbsOeVcq6eAU5GXTN6ymdLa2LMF1fyeto6enFlGR9D7QE0OzcSdEb6MfyldsOC
2UTHP75dUuNpM4mUBBJPYSzhLNCMfbYAejWzUFg/J7+TA3DXkqALGtBM1OxY2XTILM495DSjgW0E
y/37AwEeDAqEwQvSYZb0bJ3Ha1NRY9WSAo0uLIe9+zBzsgD0nkJJRm0dEdWOin4YdhXWv+mdCrtw
cifro2RwwdfoYbiAugMIeApvd7y9EOyqNBfcMhg4yrGqBKyWMQa2PaXgOsQc/cTU+E+hXi+8DuhJ
5o7nNI7OA99tJDbb5q0PcekCpY4GNnQVDFv1SWHzwu7oOlvp45C9HhgtDuQukhmC2mdp/gLqQLGP
Fa8jr5UkpFXBj5FMdOB/4nRdRgC5DNQx7voke53XR8SRQKRgypji6I0WFOseoJhxD6p2y4EJV929
B6VPZxHeKdFgd1usfJ9HjlaPPuJrh3JiR2IeInYOrfCLY9/5rg9wZnJCAeSQxcB8fk3ZRaop2LmB
OEZV/1Y6ic3xTBnbo1E/7MgyHgTKdjZMkKgseXBOYZhzNox/hKLxSPCK2O3jaqM9Qvto8ICt7e63
QgjWwEgdv9UbdCuzqAv1016qkdwKnDjI9mzP6oLHBKknG4hzmTIS2ecLa1ex5VdLWakdFK4DYUSR
Pg/MU4sKH4twCYUPrpPY0E4BWXIfRAxYQ4Nr8D3a1L478sLE86zCDqy3+Wis9Fm0hwLY0PRy+aQM
AoPlYjVrNCOeYXgCnUaeLCyXfhs3klYM837Ag0QGfnmQOhrz2TE+77fbXzFp+5KMARqsO05Gzuyu
7FMFBKQHadDHBosY9bF4Ln2KUceMunfUkkXqMPQzdz68l51n2u6lXlecYjzX9aDlhAAAqyqicqIW
pJEKOnc0jAsr5LsVXiSpD6ol1BDAXgmrrUBf3+1Auexmy7zGEpraYHixOkBejmDcZ/sDLLMryENJ
cQLyD6ZziRBqN0VsNx7OectaeUd7EQ8HqIXbK1I8CIyXveAkSfp7I0uZDvVlk+fIi+phvegdbyQ9
aXIekvuiQMUDR8fsNd8eXoir0/yh1Hke24pR3G+YRsfsc5a73lrdgJwhMxOy4NwqLyCkziaJYTKQ
T03j4OJYlCEN6yKAsekqIGEYmWYo3sQASecUqpUjwtYrWP/TtNrG1Iwp39sLuzYhMteglj/RCfgo
03hktmCHkqNb3HjpXfCuCsi6/SutsnZn5MoLqGWnoob5N6rjO9weTbgW0nwN48sywer5rblSXggB
Ea80KTuxyUsM7spCLyO36s/j5qjbLjathzr9GcESVJgI9055INUGkMPwn4uHoklhxct+i+abGY4t
xynDowMrADSURHWEYw8DxPJ6gxbkRCN7lMR7Ie382jwEzgKUzX4eJqS7vx9lyZF+Jqix4/VYZuMV
QrqGEmWi5igr8xvsPP5/KKCQ5HdUGUOMqoWu4cDEQhkPd5LcUsrA3l67axbbc4rG9FdmzsvaaM5z
4KecKhNS5F5vWqoG4ZGeOR6pXrTLcYix9oNukek6QjboUNWDAyGn+Lki5aWlNPUVcP3W2v2oHpXG
tJPdakmHQZpTC9GXfbBk0h7r9VsTX19oRDoJzhNDB1cwrOeOmRe8EhbjLvmZtyq/1pOwElebPbfF
uWJYETOz2dj83pVErd1mFFYfZgxyRyW/K05k8Jgr/cQLfIeLDH9ncLW2ANOokl2g9btjQ1bbmI0B
ye6MV2f5tRJ9rOATYg4nysk/NeK5XYGxLQqc3ZrBlV2KIsENnlQw63I21jA8J1utTiKznjBGJH9m
hJf/E8anJIaPdYWqkpwz9D0/kLE+4CBSP0S9q7Udd45i8A4TdhPIXO9tIVvsGOWaGPbPq0ufUCyl
+WrH7U0qS894pDXw+/kGLikU9Zu21Z1Aca2B3v2Q7OfzjgnrReGCmgsva8WQiP+JERH0Qa0H8lak
zo7cSULpUcdb4lDtTh04QJ2r6W4aclcwxai6HRvYX4BGTSymRqKvjeVl7z0fsecECm6dvT96PjEr
n5yIRVWXY7GHUk1v5+t7zB91AYjEg1PE/AifK0F+6iQLdC502UNf6YVu3v2Ty81d7TS18KCtV7PM
hJUBMKXEjecUXihLkE6HLSVIw4bmaAMEOgKPTCjJnwPOG+EIQGAFED8WJXwKr4wzrG9f3Loj8WmW
c1Khjw/b+WATXsf0D9PWaC7ek+pLd0jwnci5W4e7oXRdGza/Ny5F/ZqH96eS/k6aLaUHUEiKjCxC
wZZs/bsopbvSKVlCuOoG7oUaOksYVH1jYITIg5olD09o6hYMg8JWoPPkJvALsGPY4FC3IRb+F8Xf
DPjyBbWd2NsdBEeR/aFBXfQ9iHd9NCLWLiswYTQ97QvlJiQWOtkIXh3ppv04U12QQSYW5ldj2j9A
PaH5sgxc5U3vyDcTABmQtiQg4BlrMNA3yzDE7BUQ6XLjShNzI8vQE2rjf2SdA9oiwUNOC3ErJaYX
5+NpFU/Hn8MgmlSQ7pJCj1Pil2jdwr1DIJKZxN0dfn3fHV9k0DaqoRmNMF5PEmizMYKvcdzachfG
ODcXabGr1Kgc3RNUg2Nwr1FvKChbYngKcZjQf6tVZhEXYio2j1e2Wc08DorIiKL0cXYWF6Sc1P14
x+DpUr07KMol+zPW7GQvhfBZ5DAykulL6jduBDSiZnuJJMgtMbX3ne3Hu3cSUjOvNo9UDwdSlr+D
jQ+XrL0iW196+AHNMo5gMlv4piCUr9xk4AcAhITys1ws1zJ7XeZ9VvLJ2zGdGohF2u6J8b6Q5Sct
oU8OM9RoLPDkwGLOfPuYjP4cBNxJHVA0BUaMi31Y97FmxqL7ZSYcI6ArbsrKQ8WLxmSKR2POJjcs
/3Urn3JiBx+SAzJKJ5Oe2XSBXPRI39MJ+vnY9OKxJze+WPc1eutCFRxHrNzZb7ejjMWBlKSWYp7x
aBvWR7WUNqpJofT92zSGBsaIZXR48i/Te3A7V5D72/kuFXBrvkc6N1+GVq2Z8sJNu0Rz+F/6+4yH
wRJnwdZb7z8NmUujgE0aVyXBy6u0SLZhGwvtphTPNoE90pVactUQuqgcIY0fF8lh/uypO0X3+amV
eEpQcilh3urCzQOb0Cu6u09NyHVNwFGalZvlAa1ge0svKdYWNol4pKZrtuAX9vTtiaCvnmRSUULx
iYEqBjT83DrL9intx9P8zKbbjv9SE+cR2/zlGD1fwWkziluDOZKK2SmvWyjJ8OfzumMgKAiStM+E
RVtGb8IZo1YpJVX1jQA4o5/Njevjfwq57g1dy6PJ3QUCIPJyvKXLLyWS5xigtHP3ATWJmDTCPoUu
iajqDh/qLfV8+zUIq8XDlXuGP/o3Z7QYUiD7nE287gTK9j1RKUYrVilfVSSTCwi7IY2SZ/SfrSN7
t4PFwH6W/ldt9Sl1QYROIa5TnQ7R9uxUtgmi1T19mz00zg0BE5s/5SEjDFChpqgSeohN6Qdu5YEW
WWQ8llXrp2PpzcG4g5kis3V2wfpA2f7d6AQ7MngCMwdl2Mo0D0+jb+Yb4FRBWjwCmO2/na4WVZ/B
Pkg+NwcHgmua8rsIIv+9EIZbl2WXn78RWTEWSt0xJUiziaUIl762lYPN9lRerk5dMHzMVe66hnch
WXHtFExCkmDo4lgXjTtY0s9X+aOJKqZQueJu/GhW8ag8A9FgA0bOCqgHRjz7u2Ej2i7OVlq9tKYP
gEa+/QduZEbl0j0lo94tn3a+HS2HyyNSu6VF0r3hDV9ikwMwSSa3e/6iQs2B2/UQ3/6dwr7lVqES
ErwJAKa5vatPcyS9zZHMH1GneJGAnAMdVWMmdyikAsIhgrmiLKRvV4lcxCXVL15V4VlNluJIj9sV
L6RtsABtCUK9/dPuJ5otyDzxsTmxxJy6eWDtGLzCJ56XXvdNRVA2KBP3KA0DklOHLdOHRnq4Suo9
7MsVF2u9bViKr6xjScwuStSXVYCrwrnLERhZjvKUc5AmxEFnxUuRY22stoS6NYFDu0elIzKISXkw
3/v3ExcvBE6zx3JEmesHnO5pAR6ro5wM9+u5gqIWunl1jZ5jXZnnc42DDGy9WRc+N/ffyDVQJG4c
yX9mfMXEGb51CNOvCiWtZeKgtt7hk56Z1V9oC+UB8AJLSrombBfWq6JZSf52sdyHNZckRz2LbWzi
mRgOtQCqSwlbLcOGCRyRLNbJxSFM2TfxkeqAKZwCeMGTSf4i0Njwc+2uulCsYsdgio0CBmj1ZDyW
aeqDYSdS1GC5g15AChqmghfv5cbM253IOBRoP8hGlpVZmdKj6leoHzY0+qoGm73pxWKevp4ktB8f
1QpDxhJKwVa0vZCB133D+k7fWA8GrB5Uc0TNWlT+2QlYKFI+6qdn5SA2EqAAnlMBGAbFIIDWnKd+
6fpB+XGQhsiKG7Lq4Oq2kcDkRlP708FwCWVvL9dibYJl5NePmQ8zIhV6O+7RFa+VIVjQGu86ne4F
mTynoJHxehsZl1gbvbgylnGpPjitDwuWrR4wqoxzMC3mAsPI8wsaLE+8N1HU41+d7iHaaRP+4Agd
LbYLh0M5Jo33jJtAHBjt5KMcTz5CasZcdOz2smpm2sKfN8J67XcE0upiX96A8ra3KfMxKCk+N9ON
ol2qOV+iSvwbl4ZvLC38cvuoZ1Iopok/aNgzZwmwblk5StTTlc8H7S88I6jQR2XXVrH329lU/xXc
Ov2MEYrMNA/vXBH2st7gB+cSO4ffoORroFh0ZRREbobmIABghKO34H5ZvXNzU7R0QzIPEU9pf+hM
HqzKVGcnZSKHgtK83ewYqA5jmBXgNFg/P48pBF+ygWzW0bRM/tEobRKPmSqkRtn9/PyTSB8X8gTV
9uBqjWKPiyzTxt3C67V8NnQ4cuuRDPhFj6iXfUv2VMPIftLxcigoOYlYxHIMp2LSWo025sLRQZH9
z92dEYi9iLimzcr5O6FdPBCHHOcc8U/ibohwjSe7IHPoab0Ew5pBLl8LUR27gE3yqv76DaLer8H4
4rvSHJCR2WzWPkjW//vQye7vUFiw6xtHZovLFXTrvuk6TmM4i39tRt7Cz4TqHUBD4o5xIfq4zpf5
1B5aMTj3VrGbWOd8muu5rNOnV6ehT8jjtVcLmVniVyQe1k8qhdBW0aRdircYYLaOBGJzpel4h3eh
Kni0qNEpvrW2idPImppuNsJlXVu+PKIaPRekqOWZ/TdDPoOsBxKIHJdxRYbyeZXP9GOAItadZexP
l2or6YpeA7Gcd62esgSN81Mk+xD+wiiM6yeFwIG79BaTjNIT52R2HyIVP1phtazEr7pIP4BzptfR
dpV0DcjZsehS6TzXE7giHfK8OAAhyN78B0U+FIe7FXInWeE03hQXQxlk0Hm1876HCbN5sO14VtFP
ksIgcTIDQf9rQcYobGaHLEma6eUo/hEqys2XSV6abQICPlosOeP9DufamnZk+uB6eA1ovZeFM4tc
uPySeOM2BEIvJ7c4i8tlveHwitpHS2lNOA6cWjh3GQYibWpfYjlFF/dVqNLF+rTkngpF6Xajj2IK
ill9KwtjScfJ4n6NixVoaOXfmGrPpzcF7IP2yflg3tR/Q1uqf+RR7Y3zD/M1d1iqUZwhpj07lFxA
uu8gFdC6JXWi0XyYK67zwG4yrATfx60CMJZ0OUNv31C88ByNe6rbPYJcWEv2j6INWFQD7s5w5Pkz
l3ANIqg+BbTTYdd0E7NbSE3w3BM0roGBCwGexYoWDBHCh7UZeQZkaYup+Fmmt9793bgl+K7WGOhx
vD9x2qtuDFeDh5/m9sniueuXO/D5SI0NGkKzIxKXo2taDeTf/o2QLExRXnKJJwvDKGmjJk+6mZGR
IfzvRn6yIcALzyLF5t6EMo6kXD+z8lKhi93eZCl29OVNV+EYTM0/hELsOYv4CWryQ0BJszZkWqax
9TfsfINvQzPdTlhftjCR++TlowuRNytgjjuMARm/TggQ+7IAeDyNYtEjFt93K1UgkteIf5LLZIMa
OxnfwFMFxzDXnwxg+aJv2eUbo9lgNOlR6F0OVNwuhIvGG9pDY3nI+YctRrWFrOxQNzSfiA2LfquT
JexVqTYGYRKlZWvIfAbcrqmOlB6+WhOAVIDzCry/OTBbUVLdhDXQuWFGm9hBdhYGTJ7YTdb6xhVO
TnYAd89hsd+QpGBsMtvm+snGVpbyycNk5+7B/G+TFiD1c56VDN//3jgZvkboc6GRPTWtMlQtrpuZ
gDxYwVE6HtR4qyb8aszp9pTQrs3ch/P9CHlfTObBer28Fok1JvEh24LhNQtSutHS8r1UOYhDzPV6
X8Xfqm8oxIuWr1z+laVJscRCPLs5Dt5jnfwhROjGQVIDpMb/NwBWbPBKeW7ZfP6zSmpKvx8VGIwu
Gpz8hUPoKL4BO5C5OsgFAjXMal+hYDKvRLGg+HEYFHXf8uchAzP1h+2lLfy3CgytFvioorSnFCQW
AH/Q0TZ61gE51XO1dKGYdqaF3E3RBhRIzbZGiLlLxIAaIBY+6laXXC7+6UTv5v56sg4v0PAmm4xl
bS74gx2TgtkeTx+8PtCGEKmfp52y497N6ijUue+btbZXhzStwr69BHGFwWdk9Wyu1e8/OoBFPyJJ
eNsS8sEmssrkqSkFyUE3L8e3uvpCFACh9TZ8BQ3RMd73n4eVkls62Jo0yVZoVt/wKXioERyaldtK
H0WfkETXiXCF6mEcpoHnJM24vNZ/rYGn1btF7Vq6/FwgdVe8QzGhY/6g6kFF41vbHuUcRxrjV4yA
FFrvTxUMzy5eDzpL+x16cwsFKsnul9WpRxQxP6ecKX2F9438xPBSCoqp0nIigX02L44uO6+fsXvG
nivhPDJCInJpEteg/bXskV3eK5aWYyRcm9Qas6+gIS1LbngqgkPswb+pGS6wxcmBGpv2UoLAV54I
3DiRpoh+838QiT2HPve7n9dVTjeyjGvtlT1zm8qA6unRraOqvkvu9Au2zd/RV4+H6sEu6OfIWfWY
iOLCJSvmKex3YCaf5/fL96Q47w928txBd0plsC/SZSQ+AsCl5Hr1yvv310H6H/xhr/mhKm7pIUDx
I9HJ4ziwKifu5VMZBNOo3bJUl2B7LO3dxRmh3B32RzGMtEpLIIujEzm8R2I3cJ5vsiIAWJ1ax5FT
f5K/xDKrkvJ+lrMdkaLroh2U0iygxTbwIJgbt6cAgYc3SFvqPNfI4QEDovmV2mnWCuYmX5wdcUWf
jo7jCOOIyse4sEsQxVy81KVVUyYFuaLn4yzeBV8ACjFFPI1MYuOyD5yAzElwkvxJFaUrwFgsrzaO
W1nu9Ule00qUlT6UW4VwANC5PYHQ3XN5r9Jww7CZB442YoogK6nkwnXEKTlTMiP5IvAAQAWSN9Bv
1npc/bL3i3hRuEaY3JPbGT9Yn0rgv8KvEHJqKScMrSVKlNFLatEKZS3QuBkwevDxpYj2Y6PSH49L
Z9cp92iUffivEOC3Mz/faPCiU7b3T5qaXK43w8h3rIplZ7Qn3iKfvL+80ocmFKysJvrMdslCnztO
gYv27mrfYubko6/rCWzXprklFIv7uVguCcTRnsKZzy/QeGJ4YoKae7TXa7IkIJvOzNTxo0cen2iH
pmwn2umDm60OJjGp2MZ/fBMF2bgU1HMobvLtYICeF1QEm5kUw5iwiFmxidENtob/1DeJBZDbMYWj
hR5AzYo5ueWVk+kSxG67cChSSbCr6D3KGbJXot1TbI/nudJYQDWd1wqMsMFhw/dK9Nx4UHjqwJ4F
9Q+bd4hpDmjXR3D9uHrkKLH5Hw6ZffI9mrHwtQ3gdheCxTp0NzLm089/8WT9VRU4SKXziMfxqpYp
bsEOkhM7oY1+7XHhzRqN4YRrZCOTrBQASmo5zdiCwK0F5v/PcZOQqSednOJQI1qQAP5Ctf0jfdZv
kg0fkq0pjWQbXpwcAKntJR+ZcCXm86mFOe0fIA2pSaQSA/S/t3gvk0w/Qj2jlzuhz1XQhV60RURk
DL+jTdZFgoSvThc3hL8+zxLdlH4l9FgtVVhDXngdtuePhwZjwoWRWu7C7HJ0O0FzdHCChRLvFmEK
Dcemnxq+otoYvuX6f/LwgG7N68W1aukIK0PI/moOVxVAYibI88nuwJOpza+6VZirnOyidRKtOKec
ifOT8sPxAQ3+klJ0MU4F60osu2yfDCPH0AqH4c4odB+i7lWmQJf/kA3AnQNUsQZy4jX7Dy5JS8oR
GXp1DakOGN9rgqKlhmv8UjgqCvIKIp8BDz7pjggc7/raqvrVfs5MavwPCVuT9z8goOSCwnszJNot
sdVgiFWcsrLPIxjJ8FCw4yoNghDduE0ZAZ2Yq9V9TRgkwA+xy0CuJp0XdWtVpAS7Pkj3Z4DSPzug
WInHRzm3i3YD/XjePli0heg/to7YeDjHzzN8wBeZZw4ONIcjJj5DmISDvyJ/fkSb0jve5nIT758P
pNk4kTP1yGTrYcYmVB5vMJLsP7dwpIyqFKBG3W0JQewKKISn55zpU0KX8ESrtTn3WC6g0Rq2l/AX
vrN//owj2tjgHdDG/BblEWbRG4GHaNhFjH2gqfgSq9qAQHHdrlO3MM+Tg6leXiiWIO4l5YOGNRtQ
cSpqK8LDTxxBcGLcU1POKtvdiyiB+bEowhIfOuveewvSpRgG/F9exVpfVH1yofViDkQwKTjwVXNs
BoIHFrqK2i7di8sH6Euy9+O3vLrLdb40/zx6nHHUrK8M7k+rohAEQ2W8C+kMlQrtMDpagZ+db5Mi
AUx/Yjm4I56TN/qyiS/HI4I9ccnnrD94Uz1jR9GTWhLKOKWhXwUzyUNu63+gCUu2F/in+jNbhGtf
jf0HKk30QrW0m7v8r8NV8BWIOlDgv8/tpVke7PfBELuMehuHxlSV/VFdNWOWPgex5cTHgzHK9p5u
5RVPQr3NMtyAiNhOtGJgHsRRM8hS700fAXZfA1Dd0aRAxEbyOrjdR/VyBqxDTyMURqSX7SQeM5R+
d8hoBTCbDCRNYFEQqrk+qhsePke+ddLvh9NXnFlCwX9q0xRC13/cT+SMF/6FrS6GHzQICZQimkM2
gZXC9Oe6+ouAIhVLJRzkLG4PNnzQKtSfWaiXQXQCg4+eFxHQgLzX7nfFm2u5Q7OU6M/C+OkxZKVx
x1RoOt15I/DCPxAFJWpUUYL44fbu2jxmhHFuwz26KK12uD/PAlRyQVuMv5ZJ6ZMzhJlpILdJHsIh
zqiHm/D0mNylboBYf3Dd0V3pdHeAPOB9b2yHV6bJHwR37mfslHMC15h8ULFJdEsJXbt1J0l1geuR
eAqti0uWnDnK6/61eRHGYZ1oWJcSJzUBOh9cECgekvPHTvyWi/3KoDptI7W2HF5wrK+HPcMMfZV/
kGKoIfoulWFYTPQuc1E7KcDw5cZY21Gs9deKyvbSAHv+ya8nlrgWThzmtQM+cryXoja8MJ+OpjsK
SQjGxAX6bxqFI1b/JUPXfShegyVinak+PduzioI7ood/M4tKTID9Ob7fKnccEXwVqASS7zCTczCc
A+vtZITpYuXJ2z+WyaJO0ee90sp4sIMnLJlqO5lZ8qwE9twi62ZG8hF1fD1Aqx2lWBCFIVQgqeNP
Ct18EgzVgcgAtPXFU3SowKMEyCkcuRHDeyH4spTjJ2dn4/6I1LvZUNCEPSsgvqJIcLICAlLTS6Ep
nblPq7EOyTVphuuh1bkgLuMHACAFpeODaEkT+u7ZjvsWlhPalBtK8jpIu8k04BzU6gkWn5rpFx69
N/djWJnsfkHV08Gi5NkqZhDAJZwKFh+rVzLwh41f132iiKD9nz65psImFVb5JGvZFHzORHgtTv2u
raMGYQHDwMuJUy5fyWkwLazoMdjsNjJiPyVcb3CPfhAgEbo+Ssla3uf9hsVUN4G2gMpqDHg9tWrk
al1oB3vwNO7xyKx1yww6Zhdd8BP2esB7zkmdEddso8JQewz66SJKLo1S2I2o7jmGBi9oMqlk4hBL
rKVfG5OntT621Z1oYdlQboBQ7DYftsnWio1tITzODC7PXz6PRbd3q+RzWFBTJ3eUiP/sEHXFcY3+
TYLVXv5hSgiGSEJIrur3oUqd1bCOgszSuteqUP3TwGWQ6DaSCrSaPf0PhLFtx00aCFm5IOVCwuHB
wzsUbr1TWpKkH9pLY7N1MRTWlvmPNzzGhhB8IpeRzs/JXchrB5MxUOoIh0MiPIEmEwBb9pNAJP0v
1pA5Ux/u3NDlo3j0STtDTbWgH3xGbctLfteI0BTjFU7l4Uf56Xyz1rxN3VwFq4VZL/5owiIzL29p
x5uE6K7wSq0vNgqxCxyZkX9VRGA/BnAoPy1SbK8JTy0PPhg5L4mVxb+ZqdmEgqfvN4MMwOaNXxdN
hWXrlbUuqjpmpLGUvWvZYFm/75QwZVJ0j9ylXDC+1O6mYHPZthNPovSNDHDCkdAl9U7c+GTHT6qx
oKzCxL8KRRU5a8WxM9wBspCnnNIBskUeJia8OgpdpxebpmYTA1YPxsE1iDA34ihSD9PF9TPtjyiP
uDnVskTQ2jgcBHG3W5q5Qs7HKs42LN3AfuCv7AEL13SpFHthZSHAqi6mTr+CdrpjcdUf8YgWqTPM
spoZGtfdkGaZKr95ftsvxzNPHNocIdBOKZH2ok1RBXWutcL1qvtwwjw5xi99/DMR2X4/pAwi/69u
2CwmlolWm01W/u06DV252HYkQ4NxSioJVefbF0P4NHz56NdXgltbRqjq2W09D/sci+YO7k7gnYpP
wrBrFyaLJrTj/sMgdi2lEwinGnc3vlCZSl46KLfbBkU13biB7iG+9N32PRANv4bs4vCvUqw2sK9j
+X+wrpAgnESYHRnBBw2Lb/+hScuCSV4J4n8k0JpIGLHna/tjlj3ds46vTTo/vtPsd2VOmtOKN2z2
tgKK5Z1UuwwWaUKh4+2hphjWyW86QbmvzWzPuf++6azz5oEvZbA7KD9BaNV7KHHXzHrPQjv/LLKT
U2vQlJEBfyCqB8q+WtkcszC7YcaRIXHv0so8N7Jurkoj3w+kUmTmgwXZn0GPbi3DfFONfgUV8UDp
50w/VUvN0QboEjAzt69UI9KWioEK+0h9ZvnswiwoQEw3ogrIwi8mcFqmqOEYfREUkLztntq7FyP7
CZrPdT8fyDa2eW3LYicED8NdUzf2Rc8UjzDiV6aj3LGxhknVRnARgwIhcfoDfLFPp/nA7PZqDgTC
4fW1v6vf6F6gPHvgCpfrkjvwJfAmi72QA51t6AiWcIPmuUeflM1IhgWlsyAPKxwV0roRzYbYNSVl
yJs9m2jqc9coacE0u/jToTMEh6D1cVaizsU1tGexvGX7suAi+dOveke8ypjtsfygRmLxIvqvwAQl
cE/Zj1qhM573agu3I6GEtpTP5WT6OLdBd1KMx52gHTgaP4yEAjEneedpqcAy6DIj3k6/YkLQCmUi
4WmVpMh+jYd1UotfYJSWaoSg0blKwJXoZkLlT73JRPYpOWGIja5Nl8N3VKnZjd/EAqjpuLEx9OuY
UQmMe6Lq76AkzV7KrJOJe4Y3DDYmzrvDk8VxW9tcOcsEulrMvRr0lWbSpOXYeb9tBARbzUTyicbd
Tsl8WtduCHqPyfj7wJY9aFiOztFOt+KJmDlrZWwhjMyTV1/AgM1RyHMCWAIj/gP4Zaj0w6j6h5nn
z/VsRDeYi4Mb1AxfDmSjvY/17NhSYxuvLnD0q5WU2qXBkwmeZzKLbrcz7Lc4+vBRjdwVUWHcMy41
rW13pH0HqcsTpUTEjuIAfCpB2UHvdpXZNMMKqkDL7fWqmCVSLmIrfEUKq5KaJJeRmZHKYD9PAY36
wXyYJbXUuYavYqq07Q7r5mkqNdVTAuT5luMvUFRDBH+hDy0DZDQiaQpsMwJxu/ebzW5pk+g4P484
j+uEfzwXRXMhy5Eb40Kcy9z1tQGwLAK+hBoo9nRCH9yUsvSlW9W40Ev7LmbEn3W2dukpbtNSZqa8
BgsJO+dl01XNwWJX/LZsCzVxLYbD4RuPCvUe+Yi1xugW1M1tEIQYkREdu2BtG09SIeM5iAPSG/td
ximoU/3UOINVLX6186ijwOML/DYDUrGlmeyF15OQxvaYQ6C7GYoGBBOdxc0BNZomfgRMnBjIyJzN
HXngSN9joEBev6jp37DRglovKA0+BLQVhYkT/UV6jES96CcF/spi05CpKUnswCcav8fTIOa+EOm1
A44UerZLR0Nws+Wx9XGA0T4D9ybFNJPg/YUif1TZm5fG1Sq1u6IdziMNWT6tiMZkyV7pIHE4YexT
tCxstGnujK55G0luBWWRilB6g9pBQXJzP+5bFub9qHhPpXe6TkyjNA1/csiUSkrZyM0lN4P122n3
XN9AWgwQWFr1QSxMe9+76XRzGpKLYrrsF166GvHsodFYXKRuExF/u0MC9zLA6yW1rz1VquOgPaCK
q1VtL/+62gdbt/4IUSmUJ7BMMco022JfZVImAq0M3bHR7l47gfIiV2LgfvIcZBaw3V1gQuEofTgo
m4RsTL9GrNrmr7IRpo+1jr9uyDAZgLXVPpsbFPQ0U8AvGJL7V7jn/49avLsa7Zd/wjRAE3Ko2bBj
EOV6CqGhsMSkn3CXQi5Wlh+QtDh7mxIg+bVoa79bfwVi1Rb+kUFmlFW+MDqyEhtePpfyedEQkg7G
kJUXfmdkXXe884nv6bCpb3GonVFNKsWkO/g1U53k/jGHcMftsqlheZ4ij0hwjdTDPVkIzsn7VLDV
yDxeyOGfcmzum1KFC7prM0mmApm20B9J4uLjZjxpoyu5sQEB+GpZwwKSOjb35tPudMV3ENBVP+JF
jGPhLx7HQuXoMLp7E9UEodLHf9QvA9OGxtPdaXYuJKr6RB0I4afQSV6FZmAZf/j5+aygLu2IlosJ
Zlvonc0nOS5lbQA5PdHwSTo3bzEBu5dX5y29K5/Ccu0HscbjD3nC1+nTYVHs5rzEnpe2UJG8e92l
O+mHR2zz1qWvi4ztKoFDuUryoW/Z5Su6TxQk8tDZh00I7Tot+urRVkz2vGowy0wrmo9/bZVpQdZG
26Z1/edJ9y6oSv2boae8dHTs4g3BdK1O/JzS5+t97snad7XQARgv44qGROmS8yKYofQ5DwLXKj1x
ZXSegg/EZHll4koVwjKy5TMdjBpRbF2S6ToPbFXSL/OOZrG7OYvqrhEdn8bX0DE3ibenUFGkXqUd
qlSEeRR2oHonDOx4+isTzbNS53Cyj37VVorefLKDbps7ELjF3zt35/kntaZe9pVYJ1TuaW1HHAzw
GZqWbOxiv6+sAp12zxUb6Ya/OBx1zQEaINKcyltkCP5LRZbWLw6imFXq9OpQUfhDzFtniLXAePae
vVKbh5UieV11ZVcbDqk7dsc3lAQ/9l3DmGu1VNA6ojLrI/eurdhXvWAwSaORrIt2p8ayEdVtGgzY
jPJaEfw9SN7a/KuYQG7OdOHPfGGsOjjWo03KOgyVaZ8zxe6Vs0IVd2cy1+u7giiEXFA9FBWn3YrP
EREIGQtX5hT4I0YU+S0LCwrF6DV2aF5Ab/yDjvHiMcVL53guYcGDqpUp4BlTPVNKwBywXnKGo98q
TNyG6HiXJe0ooJlL2zoPnTJr1GDUsvwIAYlMpfW+Y7l61aTTNF7+c51rXAU6hCvknm4D/aCChvyh
xFcZ17zdgTKxuYTpTimhgWEUZjuwWLVLp3LPaTVxt+yTz+OkyyjMPOyfCT1M5KCjAQGCJ1tMTG8d
LPk2MT+imxn9F7C9LzQQeS72HACIeKn3kTfktkn3M+BFIzewQigw4JHYTw8f7oEjlRtSV/m3GidI
aNdOo1Qr1xkxDrSbyc2RntKrJkOjKEqkKL5ES4FhRNS4XA2k5cRFmqPZyM3OTQguiDofp6vYJ+Bq
XvGrGIecPOYFKCPYBafclJyPTj0zxeCXw41whtqHX8dAG0MQZYON9jSq6duP1Z93PrmdeniWh7Cr
vmytVGGKmZkWncC6CgYd4/BC66+X9KG6FHTUrpYO1RlKVbvN8/34y0Zkzsu/9mvdbbcVW4SA+9fz
1tAZCMk4RJUA3tygmVzr3jS1CEE0Kvdwus1AE4KTyJljvHBs9xxoLoLD+g8OunE4yP6U+xUlVopF
OsufiziHR0yBmMavLQ0EUCwev/b+STf73aLLGTdyWc7sEnW1hJlcRyDVb3gAYrYUidL5zFHGA6H7
pIU/sclYKsFWOZJGp5gjleN+sZp73wQoH2AlIgOrTLqpYK825rMRU/mJoD4y0ODVgCTxFXl3HZNW
zDHc2SieS7n9at51FrgXX3favjCudbVxYb/XY5svL8w84/q/QnCmR/XulUnULZmIC+rKaIRz9jHT
n2FwJt7lMDrbBHXEBhV1Y2LSmH50k4q/jlYVSLlBojoNV6kIHunD8wvDlQ5LFlNklfUk83J4C4iE
XOwI8x4q08hVK4mkcTHngGaXt9/zFX0zZzcKpA5jaXOY9aZLWmKVqsPaG2MOHFpLauJgs/31haG8
1hVP0zt7ma33lXrRtTQFXIsZrOzKrC5w2liP3LhnY1dMh7syO5pJbMd8UHZj6IlFcg9qEgdS7f5d
orhV2tAOeUqzccHnm+yjmFxnAVsL/E2Yn0jHEagxmuZvBGHDSJvG3SG+qiuuhH2WcB7BtORXZVCT
+RgfFalLYpqLUlpMV2yp1o4ryEAeIuZ/qcPDzenKP5gLUsYkh9Ab7llNvwnp7Rj5XvHNOHpJT1bL
hOiA8rxZLGRPL1t47cgfYBHfRHaBVhFliQWVST/CzeUMdgdwlBRVTb/F+xxOxTrKW+bR7dX+azue
oED8MJFfstrP7Ds54YjsbhxnVumUb+Mn7096C349mLj7EiaXi/GLRYf/rMeBU0MPehIBPsQTqoD4
90gSa0dgc1I+85NDYNgEwoEElWeK4tfiI6TSO+C87oIAP4DOjI4Wagl3l8S2XJfJWAVmgC7iaa3D
0Tj/yEaS8eA89HQvBc0W/PnchX0cIv+Lg77/nUoLtMxox/Jq7asWRZGVNXLAjHchTyZJHb6+d5lu
wlHdBCiSyjm/SVL0kM4lY2oT0kfmyyLJGVxJDKajBovdXIlencb0Ur3M8ir1gMXJ3j5A8ng5ZBdb
WSKERfCoe1loNqHeqgFVPQ9dt4dmGqhqANQ2+pVwgxbFsGwh/q9gKhboi2B0maxXZb7MMPaJBpJd
bDIWjSIIzTJ87tu5lDqEaOHht+ly55HLas9QficSTx6rfOo0hTCHPrqUy1GEOxrs7qTcT6irAYNJ
TbkyDyDTO3vSY/OepZ26uqA0OqgeL0V9ode6UNysxoTK5Y/30rocayZqiUkqvy3wr5MUuPSiyW7N
ZHdRDryAulXOYokLeui6PSBbztTeTvzK5ReNjY/lzRze7hrt+RgFX/cVKkAYCWmLoAW5jXUQ9z2M
f607Wtl6KV7C6Jp7AdVReRVpomni42gzZ7uDvXUlnOaDjYOTKCnjzYKx5/MCM66860nOCvq4jV+r
H/MAmDMoo7Ds4y+ruEvhMJC0nfW0gMVtFOtnowR72bfqgn2bJWBxvvwtYe92mEFF6b+vkUUBC2up
op/cA+qHXpToINFooLyWm6vg9Qez32JPQ2OZAauZpkjbms1XVBoxl5rXolpzuKhtUl6rqCrw5dX7
wetJo1oeR8XITvQr9NvkVFwSd/BsmN6tPS8oYFW/VuavWK3TLbVH35Bs8alkpBWtK8/xEaQx4fF4
rdUJA8XIPH0ho6ZsTvLj4o4HJkXCifx4l6e0elBWyNmN/hW6NTgQZrOUvJ605aTfH4wkwzwfVNY3
vGpnqEHAZT8nNNzm/HKyL/BmpeNwYL/W3AwuTS90G/tPHxOfKSMJdpj4ml7LxN3s0kE0MurtgiXT
5/wUYS1byph3DgDtChh+/nMAkRnJmXnikl2rE0TmCLQo9SogSLy/L9/x67XI9+xpIx2koZIeNt+U
bIMEHTaHGrRT/tzaV53AVBmZHpHPVTPR+XVswjzTVz2+nInNuLj3k9Qp0328nJgqKdf7oJKw4m35
kiOBUam4pmhQ+35p9dHFe/DVp089xOdrnjDsc9ybGtSshvQC/G5NHA51rYgVyy7usbQ4sYyO2mbr
lSDuJyL7AAEEfB1XDla8RGBK8Ff5zMELYpfFlyZE5JTuVwbk/PfI6CQFMdF+Dj0j9mPK+QizBXcQ
vde1a0Ru+uUm4RVXUHis8JwzMx5+ekpfoDp34KWwtERhjmA2t0LiABrF1JD4QpNBTJw/lTaWlBU+
qNd5zv/xyTYMXP2i70Vq0GWQNykxtLvcuuY5tSa1WMGagCFp2nR2TRuAJqGlhTtVUb9Zpk7PHwnn
ABuq9DignStKa4XmfMHd9sHVPPlIYakZ5TGVUdl7WnbOoI6f/bk9axnaRKkQGRpPRDiWRMnSHwYe
LEjqLaxdMhMJJtWlZZoV4eHO0gh6fX2yXGuOUj9Z4nvg0fd6AQc1GwaqpxpH53vWTxxlx4jfNv3p
Y9hD7z0VkC5tmc1M1QDBdtelb9qktMMDaLEjBYTWhc0uLkRJBKYO/DVsPsDAEX90tBuHHhNDa20o
G7duc/mvUFKVH2nCv+TBpy65kH/VZAa+jf8Rmv70cau42iYky8GUjTrb364T5KFoFcefkq6TfJd9
VozAvvoJ/0zO6J2UQHcLuZ7D4BjdvhBOZ7wQmP0j9bfbuTTaaDJxioW8UGaRCQ/zkn9nE4RwzndG
SCbAK6xUJC5BcPwyUNuiid4cMyelr6ZTU+QqZYd8J2z+2eymRrhQbhu9FJiNsPXQRC4xUiBNAocF
1toNsz8W98IblFd0+DUNpP+pDL0yH57QGWLWE3VzXCVL8njRqmuRRdwX60Z5Lq132stjaszS8lyF
2Gssm6jbKWVT9pW4UfUmbdYGHYWEulzQODPxABeJLwJzhZbMiRyib2CTbzliZesw7JnhyRyI3HX2
8DkEZrJv22kSkycBQBoVbuiTqG0DmNbTo6xC/1bNWKKY1nTYUP0nlW2rK5yLxcBn6BPS4FoJd7wd
3ie8aLhhmlR2sQKbwPpo0iwqsDQXqIWO+6p6tQGQBBsRMS7xwkzqAp6t1VKWZ5zd6gAZFsUA39P6
gpX4BDz4b/b2Oy6mVKSQr7YOIosZV0mSy4k8J2jS152Q/tfLqAIIDv+bLV5yTJaqvfR7HqszgJwJ
e19VWeqtgx2TA+k4e5ELajAniVz87bd3t3qDqTk6wmKTYoJrqMfPsfFvXh7hnnykI0vxRlooU4zh
L9+QocvXstFg5jYB00sDbxJXKbdpYg0UkZlzDFGlwL7+5Po1tZTSR8BiRFfk85AbTlq91kSKeSjw
t9+LC7xCgFNtJSBSLQ/8l3ihzwrW4+LyNO2uRk2ANtlw7UEfmjsq0900L9oS3JGBoG/nE/lvK67+
PFCFKr3AAEKQdk6ItRz/kfqcqEfAU5Q8fnsNpV9Eclnq0oRMtp5O+8kuWUQcOv8DlsOLsBnMMRL3
4ep3epxl4wmVfG8ATXXTmVUaRWUOW6ourlQJyHdRn/O7eHf3hdQUpVcFjO59rq9mLgWPpr/Pd4SI
Hk8/UI0j/5cBxAKBp51PhBXHr6f62RjHBwgaOyxzhToUj4VlzAZZfOkEmJlR2Vlj9hs/1vLZUNFj
No/RhoJq4+GFyTT+VwKxOHeZJkS5xoYtuMjY2y+mkRnYT2hxRdSPRG7krAjmk06On3egi48iswxs
5pn6iQrsAU8+mnbqnep0LpVVJkxMdbO/onPHv5ij6eBHXgOjckycfE/Ox0EeFL1HgVh7/iAPdYRv
FIVPGmfbzSu5S2qwfoi+5cxkj7QbqfEU1tPSyYSo3JV5ytAMu9pjEC0Gn0wSdqa8qNNzmvmoG1jc
cq+xbvFd5kkQUJjdeDugmkoN1YpWPnfrytJcS77htbJvp99lo3viRIEkfN0EBQBLl0DXsjZdHOBr
ZNhPlvz1M9ZtBz5QEqA03HFJ9iYejAm+tCq8f6o1v4oCnlR425kouDNxrAan2GhERWnh6MO3Hcmf
x3hir8w5Lv5XfkoR8gBL+TMPeVHbtfWogsLU4eLVaw30XEWQaB+TnmJZ7TqQbDEOQ9fijpQjugXp
B4VVNLcscLHTRmcjHNj1A7fIWoeBg6aJnZ2SlPk+9V51JssskF/k4iTNoI74DkE4zE0jvqpGICvt
6onLuRQdRl7lM6IDbq8h+grK8sHAYO6mAVVzw1SdrIkR5CHN2rn/D2qsXC7ftfaJtQgSgCZ0/lLD
BW/b/xTOv65bDwSfIz8X8+tVUpX0d/rlBjWcXjk4YekYHD33GxqRr3wX+iJw2yHiOTRTi9th+8i/
vgM97BHf/agZYMLAozSw1GKv2kpCW+f2wL4AsJgKVyve3D6gUOyShOBZHQQYsIR0YxHm1oMresc7
TycITaeUUIzs5ZyFj027pH5hvtQzY8IVlc+MbWYVqLnDad8h+lEK488mKNLfBkDGRukCNHsi2Zo4
fbyefQKEgX3YI3DaXOy24B4oGdMVq1D6VaAM+Ls/Z1HrWS4ApF0oCEa0FLGyG51QBf/rmQ9hFqfa
54urNTKwi7Gf5gHXrsYyEUHZx0cEsSV59fD1MSk2BJdfbqzvojZGySqwvjbVESqkX7S0/qVHh8LZ
NdTC/r88z3dHk18p2NSPrfXHTK/YRMJwowxydQdWL4CwbY+jChnKYpL7w81YPvsq+Pc8yyPg9dmS
79YIOozSnreBGuUev05KhdGwJIpuo7OYZBHtBHccXVx7zzR24K/UM4bbRaHRbJL+bcSgXePwiSck
cP7jlg/PvyjDR7JQdlMSpCm45HN4TkVNje2Y2lk5nDJZnr4r/5f6NqWKjYkbdSFVAqp7+nr8QBR7
RanQkQLgQhw6N2IXpNhoaRQtA6SR/g99lEqnG/s3PG6cKRRx9KBLhPnxcY/NOxWQVd75QzXu05fO
/DfbIq8/7MfwoNiHxyMuCaALKOHAofr0JLOUqMsJt4oejB9BZmRtzknmvAdV0kKRPjkWHHMIXzmY
hZQkUhhyjclkz5qCW75kdDHNJu6OHwnNZc5UWaSAJ/0e/eT3N3i808VHwTmAwNb6u8ezumpnWE9s
BfB0ZhhNN7ua60JzlsKVvwZUhmUTHl0b54jFM1Z2LTQeB52ErT1pzE1xBcfMawpvM2nT6G524tEi
Kp5K5f1QIw/oOujo8Pj0y/xZzi7BzS4JrhtykutNYsuxqRj3uwUY2il+xRMAYcatJWOSAXKlbEuH
OFIdyGSodSUWfX7Auk/SIRKvjA/By+onxWHpAgFzg9/Zar1mLc5RpXU8Q7CmHG2JRC1v5m7zkuU6
m01ZMakhluZxenq5ydwKwj010FuZpjDJRpL0tPotT/0qW5vOIXTWYjpBODadR1fRMi13vgc0mYco
x911VT10AtLPXvI4bi8xC5gPsTD+kvMTEQlGxXxjtVBruuvc6eoZ/V0oZtuPKFPPkUXo2eeXgget
Rtj7HC/hLCbRo9IYSpybUHHi3ZbHUw8x5/DNdp8cxoS+PpzGVgkKhyt8HjKi7grCLQNLe6YodI9D
ohunpgla3ErDqiYNSWTqnn5z2ddMpyQHV+VOc/IVuXYyXcAh7bzvC5OIEoVxwRhTSLGsLHyynX7v
VGllGr8ditZGnWUxwkMUjdlpohLkvsDX2ElEM3jtTmmRJgQcnR6Z3/efVg3Jlv5VPyXQy4KlnhFk
fzrhKccDQrV0BxgL15S6IJkVNjB+4N5PSOW1quA355wvDQJAv+WdoQVMgAffjQkoMzdC6c/52mJ2
AmmHQM3GfrzfIIKxj9TBSMcxz5i/oWQG17OZh4/tYwjh760TkrZFl7zuCxokUA0yDeNBYFPsWEM2
zvmN3wQ9FCQkih8iQjGG5QfbVEuvTZ3/2+x4IvrMsekX162W+b0GXD4ZdjI0VYPvLX0Cpn+jcyBY
WqgjrgqOpRw048L7FQS/M6S5KlSJEsmMkKbvKBY3n1X6jKKcCmvmKodhWvrlpnfEkXeEIUytN7QR
j9qSomc0tLmzrESNiAwJhETIq4m2rHYHdjvpTxcmZZ5O8nUNa+QN3ePoLHiHSr8IQdHduWGj8IWh
NixFYwmu0YcC8te7O15JxEtTiC/9spjHQDB8o6YRc0tmmztRGfXRWcFJWMb9eCqqrfQ6n81jZDBq
MsT7bYdUO+gmWdEEI+9ApBRBhH4qlX+3zemZfI2Pk7gi1zCPUkuq2Vj/DLPP9F/d+4a60XxTjVeL
n9N4vRwCEVr0LE+1Pj1nOXoiUOzYuaZFY2SabjkYMBAoTUcBdRI2rxnrFSM3mIUV/5gY9hyDqqbx
4gVZIyjSxamZ1xMAMePXd149AchMoGUHkj6UmO6einUlgykTCF6wKbpBQ4hUJZ4ZtLUkkKvq/FJz
Az8MrZMZVUWTaRtwY+/6LtBoelkUolyPD4DLuBX1Y8/OH/y5RfL2yZvBZheqRe+DqsDvslqs0lzE
q2EEWIAFmUrryXTJyPO3rJyXSBJwgokfLexwDooKwE0R3B76fc69Mdh6Os3+BGPIBHMR7F7rID9k
MiA7GAbnSA2ennS4DCx2q0hMaYfm57qMC09Q/00J4y8MR5+n+MYysUVjJ0ThqUsLGh2wHyBl9JLi
/l7RWaEPmquC6ukKoYGAlnSWBx8a/vfT+BUo7tCeLUOHqX5Txe6M84Bt/M+HrOAjQMrNZSl037jp
jm8bMUNCl0dwvwusz2yzemw2igDRi8e39exLSyd2iKgHHntS/UdSyJYbyz4cE7mHFVfyggNLRv44
hgQea6rHCmsZseaVD9yFNENI/jsnVZAZfoecz0mLgixelx8TIcBtHSV9SqVmJEUJNRddqIujDmSv
ZYYg0oyvI+btZlp7uk/hdbb4lA9gHVTnQBpzRxlN5x2zHT1kQGHMuroebkHjnN1lCRzmMxb8s300
mt5f7kKQmjYxuQ76ZgCW3ob6h9Yd/GWQHYzTrFL91fGjl/044TwjLtw0iyqGGV6Tfsw7Us7aXzZ4
eMXo4UfQalQGNJpgk8zrFMw07eo8143Z7o2HdjNVZ1QEV0Tx1SXtg3PQcJUxxbYZD5gJ2QbAuICu
s33ndJCzYMSbLEovUFKxYdr6R0flYjv2F3RcY98eZSGqEcgpUbWxvOLKp0MkFCxq0inSBw1RuJRD
4h8MsnnU7LO83cChx7eT3c1npDHR8YPZVh6MR6SVKywUPU09vHDfyBxiFfzz9fZK5Ce/v5+EhXzU
1Y8KyUWFBRDIkcviwUg0JfFItdxwYq8oOp/XjC144bZ8QEnqkAtw2/a8+LilM4axLUcRlI3QyiKK
V538b7sdp9cOplHHvyZpz38+R3fmn7FLKSEQUoEnGgEDW2ruW4XTSHdrTRpP1P+519Y7UDNNtadB
hHXrPaFVPScrWrDrytZStb4Hz++5R4AnO55NwReDPRTivv2h2o5BpGO4lwZ5XlDCBHumaHGZaObb
vOJLQ7+HuIBKVdsJIPjmZsTrL/7YOmfjT8T2kKLsqYPJELhIkDfY0/FWQEcgOhbI5sKFG3WUVG7l
ykwtmiBUNoB+9w5XpQkbQ0ndXvgQ8qNstj6LdafpgCyrOqM1dozT5dshIyLEeTORIx5jRdL8zl7b
CaAjTYTe5Q2AlQk4vuXjVhl1vXM8JZBGe/6XgDJJJLqqECxYsubzS3a3Zsi7+TDi975Pcw32FFRO
DVIMEPRxCr3LEecCjSC+sCc2wLj94qnh2vIgFQwt8/tl3JRU8zABUK456I+MeWYBfVW5lekdxELM
3Emjg7OJHTKoDEe2KG58djUHraCVV4RU+Dipif+3IY3JwA/n6jS+1e9OqJd08Irwj3wJlNP75sBT
UhDJKBG+B6pXDp4oTr3p8E2Xyz0Y/fuhTZ5FgOOUWGrN+rqfGO8Nbe1M3M3QWj8xq6bEwhs8fytJ
7HLNsOkd7wJPAazW4Qle1tKWag6gcdP1/PfiWVH5SMoIZ+oOigAhj+l8ZQc2XiQPMe26/c5YTMiH
iDlAD4cqIUc9mYGYSyJqKQrKIj6I/UFDWXgq16x+3M4s4+QG1uXwOd/gS4QiiwiN1cKGFHPqJpMG
4LyowYhrRLxNEmHcGRZ3KSTfma4dgD++ch/bxvdcN1dkScbV/8WDL0e/26ZjIXTsyW7H/PGsMMxp
jEosV75WGdih9t+kcPfag5bIztHQHqcka0wpxCPjpwhpuz0lFVfC3Tld1t6CG6Tg7D8XKyP5Wnxr
q6uQp5oDMb9lYRtDk5DOzz30n3/ffh1zD45ZI/p0BFXcdQnFMSw6DyOVgeKLgb5DnOnfi4yk8nL+
Gs+iYb2sVbDty63BjcsXpN0Fly/lmkKiekNrY1sgRLfZCHwk3a+jN7F1ppWsLiIPafJE9j4hzIrp
XYDTDW4vWkRubYknYQhEFzBhDDpr3ykYVZh+gK9Pa9WADqF6vAyuPB7crknm1kM1H6FnFZ2ay2MG
nGpvErwVwqbvaTo9QkMpV5RRLT9deyUSSqM7lT5whTyikBVh+Wd9MzAJyNFDuVI5ARNurTViw2PG
vedAMlKOcbS+0bxqI/pvyPGBHAd/9wa4TXoxoR+f2RWdzbLzi+GphvyhYqhNvCDJFWCGy9ZCqH4S
bbJkUdbVw/D+SQqJ9V0ZCppiiyJ4oDhwtgA+S7J1gQ9AduZ7hm4okX3gYZAMnyUIR3N0+/xuJ7t+
C4ZFtEGx2NCD1kvnUPjajqEG8Uzt/IySSbz13ZQLAx6qD62UqL2Fp3dmhzZR1J0ClI5//D+joIjy
0vbkTJ7/HvoU5izZyqVMIjXtVOXtKvy0stth5IicTymuD96NS3EN7K1WmWWKb5n4S6Vva1dBYWFh
rBkuUXv8LriO3pbkqsWvIgmJQUZimcsnG4aPk99VNl/Qpd1xVLSnszNkgOU1rdimfyPfEPpf4fkG
ieQSw8eQzPcvhZwIhDaKcnKrv9Jh6tYTX/6jKobyrJqXhYTdT72Z77m8cgDp7FrNuez0eQny+zVr
mYNJZsE5d6l7s7ry8tm8/6n+l5kNgv1yztVSQuuJxreD+J0VKxl3I601VH2y5PP3/FRwWb6AGf7o
KxDkJWh8TcGEPIUvPdW9xoMtz/fTMLUzbm69a1Ir4kCjarx7JthaqAAIN7vL4ikeqUzyhUB0H1DL
vu39AFDhlXmpjKfx9bv4g5aa/rE0iNirxrtx1bcbT0kAEhFgAaOs/5S6V3/0vw8wnhOCr708MCaU
SWH/GEscbs+7envJCn8A8updAzO3TXNDoXkPoY5PbNVa+0b3GKzKAV0rAT7EsT2jr/iy/i6p4UxP
XZFSARXxJ/WixLFHPIIABlfejt0Z8CNGDfyIsWmLLXfxNmZUxtiWfOpAaFDUCcnfW5xQG7Kd3Pb0
SUvD9SkN7SldnsWC75xZ/zkqal7LDrQLTGI7Pz78gjIb+Qy+HgVUyDmdafynRLqCML8GDvNtLZGk
mPPLchK1Re5mmda9wzP9yClKQSmTY61grwUa4qhGQ8gUTo17eq8J68Fl3BeK5RsPOToZWVDzw8TG
LaCLuf+vJiyvumHcbLS8Pe18H2X0vzWZ6bFMWjglJEI/O35L9L30vjUXS2hqRPWTdWss8/lERXHq
0J2cRPnomXpgdWB/S98S6wgDGiFcrp6rD4yTZcvHfGKUgR1ck/RxYiKJo4Xt1PvNGBdGkSWuntJm
efftjiDyUMjrMPBSLkS25osH7vH7LDUTtCJw0gmNVbLsM4WehZrkv5xNY50oP+WSQPqtvsFF1NNa
t6doxQ3gqYKyHkdsWBDcJYGj2J0tjNNFYZw+XRl6KnRhwrMq5DsxinQkVVcuYIdXEkhhhz7s4aZU
8ajweqRgAklgxa4TB211C76U2YrUh6xuSZBBhDsp05EYjJ7arGlKaJX/QRG73g9LBgNjO7RIqiPc
QzAA1Ltq6sQA0P50uVmXNyP6Ei4BBcBYlh1hWFBQmFdTzBEOlCF5drtD/sh4DyGFL8kNhzo99dL9
3wnE2RHgLGVSyPg/0phmIa9ky4H6KyLeN6p6Gv5tHKXDieNsVt3/h2MYrwlI7eZSI6EiJuONf6Vl
eM5J60xdNsOxUWXhp/HbU6+E9ZT7iPma+IKo62XjT2bBXOTtShLqiqhULBRpkq7BJTThlpqS2k1h
j8MYGglkfivLa6MWOCG0GeebTLG6lLJJ5tgS6Cfpl4dFenOQPHc+H45kUEazF/AsjRvPhbSbKoUr
ljP3uu4CMVSBBkHizXRMiZt1l3eDHPPq88Ifl7cG6wJOqMfOaEJFHt5LSE/2WKQXNTQ68UHbj0yp
sli6zThdFc5pcAJN4LEIhPEtDyc8L1tmHoY832W+oZAJ4mDPqLwSc07+Wlu+U47xabzkdqTqI2QZ
ZCfsFR1r22XL25lda+f7nbko86ZltnGfw0r1lAuZXeOBLlgvnlRokAEcbu/h03FcMqyayQTENRH3
L75xLNqbs2sFKrreSIoz1UqfD2N36IVwJ99/UXzuRbLjygGTehQs2JR+9K/5778jypSyXMUkbmlS
HnhTVCgoAacKKpB5OSiJb5TFcLtxuJBfQCL/urL8IDr3LFggEMTJCbMf6tMil0NxEh9JEQxionHE
QsVzFFysAQ0g8Zrj/dE2CsJFvWeM2S/n6s92UkJWf0hEFOMtoSXihG5uSzlOZwsxTH84e57BwVQ/
I7Eq/oyvJpoATBm5nRfVm61zmSISDuJ9HXrH3KaiQAuaIRGCAv6ruSrIEufpRoZXBHV900iswfjS
Rh4aTYC3kLvKFekxyjn3Ml7wNa9tzHc7851T6K5bcaTlphOH/OH0zEy8numw9bRQn0t71UlyoIrX
RlPBQZEDbSqOEi26I1kusa+NfIqIezn/S0jxXzcxW53IMfgaW5deuGiAXuU0a+lslkP/o3iNaQf3
KAPfHyDBfkLX4+3qHy2fZ/88XdVwjeCbyKHd0qKNWMAWOe9mEK0mljKhvwAqbNdf1+SBOXpxbpLY
CFloxoULKoYN2c6WaUUfTQj6dg7FOxaq5fHuYoyf2GUwElwaKCKX3TLCK3xHOU2X0f6iffvH203X
h4N929qg0of8ZHW79i4jIsUTualrDNR0QOFJ6uXMp/GDRacqHjsehIuPSmRjHXPwqVxFs5csXXfv
TUTNuDRtXFmIce7DT3oHeBI1YijvbivGLN3EPwiGuF8Y1bY8p4AtPZuY5MNX/stAGlWC40GuDA4/
licD7uTwRE42JQSCJbdHTW9ttB6Q/s9duzsbojj7xNUGQkNUv89RMQtnQb4DXn+/vNe7M+cmKxns
zV1dmYMhIg/Cz2JAyDmFZc1GRFXy96h41kZX2vzWFVdtrzTRHbrBgfK9pNl2vZU3fsIzynbD3W67
SHGJD4RlE3pSehTYjD+Xheyo0wbyRRUBCkd7+SQKys9ONFp0ERCTUIHAtCpoox2GQpNuHoqBKRBf
xZ2gqq3ahPgebOL3KkdYd5O777MVBwrv/mwswPMw0Q2sDQTIoyz4evQTXdH4FaAbLG7CDTKSQbtg
oJ3vCKrUxTg9LO4d6x3GQ8upweU3VuIXgezDjYOgzEB+6+QmS+drMak/CqnnkMA4B6oUZT1jvzyK
clIyEPSBL2vdZ1lEC/fVd+VnJ1LDHRQ51RTfq+mL9KVpdFuQuWUH/L+INbeOSmCwe+XBiKPRq8w/
hGK7uMcl2/8hp/jwBbkNBvqxtZYhVAMbiMPUNGgdl5cWCHlE3GaV6GjTlgVUsUxI70I6Kw2yUM8f
yA7p86B2fNz3I2e9K59R+AW6U82KNkPGPsU8hkDVzoHqx4+iJzbCWD3KdmW8dlotfjJXI6xyeg8E
iYNFP8QWu1Pv5HnSRbxA9UG+5OosYS+gQ+eoEA2NN/RVqZpOynQ/NQfMnBr2+rtO1pcqvQZSfZes
kiNWZytvHGyJ5WFFafCIOeDRGetnvf3i513L5DOn+vvovc8woWPhgVbLyfDPFOFi6X+LSIxBa1q9
Ya9QSOI2AmyfHnUmDmWeCrYHMHUwxv/SY1Qoi5LXe0UDu5sabc/XDhnbN2dpQNsAewgsoW9Klw4g
fOUamw2jncV+fqgtLzsAltWlBUqrCv7ZR3G4Lrz607yFn26/RpJaw8PIsZVpmjUSBfBdH9w0BEWk
B1Ge69r7NVR47Jx7oEhWDA0SRBW7h0r7XUYfVqr/Xm5yIC7qp3cwGseF6cwxpeD7gQ4DWC5wZW+k
0bTYu09gfr5hp4HbDgfgeBnNbxOsAg0pC57dmL+bcPpBl0ScVPBxp3L+T9MBrGKD1Igc/OgnAL0u
27M2qdbrqPUPavusTqoUTjj9IIV2L5tGlzRJaEOgAcbn2sCjxUzwlkf5f6GrAjYz2RA9rXVGa6PV
VXsl7Yp1zvknpETzetIQ8qUs276OcMoGiufNkZBxoHaE82CQYyFu1NJx1/hszPucPlLjz1xxRHFz
XKh8a4Qz5zx7JAYRvbO6ODWrcuE9DW1ayZ/zdLLQZINvoQV2KjihMWADU0lT1WjjkJuCocA5YnFF
jt5VF0Ekr/wgCs4fvTim5/W3TCWWvt8j6AUXI7J0s4bTBOXYP5llgRu4j++5RrzQCJe9cHDbxxNP
BHz+6mW0BeBi9vi704KYcgeDOs6y84CQWg6lS053xI/9Hfd/WTHyIy64Rv23LSr5236qAjmwlWUW
sjC2JYt49nmDd+BAms8FAN15986X8kc8aeM/aX0lTHXtrzdy1kjOQF9e2Z5aLi+IAY0eXmzZXie/
A8Nvj2FCRZT6WB2sNZW0LO7xUerR9TXD/g23AsQuAFYsslZG/MZe0s5Koq+UMHekDF8uo9CJqk18
hgso8jwu+fUaphI/4pCnDBRhsugKr2X3ES/50ptp0KmYghLQieVBq8VYbdiHl8LXqWBuvoqMO1zQ
7FHNlCk1l5Qc0fJLKhFZaLMvA06RYZPaECnNNwTDEcGntLsT3K3i1toZwTaeDxr7Iyne1Rv+b5zT
7VO3xZcVdg+NWagCNjV4Sxhl1kBcpiO9Hyk+faueZzvJfGE/h9Rwj4l8n21DEDtPFrfi58sHq8hO
NoN7o5GGXL1iOV73V229j3lkSZELLQAnqP0rSWrHS6VtWUqlFptt3CVkRJYk+qeTBuZERlnrp1om
i9x2YrWFymLltjZHlUNIXEH4DGSUNQXMrnUneBUsegr6WLNm54Cjot/Wiu1CPrnJhSMwo7WIVZ39
n82AoF+4r7tUYddrsNHpLAGtWqUgo74YmXDEClATefCc6dzTLXqWrBPL0J5+jGkWLhwxE+es3Nf3
OVucCfG8gk7BqX+VbiK84BvLEK7bYERhBTkCXUb0c6+BLbWwMjQmuz8QL9PKnzKtgxEFAbcFN6qZ
EtoEzLM+NAPPAa6TlNX9OP0Ro+PFjT6BaFNdvOl5UgYwtcXa6saiUY4G50wGPE8w3CV3E5ZE2cwy
1BvukWX/ggt6aOg3+o2ghTB+JR+fn10NQ17oPzWPr+r1o9/3n/ZDo7mHOYw38n6S1NNBz3n+NZZq
CPwRrLSWonWzgxvTSh/jpsS3RER3Bna5nvTyZEZ00ADA8SozlSJUeVaih3cBPeZmekYqHGEIh2Iq
1YUk39hReowICjwcs49BYMMLMw0C3WljInuOPRbyvZhokaJD7z3/S/G4dblwtl18w53HqsQnXhBn
DRZOC4cxA3hHBPDuQMnfywBoYXytfQz57xydvqBGXKs5rYOs2VVKDC4zixJcfTxMyOvif+ye6dUa
DgwN5vBbIBZxXjVRbdZ5Qd44OT8nXnw3uA+KNeaRryg1nPv6uU1mKyTMHtPywUA8UggG8DcIu30q
8dJJLpTRYVzRu6jk+k0cvTimb9XDg7qAP8zyx+CBXkHh59agJg+lFeLY+JkdvFv9UP17TltybZFo
kBGaHK5babqvnoj2IQ+aSo7QhCduF07KdPIoQxOvuwpm7AQ/SjDSXb939bZLWUW6/JbikZjA3nAX
FujfEBFE9E2g4s9AyqyTzUetxI9h3YNyO51bkx4RekU9pfYN91+csU9xqb1wBpdjbt27anPyJsUO
6ZJnOZS/ktS9N2h1VY3S7fnfhIz+ayqsYp07Pu9AZRmFHbojxj8nCajXxWrHT/4qTy9xo/PStPpd
npHK4yE2KrnuewrfdSUnjjVCel4uNwdsf2iAcB4bxelrrkeI9zXj2eueCx59TLiBlHFBRVQgbUF+
m5Y5PNsKx070axPePpSSfRZbUZ5D02A83HqkzwIBU9EzcFDsV8MIuEPnc+x7gG9OI8v8xBRydcAX
HS0xUqlp5CtESkZpWGhwvsp9euUX44ce/sV3YzOqVMJBcKEkZaz3b0jfC9Ddv2kFQjSEuBCyVXtJ
sZ/7xgJ/lTnuMtMLJnyP/eXEVu/AcQHog4U26OCGGmW743ZUVyJv8126bdYL4P7dWOlF0Vl5oA85
jR53TXWrrC6i9mkaLyk0+Cu0URiHswsV0eSCBtb0ToXn1XOsDdphuyx1/4P6eIxJuqdnGJ7qyewn
GosxdpJQsP73Lp5dfUGEFkTSCsLLXk1chcOzZsgRbJxon/AyyFNbUaQJkuo/EpZ3BJv/FnOuS6qO
qTmPVGZtIexcXPvxHlHEBCwvWcl54CXLmzuodzRRDlH+F+qe2/r3H/Cx4FF30qYLt6aCL9ohEH7A
Oto7eCf1TdPiXmioIeJfqiRNFFqkAOKH76+lL3VT4l1W6JE/GevgxLUnr+lWi7gGzACsvGPaaNjq
C2stBvU4d8efBLJ6STE0ZAh09wmn5CoHUUPYkOz2QspzXWY1yQWSpL4iGh5Cx/MAYY0io2Cx9YY+
gGc9XpiUyYZ484HOgZfILNDNdLWLU2TdA5YAqz9HCEjI95RcI8DKvgWRtZlPiu3zySthQUINt4vi
fnYCRtOqhlDW2zfVHY9bLVyZwgp5RlzOqVpYI9eGDEvZSxiGIXUrwgus8++aWLxRcuXI+cZhNgvh
mQR5a0VARVs5lOLHCVv9jehm4cstKvPpLtZCBVlkX0yq7+C+1/2aCG/4sB0o7LsYGuyXs0ZFce+Y
eKfkxdijfvE7RAqIO0gzjffKLlygfC1cK4Yk/KfOxTysQCsfQ/WLVVeLNlo3fqPtvw13G0GGBc0f
nlErKjsZSfDK4tTc+vGs3vol5rYvg7jmw+uZ6do/FrOGVZpyirK5CEZvjmcEC+JSIGIys2wXloeI
16pNskGZ8jvt11pRr8YKdtRaQEz1MUelZyQosqo3sCe4efImNqn89jZobS44TLOW6IYjV/UNrxOv
IvYbJtKtsaexV1sff7HyZaktcBx0yV3sc2Tqxpx2izDog49EsskEY6eF6Hhk01upOQND7ipvnF2N
1wUWJ2ftuMBv8MXAk2b6ibhFmkhjbS6e1SJpuEhOUTSd7unIyc7/v//dbMCsmy9U1aX9KYJxzype
mQKHy/g5v4458GXfwkOSnyxo3eg0aMK1jAsPzRDispGrlIiAYDyVBaUkIK+3yCGxaUiyHwKhlxFb
fbAcnrgtpLHesvKM34xuR4BkmDu19hixDGmh4QF8R22SDTvXwh/7hJywPQGc4DCZl+ox9xP3RPGM
pXKVT3RV6u6CCBBxf2+5zed5bp+/foccC97Gdrezgbm+3n0jbBPFq4cs4Lt6IHw2EGAzP3vdRF5d
DKfXNu7cWtPEUgm0PT2ICEpHVJdNmy/tTGYH24dHyLpqkEJ7xSALPv9F1018fbYqvbeVn2awNII1
52y6JSBRb+PLVZz5/DZ+o37aqFcBGSDp6rknqB/+i+bNRNNm7uF18Nclk+W+mWJQSAJUVdCZOgTv
Z6uxPNRUUgxNxUdQ4sgRSqSarw+tR5m3l6hXSJ6GW0F6ICEIrMEFK5AFPmH10QfeSZKvhB8W1tvB
EMKHC3KuLTdWoEyOr21IsUegfjQN29Sjhg17IaMmm7rttkJuYNGtofONDH3k5g0tw/bxc0h7Jbxy
Hd5JG06Cg734GnYcLDzcE7O5cYQ1tjiKmqOVIR8hR96QStUDZCoNpeBcAUFYvKefKGC4SismSkAL
pA5VUKHbrbnoP/PYUrbzw0/Ipow7cc76/E+ULTJJnq5pObGjtkAPlzJFGFdnYtP9S5qCFvrDsZ0q
6iP2oDYDGtmXbuABzQczuoRcBpRI0t9BvDjPZHo7wIhLBQFvvcg5Uy4VLZL3416kjRLC9H1VgBMV
3pbkSsclL215T/7697E1lJv3HKTISRlMjom5MxCXvbW51hye26WwVaJbAC5EVKZeISQeYI1YquoT
axAHzA4eHAzg/jlyvZZR2CWMPkYekH8Bwoveq3OzGz3gWUT4dhNG4wHoWazDAB/hArmuTUrU/zRh
uwnoLbxO0zD/QSsADEz2+DJ5yrDwHFZ55DWsvGBZvMkFTrO+fGcNxqsaG4EuogIf2kRFNdcBtMhS
w/PH8k0qGs6C3pHmLVCRKVAhWsBNPNYOCN3e7y1DYC2m/DpvE6/0Mjlt++gdrqsFH/J4D+CKRpNC
0VRNUQ87CfHZY2LHHjgcTvktjG6b47nR+baVQIzm0gsb3LE/VYmVNiTH+xCfq5gcKK9dB2l3oEAs
DC8v/gEH/5Jgsayz6T0zvISQ8TY0TahSD4VUi75u+BoDs+HYrBiABMMJl3AKVZ9svTq+fLIhEWvN
A0W26HpkKdl3AIPzJENzrCMwZmwBnm0potL4JMAA4wZXUCntNpfBoobPyUtuR/ouV9NvAKnvsmEV
hUvQsdLjm8aY8y11x175uXI4VkKXVYcsS/sYH54c8wyZKM1ezUIIWorm/9oWOM8NmTJ/t2XOTzob
CydLgQ4yp15DXWiSF1LI5n5OioLsd4l2FhTE2GVMzPLeyMZJZsovFZM0BQa/SqXR2xZq5jN+hR7b
/youQU6ymUAZF4FC/9spysRdrx3RwIxW4g1kgL8/2emHi2xmYBtRkTyM0jnhc1llZyg4kRNC8QH/
ls0jV2fA5tUKv+b8i1EU40qQ3V/wbmDW5XVwmTgjPAO6Til341OMTF6J1BbZaTWU3dh15TVijKMx
fUOwRl+aew08fMEeupy8mrFtLu222duvYvVrCGZ9+bI1LEb/V5MPdSWW2stCizM4jNeoubt9Y12G
6aK1A7jAUosO9omQzGivuxJKNpHAfsz1iEgAYT2qQbDwIf+8+f1q9IjiwNVj3ju8wgD+LXQ8DA/c
7AmrL02jRyP/kbgtxsIs9gPIXz3fjKAh19EywxXQyhtwQjmROcaTBZonsJIS5JHA+2splZ0QZ/MG
kwDNQUtODbSAqcAZGjenBvj5YNxMVA+1elFAlw6zl3XlbrLMJg4p09KpJXzswRJlBu5yRGEGEp4r
Eaqeg7OeTcbWETNwP9bysJ0GO/nrJXE2A1ml0mg0a0TJVym2yIwPDncWtIvM+FYY+PEjPyzovgql
pm4UhEO6t4lk4RYsrxlndlV6XuQdThl8XnF+V5fWXH5Mcccf9QXX1HK1+zDC3kbuTdDGZJL5W5iR
MBq7Y4KvzyhFiNA7ek1BcA8aj5236SHxT6Es7dYDjdpru/15tvJS7v8YfFagDpJTzpIxu3Jzt+w6
XDRuNwxI9Mw5VFG4eCiFWwDfdserJ30E5ESS4unwnVLDdrdvMixborTFGY2Mqq5Lm1iYxIz2jYxC
C5iImJt7XMtIzyuL/JKbx/dXcUR46RA5T0+/A8PQCIKAUOhLo9dgbWp77gNzQHwvjjpcGiVWAXOH
ADekDaMyP8OA0U+segi+1kHF5IjroSwHEdwLwdxqbofShCxpKdJ4MNHXR6+YLeE9M5n1lvPMiljX
22T2yFecfg1TJZVaQKk89wYLt23/XqGgp1aNPe79i95ZJdkVzKX2v7cqcDXuEn6pUretRqXDYFiJ
HVjTT6hlhcG12EWokdxf9WLYlv9O3Ojvix/+tUcjzdxuI/pAZnRlb1YpAM1X/HZ6RmEkQ4hdf5gj
l1MzQWjT7bxJWEC70cegzd7ibfnSoYOvmwVFxvlzByzvufxD+fLpBH3iK8abDY3ggCk8ELIJwpz7
ICbBKJcNulIbCq3pL8bpIWpSaLRAUpKy8hPklhEzXsioy67L2HoI7A7Y3H1jiPIRNp10em60fZx7
PkEeGPZ8iEgJd6EUPwDjhxIZpw5RB1l5xd8wHdvrTT5msQYKUnYuucXes2+V8tf4nK9jC8dihPV3
HmcG1YaNCoUCuMAxZ2wluvE65+Jwc5TP9ouHc/EX0h5xRli6Ml4xH7LNcTymJ+7dLtJEhDpKk8oa
0YJa6U3lIqT/gQGIyu7tZ2jZegK80HT3NY2xJVFMDiZnhIdKCIvF4GlYpFQ//mxKMa7nhPx1IY6e
5nkeBjRsLY/OfpDCLwH8jdbY0cHujioxWuewkELOKKKLa2s8IOSV4Nwb17/BJrtE59o5h5mJC2pD
KLgxagpj/E3yumPYc05g9og3MriTv4IKE1ss1gpHoetU1ooZ2iZen+/LPSFF0HYuH0yNxAnnzwx1
kgo2jcJBYe9LkZiz79RndU5Uq28Qor+7xnLweFxfKFOhFc9+PrnOpQLsm1UleMu0qnhSHTyvH+Es
4v3RkmGoZVqvjxXGXtDWjC+SjaBXMMqYYtbQgJS4pH9u+28yeUWcdcDC3G4/z8RzTDL0A8xlicJR
B8uIRl+fd384AB4sHw5CEtjy7vKawzhRdJCZW639QpLQWnnNE4savK+3eU2LQtc78/MOtEMmhC/l
hOwLy3uin7UE/0f7m66MMUOPye8JrxJ7/6f1k4TETm6nZplczxL+5OgX0eE7ZvvIj71McGDj9hIi
Oa2QF+vm7wBMiFuCkxSaKugg9G54cl0ZH7965Din82Nne3vpaVjGoviwOx1gUgfBFa6HkcRKGSSF
6C/9XfJqD+9uEgJS/AFaOJFvMfCV6rZ9tzW1i2+SvmRnZNjzKaQmsLe4Qr60ZNPUvsqiiA2bpt/S
3zdtng5tYoKLjar7jWOkV9O3mW9mokQh87aElB0IxtVFn8vxlr0j6eMkkqVpzNoc1FhOdF6VSmyS
YIeD48EQ7Sory9o+7CmhEXvxashY/sW+isboBOvcxjLMtLnfL7EnJaT4YqjphzabOivw6eHpCbHI
M4VQBWKPeOyBYvROPNoe/bK5x6Nt7KYlxmVtQGZvvHHgXg57luF1U1oVUmNGo0movcGNfiiIj8Xh
5hqePLKcWTotl3314aCG2cPHDZtr1F4KFNZdbSLROBnaUUDdu9dXWtJBit5V0p9Kjk9fS1z7BvmV
l26D2g6kziYDTZ7gYi5wxs7eqUidSXuyR6fhkCYNEc4VlWzA42bxWIwxHwEgsVSpDChH9JGv+WHO
LrrWEW4DjALWUnNiCLQOAJVqqpRhCHbwqdsCHVzfBuqQZY1/SeELj6oocKiRc3P4Mnwg99D5e+tB
j/30kJNqrSzZ82lxMiLlpJnOzA1p88o1PhSMVasNYC8V6oDJm90VpuoLNnLj3vP/sFOch/xPXOH0
jrHSwlxRNQ6Q4ewq9UNa9HSyKGjIF7H/fMaKqoGqc76ITHKpesJ0Ob/z9ec6EkygTcefAEQHZdIY
f1nMdhKRfbhbikshgz54lBkLFztPoxHdg6K1sYp4B/Lqb2vaE0cxXDI6sg3SjLWVw2fCFs4+L5AR
LoUZWiy3HtU24viDoQW4hj5iBy2Cl+1h5xVjSvrRyizO2glA54N8FS7er73Qr+0wuXtN26m/fizF
/k27TDff50ZpqUpAXRNmJR7QD4mYf2fBlO9XbT+iPp/1TNg56VRZC9Z/1c0j75BX9zoxlfZVKDjs
N/offVE9z+kYLZrMcSk6nF9sXvphcumT6V8ZPcrDFNebod4JFPyphgh+3cqtJ6sqAJIBX187u3l4
VzFGVDhgrA5zuM8XkpLT6t82rnVGKYNUPlZMia1qwJxLRSCtCOslrV6QMM1bfx8VZaDBe5Gk0/Ow
nbPsl8kEx4jsuPMYuGgGCYe28jBmdBN02ot8CSiIuzLv+um9tbSkkXGSEToQVVTcYZodqV/YfxGH
5uo6jGGT/GBsTvKNZRIYECMJz8hR9KgB0kV7j149Nk82X4j8KFCRJZTw2L4rBzCd+2y/e2fmrYge
SXoY6nMGi2w2+uFtWDPwEmTgtjeVzBWl7HkuGAV3Hu4/OmPmf116vGVH5FJWDZK0H/6o12cf6XvS
VyBfFclrtd9/P+ekhZ4cR2oZ6y9eQfaxQEuI32DjXCqcA7g4MzvXcJmq3ZqswgKUsy8Z3EW4Z9l3
GvXDAVs4sHdDFJt+SrhGTmfQn+fsEd+ehjPtNobk/zRtfSAe/sgzoOInF58Onl+eATuFIdlE0xo9
g6SrBTDGyAIJSe5qyziAuQ5YMf4GpejfDw4SvHjG5u/EJZSPtQIYlL4ZLiyCSvEj7Qo5bXXM5Cd1
Uwq3s0yoC+227qHvT06tWJrVGCCNF5uh4eVYTRIcUF+Xu/cQ0uGH7Z9GJtcVwnCD3UJWLiozykn4
2N3jLk+77rQlW38JR4QiVpLa2u184P0JUCrq0TnQbTjeODhlHEBWz2PdAQVx0IZ8CM2epXBgH6RM
3xap9kky/DFlh/PeY3sbbry26xhRNPugmuqT3HLsjqX7FetTjO+mUola3PCUZQk8D91fkZMYtKPv
ljlORVIUDUIc4QsxvqOz7ShCHwbep3tmCGG8MUOsU8UxWq7KHK3W0owzbfjTZARS6Fj9jV341C/m
uaeHQNqGgqO0lUgQyBFcjNsjz8wzVmS0j+xkuDGiwoyUFDNYc1e8zSMyOMMCcMpIaJ8+VxKXfhEW
PEP7vpaHKL5sGzugb/6BYqROnTt1SZW+WioQ2pjUYcMFdT7MXAlPJjSrQh2+Ku7q1IlWzAHCbb92
BAtVWXJlQ6GT2f1teBJAXhZEqV1uQBWWpDVJHAUBaAyInIKvMd5rhfmQ7q2FoDV/2Gad5XQ1BKXj
hYKdClwWITD0k/g7n4C6w4uG2opJNdiOGwTVjiYGefUHK7H94THc8oBZQWLolYbVV9fBuhSa5X5g
p3EeyvHXsJsJ9U/fLWrv/ol9cJfcmg+WvtLbEUxHt6UloCKQziTi5YEQBjMcWveFkEC+PqPV4w3D
QIthEgxixN6L4iw25aMdwKYbxiNJ3wYTM/IhCv7ZqEr1mbz83aMAvvaCYoAZ7glcm1Bw8RI3B2C2
fEvMtcV32yg4OrxbATOMwWJdrPqyNJFsJy38XqYdsD2BQJVvtP9vLg5rxUxxZBx0cQGkVp0oehmy
C20H6pjUnVQEbaU1Hg6FCbw5K1715tOWDDPHSJB+I6wNwuxsFAzZP182BSfZgwMMkaOORGC1/JrI
CkRul5GuSAOJXoxgmwou/xqSrIbHE3R0KK7ffgHZxk8tyYwsrhsxh5SAtIDfi80my+saQg/4ut/k
CICLbC/zspYZDJ28YlF5eKlsTGfaW3i4868S2H/6lipk9PnwE4hY+1vFFKXdAN3LmGFIuCH7i1W3
DDUnDxL64fOLnIrBUKYF/xyO8LNcr7iUj1q1fVQ2ioWYF+6+nbxK3aVkwGPGFWOwVNg6E8oFpTrC
ksocrdyr73mGUiBGktGRzs99d3D02Fx/gjkNHEqHFRamlHtudjh2OZ7sHP9WBOpskkR9QhOeyGTB
um88T+ZbKSAW2nLz9KEkCosfW6q6Ophrdr/Tt6m3HQGO1nQe31wpTagkGY7SDtSrOA1Yjj88mNBh
tTe/r3eOXThLahub2lxtCP3i7/aCjChfXNlYeuL7LsLHvE7TpRQ4qNwMeczpS/ZD19jiFp1ibypR
SHUSIhB2+11dhRg57uSbePYcsPoCljnr2RHwfWB1SnLJ8tcHuG2XqCM0dBnqCeMqV7Z5ukjRr/Va
wR0IzAenUaiOvwGRGYPOhXPRQIiEqtdqT7sqZomCGluaK1xv8Z4G735+YLrmFJdWGnKe0tA1SN40
+gCGsd6IDlwHiKFcdmQuPNLyTP+ChRFrH2MQyYkXC6kwnlZxA/ugPjWbxfQKjIK/4zHAJ6qkZwuf
dqDBT8URGvgUyk8F35UkYiTVWW+xkdsjPrG6C7GBGvvynop9gBK9xQd/dQQUx6XsHW/tCVGnHM5Y
5Xr5GRU2gzSCAL/DUOtEHE+UX7dJ7Ir9gbMsWRNj/HCXWSQqRkHbQsMfsDxxi6xDVElsLJaWfPdh
DmpzOwL5r3nihyTkpTTkodMivdcpTKRTG/+SS49cuUd9/4m2d+1rYH7UIVwi5+iAszoPt2OUE96q
4zchF7offBaQgor1GWDKuPJ13Lo7/1pk3GQc64sx4aYbuc3WzrKayDAF8dy+2GwnnUsW0t4snX6h
3BHtT+ypKsqnnf06wFgDFy0ZuZ+QViV+UzfBI/6vNCLMKtSTAgchRf4jsCw5r9veCk1ub1PHREFT
Fpobx0XtpTFH/63J6D/RPFOxO5X9V4dgJ4EEAeC9U+e7XIp44HV9py+ynwi685vjhp9xbAl2KYnW
85rXFhZEuiB9as5UUUCoFStFGDGVl+KcgpFA+PUZoMbVV0fEk/V6OgKzrknCCZd0YaXz4puIc9VV
ZSkYoO3iJdsL+6rXshoKBHXveP3tSWaTuCK2q8RzOAEJjQTAnFnq6rKEiupCKheMhT9GCUr2RzDc
0eX0HiHSj/FSuFMFvCm7wl1yQCzNLxLf1EhVHguMyX9kDb5vLaaaSuiM8FHKwYsteAnoD87h487O
pGFxYLGyuq8cMoqEZj4Qp/O6MZz1DHJewceDH4sf1os40CnPCCXFkvL27AweG5VEpBNqUTEehnIu
Jw/45X5wV9gSZyGmpBjPiDYq8JCSURRqINWNhzOUkcVpETXbX2xCCgUwWczRElipQFCaeoPmovDo
qQXgCOwd1d+Wh5OIWGmfd+1dIuxrs0JTH7qn/JbvtYEolsRIz7pCx5TVl6P8nWmXdVaieENgdlpg
4nyfexmG8aBBbzabCkPgV00+y2/cBmNPG021bjsoCgq9JFe2g7U/0Zd2n+G+nOIt0wYCxe2V6wXx
ELirk6Eu7580XHh79zGIPZlESVDsDxMDvN2md80zwNkxIHgOkhZgCt/GodZKIFK+81mvVg13tOvt
EhzCZ4zOha4R65Mu2NOFDGxLBaaDI8YpYwHIsdCUIAu8pLU1SQTjAEbVINixlCZNtdnn/MnE42Ko
ZJTRofynRTgaLGZqW3QLLY+tG+B/kJdhYnXTWzwDmPXzFvtfhL5j3HQ15nrQCqfK1TIsCIBZTYBN
s5zGHh008VwtypYeIcIvuMkYiDEbOSB58PIt/s//I8z0ClV/8Eum9T0uqoCDTODwilbBX9Cuwd1I
fspn53s3L29QgamMwlsd7O0ChuFX11NtEOEe7Lh2XHivuKUJzFra4Kz5Ev3a5QVazId5mCVOPEbz
au7JxBacU6zcTGMkAyJOgQG0JF8IfCfYiQAauaTjJ23WNHDOgydR7IlFzKKg9pHrn7IGtr9gnEaT
j98MZHpIUhFSQYfaQsYz3L+BhwT/ByvrSXG0rFjJPouSpOZ8+gjOvpj3DbH/zTlNGCUWqZnQ45dw
YQAQEbJVKDd2SDooc++hpQLL8YT32MlZIi+t9EA+aWUEHyfJqT5MrJEAjWbJOYqxH1p6twV2JWgj
j3jSWRVP/5NA8oHYXBy3pjXJyeMiT/Y72eGHMhAeIY+iEHGIffuQnO9RQxngEpYKRN7BjSfDkZGY
AZeUHb2aWS1nbnabdoGb2gkJ9oMs4V5LLXn1whEg9L/FXeDMoqVAEtbnQMOmItU+Wh81ni2ia3HS
HEO3J/MhyZI/jzy8cC6n3xs8ToDWkczkEEcAJ/92Mu2uH4MEnwGpPEMFucm3keJrPk3w45taLeMU
4F2cz7+mQsE8SnyzYuHOcNmvX/X18YjE0ImePu/OwzoZsfKqIhdSEC/nRBArNkIpXf54dkvH9zUb
0nSRUXvAGs0Rh2YewLSW8TmHDwRbFZHKNt3DNUdmH1Gru+lMk+DQ7KzWKojUByu3nspgH15Ro0H+
vkUbUNmO9FUPGngJbqzxUkFjqO0t1jTwy4R2iKis4k4KuIPAWYzChJwj3QsHOhdl8MF8hz7kdRoa
tmdlz5C+u2ucBY2o5bBPDSsEb4A47qxK27jXzRnRxQlzYKxTuK4jrAslhwNIyauC3XZR+HCvEpPb
JeHWLNRpcxipeduXiXJVNHER7vc4WwCmNGCzGHXC/lHQtV/DaDo3CfEzvkJaNqQSH+vP5VvRGRBZ
ypu4LYWkiNde3aIA9aet9f34y5qX6+KBqSNBXv7H+O6Y3Z/3p/bOiwyjybg8B3aQmLS+g59Tlm0Z
dUwfLIJjgYEi0mZNAWY4G5PqaGiy1J0zh3WaJ2oQOVbJRf0raPZbzOgDuAP/KzmpLwJUZ7gz/GCs
6jNFsp8Xjcjklav/3JRqFQhxVah3L24K3mFlV/u8SUIT9FNGYNNJzt9mD6A5oITq82DXU/q77xx7
JRe8ZPH/KBuhzbBiu4ieA8mLtu8Lf3z2XquTWWO74JmQUTnDyXp8nzUNrAYsSHEWyxnxOhhtjUEu
rIBQSFNZpLAnDwEf8HFxRxrXmj4xM2fWvc9S8P65JqAZIgS6FnWMC1rtuT8SqirQp8VJWn8ra4EK
OguMUgo8i6kldVIgd0USq0URlboAwxqo85vLObrMrbzZu8VCBQ6lYEM/JOmE1pFJTkoZLFGgkM35
5NAcIKfw6e99nJEP5c/MsoMg2e0ApdKAFZLr5Xp4xQv19PhmIyj3AvijQZSQUB4CalIQYrMz1i6W
ImYUtRkajEX3FMxfV9agm+8pwW1/i4NnRCDVZcCs+t1Fh1KNPvcEU5BzXbPdMM78/zbK2vNKfwSf
DYuJsUjt29BeJfOBCSaUorFqk41KrRTKdSLaQS3eMvw5OYVRUP36VaWNNEFwQjRcHzcKbiFd2rx8
u2s19ukj6D1I3NayZWAgTY6Y4vLr4be+iA/az36KeTmk78c911ksHUrOt47kSNKZyEQ7jQIn9R4R
skSEmBg8a0mttfsZ7Mr/RZYAqRAUR37Q4wiFnJR8XUfl8/LMGhsFCqT60mUT2Cv24u58ioWVTBM+
NSVOKMJ++Lh4akFB61LDx6MAwsBLTtVvb76baEh8eIfuF1h6Z41/jKLnmoWqtBHEkS8R2OL606/V
kN0sMc50vpJGERLA5wjiJljs0RJr7xa4QFS7zw7ZYHFzm/Fu2HAgfIK2SIxxbYGRtEhgwkRhn0Ay
fTFd5wdcbc3oG0mVgh9JJmR38TXH6B9axdQ1Hy/7Q4TbSY77ZQTaTrD46nqKGuY6lEWFdXiA1EdC
nFVRTZ60WSHoZDg/zlUY+65+OxH469dvL/Z7Oz/qdygaFfvY6+vRDZh81hNLmhib8ymk0h5dwN1a
ekuDqPUjEO5ALRv/52+AyuX+0/luqCnDFpHMY4gWKenWUAxZAfrV6txRNTNjUvVL3Cz+TAzfudAl
RJEh+NsWn3Ar0ngSpTtye9ca331fIhRzceTUdcOgtzUeNIz/rjKhFSvJ6otmr5jSaTBj7maFJx6t
6AOQuwAGr3/rMFFF7FtqfnkDRCQ030ZkqIOT8jj9gFRzBoBGcWhzfO5dgomtyHteyoU/mvS0g+cZ
ItUQxgrwMI7vupR4tF8wXIc7+dfn7yx48+Jom1jcXtYOrshpH/jkL2rF8/UL+cHhpCUUfs6ZtlOh
XFIUk3ucWePH+Ps/DAHqgtJY+6rlTHesgqbqs1cW9sU/w19aOBaAW29VbANl93BYIhGuU05vleDT
/MWuUbfF8i2uMDhiWTZ/fG9H5qMeJTYWoDFT0ItD/lhWxAjme9wZ+gxQieutR3nNfa3aavvryV5w
WPEZeKt2kLGilZC22h8NhTMksDti5WPBcDqTOlrrEXFi1l3ZAPSANMVxODGB/14zFgfrYJYXDvTr
YoDT+2HWDXCr5TyZErIF9KZVnO8krN+/XM5pndD8Uub8PHhHZ9qpuG0OmzmoifM5VC4VtxkzS+Cj
yU1gIUFzn0QTyMVIWtkyQyNkrKO4Ztq8sWPth5r2/OKI5TxBB9FiN+QaS9whRO+OIXeeaTqmBiUk
dN7vh6e5IoVFcJ2K4BkAqfs6WbeGWXIZWHvCh6atAxnVcM3Iw17Bd8KQhqKE7dLwNx+HLhp1pi7N
cvctATTTWkTR33oG6sweCj6y+2p+jqjEUalMD07hCVmXhVypuvOW0SZzDCF6KjJL+mIjmN0qiwce
HbnxplaV8RcH7xDVL1Hr6IM3rrwYwqPGZhjF8+VMeTqZNDPjvUN4tQG8p2HPzOHVWiOn76JmBciL
MC3D/7L46CVBSe96zDKQUldkzwAtFVAB2AFFT5X32qGqakKtcb/2UhmK0/WfH5IFK6D+bjFs6SZH
+cZNMKoFdxTLJy3Bl3aKabxk8iQMSVARwa48hbUR0D0PXn+uz+Wwu64gKVENJzPtRBX1XyO6nb4/
hxuls0/w4Zdg0aosfPT52m4cJntG61UnfRkRyq4l0BLjNLrn4auaX7s1g12u55WmWkK0al+oxTN5
zG0nMGs3QBMHnZgkvYQABCPU3L9K20mDmR67RvN2kB22BlvQrcJhHw5JXOMteIo1y5BTB59/sf1V
Za5NcwryE8MVUzQN8ccU2Jlqnx1gQ21AgAcJ/nJqJaepaQa+ipcyJgPTOskbKC4CjXE83sXmXWrX
B+on3WUsAt4tQ8qbJbmjiou/VKUekHeY1nJeECKg9gBR6uiRX8hqNHUWzNljhYYrPXjjNkeYSmwl
Zwdbss0pIRgnJxNZTJhsPpLQYJIBKPL3fKZq243f+/HbSYhWy+ix21uXPTkdXih6bs46Wy0EleOH
1DcUfI7iJW/dU+jdWDHlXkIHtVVM0e04oeDPpNaL81u5TC4M2pWsN2hRLBinPk2IQUD2cZoPV+Mj
dLkZFk4Ez3LJPywa9hF+A/lPKtI0Nnl6CsCCGi0F1vsPZmrpmJz+Donzjitz17PCPqaqzdbnqK3g
1ioOyKdHgmgB+geex/c7wczqMwg8jfXO2+g+pU0fSMLgx6L9nZmGwZgEyoN9ZnjLLir7lbsZ4poH
S9xiZg/yQ6Z5Lud1lMuV40kAnxNjfGLAJ+R6q2w32AX9qWJVLjN1zh6GGNFGOSowy3DIuD+OYWfc
kegvlC2KcgcErZA0unSXpj94fgnVqg64IVwv2GiNpWOll6uA9I+H8m0YufB6T/yMraMmzlPJ/4dK
GwwGa4F7lw5L/sby+qOAPGyJ7TlFPC0/oRUGUOGzSt6tWvZqgcd7O4mOqQi27S9DoDS+nCzzcnJM
Lv0HBW6CqwlLNysaY4SOY+6xJrz8CtD5Uol3byDnLM3Ic1K9n3+8AJ+CZtEptXGgh9kCGbY/7E2J
heJdcFN5mpRsMKFbnIncS7exn+o0xls9EeyZlDkVpcFLz4JjtE4gHgt3h4DaEgFvgfGElv7686Ue
NRSAoNO6yqal+k5I/LxjvZhli/gU6oLpyGD93K2FtKQIBnEts60KnKmVG0Hzaf6z07o6Uwn8zjMz
iheOmfGvrp22yklRsS2jYYc0cl25Nz4AyqqYBg4ejOwRkQl1lp3mrgz1/6c2uNdwr7YpVouD1cJo
ux80t57aCMRBpLI6Q466pbLA+Ti18iKQ5L8Bpf2itvBF0RQy+rDRr2e8dwNDWI8mg8znz+tYHeY0
ucDrZVYVfrfzahyY8ppIpdv8qIuwgFmd/i/HhWIUyjaCTQC9IQNvx32quvp656oA8KYgvD+cfQPB
201gBDwUr5C/mzZnfI0AgEQZ3aM1dkL1ryQVeORy8Sbbp24PmzGTesojRSnWUmTOGkVfqXxOkwgZ
pYC11EfCgNJFekAcryAjrTAt7x2YMuB/uAeqkvgjktdgzviAqxDy7G5rFzsXfNMFy2ef1KVDhKxU
qnroFigBeXHc2/CKZgslDdeEER+2hh3cTFGurfhtNQPqeKKU1z0HDA7tbeNcprwnOeJGFwH12vMU
6gzAOsme2EICcljhWoIJmaEQxCZKedBqJEjmJ5BZnS1YfvrUMzRJvzslo0sdL/KoRxu/4YgtasGb
LdSuV0AQqdQezi9BGVo37DghsHnRGrM0yeb1xcoOKl2RCfQWquYHHDmssrSAZ3b5tX0i8X+jJQpD
axPYunFlPRf33wM26STeWkuQ17pSKJDpw2uks22KP8MSGzHoA0jvc/+feIOWLoXitSy2xIimIyEt
WKfewYeWEMCniQ1iicP7DRwnGN5VD0SLbUrTiUQfYXG8V3MflEOJRSgnONxmeKDdzvnUSCV58puf
lAA81ThHOFjYcIYrDzXynjxIwnV3K1RrVBKtpIgk08W+fVgWhpfKS3S2fUYlVkCXcvuU9zh7q/UA
vnswNBKofBWa/4t5XI7molZsZQF9NHsNdAA5+XW6hW+tuNT8f2jhS3f0fKQ4p6N0BYG12tVwMHRp
1b77psxp02Khd6bbVaWZR5b6TqmEgQkpfPpK+p/DBlFMq+L4yQm6dxR7XQHoep7YFa9MywDgnrp9
jvAqyrr9DQqyEar1SoMu57r+K9KG/xBD7O9ovfBB+rz/jl+QY+eFZNZegF96XoOQd5CuoWmXqDKU
udBOP6bPk4F/fJUfy3KV68Rpq5x12HZf0ZyN8YUIjvatAMw6hcbl9DJ3fTb9+FjRVPzafprpBs8P
vLtW1OxvNjlUxOp8MBQ8Xn8PyoRhKUyphQd2JbZFNaTeO0RzSDYg3YwV96ntdK/dVajWqDpvJL0T
Z+S023xM/qnX/X1qprha9N0gXe0mR8G1gB39412TIwl/DGnbTSGQKatRgmD4IYoy37D8bOS8mgIq
6e8DWj5GqnaZf07yvCvAHUTMPMZWxBfPcT3iaorq38CI9eWA1jyAsiTJr3KqsiKH38wY7wbvXwOD
ZrN4RSYln8UF78qgbzaR7jEkfpMivyMhYHjEySk701Yu6vec9K4iroN52iH3Y2/xYVMVw8d4SzRO
U4UBijYP+Ub/HfFFT3rr0wf9wtd0k30x7QzmXFc24C1L9Oi7tcZ6gA1A+2RpxO0269aM2na9ZLwj
/drO9n1DNnV1/TwXJbxE630MW+Z+7heVq8AMRluP/iwg+LbP33niV3uzXkYlv4GlpzqrcZQIYrWT
LvzPTwO6LulFCKvlajNnITsEmQqE2qe4QdlEz14r9sb8TtMZJGP0LuiQl7aVew+spSX/Rqt56gGW
87UHJZtNw6Z3h487YCSCyaq+mJx+al9DYtiQ9hrkbMnaJGkciHs5PxNA8WkIpNXklJ6rl9NOD75d
ySBz1Xa0uSzuy+xQnynQ3Oja0L4/dGTJc7LhWsnrzdDM3CaT3oz9j2QPZD9YzTZkz9adl1/cCWUJ
QLjv8tx3dLN0fO8v5LYO4jx6gx6e/IBKqbMOVjoRQ10vWs9m2PzW3fR4BSDmFGty6eKeVWuNLLKd
oTOasM4GXDBLPZrfL0TN+BXXx39unpQ139Dvec402zsxGH0/wXqYAoBBxwhzLFuluXHqfTvex9TL
R4H0N2oV7ZP8atiZZpMjfaBZMxVtUNCZVBldNTc6DCKO3Mprc4mFOZ2GeAU8s0vopCC8Is71i68M
KwAAM3ObV2cK1t2fIglGyNjpCqEB9fM5dPovKMls9+gvzFgWAlUsj0aErhoe6ZisLodWkerXfnuV
JvHwlbnygGp+uluEa2bNQLWTVavGkbCrzpNTDBpdB2AmuMjPULFK5v5U6x8oV/q9YBx2dIwvSBT6
EdpFgXlIJkDJIwFvRSQoBjyGrLv52hoJuZKElDwWIAALEJ0DlD4JzhyRXqrah3HlF8zyfOZUeEYZ
8ZuKChGU2t7oAtyjKGaTJ6DVGznkd/r1S+pHVTujQ8hf1FDKIHFpllfl8YuiDTqgVFxIkmm9OsWX
PXHHiE0OG6i6GcLZN2Uus28jGqGzwRqMDfZFi8MS4saZQ9s8G/j1oOz3F7imppSxjOWpYg0ZhrlA
MtS5E+rtEqsHQYvclrR91Po6FL003V39Q5KSTw4JLha16Ohm6umR8o0UA6wu9/z5GqUbT7aXuKq7
K3bN+fwovqF22dEbTUb0z7Q/m8vPEQ78W04jQ0Ejbkp8dtGVw+rxxu/HMw4bVXLLtoBUtbA81aL4
5kKj85ftRPBS4j92GpkQ+TVQQPbdtZyw5ciWAea7UkqGPC/2oHtfv49joyvHI/Z+shilx9ND2ggL
5y06AShliMSQmmNocVsI+goXQm95Q/oS8PqjEyY/1wKMu5GVpaKyKYMGHXclGrmO1a/of//suP9K
0rBOXASHfXQ/PV0W6pUeNhCrJgm8gNOBBCSNTLPT9i7KoSLeQ/z7BYvGi6P503a27kExf8fYfYZh
H4I1XMe8822Z1h6L86IhUTfbYTiwccd+VzlSV+2kKWTbkMa473gdv5MpAMRCx0gWFofaVgsYbfXi
m7fCVg42rotPyC7ems+iux2VvyIofmEBMirJLcXqbU0jVF8AaS5YHjJTSPC3bhpvSNSu+9NiGUWD
sNoA8ME84xpn9zzhg0jg293eU/HAAjnDTvoDriNOzmWgXRVvpOLglZBqoi6kYHriuxcfNM3gCxyG
VJHXUjJlCd4/09+zjwQr7OZtgo0j90mbG/BrcMzAyl9jksKhE4/wRy7z2m5fc15DE/DPH4qELg3I
YGiLEp8rLCSRswRQ/GnTNDcqMSdPmML/pgyAxHvls1p7vhwD2j/MXlq5QIUVCzWoKizx0arXNb2k
qnlkQfMDrsuYm5O5UPVogtG6CC1mNslivCKzt38o8O5QSRuQq/cUqsppQdACsHMCmENZfOWkRmuN
3TS/T+CwkVjxpZLuUtRsiIBWtk+nwkQ6JnKU2GFp2MG+GW8KBL/m179fX8Dz0ur+qxJkMpcvhK4Y
8mzaa1Y/eG3j9Ip0Vv4UzKbSxbQFMI0A8HibW+atI3X/WSjFTgzvBmysRDH/hatl2dUACg9qmj4L
aCNGM1c9ZUnseScuOB1LzkyNgyJE2rPsnvEtRcxVrV0NzLKH8UV4lDorsNiy0wYIIDKxI7UCwtmK
7lrDblxAl3NZS7Uw06MFG7FlgsRZOqR9y/7ae6tnQ+cUwiRyV4ZqcPv/6ImXxSSC7/T3Bs992pDi
TCaxn14VEOeVgtR6uQX3jnH7dqX6AFETYSFX2m2Jhsro3LNOHw06wTqYwWOsCM8i5AII+kgssUJ+
f2hbRyEv/dNmkd2Kfx/UpD25v6b+mTr7UaHQTShkCNUQ/5LidxUCGIYphVofbXzp4a6rqyk0e/AE
AW5atDugtNIW9UphwLjtQJEEvVIqqt96PcwOLjcpwZQCHE1aBLKto2xOmw6KO6xQyk9E/6jd/u3T
tgywKpD6eiIX5TagVdKJRsmdIOBlHIRUUHHTKjyE25mcKzWNF9XqZSR9wfE8NC1wE3fuTEgKrLQ6
IM2Dp84S1JpwYFaVbDqM6vHv56lCaFt0WF0fNE2ZdkiOAHl/qxxWfpV93D/76+HMqu0V7Ng8OV+O
VsCcy6tXAzIRvE566k1AHu9gNA2+geWjzvi7eKTIZzSGxwAikrSCnK3+UrgOluRs44TfIeBm5LPd
CAYXOBwTYj/pUHI316ZnTde4T52AltpFzcruvSEhgueBiYl8wLrFjNksMA/eOV2jVLF8fDWGQ6fc
DCVAiyvoTsz1LbmCrcAQvYaPZ3jtywdHOR+32JztgaF28z1gfCLL0rwRChxdZ6D8QQejA01MZ9SX
ULB5s9JY74nzecFjfc/Ny3HkqZae8rjlelEQEdBiTBTof2G1Is9fEG77LjPRPpy8guBJkuGXtSM3
GaJZQ1+Czhq/f3z1Ovb4BZYvBLuk6FWn9KVUcEf4SpPdMRPxVFoaz89gf3sPpitxTD+GcV+Od9vN
rjnCeTNTfpWEdgAjro7NVgAZkfc/wrb7Mh1bSw1ylOee/O6M36VwMVuHH757a9Cl4Sj9RyPnHVjJ
ae3kmniaRkj2w/f7XAAxGomj31npNUfCwZinDmETXGT5Sv4JEl5k7TVp1NxMDMPGffvjllj+YRSY
8PW+HGzI1EHiKHpnryMiwpdfvMW9WHIcJ6SoPaTBSpFYj5E+Gd8EB+ceUf3ttxnxbsJW4m1rO2Bs
CQw9AMM391pKwfIvtMd3Z6nsPEQ3NqM+kckYu8E80tMsN6xyznOy9li/cscxuEjapYua0aDaQA3t
BG8JAvfJwPwr9V0Guy6ckbD467IeGcpXHxd2qe0QL0iD2O+PNG4Wy3gta184llu/PVCpZSQaODhC
I5YLmGucs5OkmzMbw+ZxATx/8cP/PYVhG9iWXdo5oMc9Q2Q21LwXRXDLaaJiPOtjCJBulhtpvG/k
Ii8H4f9L+yGnvfxOUod+5ny5zBqOQ2nEsF+6dDw7XBROEpIRhpEwGcjslRypMW9Twg5GjR2RrTkJ
ylQmbycTmCjV57pQRsT2mfpwNSmZSLuh0Jvll0vZCp/SCXvM/fHhNX40v/d6ji4x9+W7GLkm1Zvc
oWQ0KrD6VOmymEGwTn+twI1WBfhC4i3ilgpTurPTeX4kwVTqejGaV27A7jP/60X4/e+zD4QuBlh7
cykyCvsdQkddEDpmcvFxxqqviaKGWB5Gz+7u1k45QIjICFXWXsW6rr7WvY+SUs1WmDOvGP2W9pTD
MrZPnfEw+S853/LBJ79uj7BwkY5jA8f528SRZBznt6qp30MpcVPF2R97q+dt0ik63QgLiqwTD2kC
ih0DHX6VC0gQsyN+Br3e8YjYlHmD0RNabt0gl25WW9UIZ6UhXdSofKGfALQGHlTHZ7yVVMKdIQEV
7012VBwR7USNG0m/em7H2f8WkXU46BExYzKqni4VOm/oct7rIxoo/bjlqm66DRqsxq6rbpirh2fg
mN2V2qznCEcg0KADmhTonsan3g88M/XBJW+0mClqrAQXJNACJoa45g9Hzsvt/uS3MqD2ifw6/U0M
4gIzYQEbC9Ghf5bo3hfohsZUqU1YvI1jeb+so57O/TWvzArJ+XUn1D14Use6blGHx64apHXAA8J0
7qakjaHhVteft1cdXKv50ybvaRxDLNieA/ekrQVISm+OjtyQ/x6sBqOhRqjb2hggd2IecFpDoI2n
oVlg2/2RscAwA26mdeyf/6fty3IyxwL4RznSCJqghHVhp0QTOdGN45CURtYZLG+bw5jT3opNdB1z
Oq6C4ZIM9iNJlzKtLsJDGQ9ThtLLvxSVAdzgyrfGWU+PZHPnxW/slWsxEBup4CXKPtoHsrTrs6IO
RClXB/W4oLxDXzLAvAoy0+0860B4idali5nxiwB8KoHfUF+oUMqY3ot7jgm2YPAcYuSreSD7esj9
Gumdw60ARkwQXx21df2JQr5IY5hAqR5jZk7qfKtpUxtWZUTl3JYEhidEs79rWssPlBYR0ICwfSk0
wfDVYFkGvngjZZNJjvCQ4lDsQXv0+2UgoslcOJgnxoljys8BA8QPG11Fr7tPI2WIemZ9zrRwtmNa
8k/Phb1sIGzqPQ1eEaFdOqyIvgmtol8LJYvk4hqmC5N4rSZq6OKJW/UwOUwJlMJTwWwVw7yTNQOu
LC6t3nRu1EfVrZHz4a704vCHew2lAvTcFl6aA6M43WoeyKYkRlDcxcj0s3i+8g5qxsz0Vi4oqzvu
FlYql/k2vApNbr4adi7LjvYioRRQWXMMlWH81JEySZr2BJtb8DIvZqx6R6dwTJcba7bpjdqWTy5F
yC1TVmrXFrjm/0RkgO1rVaUGg2tdkTgsBgGbw5ft+bg/dw0xnBkr8NapSr3BTZ3vso9vcoiPFO5A
qKX9FJN3CQRD1uN1VzePMlh+JB7HHRewQzUs9SAmq3T9nHFxJnEdqGg3i1XxkSFbrKIDuSbKfv2C
q6t/v09tBOyaatULoHzRtJ/fRqdi6bFLcFdygavKupKDwTL8gg7+OENe3B55uUrcoPNviPniolyT
OMR/GW5b63A4BrL3RB55gfjPdNy79iB2rhZmpgrRd5CC/tPt6h9EQc/pd9QV3WOvEhJRN/BjM86I
rXxGqjz1p4wXg59MvV5mOpOuAYE/TUgB3VM7OGXjVaJ8NVHRQDQ7Is1XrggBhiwBk5LfePwSrtps
2Oa4x8wJ2+1D1keGXkKcfcxYzIjk9lC3E28pejLFvukWsNubhGPx1D1Kz23sg/OnFYKY1t/9nWV8
eYofAcebk8H/fg8xUhrH7tlSNQfXQCwnHIASmPi1JMhmU7AVSwB8E46fh6ail7sRp9w4lcG3HKru
7BvgcHWuHG5n5Xxt2xnsLDKikePRAKR+o/Ns417f6gkxeJAxTl346ieJTQfZ73U+H1UtxL62djOZ
IhBzDqhwQ+Sye1/3sFxqdtaKMghZz9qu1wFiC8M9kzzWF3naMetXzPnzvJXwkANPaQGwG8NIyXfe
BIRC1jxVcCX2c57vBvF0Y7Wvk4X1yrO1xwIhNz2VFkBAxfKFUknR4vK3Fyu+ipEPGyvDzSUEIvi+
+X5RA4/pbGS9dCpE7IqnLGpWlbqbRrtwMNt8oEk5uuauByRH0mrq8Botbf1CoIvIxKoDsXtTrOHF
nkrScJ18b+EtgUHZYxvw4a6ck8n3wk+dmUlj8yfWhQVi29Sb5dpzMxqXuzQle7bBZr/CJNaoGYrq
DAeq4w81VKD1Umo/d8D12BRVbpIFdzfDpJANqKkRPQB89Jre8QYrgC2J7f0rnOGNMZ4etXbcQSnV
dAV0Jbn8xz3DKbYWunJX6JIj3rlPRa1px6JtuLjy7cWlbIC641DJtCcgYgPqAYozQ2V5o9wdIlyO
x41vOsIfpr5uaqB1vdMGdx1ikSKWoz9BZnGRj4MJZqW98raPf8rNLFBFD7yLl1NyLiDEuYq+DlRW
43ALkb0HBEVbPo/ov0kAfmOsh8DjgsIdNy0TlNIIj6yMFRCrrk5jiuGZlDBmtJo8eEnPukzI3b5i
lwNvBqXeXTK9EROW5L0Wap24jSL0uJQHjQXUk1apNPTvc2gIF4zcKhNTfflrjDloGMY4BXfJmGBd
6pDwQBwDKo4qdcJh2E8EUwJlIYr2JoEpQvcFa8ONJ1CrA1MKg5V8dJW8Zd6B/SQJIW0naB8j1FXo
yzyAdeMI9Jh+CM61ikSqPb+1NvZY/2WaQm4q9uTDNcK1f6hDpM19647qmMFNncI0qFIMp0veSm0B
MNQtWr9dl4qcqeXH2MZ3Qbqu4FFiWJUCqI4NRzv7/b32UkhKXLPR6G/Zgoe/f7+OELAqAvs5iNGf
xkpFIN3KiowsVb2y+vF7lfvtzBtOni9tSJ2zvl9JvcxCx9mQ0OX81Oee1D1dO6I4Lejq8F0QXFq5
//wkONUtxoRER455kISFQyCJQNHvNlUOVRRSJ2mXZb0D8rIpOlD6dvkYQu+dPcBMhnGnB0x7kMI7
tcvoPLA1ZWTAoyNfYxMb9KUwkjSlx0VNUxoXhYnjJYSK7fddT68ZqZl2qtS6l3TThpQIgGsBbWYM
tzDrEDki78igIK/CIfP05YLgKlk/NgzoRJdfWsrgGx8tZRmyo5Z48iBw90itMDEqYxQIh+FKthcT
ZWj3+SI+YjLg+AMqCF0G2CLZcsBps+R7UUpESY0FTRvp+DkUajfyuRnvrCGnnKLy6oJjrPnU0/Cj
e1ZnEEaq+QPUGDbRgz1b+oeuTQ0SAis4sXK0aDeH3snV5LM7UwIKXbwPcWy472b9Betp+CDHE57M
gU39pABbtXPHW1FlLYLCXeKTl/7l0GxAaTJ4ujH2gxnOXU1ujTsqAiijt7wFdJc0/a994bwWNAFb
4ncmWnsl8sdQNJeXgOnnOqxuRnfS8M63tc0IGGz+HzDHTJln5nRLjRg+J9gqAxaFIdom7+yX3gk5
hU7N9TLatlmAiMmGjPU5yhWir0Li9IoGJaBZXt1loSa9w8D4qHAgQCMLkgrLYGt30uDhmUoleIIa
8XICYtvw7ReB5CQuH4iwHJxv825XJUF0xl080b0SsL0twOtyHI1vStP4g3pMxlaZBNLvx7ahCSE4
EyiZykRl4aV5MFYkQCEa/fy9GhbzE9UJ16B0S+jjnWuuvM1QisZsbRpuRDNgvBhj1iBTyLHW1ngW
ETgbH+/E5wQwGQO+Qm/LUBYBobmxLe50gTF5riK3Np3mJ23lzM76JlUugJtphtjKVnAEfHBuB3zc
jcPNBIPfNBaw9hbg1eps4m7HARboLStoVkfoiLCAK8VR3m5qScqGBVWoZxgSpHh+YL1YywtwsvtG
7KQ73Q9PQtzZJs5oecZpRRz/ymDZ77WeCzQIQOzcm7HoshseNhhgYeBSZDKt0IfcgmwqY6Kivykg
vLobZI8NTuLTaILbYwSUaHxSVJ97bAsTPFCfM9qCwS6X8eI6C0+p+cgqBwxSq90B+f+QWTuOqNUK
/B0DuSxmwqSYc++kgK++HPlmqJ1nzKzIegJWlm9ndg7RbeXtVGWlmzdRdQ8Qdc6gh0XLltJiy0N8
EmxDwtGEV1vt/4hudCcWk/R84tqXpXDaYXYjHCEC6jlhJN2Hzb4aYUVW3NxyUEMJeP64DIGlxR0i
dBGThrsUp4dKAettLYgeWjkGKcFtJM7BbsDDlb5YGGJanjOg5k+f9oNB/JxMwFwAnM09lK2uMFpv
XdKqeDPy9hOA358ciqEur8sDnZDcKDLqUgZ5CrzpzI0GoKFejwC/trTsUDsSwtSOpcKowMHP6ONa
SO3fx5nn8L3d1g0os2XFmsXMQGdrXkZ9NApLQ9fJpJxYi20m35i3SM1GDO0zVoOnWc+4MUxTt9nK
q9mRuh4ADiQOoBYomewdzu23c49li6/VoKczfQl1oNBQbrX2xCkSC8COIy/CLkeK0pV9veAvzBpP
e5v5jvPfbR2h4BZHij4cRsYJPCRnBVThFyHXUxVvOJDDOfHLse589TpD2MCpAlMJZ12wrJTyIbMD
xbdBEDghSVicbIiO8DnEtsxFO9qfObUv1TLixPizHQidImgZ9EZ+zHjLOQJ7NZSZgYfrLBUOME3u
YLHrY30qaJJZbcdSEKQUOVem92lxPE/sybEnu70T1T14K8ZIfkvVg4D9JF+ww4wykAIqo9WJexlf
m9QYwCEmzZBUNLbFUnhCfqm63ipEbjVxOJmkoFVO7mjYDcH9gBs3ObfU0TVABwwuA0Us1Xz5VwSM
HwiRjRlBuySwgA2qyoXroavRhFmVF8ilc7fk55tT8RdDY8zWMx8pboutJDPRvSdEwyQSAfsbRePn
RL09cflYDuSZW7VTJoKySE69WJHaJCnnZNcroiCUfSbKgpHXlHVZ0h4Gi7bIpyQIMpeCFDDHiCFx
0qS8DjtBHbhPmUMjcVzvJz7brKBc7P7k4Ny8eGo+l8iENo7oGbvhkCJla2ECrLdV+ncleOZYyMtM
XSkRzRoeWDO1NMcPGcEprXkKYzysN3w2NbjA58QS1TPR/QIqxXmHjTQQ6vkeQSBqAl5+Uv5N2Sc6
fe8jn6dpTfWCGF3XMbnd4wGrJnTuM3wk4MVCIxCekbZ56CKVE/A5/Wu4kLLmcibfirq8rSeanKAD
LCdqPFL4Ytj3I8unXa1tdQDIqqZTbFG+epjeT0H65GfdhJUpL9mfUrMuJFcFJyFFGSvMn5I2HMLI
At2HYQBYLuqg+IXunFPlzphf3NGqMylJjvy04qH7E5T54WsDbeE6BGgVG4ZoPVvI8AblfQ5vRUKj
5dB2wvYKlAg4WKAfUi5MD5FxVY62JFp2COTkBImVH+M/88+IDf2ZHN7kKXQd4Xzr/8PWMtV+dI5k
KiVEFrdew2GIHnvnFllfS1Gv8y5ZCmv16GO1lb4P4eez/Tg6Y2PclX9UiUqvb8uCwKMFNhE2tRtX
UAeHCUXgvqqiCdCeqP/iAtf5/sjOXrh+qxW9bn4hRP8dZiWU9Hp0BEAalaGin2/Vk/CUKy/KPjmE
XEV5tty4lb8uPMbYeOBDFEzWfHYMgglJa987LqHbFCXxqDdeE8Np3yb9uVOxPlrqo5b8j32UFDdy
J10O9uK+0/AqtT/n9E8UUAkekys6ScXdgxMr54b3oKC0hQGyA2gREckaQEN7YsBlnX2sNEwZKO5N
+qjWiIyNP6kGPefKaNT9oxuvOSuzQVw3Fm4QHnSQRMzhlm7sjB8eP80Na2K/rLfoG+A/ZO+ongCM
a25H8WoGVBYTYq1kCH5S0HIY3iyEbvdx+YsceO0JYXBWlQXSqnQM9qytiQ1yiSzb/V5VuOhvaLA/
vqgM3W6ZJmGS1eYAdBmShSXdZPX2BXBtNXI0ioOf+9chXKPw6lVZSDYXi3E34j2Ahz642hQDV+nP
p6S7kAnBnfW9F07AGJ+uqpNz2oKSOfGU/ANwJ5xMw+RXXsZCcSLjxgY4i5lKb7WjI6S6EamgejUu
aQRcuB7+baAdO7FMRI80mnsQg8hmdDU7z+x7bLruGBZJC54GvkMT4+FoW/BHX6vcXTvLVWz5ruMU
PevUL1vDILBYXokVz66yniSOqlO9PB6hY8lv78e9VnfckuBSsZu00tuk+Uit5WJ1akQ2XUUlnM1o
bIRY/+H9MK1K/U14Tx1gEgl09lZyiLqXselmV/83lSbj6KTIo/UUZsI49kXQhheoxHus733sEYbM
JfyNYCmkNDRJz+Ggno8neeJHSRcNYF7Cz7V2MZ6brcojYZh4+nrXa170C8CgaUfYupTzKplYdChG
7mSVTbwFn1vyQS3YlChqZKaw8WbmUwVI2Kl3rmvBugH60wnw01qlx8PC1R+BnUNyC0o73ImOwqpI
3TKJOkNY0pKUOSP/LIZ307iYFvHSyP6ePwsecpoTWSEgfn5hDPzBgPASeJxEnVmrMgvaypFhtNLq
rccJgxwvkCOPPy2roxhGhjYaFl1AkvGTFHAaObRsxVJj28oHnG9n4DA8Lik64GVWOdaExuQRso0D
bTQSolyo0LEPTOi9l18LKl+acgRvzJcZBfM33Mh5k9I7ARiirEkJFGuftBYpTu8Xq17z07q11vsh
vwxD2mXnl7rMDL2QjcZuLX7tGOpoQPw6H2ykcL8me0B3CHRl9uyxBMlbZclEFUhexxgcnaSbH5b4
NKlQCv3xoJr8blQzyvewJa4qp5SjVHexIUS2rx1XApRSqoMhxEJET49ATojD/pqleEQPR+GoWp0+
Xaqc0i/+ke2LorlTGcWW6IU/n9nqBymkgYtN3SWeJTnjhYoUKK3iE5Emsh8RRlyE/F8usauvu4U6
DxESzk4qZHF0LdLgsLPEiMUmvQXKPUYAfivznz8buykNM6Zy5J9n5nV86bnLRBd0Pd04HXtgJ5st
Sz9icvqVVPoHmthUdHhOISOamvU5/ekm4+bspTmcbLrb0GSKqmbppcfk8USmZApXmMzJxNu8Bb+j
4mOavE1DGTJN4+gEyZgWfl5VmWNDCUiI5z6ZMuPom8ki5j5kFXcNMvu+daPQtJLQoUzOZDzTS9vd
Sxy5zHrXXugYQEy3G89FbjacZGW3V/HTWC0TX15WzMJDfkyEsVMNwYO3afeEcRuHleySw5/CxLmc
iINw78WI4govVgF3hk5Vft9JA603xQHt1QTVvhTDQSmJ5dAaaemO3SFKIqmXwH8YjbrGK0MGQLkm
Yguf9csWvZwrLdW+3Dep0inpivhqVNwr2gfOMvV1FSmp2YbDLhyJ9gqFf/IFf2OqB9oHhxwCx+3B
JExJBRm5xRyALIrsfee76gkd4z+YvIv12z85et3YhlCMQM/RE8H+Y07vIwL+da4K5piPgl1WP6r3
wfTTvYOnDa7+UnZAEvRcgNgisV6nuPkm6BF7HWXG0gJdDE7RRMmYAEAPnJVpGdih9OkzzEpgAHNW
tqf9MsTwxhY5g5Qj0NYgsjW9r9fJToFmBRhozdOn+r68rXYuDsggJU2k8iUmE90o9S8vNi6xP7MR
eL2o2K3C2TILwQ3/jucE8w8GsRx+JFp5RCZyjW+4SXJdXdtwvbP5igw1Po7sUsVgAogZjxol1RgJ
JL25vGyzmhW20dAnD/IkG+KtYLlnnhQrG7yjqHy2Dnm6ErTA8IIrkIR0XRAhog6p5dPKmb8OHrnO
iXvU89/LuP6zVOQ02vP1fJ9PpkymBLLoHsn5GHdwLU/48t6PL8WqaZYolT3lXTUldpvtcGD9l/A1
V3vS+I/THQkdLT1xuSg1bVudZljqoNiKSLULnENtOUYqWqZAw2gYpiI8vPAV+4sYhS7jRBFrO9wr
rn78iJ4DB9DCvx1L3kzyFK3MDRcCTNTwl/KmugwlK2LB2ipnw+TNZIa0FiI0B7CwMxjZrTkML+kB
8+m465zEls8hZIXQFJ4593znBWotuNHcotaDvjcuLZX6MWTm4PzkHK6PI0d+C0KoYnEnHPdDa/8L
lcZdmt8zLY0vcSIom9SZtlxpOP69sJzzoEzFKIny9iLXycVkuxrvlFiTawVmuox5UAHgOXPA0h2a
Lhyh7vuhvvAyGEnZ2Zbag5pZwNXwH6gXIP3LetGWFFzs1Rm9wz0+SQ7fpZZMo1U41/769EQEaknI
oc/f4os4hVYYfltKnj7WDZDMjuywothYyxW7srITgbB8zw1QaIU/gVVz6spEKg0/Ib+Yskeyl/aT
fX+QNHJG4RCpzgVoDk9a+2+A4sbuQ5uvMBiqoVQTTeH/HgxUVHuXyOUPUQubFedD93c/9fVIi5pT
eT1ykFzwogWDPFKp7n10FFrfKdxAQVWS8sljNbUn/QSf16aIMdUMn50JtIjqWCkFqYiQywCAMbPB
s/ndJ58Za3dYy6Jb3I698AiKXErqu1VwIUjR2+7HqSEb8G7rcly6ieOOiCjbloTB+AP2KK0Twenn
rBO+QGKsfDlDA089Lcena7LW2LoBJOV1l9+W/oQqvZ265A+tlJ9c7fS2J2XcuC6jNwkG2Di9pKre
7OoDdHE+32pEuGhX9RCRXY3wGBZxnYY8SRiTXPaWHAm6B1WKyU1CO6nW+uCrJwzJrYzgZ8Os5chj
gyS5dNJxoXEWDnhm55C7k2T4WJGFh1VjOGNWukagvh7jHuUKQ0rbD9ejoei7upekjjMBwVWUBR6g
ntW0Mgsw1F2DkxLVJRvbbPDeNZHpfYH38wolrOpoHvkKAdzNi4ZdGUJFGYYkgh9kbogKlKZOVpIB
tFRULqxeRupEdBbMmVtiawFGT462T82icX94UwD+MnEQBRuvrf13tYszSQNhtQ2D7U/PPS4oDsvn
nUBTLNTv0SdLlo+1mCfUDgYodEoHFkdbWb8CFojxGVDupveT/UECwrcw9tlvyF12IW0bg6jIllDN
SQPTHGU+o6STfeMMgVf10wd0vFnM67I5EKW1pZfGyb+gK2dZ/swLcPIZzr4ZvM3aTZ7vFGLUyD41
0/6p1hDB85id4//Pv9ivTppQDi9DeJluIC8JnPQEfde6F9JSr6hDAJQyCwAcNuDYa817T0j/adYn
N9xjXo9SweUJYzHKX20AsjN8wqPMkcHtd/e7kh4C/np5ZssceWjX5wVghbd9vZcYVuELWKhb9vE7
tedITugZLmSu0L3UCtsRSyCra3G/G9zwwYdbjjilLRDjk8tlzMlKG0bTG3YZi2gvw3RW10+I2DV+
X02XrjGE+FF5xhTVEpH/7FeC/aeBYJNMuXzAnnLwHRhVfvuz/iFqUpBBvDMmTFwA/k0MjFDxVW2i
k3MBsuq4f6+NTgmVzDZNEXGzBHMBAMIQuyvjHtXWBqprHRmixQgSpVctln9cNPZEy5Zxjb2gkkBs
ITN3dyTyJXX3IRmRj9MvY5jNI5xs09N8nuNEQY99InNNO8wS4SqkBow48h5d0iJo/FFfiMdOknQF
bWwThJlbe3zZQyr91FnLGYi4nwnfX6Xwq2E+PqkTTiQo/bYpJwiRBujzFmPTpFUG/DJy+jSHxRWn
+ZQyXlf1bgGwlUUfxlGp/IqqxrxJq4QGJmEX0y9DbqW+H8mdq8f+8VmhlN6yTe80AJHWcXu2fTSk
YsrheUJ/2j4I59Ea3X6dm0Pg3jJsmFbQ3sVf1RktSwyAR/mVBZhCaPYPBHKl7jua6lz+w+fvATxI
ia9Ldg5Fg3IFZt4bWSzPOvWuir4ctwajbYBvuI53N1SWfnmqzuVA/4EOu37kNEZS2mlovjzGGb5Y
0CyRw/6ZmzOXu2nBA35X1iyAwWL4liG+goSRedvJEybqQpknTrQ1Bf3Ty9XcqEiHoCj1gxoM4dyF
LQ+wXelZvH4pPlsASdkQ9Z/h/SUjSOIwaQCzMXhLg3W5ZsaAJ3LbSrOWCW7fZoP3lGRqzs8UErMt
qNJwi21IWnNVdPsEKlQDH++BImkqu2VFaoW/FrE1yqgDmQgyofVsI/oYFvpH4LzaKseZVGLubq/C
jHu8tPbQguauNnw7q7flwAcYl8G4+922ZvGIp+se5lXK/qiF0cyi+OnVHp+yaouqNim5qYZv+wYH
HanMMO+wHKt59R3atR0RSXmzylahxCor97FLAMovaKw4gPs/m4d7yM0VQZSNf3XmtgPvzxR5qxIW
6x1Na5/bjI8o8dJbBaYPCmamF8jYoztx9bEiOaZNRk+FfiKhRrNqlOKTpiewDdHv/R9Uiy1KPZmE
6yohuKpXlgrpKdapGV6a40JSIAeSUfsJjhyHczLi5PRIlAEdmQTUIzEiTHj9fWQAWEgPHqx7krYQ
RL6JgsRqNSzoNnB1TY3iQ3/WOdg3f5+Ak7i4yK50HW5Uy2h7LZunY/3ijLisJJOZJqsIaKDmUzyu
gfIyNSxVf4aiC/9CaOFJj5dNbfVQ4d9JvvOSzOr8PzS5em6DSxJSMoSbIs3voiR8zGXXly8mz27q
0Sl2KUw7Lw0N8kqLjNDTCbU6Rvffc43T0lx4afmY1XM+GdGyDCbLLjPoqqJznPmWsW7tPrqcODM+
lJ4z1fOWBNCm9qhOLmGN6oCCvAiTdlBhq5L4MSxxhomy/C7kHvBuhImxBUlgR11xfMeB6ENQJVsJ
GIiGiVBBy+bVRpc2L4kgWcWpjMrzr5V6NSjWD4pR6ud7HA+yPH1u9pr0iUirsv4eCE/6YiDHgaAi
5LnKpy+/67hn/dxIFM0rRa7KVITuw43ziODVKWPWdvrYrAB/i9KEPmB9AF2TU+2Ut1OekIB8pTGf
dc5Rujc2kTGufmIxCYL0yqEdyPf28skHBQB7tvdnGLxjHN/eRaJhkc0z1tYmeFnzBc4YqONqCPiL
mbJi8e7xOjSMSP8OvhGEuvyBAyZv9JR9H+hyPsKWk8nU+nFK2sGGcUXTS/LeOb0kOfRWK70e+VDh
zdL1TzX24nvMdprJJSFBv0nhcljcCSQzK3L7QTiPkRDOlNkCYyrIiRVo4I2Gh8+mWTmklKk5Owdl
82MfSrJ+Z11fLs0+WBq57LrRmWiCa3I9Icx2yJk/6EW7mlvq+IA54xY1Ji94EFRrD4dlOotVLqy+
duYYfKBAB5oj3f3cWcPvavx/JkhThDeqw7cHoDMqXlyoT40x4WMad04c3bDaP3PkiDMzJcJ8r7vR
hEYFMwFfjs1mbWlDi34QSjhat5c0gIYPD/jCgJSrPKwNeK3g+Fv0gAU3Nz2ro3yCT5B8OyiZdAfr
+kouqLOhe/1j9vZ8sYjl/T0DmtIsqUB9+05EEIYgwowpKjdtWW5R3dz+UvqFB/hmKHe+fXhJ6kVL
VDTcfVc8tpQuSEZZNrniv4kbiSPZn55xWOwsoTLVVj1uCjL1mDJOSox956B6Be1ujR1Pdfr8GF4E
oA9I0JID6OlnIbXtZ3O0EcRmyIatqQKV9MgObDSgOPylWfbSn3C1qfgC8CZRMQ8XIdz2BiJJFI5J
vsPhC/cREZFy2o0wtqrbM6h4M8f0AX1zSmUm0aCWBP7QmiEOAGeEPMOzbutu2wcaqKvMNMsRbhpp
0mD5j32ouQGnJLwxNzndoize9ibqiDhinz1mQMeQ2fpxZdIwJsYLmtQsMSmjlmRvH97oI6Bp6BJ2
Ifr350N0qbjdofGGvVy2QRJQlwDiARcteAQrCuJjw7mGpFb/mphM9aplajdydv7qi08bTQUwFCMM
y3jcG/o1/zhkMKOU5bnP0Tia2+0NiX6YySTacdIaJPPM8fltC8ak3Cpj+W+xgUw0QoQGgfNvD12q
7n9GjHZPnRS4RxkYrF6zTQlAJJ1JNU07rEjFwn9+j5juA6VR/xjTkvPbjsQncFlCHDTI2ZoHVL/b
IP53UFpebeQbfH7M/1N/zRneUlaTV2hXhvu6NSxHY/59uRMBpikFYXxRmB4kHAwwGtAoy39SJfA6
ld8HjtpiK6tPYLU3sT/ZPcLZ1YJhWhQmvkI3lNiAAz1WY9wy8u/ZLjpCdmmmPtOrLexssBS47/CX
IV9iw20bKQcTpfTmziavJ1WrGbFfwAUCh5ym8BV1biFtPjMfcMgRzKEE2LvEQG0bkVAI0QbgeAY+
6EepYvv8/egShA9F7BJJPVD1ALZOLxNWFFwqvTkRBGLBG5qtpgrATzrW14ddL8h1DHgf/AOkCV5q
VaYYXv2be2StSUGbshFrJKHf+ERwGCRzwHAcp6T+zi276bibYhS5ULkE0b3TjhOuxjRm8yALMhhO
apE5W/povVUmNVVa0xivG05dtsa4T3kGqxK2ftCBc+uBkAhR2wS4lEYF0KPaRkuAzrjh2ORNBTCd
Jw3r9p6dCnbVDD60HUz8UnWGkvhh9JKdoPiXVzC/TBwRqtJXYkqvy2srCF+d8fJjQ2cvkyZLlvc5
urkoxblt7KJKqGOrNLYRXyArgD2qFn9AlMHV2x3VNdIEb7v/qUhFm2KTLsogU/dd3pK2jEo7YApa
cJx6vFiqHsZ48z6ALPoeS4wJvrg/4/AqhNGlIRsqJdI/QunTUirvA9kTPSMuBRoS15IFTngCmWVF
W4UGjp8qsNSVxJmg+ADX5trbUd/ufwQVesmjAN1DBo94vzlH3mMAkSsduEX4xMY5fMoZEQ9lJ3Bh
vyUNTkLQY6jRBXBQCzQdRCPhbsxg1syHw4Hfu9CMwve55PLYqA39PJn76IbHR3ZcggUwHD450EKp
Wxh8BapSK82rTFvGBV3eW207BVr3CIqyTJZ3zfSNXs5TjkJKp36z1lKoCSuZ8edHbDkf85P4EkoN
t7dhMSlblo0aKfzpq99G1XsLoMMSPfYg6dpjDrw74ZzTjnHvQQoc0rKwgY2i8F45KkumPHuTtqwL
Ewd2gIcGkKHKm3DxSF4cM7uM3ff4tz1o5dF5F/eREsg4s/p1NaKxN+lN+aAayotGeGCzOep4sR2v
CEEOXS1N2gO/D7gTcnAKoey4/C/r3GcmR/zVCmLP3+ZIq8qSqKB+QigmzirMEUzT/oeaBv+4tE4i
lH6yO/PLr6kJmktU75FbBiNzTjTPjVRv96BfZ/mfDbDJgZc7C/BK1Q4m1+ffm4jWtQuIqqk2lh0s
OOH98a5C1KD5xlgDz84EWjtjXb1OHB+jxvksMO1ven/b3TPr4mu5/wrTzI+6oMX/fZBF/uS9hnYr
PtWIVmLarXkjZaflRBnjPNTncYUyTfuJU/y2xrt4UgcSb1ptY8NSUXoOTS3Tm3F2QC8oPwWPiJJY
FYgciQJJ0/Lu1w0HFUN/6yJn3GM0EZPgshN6GMz6xBZjOWx0MaRNifQOlLYh8/9t4z8aCoaBGyru
+G0q7XDfSOwhS6RptJRI3bbKEe2DVBJDcwV8Gqvxt04vdaULWpz9axQN42sSPciYm+Y15PthXc8d
lhJ1NcLpDLSkAvXAgZ1VCTcJ1wgZVzCigmEF7sgR7/iHTbuFmlk47zfH7kmGQRFZ5mbl4qQZol3C
c4Ormwu+TyMefetG/t8hmAQ4465RAu+n5lNFhrJdcFTb/IpIwWKHehsg+ayBu3t/vXChJlDcQTFe
JJAZI8dG8IpThlzCjTjxdBt+6gDN0ByR8nPJeCytigTthRW+IXxf+8atQrsCrXx3VXQkyWwpuXdR
m5mY3+9EEKlFfb8sc8FqrsFpMtZJnDvuUBmZv55SycSLQTuv07rlc8gMrqmntB1WiRVpcw4UbmaK
Sy1jPj021pC4hi5XNliYm+EVnK2f+mubkMTUAnwOrTatf0e5Q1eCqvYWAY5Iv37mRVjTyHul7201
ccszOJvxXG3A23Mv4Ty7Sukx1tXuejC0w8qaoi0bL1njwN6kSGZ7iiKV58Am7PuXMmKauWfcrOHO
qXFiWap3XbP6t6UIqSi/Pq8vgi5uTJiSVVWhESBJuu0cg22t7pg12s4BYT6uRvIKDI2PK8KM9OTn
cCw9MLFqDVweJsvBHicZrkbHTko/OaBCDhVFXFD/V66W+DqtQIbsBG06V9zeliS1Nc6H+7OXNsHH
7XBGS3p+Ul+q7sBOTRNGq8P5DzqeUC5PSK7Jw5rrgdLGgewcJUgwx7ersZbAoknFSnI4sfcB+DRN
1TX4Unt0ZOdGyxd1FlmGcfNrE/bA1GI+dHWFyNCV37yinJxGcB8ePI3YY7boEdp10t6hJui36vUk
ywrx/WHZ52BFJJZbrQ9kQHXEBcojGIIjxFRgORbLlafaSUHD3bB6h+JmTPocf+0TK3NzdUFzHScw
I8mTib34tlXhlE7ptkL0KA4f6A6/9k1u8XvlIK8bLVUNEjqEGM0dNoUKQw8ZarpRpdu/9aMdAI8T
hX96XSNmj1kKKHJkK7FA+R5Dgw+Vut0itKJrHTAI7WuigJkbNMSN6AVLPs43RriPfXcgNvxqShvG
WI1Rm5vkaZcH89ZCiTax1PukLTM973cBSJ7OSw0TkXy5e3dtRHF7oJDRpDNsarQ15EQyTBIc1oaD
zG55Z9HhdLPi7pYt+SBb/LUZZiCgJInOWvI8/nzhzAKVVtjiV3FT0G14GBEThDTrH1vK33Rc+fMA
mFFBfMeCKJIz7FgzBdKgXsPmRbgku3El7q4k4HXGqQ+RynQ2RXvsgM0Mob2kNKUPMKwkI5tlOrk8
o82GCVkzfbW9XQ2UuQIUOzGyVhgagFczXZe6TzRBgp8gb3Kx2ScpbQ23T1D7QjgwqZxnwsQwxrFr
+B6RJWityioy5lzkDen/n8+3CeLU60YelTOxgiK/4J8NWTQCEt+3T1L87avVjZ2K828DKaa5vkAD
moGa9ZsM71TRdL5jYy3K+EsFssty1G5Aq5vTDxSkLshaq/lux4fPUgqta+Wf8NIfEWG8yGZ3lOMF
/jScELbIjyJiG/vvmyDgdPoswevN6C3YBNgpnsXlh4tbm0ZZocOMkNyRzGz+nXEUaR1+k9pacDir
TVekJMfynMddy0w/CLokXx4bCQuvuJlFuKkc+4HofcsKLXnmGcXSs2R/IT2pJhjStADIgKaI2DrB
P4+Y4uCsxf0SHmxDcj2berk9/pV8VUBu1L82eHpdLY3FLuiEVcV9TSWxoxCTl/EqKNef0VI/zV1s
F1JDjeJE488e9uI4eUfSL6ot/wsL1mbeHsYi9RxRPs5Wj4jNLuj7iWiv3O3AyFKO79e6lqNygzeY
pA2F+2lfCZxHG8d6vrYdbkCemXG7wwhVHeCoDVjM+YQqIfFPC+2djOVORtTsVzf0xH2Zp1PYeUz5
wwrOyrXxut2RfcszmBltxHPErqYO661KH2vPc/TDIuRYOQfWGeTfMFeLBQHf3dWcQ28i1e7ZE9q6
pLUa8tvHj44muH3fYUfT68FHTyrSr6O8YZnKzuzR+wOimAYnh/IRpGZ7hj5ky/y61xrN3y5TReFV
G0vpLWX6IFoigswOjuskHUAWucHjC5tvYc9xWO2GqScv2v0WEVj38gk2YrYmxygFHC4sj+UcIrUj
mwAyasGnqablfp06em6Ibhu7VY8gel892V1D/JJYbOj5ev+CaLzvdrysygdGqkUROiFcaXCwAioT
K1K4B5kw6l/q7gOIOTz7fAZ4oRhufwCMg3J5od5Oxph9gp8KlvC2oRFGrDMtEgbFxLj5lcVUyy9c
v2AgC/OdL9sTU2IOrH30xCf76QakQyOwSftnO1GrLsw9O2bKYlI1cDWgR/+VaR5vWWmLWzrhFuX0
kMGEhACyk2mt8p/JT2Pm37ASeRv31glRBCniQIDa1AIDIxMoLRFGjSzanTWQ9JiaRoStHcik19VN
GVnfwPze4bRYynwhccIM7opB9dlAYH/lvNNRJ0XUnovgO7scSpek4xaht0IUtoyVNUeY6kOpYPAQ
gMHs+U8CLaLSA4TCiA+Y5at1GLCZAKH4pJ46iWXkI3SIsH2ZOVnrEJOMq/ijPxZOCr+9Qlw1isfa
ENc/sT5zgqbCF/gf3jqTLWWmXFjKMfGAABb0PcEPqrj5dSUV3OyhQA78AF23pmEikKkFkrJqgKJQ
G5N7osXrrSSzFIqiNVPfxmI74Ge9ABLExqhjK1ZFIp8SmqCDeJ0yKjWo2ekdcaV5sehVm9YaC20T
WUYvVIy3YYqV1llzK4CQ31JLgojx42GZNBsWTRzS3RHwmgBw8PUkyvP7VeCXuXaVMcWNqEkqAoRW
oTCZGubuFqMtWlmM4O/fTQ0CKFT9V5B9ikD4GN3byMcXqY5x9Nm3p2V9uvViXyXA93HbE1WhPZcV
6or++p1tVR1Qb3Bn4cCOXIyYEEKtj1Ha6gZM83YYz/E8lNa9IuvTcK5clXwIrZ+J+EcjjsITWE61
4SjN9XTdHn8zBi2g6vYvsVIGW6t2t8lwzpFhGIDRQto2fuSsUOgiVtOCxxNj1oFcbFnUKElVrfN9
M6myDN1i1cH7TtlK8V9S0SmpV2RZ77FGLxUo3Hx3QocMLv3ATg1oQKVNsvVUDFOL5mv2v3hP/L6E
nECrgg7EKHj4vuACkxDsibiK9/FUNRePlJK7lZaDCapZRvT6st9NWwYEFdI9RDjZe7mZs90XBxqW
puuLa33yQ1jD7GOeOxK4LD+2eFOXlF09GRBeQOaPOUtDCxCyJ0FqPavp95a633H9TK0bpFdx0+zy
fasht7CvJ9f2ukJTprN7EU5OthV6hflcpOVqXbgNJnl0OVaEIw9MTGJ7txY0NxWQgLhu3TlEphF5
J6aTTQv9h3xVMCArnOoVfXXESBKZtiV/82oVmc1Y70WCgaJsCUC6uRDIC/0PuJhDvUkqUnqJ63G5
7++NHM/hflIUWWAt694Nws72Hvqfwy7+eE9ta9+NwyOO83UlylZI6MiBO+DQs1hyF2a+D48KXAds
slbOoANWhqefjtMswp+29eFSSugZGowXnAGOPdvWr5jfOmzlnbEjH9ePnsb+tIQ3vM9xak3a0FO2
qJgq4coHkTvFixK5oVEHq7J/VVfxoFRSfW2KlnN2NH5lSxmYZ36aTJ7k/eY2uz0FjGR8EiA/mTLJ
5Z9YlbD5TWomEsuWs6AJzjF8K+8olHj8+AbVLySlt6SAcqapmnijAY29F4o6o0gZkINNxaQErEq+
GLwnIwiqFISkIYl0PiImdVd6CnLACrwWUOdN8zC+aybqETHyYaZonMswqDErCtdOABhfAOodMqJ6
gbgtgkih60ivCzaRXxiPRKN+TkZD9GTC7WTkHesIS+sxYtUVdgWWF4d+SovvBiTnbE8tB3e4ruEi
3iiyxjgeDApM3WM92ky2Dlw1VniRM6XhpE4rptelqmM5Y7VZmEJEfyzGKU/Yo7Dc4gK2nI4/PGso
kEzyr9uCsQQylT29T9LQ6/f4lmcMyp2/ng0PECM4gisiBjjepLi3AO7/Hce7O0Loq8+QE8V+VSGe
bOguoqsmnBhAyGVhWqtiZpvRsv3pc4VwmHnAX8+gySHfEHhlifKXQ2n8I01fP0Dq7e3TnVO4qXLd
h88e5ecRZYjsnLNUN0HCAL2SIO7PRU9P7o1W+JEat8ZI/uUAkyRsvfpD0loc5RFsuQfOs7Z+iHdU
0GIpqS8/t8Apa7ZYGxk3c8xeyxZic4Ug3Ug4VyAlPnzuEccr8q5BtOCSNyg03JZmgbZnOYIuluUR
HQUt0aZOaqILOAG4YdOVI1+bExsCqk9pBkr1cFvkzirgl+DWE9NdglyrOcpr6JuCIuOjVu8E4rYx
dh1N7no7qK+h1fiLyvXnTiC3W5y6+bm2VtU0TpobabarOKgSroB6vXzy9wcWejYR2Ixtug9AN2v6
U3iLvCITxjytQXi6y5DX5S9LNh1gdT2rsmTQTfWR7Cb41y+DG1XFP0ozP7/pZPm5BvGVlls8Yoos
xaDKIxu61CyZCNxwaLrqDiryD3iNYHUNv8mOx+I0z4941y8tL/beaXJD4yqk/vFJiIt0zkcGQAE4
Os0EWnUojGXUo/5I/uXvhCr/kt33OsLP9wSEbjR1uzkvidybqP61rPFUPY3NHfdd0WHMHjyWfdM8
APefR7gWGDXMP4wwrvJ7ToB5oD9+zDlrF0WcD+GNqKZ8qypggp0VxI5nyCAtSkEzwBqBUYlXtC5X
U4GW2qEEif1dDzZ8HFaYdaYxWoSRt/67i7s0dCD3yyxiMVAxikOBcHIuO1HV13bdV1J/eJIyupUX
GuKua6HHQza1nf20XTooQ0p76O9sLptByJfuwUXxwUGnaL0CyD9Pw4jcb6DteU3/WJ61k1lCYgI3
1sQBM5CJ9KgEprkK+u3aKkZDj7GpSkD0ymr9tytMMGMSkZPtyavhsmNrVM/utmJVLoAFjqtq7BsM
Fe7CyN3x033qC9bzC4jvdLSrNaIuleNCuxJQCF4B/YLhl4mCUqi93mf/fHjMzWWAYKVPV6vyNhvO
Lw0m3OHf0s9/dLMr2VzKxzEB/sTWsetH/MGFGaTMuDyWDHNnRs6wNvqfttrTzXNAr/oIz/iWGbtu
MmO1uPPnwQUm0qrmkCYq0NZuXhCGaox3uizXaij+jWqOcVFpoGClwUrCmuRafggd5DEmzs3pQXa9
Rbk4KWr6P/84gZVJGIpieBaCBptnr0VzJYn2mf+sP3tb2bsR0r9cWilCGWwzeQoOo6dpE3bp/cIN
5Gbwm6nFuPHLGyFqviPajd5EeQZuWW3Yv/0vSHqkXve/6eAW+RsqO8dkv04DiCQErQu01jmXGRs6
vWXgM8rxk7WO4BRW4IKtzGmtqIdEKGjb3L0S1Gq4uatgrTboLP1rXyzKcihkpHeB1F9mYZtHCOUY
5ehPBcLZpF3tgAhUA3/Jg+ZT257dGj7U9h85G2B6CGbH/4yYgbNvQWXrxTkA+smLinJ/fNA0r7R9
lV5yK64H59TRgTGV9k7jy4s67dXOSXhw+6O9XBR3pPzw/lMiu+johw/6rPgMoQydwBFDdQyb0WPC
9Ufyyc+8D+U8CdB7tTOcjlE3ZikAzr0E6a7Qt0OqqIxVSFCG9R+sKxjdUEnQS9vethGS2Xojy4Eo
I3fbuhPn/McC6em4OPg4xnBSk1TdTagvvxsrsdS6gTWKj4TQbheHVM9jDnRr0a6AeXuVcitD+Wul
DaRalkSgH6QbpGvvxattBfUzd6dzS3rIb7fKZTNnjKOPUWvSS5HeBDjioXqMaDhB+hyseTxBKWNT
n8nsFgb1a2jHGVaQnL3MYGSzOvtGDMODhbMemurTaUv8ojdjHiOqqPx54DeUtCMJuKERE3iaNsKr
h5RyTZK6AHsR9EO5KPB1Mtung/9MJktkz9dR5PceQD7BXBb2CH7HMwXtew9NLRrSP+MgGk7HEb/Q
CXWgjJNkSVSLxa4S0CLttgNIYTbfAJn51MDBpVX4GC6w/HLvSIlG6fUlUOMQDizDdnYa3gOAqZV8
3viBLaC5Ry16tlagGeBVk2zOb+kIQQmfnSKyivYJGr05cMymwgMD6Z21TUx42dsUzrd+ug40HkLi
dJY8sn+D5bukI9kAE84w4lJkj1/5g3D8Hdz5loca32qg+HHLlJzHTgkDugvHVRKF0j/rNX5chxq2
THN+8oNw6Z5GOTH3UP5bNGvXaBYqvx8GiroGh8szbQOUhlltp+uc21NC88UhqWNtWkhyo+MovwRm
3mNEWY2zL8xWDRKnDOiIlZrscl5WSYvHkNiLsWVlVDc6+wa7+ycn/IXkBaeegMVJUAPRXLMSUFQW
C44tBRKfdNggELk984VoAnRk9mA/RIBuYLgGkAwUbm517s9BN16E8PojPNqbzo1j5zQKGzz8z7Fa
iY6Bbn2eawx318omAMFv5hwP8Y797kUDyUUj+ms8UtjXUJsvb2KcJ+tszmo+8rWcXvVpe18haBmE
uVumfVIX6phj3K5HzleqM7VXfeD0RkjreQP9jvpweOp3y3GtdZYqzKNlevzNXnjXrviyg7giLY3Y
a4oIETIacHAX7hzgRrtYt6E2qDyEOUHBgQyFUArEX5ydBehvo0NiqWpEJOAl0dLEPP7B0HgZRbfb
99oysauLUoNglNoIa4Z+5B9ZEcWqlB2mEoXL7O1Jl6seNiAg0ATLY85yEHqVCF4hmKRQ/Zy4F+IY
D0FFv5sAo3SXm0Jr7JAqHfbLIG7RkteUEObXvaZ0TlC4aEMgwib6RXbrP2YVVCGWEVCpeI1071B2
MAqXvuN3hSiTVW4AO2jfpzhSqCF9hkAwBrMYYAkMuzR9JTJehXKGexbeheoSWphGZaUKOUdLI43p
18UPKei/pQ3wrhonNFlUoNnbPrBWl7xhznytmBAFTfIhSfcdLCaKfe+bX1Zs5t98qI0js5BAhCiD
BZl7BougR7yX80UcT+1V7Xwltlwa3LL20TEivBtuPs8jba/mGNj00GGBjMipDKCv4Gl9hz2cB05v
6M8t439WEME8olf/RlQTcL18DCOi2OAGbD1FI2MEIuA1YW//M7inhbfNE0lOUjlLBUvGtr4sgxiv
wo54VJpRDuFGCtfJ/bfNWzNME9ZbOwB0h69E9lv8mnSzhM5caUDL20Wj6gUj4pcx7a5sylwj0q3Y
DjMImOcuEQLac21+aKQYmzCVqvStD1MQ40Z+piI8xiF8SCaH3VNBu/j4kyAm2MXDxieR7zA/u3pm
xkVU+VHh5DQA5ab3Me4/BnRm+h0WAFrLkFvjCx3IzDacdgu/yBALF0GqB7l16gu2bSsfDYsGh667
WmY+igfFppOVSZ5va2TzW+Cx3zruUr8ncR5JZ1ZsDBnOMEpIv8JJuOEWzTFNBMKKSqUuATsTJwDy
8P8XMiLTbUtk4ScyYfgqxzbFW8aJqDS6yUw5cxuuyBti22AtWsuz9FSrtDIsAo2AwtWeMQl3V3Br
cH/d22sEF7ZgMTRc7nKoFZXvzEELAyvZ3StjISFyYtOxVGsAhoxoJuUCn0xA10AC4Fdaw0M6PEgu
Jisv8GgBEY1pb0v10NtXoMFmWVCQnPUtKuTfNalgKEftmyjBDiDOcxoSOjisd0obvOkLXSZTiadK
lyjBG8x2/MYrtdXc1uutoFByYIAGvqCkQDXsIhcHweyneG+6nppgpCubWMt1gsKtB+Bv/cD9QF7d
IVNGm8AjpRdYjbFEQorR8d/CdAxBzdSvEywBqUHb3QqryyvDvDZDAzo/GzijwmiEGiCS8zIErafW
VIRENy+u+lvCvDxBwrW3f+vx5uOiBrOmOJCWGWYFpy7sj+f/qgc6yfEt+HtJjWP/QYyPOp8hlDQh
LXM8kVWG9sn71cwdjgd2qIN7+2pXx7yUdKCp/f0r24IIz22nVsiyrpb0g6TnAxUbEZwt2az/rU1B
0ZlzMR5QvpuK3AluJB4HJ72hXyQgAM40s+s9HPeBos28dhtfjOaY2OvF35yfjjFVx+ljydIS0We0
VTgBb6rTd9X4b9XHdfcBOukyrn8xfM29funAf3kd6uYT5ZyAe2WoXvMJ31YrX9ftje56y/vgJ9+S
89jjORPjbB5vThuMk8/XBoLRRTzodfngNLafTgWtENM1KZNwVDW3lwCjRTRqQFgY+sHuEajHAD79
5hhLvt/W2Yu09R9iZPQOH4C0faXydQCYsp1OFWXTusZRfKa31qvGrhG8hHTfo33r4Bume26+Kpq6
6MYewneHsuJx2Gm+bJjF5A3Q6ghWklg/R1sv3csEjMX14It52n5sAeIoGPOPnm2/hloVa2fs5AP9
XM/kEli4pahHcRixkoCEZvGwXfWT77vxSYOA73IO55/qcR/K4mXOXQJLMh7HQYnSU6OLCKIiGTjg
vucEXBDxST880NEllpMZzHwRI3Ps7BUigkkvg6tB3j3m92kxy++Vienhu4Udoe8y/mpAFTvGvfSX
tIknB+vyfHFsioZyz4g07r/drWpE4lOWA+0hEuZx4NDT8c+JGJn30b1Zw9nbd1PmOnJHsoeBb8iO
p8oqn8pH1f7lrjFZ3yAkJJWPIgsDAzacatWp3nMiiu/CkPbE1RkSWd37HuAyNSC4hRH6KXZAeAKj
uzRXp3N0SO1Y+BvML5FWDfcbVJXPRzLjfawYX5mjQoCR0TeRV5U/UkcQDllsRL7No1XOj3yEtkPU
BOZ/EI9Ye6n6vmamWwj3B4ZMG5B7fjWc+ZmRHp0wr6GimzzCPh6Gr96DXyxeaVqkTB78AG2iEqux
20TOGqmEQrsf/GVhWAnrHvTVkmWAM5l6TF1pdE4vRiZVewInlulbJP8CEwEqA5iVERGIA5yp5aD/
sGur312NtX1xPlYpusTuy6YBgIV64uq8MqAvV073iCFWXx0J78hBts92EfUoVJrr7RwNw9U+af00
dOEJVZ+cT/7IR4erf0DZQDJAZumI4/z9KRBknX7XtqHDERYP93txg0EQ4jl/y1zoDTLGI99CWJ67
03z0vX8hpRhZntgq/LDbQi5IR7ivLurlHbkaBR0ikEOQ/nwXo0yTNOklfUMhjGWPETG8fsfcjRG6
AvavjgUFNUDB+4w2uuLTU8JdfmIdCB5ddZPDhBnfzX0m22aU0xzpKo53FWwSYsYK+ZA3ZzG9PGqy
edbD/cltDmsu1IB3tqEwRp+0pq+iz7eJeqvdE0ebU4S37cQtr6po7NLXc+UJWjO4JoIixhDAnROl
eet697RDudoRShm4Hxg6AzodwzZyVhTTy7KYnawwaOmkDihmidgvJRzDcqTRKG4Kh/3uOnXwMJB1
jMFs6dRaqhYJOs19s9WP7OcGf/q2Olw/3CxnW1ErlizunXENVKdZRLEK0Xlv/Kj+SUImFZsR7RdH
yqzM6jeOIEMQFY2x454h+v0zp8GdApb8aF+IJR2oFgagIi+/NFVPgfIrkKX8JLsS/Hy+ZTVX83di
Iw4JFl62qRv0Z4y26ZOf4LCvchEYtTmmtcMnriFTMToj/t15r/pv9moW6V8trHiWw/ZstU1o7KpP
5GExxavfbQ32TsH3suALUqXrnC0sBn0IoR7VBX71GziHtFc7Vi61kA2SEG8eszD3NLJg9Z63xNPI
lCSsh8Ewce4bkwl2PaeLp6djvpNyHiXTGrzSPFaCfH9BL5n3W3rcNuX1ro0xrKhwNdk/RD0Jr/vO
VJJVIDAUiRlK/hEpUOGWwBAFYt43TE2z5JLNGAdvBv1RUw5ZCEMFUvzFUad5Sbi9oMODgpHESk8B
t/c+UVXFWU2Svd5Ox4w3Ii1hZ/gurbOB9TFs71YbL3K1TNs31+Zh5RLQWAf7F+D/x/ef+uknVkx+
Dwtn6xeApe0tIzswFkRg4ZdL5uUlyrsrmnkDZ0Ns5rMaJuYnkR7XROAo9gRrFmi4Iw82xy8X3/5Y
JE/qLg5RVh4lLHu2saDj/fUCdLIGqFVwzWf1Mtp8+zJ8W0SmqfAlYEedtSNPyi1IsCRPtDiFB7Aj
Vgmv25TdddkGo9gsAS+VPxDRZ5kCuTEsvztYkWRHAUpdPPiHEyjXODjjDX0xKMDoTdphJGzXqVNY
AdEOVj4g7D5aqM7yG5lm+15vBpJjlgn/7rQ33lY9l97n6k+bTvsTg4Qif2cxhUETu0ZHZj+FARbr
bg+hF1k1AJ11y2qEeausCkPtjuGoRoddpGSLnZ99ifuyQsDHhGeEzzmCYXsal1TVuUuxJk+xpLko
NtkJLwZWb5uFAa/oun2gZi2KtpaimhlPa5iicWphy0zXTlR4W88k46rIzOfusS5U7takgWVxGF9U
1XmsYmdPZ47R3B07tP1d90wZHFF+AJIP2JwkUgGL2am1gwJD9SbsZpMBZIAjHPJGtmNMlkG0KmHk
1cVRlcEn3yVQ15QMKmhCcR4abjCIwHyAK98RVTPkVsF4qlgdNB2WSWe+C5GXKrr27eDfKoV0GgjJ
wRLmAC21PFWpdPRJRvgbgNYUkXnrOPzTpiuY8zMdsmGFYiZqrXW0dyfu2pljtYlNH1r+6NuT7Dfg
KAuwKSTIwPWToX60uLpw2DVfqgO8ToCMEAXSr6zS6yG84PZKopY8hGmjTiqYZ3ERK9RVSluO9NvA
zjKki2B2ktVH+N30YxsAScpu9H0KfzIovcEECls9Z8UHd0hc38D9BK47ozl6sMLuTYH2kWdE3jKj
2nvvwjhUjQBQBxrmJlKLeJiBDTzb5822n04BrlmRA2Q+N0PCdRoM0zY9RfDxBX9AWi/GCnNzOZbB
PXwNM2T3NARqvVkzTZxlcs5icr4Y6ax1XqxDFnuRutvWMTUdZpl7EOTfdO9KVaZOT+d6skGSdjfa
fETiPJEcTQWmZa2Kbkgln1iejw+sqitF7j/ydHyJ9se0ugtnHNx9yPklW1+BnjBBGpjwF7exLR7C
6h3Pxf17hlgXtnVVQ7ybBpyhsW8lr34bMHfqCaYR8vXgXkD5OwwOvlEMkNR7I7ANWt/n9jMN1nDa
i6L7yf/u1FjOuogBJg2IfDFPeOZ8SOWGMU11VPY4X/rQQihxCxHynFdUVAImTJWdMH13qrAN1X41
mJt8ec8guPwxeU1vGIHkuXOSOf+BiFvQp4FV96a/EEdG0gdqjVHzoR+DexUWPVYR0Go6KZYs0Jvc
Z964D2obojlU5lRBEaBPix0NiZv/Ldkf2CLJTrVeD918bqMNc23MPHlCefUhRVxZ7pqZew7fODfI
QyR8n4O98mx27G5wx834j3B1FJrkRNzx4z5OcgnSbhBjPsHOV2Abm4hAShzzmP7u3EXG3TyoTesl
nbU4RQjdUhNuNFOA+u6PRBJhJcJm0cNcJ1fenPl9SHKNXAwkzJsreWE21d3x5upuH/P8PE9LD/dI
f2TCBCVLfeRZN2ITK7LR7ThsGiLoEeFX0JbJUfH2CU1w5eIJNP33UsM10RfjDOgxuG04DrOevJd7
v7zaSCjRhd8IupXsIPb6IrOVFiwP9iwIn6ByiMVBmSm882Vq5Ab0RM3e+tp4k9dfMchOng2mG3rD
/9GIbBCmVQyyatZCzrow9ECVgsfurygIzSO7xsIGZM/86fYwi963+ZEHlCIzsoeN53vKwiHLYUn/
C3vp5OVzY+6jBRkV85sv1kKodBWT6aECjGIlxy9erEJjUz8lkShZXA8YqPFn7cExE+3gxUWdGUZu
atOZA/Bu0JxbkZTHHH4V6WQmhNDs2+RlHntVpZp4l8xN0WSBFuD2QJ4k6tLDbwRUA1mCFnafU5eF
xuDWd5df1JFXbiWhg/8SY3o5eK56dZfXuVu2yYOvAcme8ESGvc/CHa/UBizEvQ6elVSl6eptKOqg
pgelmXLIhZHVjlsOj3bFIdjbLEReQXgeMW9b1GtQob1ctf0sLMqOcuPDhUptPLxLykAXkmBE3nDY
pExCheQ2Ie0aBqOz41RvCsWqoOvvwJaouquL5JO0Du9jia1p9NoqQDCnt5zE9nJwbH9/ASPo7LkU
BAncF2Gb0Eo88OOMVMSoHGz5TgxTRJYEzR5FtBZjRJLsCoanoJiXhQZNX1zitczhuluzwunKMdWC
y57etOJU6NFm3HHIPMD9m1SSBgaHrBFMrVpD7CBh34Nls6rXIX6vdtV4bz7y3IJFPBqA/sz98rgS
Jm2CaFwtM39xPAbcsQHpz8f++LUU3ox3RPubq9mkiSqt24ahlqr5ymSyiueYuL7TIinNjc/hgAvI
ED2TzldBO8jXQiFsX1oVcOY0vbeVFXUJtNk0xItAXBQ4Tx+Ifym6l2ChXcNzWynCuovDXVUGW8jw
NmJIcGxhSyCZziTpOa2IRq9wVuU8Q1PU2h2Qp3PoGlUxX21g15al87bxFcKCBioubyVeaUDWdvvk
6A8cNO5K8MhjH7mdw6kOd/pOPU3YYmUwmvgJ9Zf6fNWzRwoY+XIG1iNI8bBZ0547K4EKUbLuxyQH
wmnhzMBFUOo+1misHIw1DIINqe3DI7xgrJp/mxJoy1Vm45mGlS83YepUN+qGdkhcwS/4aDWA5AfK
gfjz4cCW5GN6GaEMOOLKEhoK/EzhMsm7FHsZTYLijOPGkaYkI7wHF6AmROJUr6Kg0WMjElC7OoVM
jLxvzu1TDz3t/UOwvMTHxvk9uHvXmd9FYFd+EDEs0LeKNrYsiHM8bjmTPV4lmeDZyfsYlL22ZxnZ
CY7mK63CycZCyjD85/nJIGIkfEjpg9xrZCNLtb2qJ3EYoalsOru1gM0/NOW8TkwlfgzWKMnb+V3l
w4U1od+XHsCARSrx8tSUwLoI6HSNRjsEVrAAvI7q8jXmmj+Xid+wj6fkfpz3BNIQzSRZ5mpbNn3o
05Dz4rw1lDDy5dXyFCs5Dhw4sxKccRiQpT4IOVWShUD9+nKwWux0baxukqBw2LKRqYhAySXXs0nj
B3usFFNS5oTpE0Zx296pvmVuoz864YStXm1CyalmOLJtcWKn/RJ3gVZulBexI88YozPt75mE6IS9
kI2XNCFaPD0FZjhmMdrF5fdMrBJUTFiCra+vB5r51TPhhluh98mEG9yqyrvbtVmVXRdLaFRAQr99
vTu8JhCP2yr6/eRFgHrC3na+Ju4PhjKJOu5MI1eGf+cmoGgkM5RqwKn4NSX+kGf6N0P4DPEkU1oX
Lcl9dxLf0a1EQuiwWY8/FV0oP56/yWm4TmMvpUgbPm6L54ymCgEJgoo9eQnWiljdNBf2pCcv2Zl2
ZUK32459RBdEYcFG6ifK3FiRkzDthsR7GW4PVQ2Gk2enRLewXMjfTxynXR44X933FXGQTI0N/gW3
qrnNzF1YEEqChUqtDBRFeYZm+hK5BQSDzB03LjtbkSNJrEQCbVt5ELYv8IVyZ9Uz2JTXXBDiHamu
Gjuv2f+aBPZydzF3aigVXX2kcBvGR1mJX+zbiZoyCA21idF7e2Avq14j1MyNLeFDnpjXOBiwOYrI
KoO/JOgYAf1s//UNuDyyF0VWvYk5vPtRBgmWCs+ayFLU42h0IeDiRvN3H4dRnTyXzo91B11GgP/B
BgNu8HzQXKb/o0CfOZ2IkcNBMrfgbz5LannoGEOj+ZcXueWfHLBhBtDMExsm/7N7DA/xjPaHJowv
HVYJ3OdjQvJOxId/s55R2vj3YcqI6asLeDv9q10+gfOcBTy/k3nph3SmeOpohE55ntFybJdUY+Vy
jQ9eeEFjJ/H9PLogSvrZd5RT3bEw14Bg8qHokzl/7zv9ABPRA5GK51neNUsOCzqigaPr7IpVhvJB
0hB7ssnV/liE82N9CmTzwHUdxxTuGaYCwYRtgVr4kaSxdUSts96PIi5OeO9EXq6f8/wzpvmDDov3
xBdSmbfxznS3mgPfp6JLqnVazueXByTHKf39wnu0BIpv/gDnWFAl13N3l80oeEMe87B+wR4I/OU0
nPDl+HWOFTzAbvhrT5dJ3m6wUvjMc9XdH/VW2BAslvlKmIYr99rfy9k0bgJC2pPx3rSuPUrVSsWb
FWOG/O+P/DIj/zVoyaXJMGScwUo2lqE+IRbAxjLUOFPRysZPFm9vqEqF7Dt83WZ0ricRScRj0Eow
7rVzXSxwqw/1GvzCZ2RmWpUuq+XVI48nzeZuqgx22mFnd1Pmce/U4QaTqoHHbVy8+wItAUa0dXY9
eLf3Q1xFtQzrQtOYZWfrsOFHwqI1XofVaFHi0ADNMplEbR46B7wn+QK8PwbqDlHdB7qJ3MV5In30
eL2N95+t00qtOKzaX/UOFJ0x4MXUtGnGm8NXQnnU8uAd3KWMnywWkuzA+HAebt7jClyldTE1xd48
RnX/WuaXlHE+XsJE2A6AiQtqnNMii/e5nkJCSAScIk5mJ6Rv/ATeSSEYjq8NHTkaZIaKXrHkBeRp
BBoqxQj+QfBjhn+e19l2Kr3TtX0/8Vf2lAbd+hexOe9cECBMJcyzgwAwcaBtf9fJ8A1oNVtzdfXz
u4PgJ2b809orzMij2qAHVAGKnBsq4SUuROsqJxiOXfOpWgkDyqp8UmS6T006SiuV6oD4GwCmPCpB
4058l9y+ko4ETDQSb3KKBxGhhqGKWCa/eHvJsh/ZvCx/s8raVNGUDvp4dA8uOCGB17jUDS6QQppM
5C94+zB2bDOsQrbDQtKNLx5FVDQBdClgNJPe5BUJPUaXmBCciWPQnJIEuZqrQOESdmYE85ZLx+t7
oAl/NJbi76D0cooDrzFsmXSpK03CniejlhCnSFV9QupyLxyF/qc+4wxCoafeuKS/h7WRoNm+fyk1
gkNYsURbjLddn9LsbIDuIA89oFQc1BJYXIL/n7tcnxJ3N1eQW/sjBCPLOSpTIkJ+uhgmI5AZPKTC
/AcSZRngLK898E3qkYa4/p3Wy+OJf30Z13zTD+9l0lMnz52SoqW2AkslEXuEMfgirxy/IN5jZQTs
ubpEoY7TWnh3+frvVcoB/rflnPeH9m4Qxa+LDjwtCnOvfEVW4nlo8dFCqfwoPIUha/ToAExnN3Pw
VT3sFlKgbr4UGf2RE+jXHKDlTbZPkwmKBB9msA7gkJaPLOxonpCjriOgt8e4qC/qpXf7odDQr/Ii
3RRenewMTE58pZOODmGP3ETztZYkZFQ1mv9N1lEv2Ve5g8tt7ROLrrmujl97O8H7Rky0LpBElYfU
n6eAg0w1NnaFqIUsGmZVR4QgVSCV8HE7yrbwkegHrg2IUJ04PKc/n7BK9lud+SlYT5JZev1XZHhc
pSjWloifC0uFvd96LgjJSD9SFXhcWZiHpI3yOlH5Iu/k4w+JxGGhTaocw+rGH4/Khn0xZYj7UmAW
Xx81FNCBcc1hm+aM0qMe/+uASUEHXdxhS3zCIzCWGvQrUVst7LE61j006CZp3nPiZECQ54zFYK6X
Em9/PX0VQm9fK/OqxnNqzcATzxkNUxUfJ00IASxG/WfhvzHPBPqgXmTefDdPxhOgjWAa+oBF38Im
t8FdfVrhdTk2WoPl9eHDRNKCoxA+ZaiX9/NInhylKJknFS3KaJJxw8fBV6knVQ5nViikQAIJtAz6
3vUWUtOYWgw+oXnpyzjPnZY7fwtMKgKFiDFC+V6t2Ol0vIJ5kuA03qNFsaaeMSif4eiBlAUQJSWq
b5s6W/W8+KQET85SR1oXRTGv18mBoOFQwqUyF9lJqmTfNtAv4C9nI/zKv7KtFYCG/5aHR8rrq35u
0NI7QdnkB2FjT+2Yo4MnAwiZLNEGhQZozfR6OQnFSLhk+vN0yN3UJvcPo1uY+2w6PsmuB1l0YNVF
7wClHxEi34bruNaFH6Xr7b7MX3dKBTFxDSWil4lmew98OEiSLdypa/bX1Nj+OHowVrEviJqk9n1x
j8RWCVW7WQa/5Zput8TgDiM921uLBhEzrfmUhONJWk5HHcWZ9KJCbMu6MUSrOtnqj4JTYKnCG4y4
S+LuY5MFp/7hTAAtKVneFNfmNskNhvXbSeOFquolca9Puu5lYwPw9/yK1d3Kf21nGnXQvdWFz5ho
dVyJy/Nn8T3kedSEA06KHSA1O7JRSEXLUZq8NridKfPMVAHwZCG7qcYPsOWs+3OWka72RVPT3ZFt
iEtsoIWseIfr8pg8qlFzp/J6t/+0qhhDybcXFiowlyfeuUE38kEI18bPnezdC5VzrxfRI8pFQSVb
DaF4j4kPzXIx2NdW0sfJJmYwbAJsj98fzXL3Ki9yte6HlOEVnr/ckADPvhV0/wjNavCteBUR23at
9fU1sqmyPpA8cqFNEN/i4pamJKssoQXSE+QjIFGsSoSRPSLsDOmegbRgpQte7JZWMCF2q8hfj9bY
U+65czvEH4Nq6rCE0DhKYEEfH1ZpTMDmI8sE1yVHcCONHLEuyIJsag9xEaRwUhYuiiXJIgTQY6QL
D5h4rnllH1mfFAavmj0cW2GfyG+v8nlhUfTmw5m8FIXaglgkTSJ6urtMhPVa6PYJJUw6fqMtj9jr
EEjIhmWIL/eK4yv1b4SmX6mct615kPet0h4/QYbBEscCOSvNcBW1fb2MEILDlJSogl64YTf8cze2
1h2+XPW/y7/Sg84emNjWxQYuKNonvEOu8gZ0IRfUcmSsbXZ75U+2sXcVGqZA8VmCnYMlV38Ho4hp
ycBYhreFL6FHk86ffoEUjdVm3782WJqw3xSgtefrUQcVZmQCpeEFfrGVwHwrLRamU+UASvajhZmc
dVv11+NeX3JRWFCmNYqVfk/KMY9XzNck7ekAzuirENHU9+zThUVZOYpljHZbfePalDEyMu6Cxk0X
7IEpIN3m0VytYk7tGSgXbAPahJye0sFJOynvptoUKy1VubOv2O9pnTcMDq8PV0fXZEgenIPf/M/J
F1zq52SOzImCVwJw6ZvyBoBDjVmFDqZipGYvqneeXzxOnty3FCn1b003u9VymzeR/CaHDBQj9JXh
O+AkVjeUo1ih0gXdvPLHJbV34BGQ0R25IkCYMPJuppFUel5UqWMTGy3aVJ0nnbCaUM8PYJd31TQZ
3o4G2x0tl1XRzXnV666u5v98Q+fHTpeohhWF+BVz4Zw576jZ8o0EMrGQQk80BJtVH6JiAYHn4/xO
I7M/608j749MBpIAwHddAHN8N+SbAOEITnp2DJhAN4/IE/nKuNgFYDlLWzWh+vuVW6zdUt9IPpfb
dJqvpCehjdknGk6godkygXHq2TIDBlyRVG1o8AYsw0GQcanZvzG/id7al/9apWdWdlTSmgArAzOe
8xytuTek6R5J/Cr3rcYWFb0OkzKo6imCqaRgUiZYgPzWXQ5LRaRogqGP2h9hYZErgJ7wPiaS77HQ
0AFYJq5RBcfpy6h16lNTuU/uJoeheaPP6S13xYpsp69CkCDSPLqea/qUpKnSDcKA0AShbUfDi4fy
hALLdu+bp5El+ee4iv6hBFm0AF2pgN/akY56IEoupnsoLUinGRZAe0A+MJBhcWze6wzaZkQ0Uz1a
0B1Yd4LF5LHe5peLr5veB/0rcn6NXwHmye76RAvRGt8/CNYIzlyeuu/TRZqF3EvQQNeuacYbd6fA
hJOBP31S23y5KDBkLXge91eKAU2qruZC7g17DGBgKsJQGyu+O/XG4t6HV9Ex3bWw+GmJ5VQ/FQzg
FEScn/67zFOIzXBEq8nWKDiZOQkE/mDBVX0n//fcXoj4GpnITZNmw5iSBaD+tJgTamMSTNTz6oeY
104H8rBELqysX/cs553/+Z60PalZ7x/VSZhnT3Ep1rkinzuE9gQX825aoUgLZOQtSBqqLTbOTFWE
HzW4y8v0qCKxtSKA1aSMl1VRLcnL00Jea/K96DNrBZSOHqwqGjERq3ySLpVgmmCnVyz8mE/+iXY/
qc6t5fc3WlmnAmBekuM7N1lFqdZm+Y+SULYysy9joP2eOvwk3nS7AOzILUPyX4sydDFEnxelH2wt
cX+YB46osrwpqHZKCg0EPPFTRixPu3Au4RZXM8lNH6btUvZuzh8BOC6maw5Vdu4/x4v5K0JzOU6l
s0JUkHI8Y2elGxjEgEcIARJ7J90QNNW3t1fJaKCOBZTZ92VliunAeCAurf9GmXqoDOvBpsJLWa49
EpWcF8t0Wkuz1lVinoIRIm152AKqZRcnNTwX4pBkbX2HowBGfEYs2DK0m+ztjE2dXMdLjmgORz8t
mYljNKfI1PP9YGFiw/aVKWij6YyUKGkHpxhapkuAwXrQ6auXSbm64W6z6hvuBFU0uRl3jUanNqEp
+/ba8MXFXqzQ7/pn4no0jmb4VB9fHL+xGtAYR2B/5RzVDM6zRT5kBjt9mry4aux++x4W2TKOGglr
jZF5WrBac/Txm8Vhiwn7afVBRQShVYqw8A6dmO5+zcPjv+r0FVUcDEh2oo3hKX3AbdA3EOwkjMZz
BMxn7xJe/iDIkEbc319OfIHujSMwTzo5j8Fcv5rmxwWcOnosEvISjV6/CHl9jCKCzx+kHh2X9B05
KJm6faXBu4p8cs9O9xHLCgv0RUh6ZrxdKa4vAcWGj7itTu611w1UrW5UWqkOz4PAn7DJAgvg1BHr
XC7sfSWQ6pln4TfAmhUG931yOfwlMT7Dw90AVrYOWT/E0FPVdMF3oKW5W7e9f/IA9Fu2kKdf5xg9
Ky3Vptv75Y71iwroXzclzLk/xJ5X8/vxrPPEUV7csUp7u/XyqMr3CDTLuOahNw9L0894VU3OSZXf
2TXCklvmrfpZssJH9lFuizPRAS9ywtQnQtfjkta3Z5Sh1jNZwAX5wnb9fmzC2KWeWRXjEHzbuRbR
brOnfiajiIoKnDpYdBx6aOaaqLPaJpnljvBbv7ngnd5nadOR44HnYRQGhmXZpyurBkbByb70idlB
AAri61ydomW/QOoqIzT9zyXEohRUU+0a7Fby/XE1i2VCWZnSqsK4DtYHC+CKCbnYRtDLOwAybYY5
eHKqvJwss8FUIVufzhCUVNTR2ij0G9NBcXYM3tP+TENhmfKrvg7FSdssGVuunjZaZ5/X1f8VFdk3
BXnRZdIUQWGXtSEpBKGjMZYQfE79tWtYCd4W9hZabHupgRWGMpQvLNyq1tV1BBvY6idHKPonxGtx
XVvmfOk7nf5w6wFE4XFfqgeIcKA+FGCYAJTQmil0ab1RAkbJUD11Xq9QnHmaAXfFv6WqcfaJxBzn
xFPHbT/wrX0PV4a2VfKPFKWzPujcA4ZlGBnixRqixisBZ07H95qDJPWSOdGZ2WXYod9tUzbAK4kM
wUIUOfBCZjwXRie7aOfRpZGOeG7lUi6n7/USe3Kho7V1tSOk4wdVvhhqK4AyzpNy0vK9ZZyFK6gc
28qdo2XYJspBcto460WDlR0LbDT0Uadlv2Aga06Gw/URqz3vHKZsrW0F2vCQD+6EMz1qFp7sbvw1
4bA80dmw/fcmAYNKXdnxQ1gVOvP5dEVY2Jsil0et9Cwbc2tkKx5N0k7VXJT6Mr1fErnXNht/1iVt
vuQLJfKmQDZD0zhWhkYPZG0TQBqol4AgPoRcZq3XNUU6AZW9TH58iyc1FymRFd8+EETAiJ9B0W8H
EpobtZEJdIJonDU4/ZKdm1VQma0WzCXKl+/mviCbu8pPE++YXAJpW4nPcWsruKtJ1+7UqsMHZ4Zz
1HQ8rZeJaTx1LI4YW+4B1ji2K366rPGqVgCuWRBzHmGGT3JvTMrg+DGYC/JDLLHb/PYs6L0lbrun
PNvUzSV82hRPVoRKojDNFQEpLxPkmy2uu1mWlxx7359pe/126dicrqXFIYH6CkJGLsY1TXTA4jSP
D5UYlRPC2Ocazd32NdNQHtLS9YTESzTNm8hoC/RABTPDYLkwfBdN5ZvTi5rcsEprQXaK5IjqhuzP
oDi6Av9e9+n+Wn9s0Vx0TdDXlAL6ckzBwpEg9pIInEcwA6+n5nc6A2kUbBrfQvbX1/KZsMJjwbpO
PaSbWxV605+FmOiOQHobjn3mcTivNBowUl2cRhvVZ30Vj1nM+NTGT3wIimaDio7bGzDc+aPBb4IL
ZpSa84LCUR2Rk11PU2DGpd89ai65unmb65fdC/AH1wW9gwY991d4MRY1z7HGBd2IUXh3SQx//SYU
nkzvjy7JAmRWZVGjn23l6R0J0/oCaAggqx0F0A6PnBc9HE7SKTQY4zHLgYJAmHCTEF/6MJ59JI8h
DAuXy6uyGi1lxnFm0iEc3dSzWyeyKuyVCl/5NRIqqBpspQmnV+8JtFDGKKuLfWf6wbyE9OfbFOQE
Xpb7Eqrq8icbaOFF+xq3vOSY1fg8epV45J/H8LiaB1qNYldgjN9QbdFu79CzBQgLAT/gy4C8y0L2
aZw7og4AyYs8ulsbG0sWf7j/iD/cp3qQk6/695n6870SVcklAIW6BtRTpHl+7Q28BPbEwXQ/12sD
3/slT+AvlD5fOLwt8y5i73I+qFL5JRhazwgyNBuMLIH/nu/3KuDPPDS/l8v8dSh1dDelQt7ryVBH
5OikuspeSn/SyqSwTf5BiMqgJUA/IAvLDOUHXE5fMGPmUYx63JnfMqnEVl6At7ouEITKnwoZH6Gl
0mL6jRujFGXhfuN1HXAPGvImPdhyBpTJoeV+sEtZkIH8VWUf61bm+qCXuEfciPjtg84QusJZhYI0
fjXjrUPq+sTNnVvmQjRd3kQvcy9g/MZqbsGHeBW1ZkU1zEkR46rM0uGB7PoVb4sDzWLEVYVlEKlF
2fxeN8YIQ48ea0Kyf1I5JMr4JsA/ufwTCY9EaXyvPUq5Jqn+DeFSTfwyjq0QIJT/pZCqszY68EsJ
G3TcU88MDAWVqfAHpWSr6Km7EOTKkOcwjrOqVRdy9Ge/OI/lWW1iNREqgum31mNL6tlkwBYrq5m0
Kw2wW0yxVUS4cGroxBhhf2RbDqTsRabY7aOETmd0RB9p/37sJ8uAU8JUtjkeOe64wQp/s6yRFWMd
JUmHRlO71xYAfZ/3einxcoDU36skNT3+JubLbt9aLjw+Ei8spS/aFh+2ARZfygg4fSHMPhwgbG/B
TyorrC13jMdwRxqFhoRnsaB+jYigcwUVf8veHffz7FI/gQO2hw+03OVlk8jMu4L9UiZGqWF7i24B
+uAX8eY1LHHMMYN09LLAwxsaBJaZuCSI5fxm242d+0twuB0r85HMTYMb+hGa1GmnRs90OLfAXhyN
/MzvLJdGh5YjU0iqN5Q+0/xYuFizSAKYbd/FsXJ3bimvw0hqmCobKI1vYwsDbfQPIOkVmahAxi2N
c3pw/hsUFPOOeG8FiyWGdcKx1wLMz1oatBgYqq/rWYbHxw2ZTeLIvZ21fiyxtj5He2dOp5jxJKqh
79tPd2TchvY5yOFm7CbNni2Y1N+qfR2i8CEPWqlWPg+2de99fwvtoF+HVmxaAQvHkNRSJGmyeoAr
bkD3ysD5VKAxBXP5n3zpxyecZRbgmOniMJWc4fE9DiLzFZHa9H98R6jStYdXiDq4Zf2pz6BvL+yU
/nP1PpIMeYwmgeIqlBMeur4Df6h3NydIu9TCjmkYCFfJSvB7bB3MlBv6i4c/yOFAG7iQZMfFcUc2
7pjUZUGG7yrwSdh7sdaH65kNszJDL6ZwVh4pCzykxEctDEkBw8J+2oypmYFpr2KuQxwsKX/RslDv
gJS90WbQhdocY6Ahz2+MbocX+NxSf/+TSHCaEF134CQK7xI9yvk5GT6ndqfNHo3z05XAgdwhTOC9
7KFASL88ThE8GbVOHiBQoHwLzAgLxjAAwWjDKlian4nvF000mQOXb3Kws+qARtpCh+b37wlzKbSG
FkaVkaVF2JwmnfcG77891hpkD1j/cztv9LVY8XhyVhOybZCl8tSOd1Z76PDjldbZKhnc7kby1t53
ICv6CY6R3iiz2G6mvd52HQEc5u/b4oxNy0geNaFMJ6eLxeq3xkHgRefjAn5jrqLdgQVTyOxYNl9l
1XckUq3/Cm0TeMlmAAH7IOVrJjrHQo87jm3arN4e70HobV3qs4PRhTMw7GJzsQhdVef3pVhAJbds
t4jjixAdMptU+IaqeWGFwTTP/oqAX8eolVni/wpNkE9DhXmr8l4tK/+rSVHxivmvI9p/PFl1oAoK
OieaAQ+exEdEj4+ZX1J/EhxiyPmHGsLU95FdCh1wf1uZcrLnED05p7JxBcA//CZXZneswiAC2qfW
kjf67U16MctTXBXh6Bludf+Jwlg7nfIhnzmBbFCCCvQKnlcvJdSi2VIDx0gvfZXWMA2dZ9jSl7wp
TpaeiqQCkf4NigSUTj8HWXVb6YNL0ybdAiDt/XKhUl0eH9axCAnvoZFCh6QnBI3D+iqsgHfy/X6t
MB8Zl3Q3CyXSR4axtaMtvFxfQepKO0hdgqc4Xc28Rh5soF75RNfU7arZ4z6S4rSy9a7Uu3OYKYK9
eCpjSm7cBbrPWB1AGT88Yn5DS2nc2UKqYwU9i0DGivUAj70ctWWlaHex00Q/2QxIAa/23cwusly3
18dGHGtwFldEmbalSNVInlBzGMN6ATCX+gHINYrr22bcEJ9BZT4iiFCda4iGG5m/om7qKwmZ+0g8
4oEO/osxKJNYPLQFZ1aZdYLuq6INrDU6qTsyOXpKISxhypd6+BOyitxh32R44R1cOHe6aqd7jbGy
M1rrtE3GiAfs6iz/D0Wr8D0+ztBTfel2lcCtxopdo3lPc5QfAfHXHN7HvGjih91//WUPBbubQ9CC
tP16FtpvOH1LAEt1yaLEbgpUt3VHWOloGuR5+uP4TP2MxPIc2Z6yTkG8pV81ju839PBS+Ix1OLtH
vAy12LTSgI3LjXk25puLheqxcubTv6fQRI3tJSmXJdJfSLcOcvyr7ALGNBWn/wWUqPmpji/Gztp7
2zZWvaQG8NR0XCETpQ8IBPzuHJNTQEhRYb4AxgRtp7UZZBdCEbw6iZOvq2zB3mtKWPGGCITuw2tk
md09/ZCaech7A7OqcUMDJEkWZVZ17OpqKG3FdC86hphCndn660Zx6HcFMWvSaCJYWqp7JzYjcfVQ
sPX5UTd2TrEBI+G1C+yr3ovkvDCLanw5+Howx2I5pxoLODQyG5cjWp6ptcGBRV2ZYHn+J3Vr68IX
CmLaCV53rCxA2VtXUznRBHdvpl2vxmWr4Ov2Uhw3JmZpXlsnivGEcS6uRS2CoRYDdv+pnAxXQ5fe
V9pP15Fl9NGOaiOr40PEYEBmWzFtMLnqMxTexn9z6HqxAUPiTIh4PqTp3q/lcqceg9p+icgGYEJN
l1W1wrKRd3LGGSRXRSspLo+/GbFvxEw5mhBApkz5cjopa2VogMXqvMB7Bj7Tckr8fYvVKgnIe8Od
NPt8rir+1eVCo4z6/gLo1xK7hvZFflijBqHmfqeAu4Oth4srKR+9xLPico6ZS/aqjcDgv2qk6IwJ
hbr+TZKujpdNGC8mCzf6erxdhswPvqqdlJGxN/XCm063UhCXH/BMJYWicnQDM3+G/8ONvgNFEsD4
+RwuQ7QmzjrXWaAXP76CIcRQkmckydvNGC/qmuqFAq19k8VzVNiWViBcjMKm9/Lubx4yyJefg5nX
W3f8icwC0oy82XH1TDaVeJ9Kef1zONvUitVsbDbRAAniFWvnMfUFjI1IpL3qjWeg3nYsInVuWV8d
wU4Axtrz8eSnib/j7vYK4VM+cVquW9JBJpCOfvGK1aPyH+39mQOED3MMrs6JoZhjq5g5oyasgCzm
F0uhAqK6ZeaLtw/v537Cu/A09RRbCLGVK3sPxJDaEPwqTCa4daHLnZ0WUJlUfyh+ds960DqpwrMx
lAsbr5dMUG1jNHp5iymMzEzidE60Q22kjjdlLGEtJnENr9BMlieOfqdSjcSuELPo+DEbYk5mbLbR
EIbIzAHg8pcUd9gVxUFZ2TDZnfaXfg4uyxUGkYqlIb8ZQCuyfdssB+G4tg0Zp2HY9yoRyZe8TzNM
uOuVbte7jWDfl9CowIMH7SEH3p6Y2pOytUAYLMUB/KkeFzdc7PTI0TF0XuNXQRJcR0EHojffXv8k
BgCe9MgtIuufZ3u+r4h8CvxN+3GNfR0qU2dTQsZ8+E4JXqk37yELjuuFxoL8Aa8yXfIy5Y3uywYn
qZQ4UQuZWY6SYz8NYoccLNBpIhtcEMSS/KjHJ+9xM0CPHYowip7JnebzJKuiRW5/1jkKPDfStYOk
MWMCOgEPGFxo9Y1e4VU6ddQ2BTb86r3UQW0A8VMRMYeom4mwlZ7w1k/IyYAPO4TstO3qo6AL/mc8
bG2AB3dczArCJruHMHUyATf3pZdvDFAXpMDGDesxt0NUQ3C5nxbFWRERQXZJES0hGvcwOfDJjVao
vvxxPgs9O9oXdIKXwbvAxJUm3q65AC2WLPpqkFs2FUxoJCqs76T7qF0pVZx0t+MaBQnmJEmlkNAV
RGOrwRRVZ1V2x+uCvp/naYEiRz0jy04LyV6gmOmhc+ryAKJmsm1BjCK5YT56UMnBnL4cC6rgYCy3
VGrMo1UWG/yRzd6UNlHAEZAskzfOdy8Xf+hCExS3tt4088fEbYKRPThQvE46S0sVu2BenU8w7ORS
XvlyDWTEaWDf6AfuhyQFzVb6kz/PZfuh6BwyqliYj4xPteBWsQrwtGIchWX1VcPiu4pxOV5YTNaX
F474pMJjwK6FMinbEa3S6pmyAGY5/AznBss9Ra0UUSbDrjTT5Mgqxo+70W2AivLvv2uToCS+QAXJ
baejZQvRfJmu8QHrUSKU1IFc5NfEWLLBs6ZBO1MGNPu67KDmUQw0ZNdMuqwQwAe5BV5rR52wClOv
fgq5OMh48la/5/z4leg46ujA19y71EKJC60jPA+9X84J2Ejya/h2m8K967NZ+Jv2ctwWEuR5YfRk
eLOaz/ErWaoTLsJxXzFFc47B9szIk3SV5aZnA/qcX0HfLh+xSVx18A58kkRazlvDThl9bvzgml0A
bJVRHn3p8KX6D54YXJVwngMSPdW0bu4HR3WttjvQNCBvOOGTF8TkZgXuT/zpElLsX6ZhEk9u3rQJ
PSWYCIoLvo0dbYghZuEWLms5UN1buf6TR5b4nnA5+OgcqHnp468mgIofWe8akpFgFNkQa1VnanBH
lxoZ98Kiih87pfBYMfkEg4nA/UxI0aglYE9PucMl0qYcaOtMCRnLBvd6+/12lRkMOhQd1Y91xp71
F5BxZ4l82mpXBgJVLLP+z1mGMkCc6DXBCnm7lJ612eiH7s9cGhVLRLOgdwrO3tMwtfjat3bBmChq
/3/bXlA/wVHFC66LaKyuEhV/iwl6FBSuEsbKuFRsSzyHhc5sb0KifyVs9r/eDX1u4Zq7ve5KYfwB
FqYQfkKPTKLioHHWzddgP7ZXIvg+9O/evCSYI46uPrDCDxXYd1ypAuhxXqm9DT6rtrmWsH98KdYu
cTzK+Q+D3cBaqGb+2XqUpksZ0O/OyOb80OY/8pizXMWl99h+ESjSaHxQpGGjXV6XSM2vsUR2bYfz
kNZ0VgQFeUD0AAy8NjhwwR5WoQXb2ZOz5gWOC+QGVcWhesnODegLGw4PisjKyMZ+NrmWJQZIy2dz
yOBAOPpxDNj5KQjRC+2XzgkgB9WTElKb5nmJFswtJneUAbL5+ihLETRkVTB6QsSBcvQWizTXU/Lr
i81W+yFpHEsRdCyZmCs2nIsilUXq5ffqvmjzWCjvgqIeUL/CWJSsULSIIE6/q5nta5MYpX3uka8H
5ye+lNN2wC4JkS/Dv/DxzUCfhwJ8H8tDaqCR/sbMSfaEyYa0RUmuXsYwlQFbWAUq1ftcs1OwR1Y2
KF3jeK2GAxSiew27G1FJyHlevifJqOJG/J+KBIcQJxkYGLkArTXgyZmnFOtlV8XwX1pov9euPRyi
J0vJgBAfpBi4CVswMpB09GfjvQxVaJOM3Begk/I9rc3Cvz2+Phb5hjMPQA8nel0oBk0SY2r8aSWa
t+U4Os5EcsLeOVY9k6ve0jU5rxGuch1zMRt9wsvM1s2rsARE9oHyqSMIL0tbRX6BcUe3QcQ4noF+
JALIMwBEwIXvX7HrltYOwCUGfn3XaJiTVZxVTmBV7odzGCk+u18yoEfLrqlX+jkgivlPSTWsZ4CP
edBOZiDjcnwu1YuFSb6Nbzln229HNCcKDt+HvZhegV+vS4k9xGXTC66fDJVpIvIwKtpR1UZ5+WG9
9/M1HoKSlhy2/nqk2Wg9elA51mnAkxjt2eafoaRbM98lwZppWakJvnfgplYjpSmX6RY/k9thNrOV
Qtp43+lYa7fe2M3JU7uZzAZLGeQWCZk660p/W4UAYkQTYWrRKefyavECpcj5TvLpT3DIVRikFeUo
KEeQ2yjfTy3VBme9kzaJRBfWezpYj1Zq3BiAEsB2bqZI31P0SV9A1WX+9asxxd+mHeGgZOSIS0p0
auTKCHq9Td8pXWACBD1wiFGp+3cPfyBmS7hMYN7L5c1ZgoF499bCJt5jLXOXgY0rnNizwnH2z4wG
MZ+d2pc9bW2kLk9MpRJjB+1RCOMSRuhdJctp6wemnHd7aM64iJc3WozPu7gO+WylQSu9jC9xon2F
451kS9cBkZwq0UPpudLICnANVeWz7I637cKnzlg73FrgJQ3rUuW02D35p4cAzIvb6L/MRjhHxHoL
S3fgW2AUu243PHD9K8Wwyw2fXnnIGPdcSywqU/1T3wElscsRcL7nAHA0yW3ETQlhV1RlYnKgp0vU
P9wdpByUq3xDKZrR5j03vYVkoMCOVds9a6ZtosYIlff+UYeELSb7xXz7vO9n/uIMkE+0IE6nWl86
nHhZy5h43XZrthOdHeXIiARGyzn5IzkoB+Dmd+YEudkAaybsY8p/HKBUVQ8MPvCqnBRli5e1jEzk
UjuuOHtLkBqxDOoOtUf5kXnjV9wMPHeP3akje9/bj9GtvK6JrI6Dl8CeX6vRL5hcpasaJtQzsEkI
KUHyK48cp0zQ17bINw6rTyrY5br3dmMPhWBTaCUOtyvXSGIMqNwAtgVCVG1JortTiO1jT1yKnXds
EEmlNQCFOlJYKmrUSsXL/MTBVqp0YT+HnZ9Ny1tdkXwyWgcPLoA1M4XVJ8KuHk1505ZEBYasrG9w
dFosNYy9iqiWZ3gXrp3dkcXOw7o4sy9D5T3AWM7FL/DExwgbTEm8hA4LSws4p3NyOtpmNkVWs7Pu
AAmd2RT+goXpx2uZorMQE1P/IZhpaVHAlkuqxumicORZ867AEs4Y+XlReN7o30iIXSbjMysd3/uC
5VyyObB+fR52eEsLnX8ZocRCXLZSEIOtNMl3DrsqkJOBQJvt8IIaDCk5IAwkT6WgiCygIQU6GYiE
fhdjfpOkV2sHE46ozssipYvMbRXFzw+3yXVf248PitJWW9VXovaiUNUg13VGxLjW2IFx6rY3m+3S
0EY+AMjtFkvN7UWpdz3LFDEePPzMr2kMHkOeaumYKZby+pkcB2CgOJeunZiEzYkKpd634huqyehz
Mp6BOc7uF3+Ha4soZjga3xepfjawdnQhhxrPBfUxrr60GXkriFBj1IzI5OqyZp43gGCQUxdXaPhA
LFtJuiN9bvcplUnc+wM3MBwxWuU6zUX6vqiYe+zmXavU++9vhAzBRC5xBUF0X0E2nn1kwA9jAx7P
A3YSPOzL/HKes/Th407LRWS1OUg4Z1lA7Wd3cSRLfeBb3Y1vPoltwVq5A25RDYK77tmR1z7jjPAM
sDwooIx55+5XafjaqDReO/yv6jSSv0urnDlphxvenLVskl5qZBgeRrjc59N1t/vFvwhUmcnKfV7J
EaU8MYS7K8sutDt8OCXLfjL5QlhzDSOG5cRUxx3Joy0dgtbK0hUixqr9/aSTL3GdyqpIM3s/mjxm
w/SArpw74hY2kzdi8Bgzb5iZInraMd5xxzW+cwk6NOiqXmN0jIY/WGzL9yPbY5soZfx88l8jyhIM
j2dN7B7jRdkhPJaCJkViX1cTJnL/PhZYTu1tMY0X5cucYnylALYImQskus0aOvXJWXEeYIf3q7qV
su5Yhy7mMsW/FuKk2VYjl3W126LcBxy+ydjPfe/6neBN11AuqXqxa6trfm6aFESb5ZceRn8bb0jW
SMUWpPH+3MZX0Urc8v/ONRQ+2Qsv8YdT14tzcvlM+QPuweqMP5r3s5rN+C9i/Yq9JAMteO4s8nk+
6Kd6tJAiCcnga8kb4KHNNef/VEdBIOt9WseNEC/R4GECYAkW/aSLZ+FW2WKfKKVZhe40lPcaSTZb
d8g0TBv7P0C/g02gIjl3sFqv/mZ/aAe3KzTKUP2iIJoQnFtP5TqjLzCXV+tgEEZCwmqh23n/KBfA
O6ZzCSaUl/LHgPtDHuzWcDoVGEjPPyFdPNxI6xj6+dGvu5zuholcVwVq1Kl0+mPFKlEC/et5CU14
jKpYk2kNi1Ml79JeOWXp6Dd+6FNXX9FK9xfH3yh+9nJPEJ3RwW27QfQnhMEymNom5ZcAsl0T/ukc
qM8I6484KpwGmd/PHtBi4heyrVTRkI0hWybJk7wWG0seuWjbs3jcNeqKVjzMxViHBPY/5QsI/Oj3
7WR0DoaY7bLHV4R94KZu/oDwrtg2Dtc8y+j/wk2OyAZDas3gCP0KK/T9s9aeDZenryKbLtbGmXTz
kpDU9Zr+J2/rLtOMMxMf7bUwJauGbMYUEqMEy8zDlpmlDJYZ13FkWCRpZfGvnTSAkPgj8TdfUU+z
qDEn+3p59IOe0Cb20cGAbxaZ4Uy+D2JRh7k0BuKJF6nwCf5popt3PQgSo36sVrh7rF6mFlCuEcFD
nn0y6CbhWOYJXpOar8emlML9jq8QNb4EGa800B1Y47KVJv4TjmfnRUH2q8/mAuxbZrurnCZXMt9/
MOkvpIS953yEeQObcNmyBNxTlNrn3Eq/e8QRFeYf+2su4hxyNEkmT9nlfoj1mnf2EgfyA1TJyZm2
rGndGDVElREKNUBRPItwEUgSHcnr3LGaNoRoKPAW+otK1mLNi/G29lySnCSpQ1s9UsAIcxE63n5Y
XfEvkNxrIHlYSvqmbR59e6FIjZO5bruD4xPRzS7iMr+NHVGwUzwv/sqRo5WCdpAtV1ZSrU/9RTNp
72y5zRk17OrV0p5QWBnvjoUzEmmJXa0kYClcqu6RyttT7GUuayLTk6KJdqAnxGRwHwVTfEKLUYd1
YIZ8tFg1uG/5s2Sr9gPDJpWw+4NJFRQF9h1B7Yp1c7qUjJfQwwK4MKrqfUjHbuyshhJ9w02TTKfk
ZpwtxZOISkll/8yxhsdqFnO48maz+qXJXWq6ayuSOPFOdG6xi2l64T1XJSWYb+5Yc6mMbwOnaNBw
hNV5c4etl/GXKL5EpkjFZWJ/UMxF8KSifRa2OOVncbp01yyk1cm0oTLCqiDcyoJQC0mnezREHUJf
TwFe3bGUV5rKX+IqDFFVh7fljPLhuzaTkIp5pZiZkNL7ArzbYIkMSMjFc0ydJoSkJljZSEh460x3
27badxtNYw/lq0jlRbN9UtAHMzWnPaQayGKFhBe2iDCb2P0mdEzokC8psYftlVvS/lQFqb7xvanF
KD8KBN1+AL5KoU6nXi6CLaa4YX7YQ1pGu/Kc8IqRVgahXR61Fcvls4v+NpYtSFAqeG+3Z0Q+/IYB
xVT1U+a9ivrGTmRn043koyTWcRVWwVUF27CZFle3GZI3q1ZZre9oZCmSEZsf8zwJDrmskdOsr2iH
9bJaHELjzOC3paWDmeGh+R+uZaNUvs+m9LBYCyWGHjt0ak4A3lY/2YWS1BR5KIL80+7XY4aCB68x
zKG8Q+2AppB7NHdhfLDMWMN+awlnj3FZoBi11l8TTdzgnHkLa2KyCKX5WJJvDDPTEv/w+nb7/9Kz
+EQetjbpOJwC5xOrCaAcZsnRnB2Jai6fCEiskSYGY1FY2dpnvm/gBNArAbh3psLgImZP5ZaJ77H+
5i35ptMjQ45AqmbRI3+UV3bamLLPkf4rPguhxo6BeqP3FR3qTRLijSYZwHQ5MKWRrmudj++i27Hu
eTJLNNsQyxL8rwsD3vRP8mr/rkAdNC0z6IhfvehDFXlgkfOhQsbdt08GJAdUBwrGDq9FvkEdNg47
PbGKKHyEC5Qw3ruYZ5fLUe5+cshIw1eqieMP9U8ryqcCoLEDalHx55JRMwWCG+G8h0jktGV+9Qtz
W028TlCHzVD5Wm2EhsIDCNeZAJSycHQMAGsu3/6AkUD8lR1wtYnhdywRnwZBkfJBdQ1ZRdK3TVlI
0OKdQqPfx84QlCTY7H+OO+PXEXuGkf98j7zeGK5fehppBOiNEHA5Azp6zCHpjaRfHOCX5DGGav+J
5+K6c1DC3jUUsmyhrfqd3KKVkzBrtJSQyI3X9F2kf+2ikszVLPBGOWmR2sav2LDKvxh1z59O4AMG
K4+TuSrlCK/A4jnQ+oyj9k3EX7DYIvHuOz8bEt9CDE9CEibaSrY1yTDKCXDlCKP2ipkAU4m5/waY
xTRcTniLm72PRCLIZyDcisftPtO0YOnew6XJgwrF1052Rjb8Pe49reYYUbVm13zM2BiSmF0jecsI
/4rejdh8bPlD/FfiIrCs8dhxFstP9gmRONStFCekrNYtPKlvbYd8RAqdCBdBDp5Sozw7w1yySeh6
GmTTfM3XCRiQwaQIoqRzeH1ZzyEbOxabWO0qEHKEAXf5ECVJS//OW3+K16UMBVbSk30nGpfJ7EGq
Xo3ccIYVzExkLlnPuu2f9KlrL16PQ1biBw7bB89HL1Gy1iW6SbWYKRvKVpO/9ulm/wa7vHj0X8nh
3UWPbsX7fsd/cTUrIg3LY1EObO6/CxfstQw49NgzWAixHwpEdy4YlpxWvhd6y70+jA+dF0JCjT9G
oVzlbHVz95nNHFizlXLiQjUOmYo1NWN3euB2bGvqv/mx5NyPSDFIgIrr2FH/HQHhJXR9DECIcM/J
dECITNo/nCaJdfjeLR3SVRHhGlkH/Z26j6/s1HeuiwoTvZ/84UO5EoDzDIu5UvJIu798wkSBSyKJ
JkqoK8XNgy8Vm8DojWSPl4/AZvjPbFUyDnnBmQl2XOEHOeBThFcA+D//gqaKkZd1ZbBVuERjBuGm
83EX7bbcUQW19eF4pMgRAqyKB6nJRQ6hlVYLuPQDRBeTWJgvvmOK9XzQbU/HgB8ynSeXiU56RRxC
By28gP0fCW/bLQyp44gNdjS9Omy2MA1zUrTC21OOW8Gi+QvzfP/hnNbXlU6I2R81Y58tX644IUGl
bttsXA+DJWND0Nyjcj2FuIqgzs6KeqRHGcGkODzClbhL7f/EaI87HlBV6Kad+XgRxOc+itX6Ah4Q
VmtVR/kylb0Vbvn/2L7IYafBzqY0CUecGDNsmp9jzVxXxn6o/GDtS1jqoxEtlM2QY0tzJZ0IdVSf
sXipAikhkpTH9slt22A2o7RWaksUN75331o4EVFLuHAjbWBRKghdNRHATxUKeNgVLbLorELjygl5
XCtHcYVp4NYYJmud1vqyeuT3pThoesGX4RBv8eGGOIHOCzhtUAO8txM7iwLRQB8ikw3OQEeOS5Yy
D6zerkV/fgsbxqijYxkMC3nPnrMzAMhT19XQe4W5qykcy/vdMhd/YRCaDoEh/K0kCfGg9Ys+1kec
e5yxzGJMdpfYcmfy7fimpRMOE6PWrMcdnT01lIPAn8X952J8dVvLSNWkzyTYGc/7OXjeyHNc73iC
LrcwUM3ib02SGrFJkaczCogYdA+syiZLSig4rtsa6KLUvB9Z1r7jHLdzPxjw9cQvKgm3dTaIY734
gB7+x3uheGhmTMxWxZEuVG+ATc7EnbAMplA0E5Osqg+ZBJJhdqviEDHW3DLKWiMCH9DIxUApkxw0
dYSLHLMLeTNa/NLz6eiP4a8XCrjbChkgrnOykgbWEaDurX4LrXj2U4rE2Tdomyk1nRHS6z3DdBip
rIYjhTd5INS7SGhsrNdxBMGxXftA+2OTGaRiNKYkwn38pY7ux/Wg4jql90j1wcKNfcFZ2lhnRKlp
W7ItkIYCcF+ogrnmV1fjzIJkv6SQaP6hkK5kQh05VEB3hyAoRURBjWae35xqBSCqy3tDCT3gF5gA
NOXK4acLLJ7XZdXeg620JR4RCdRqBH5jvWJGSygBIbEMbYKaaEsoU4pZDaB9YUgVvA6Iyt6ozzle
gfruTLd1DiVshiNZUPvlDG4hvtxJN+2bfHu6PrCC3ziRFvh+vS1ofjC8ZX8LP6OeBnc1wiAZbg1O
xxC1An51BWex5/b6yWkcwdsnNtYfvogc8NKInNJvONR0WjG5kBKatK+szZ/rk3lrYGt4hzrFm35D
WsFg5DyKVY15lZODvrzg9ms2PvtFhzk52REXcNohG9CLfk6g9sJsnFGAugOVkJKICsSpwNHxhNJz
YGzp6x6DXPjtgwWn4Sp5NFA6pVKSsqixLJOMNkNcqcsXeeTK37QsPMpmgOjttkXP2q7ilCIpwL2V
222ML8I7Vipx7MtDhg6IxxgSYrBgXvRAqoqEhm0V3IwEEuLEu42z0Br+swE1goTJu0YyQI/evWOu
kn7d8Ge9pN5ssH/T3/+HL/ueoEnyqgX+GOPf3UdayfNQB6Er4YgO8PAcTL8XIe4aINNqCvzt9s88
lTNvAmFderyO/7nf3Kg6i9Yas54v7weGHn5gvRq5xdUjLLfX/sCD7I/W3i3MowLkxFd1RaaLI8Wx
Ky4axRvmRCsueokfRP2+KCvq440dtJuyPai9lUdHNHQT+qvThP8q/TEdGOMELBbklx8uzanQ8QA9
6/XerhGWheWqQGkpl1vFae1ciOFm3FYZVkmYziI6CBbFpYPx+r5u8HOcAcsY2DbKbncX8i8Cxr3l
A45Hme8dX65f/04iijKyt64YPcTORzh/jP8gpKhwnHGG7kRgihkVw9Q7EPu5ofarQzaWc9i2eMlT
WXDsnuDiOA1ZG7kTIuqhYk6WLb6BRWEzbn1tlX0RPm73QeBqRYKUCnvJWGvw+x62FkrIr5io7cOX
qeSYaUVOi/82U7pfx29bWOsOwNwBUAU+AOtYiks9AeEq33Jr4BLcz6lF3bZS6tdI8Tv4zec39taA
rtZc8qqIC8odAwrN2abA1RyUjAh8QYgLbr4efvL/M8p3PxqTnuADmlyLrPVFLZrCJNLHVXllFXk6
a08L7HVsYoO/tCK7c7DjCqvialVlLyK/Es85U78MMesZ8zvYDHbjpxavj0aF2X3JwM0rEaPRDTCQ
lYqltp0dkd9cPQ9EeIBH/0HEuuwoae2CVwOhXWyHqqLgceKsqILBmmfXUrG2VOS+/5R6JWKaouyK
BPHRccpfSrVolX0p3tb/gbphXzFpEOLdWHWhk5O+jn4vYwdf0Q+EYoRcOCeCbI2kUKSED5NJ2RRe
3unBrjaFdk/RUwcuW+jJlOc0Lhk7/eLHJYnXlpnDGKDpUS/MRIpzp0GWCDMHAkbC/ZLORnMeAknP
S92rjy9bnLNmWonA/UUOPjohxwvKGu0YHtS8pRC2Caez8VcFl6/GGYx3dE5cFYCiAzGXdecFFbLr
J3SjcAa6NaXSgiazLEtOEEPUa1Le+VEd1SglE7fDDfrkuKSYMBhl3OubgS2lsf4FeHV0XFI0RhKR
Lhr1kvx4Rms4aA3uBNctsbOzDMSAiX+eC5vYZEDUJIY8sCw4cEnLbqEAOeLOPGvfPRHmClvHJn0d
BMb4GdLOhFQI9/g79TK+fvF1nIdpIZ+8X4YRRiA+VYaWvyFxmy5yqejBxaVAKPbnMIT2jgNC0m6x
yYCbDBjksvDqDccYmtBUNnePI9qyqstP9+XZsk8DSzl7Xg7LpuQG7ZPUSNh/Zb2fuQwn0e9T8QnT
276/bjzmToLGmtDpurX8A5IqdqxTNODGs21hWXQvQBn/mnWFQkbtezk5ZJ7h3bKSqvZ973p9VKF7
jhKw2PPSoSQLdvwLjVQZFqadhZKUq6ceugRPJjmtmJqCUE9PJt0AXEfhZJNgs4fvAqcqaxspjcTg
KcWSKC/g3//MVddRE5t85byJsgpr8fzZp1KAt0GmEKUsyA+fBEdAF6pw1iWBGF3tTcP3z6MB5s/y
nyQav3py0e78RIYH2CCAleXWLS0pCW98GISfOJVtLEcm7ulP3L+Oxdt+B+REn0QTNEiRgCylt9Ko
I4MqnYOYVtKMxRwdMxZKdSNdnJPR3k/Yf07irNPA5S79jm+7zJ/C6a5wFRiFFlJaegd247KqCKvF
TWeAJD8ON5757J1u/GCDU0kFQQLT03CpjIsu5XQZS76s4m/dcMn2aF/35bYSmHNAGyPMye1cRote
C7fSIxXfPNPpzzZN1gLq1pSQ/DNfBChAVsJalfp1nGM5efM+X632EPBcA9BcqvKLtt3HhOTaDkYE
GXXJY8gKz4d1AGCbJQX6NJjgeFd54FaBk2lFHg8gY5tfPJt5WWvsR7dJqXFFy5L4pjP8InFKNbST
t/RQSrfmaoILknG+TTU67rwTJ/Cjm3tDN4i1pCB0Uh1oozadxIyrJpf3bdVRrTYiK0iIvqv7xqCl
xVAS9SNwVuccTaBSCMA4L0rfBqWNfpR5b84KXnsuN00VMhaEBIgDomJOuOm26v3D0qArr6zDE2aq
2qa0RUJGvWIqal7DT/tqTQPVKEUhYQ3rqieSBLvIggPbyfWH3klXg+r7DvXfgV7WQQeiORkavcX4
QtcqWLaZZnZq+fnjQfryXXcAFDbpvdSShqz0+FEHUYc1erhwDQ1mD7kRRebaW9Vh6CGnJwuvGITG
e4U+Fy/jPwmdPkcYxzz3RGd/1FWtJq1Mi90GW7sPfQXNdUjuJ3Ahy08bIp+gAqM2E5fGwEQLZL2O
zPBIdHhk+KcuZimzoiDiVjg/zhfg/GljtHzptFIknB1STDeL209ZPUgD4Rd2SavKhdDD1EFPs9CW
qXQhN86Dkytq8AqlLhvKRQkmfsJQZmwEerjqGElwgtAx6rQhZnmz2775OSGK5DQp6wnY4GdyCs6g
bwBC81vso7n5irYz8ATDiGZtJEKXBt72zCvu4JAm24ejZlIw7eyMV0zJ+FqvS8hGDUy3y3U+MaQr
TWPB2X8KH3lX8vAEnHBBTYykXzydjJArjT3aAuYI7O2VrTBQOa5nr5EYluXzri33NXh95JN6ah4/
yzjWHlSuE9+pMqBiQjboi079NWNzVRLILjoNfGF2yXTcGFr3RnhyjcUSLPjUhhr4DeF1FGLBoRWM
gHMwgwZqBwJiyCR+h3QlSmot7i4M8dbh+1ktCA0qse7QzoQHLN+nXo2JT+1BOLHNBxrO/VeUNtkY
t8Q3mfQAfFEP7/2zak9IzS3ySFkbNNic75YVachVUymSyUT32tCBshXPBvxXe6qtCKm/SIaE3ZIN
T6IXsxRluLj+RqvWHqC9/V8Cgw2YR0lERkN/75B3bVvzwRMFHery/S31hLIY3rOI2nPAvawz/WLM
BhAGJLK/CMBrlKics0sLH4VHYIgor0NoIM1uCkwAVGpRO+6vsATUGi5iOa/7EYl+cGC5mNYKun0E
p/ShAX64nZSmSuLUsaFSx9skuK7ePvx3BK6rxzyZMOU2C83kX97914d9yp7Osgm5XpkQZmgXdV1u
PIs80JOYeMjUqpM1Quql1bnKa6ZrwpVTseqmoEu4NYXW4wQFTmBrUIhqXk9cgzi3ntvvRQMVCoAm
Tnvi6FhRRll3afCiz03fHYbTzR2B0lGhWKM7QpV541eYfyyPaF7/C3paVNP1+aUpAR886qTJSQjK
i3bi5FgVeGYSODlr/wQ7tk8iGHz32gAdseJLbj5eowg9NLJ59ZmEqy+L3rKHNs9mmblp/4+9YKZo
1jlCOqUjfsZU5d+Nt42fHPVKad7UJ5W9T/awr6D/Apxwhg2MuMzmscvlc9JzlH4iusImviuTOXav
Io9jettnbj/VI+x3W9lsDlMSY6sEGPnsnUm/mHQMISnGjhJxqtysehCxLj08NU0qhTwHJ44YprR+
rrgxjIRzw3oAe9Nycw+xvDb4GFKqYtQfT9n5ILnjt6uTcaCvS6WOgP/2HmbDcwCFeQh6yrGT3N0O
XEOUvy7wUKZj0z5i30yTLnrH9iusOH5eCH4hiPjy4+WP8w8Y1XcOTKhDkIKdS9jFD6v0jGkHm+uf
V0CQYx7Xzo2B1ulIb39n6vp/q1lGoTX7ns5I+WD9fTgR9F1v3w6Egg73lXi9ogmyBrH2Yu8ozS+n
YQBX5aejTDXTdJd/iJPSvYkS9HCOYhuL8a7pjTICkHwK5bPl0Cw0c1/9Wv4RwdWHWjs5kaFy5/f1
Z/NMFxHzinIHGvbRo3Kqu58VXzMIhnvwuDUJ/B4MLPqe3rfBBEBslsHMkgvU4NnTZu1eNpE5YN0+
w9vqOS5U46oEuF0g41sLkqR41bh5M5AtZ7p0jB7Zb54RTvuxGjtlBjEHnvu5vcJTZ3iu/b5yrEd5
RjuIsf89M9IFcIB4ZEitOSFUh0j9Xh16gV562F227azmGCwv+8nrwRaCR/HnhEZT/DuplV8agykJ
Gfnf2eTMLKxYAZ/wrUxwkZWBPeyvXRDM96h9WvDY/eHJTIC+Lc4Icn3TCHSw+f5mEMjJl3ELdju3
S8niB+8gIMh+POgRWQtmBySobS0yUGBpgww3bj1PiFSbbfXcTEuhs+D0R1yAaXKk58jTwPfShuwY
apItxyTZYeLvdYwQt7XSoAizVvxO5BcDjxipeqfj9/K/D4aLDwDoxYBw6j0ZHdrsnq4zKZRnNHqk
ty88vkQnS7uyiJIWmc2T83pl5wCFeyF6tyi1koESlMdzWNBkOvZnWwW3qxZaa9SpEScLKyZPnDHX
7V/G7RdP3vCCOkNqK/hB2x7DAvYEeOLuU8CFfKkv5QGDK2P2SdpL3Av+v04QmiVETwL88eNOjd4a
2KiSB5ea36uuzgV4db/NFxRl0kWVYNRqswb+t+qSv6U+8kwuBZ57T21entG/4pXt0yejD1x4iv7E
4yfUEKS85qdgswdaEkteN6zXJfFWC41vag/LtoEBwCxsb4YKjO7bvnwZuzMtlSZXM9Eq7oP1SPvi
r/ggIX3edn8ohXhgcgP9IukV0G8bzvJHRgVfRqLXWk8C7gR/apEQ63TGW6k6SGeC4E3A+A9ZjZAu
JIsGUYWfsYJ9b5aoGWZ79T7YZU0140iLCT4HT55JoQK8AMt27fD+8HbNKBy4QzU8IfmjJoT/Kfvj
X4/YQbLbNS+CsniJKkLHIckkHT4SPABvEo0c/E276wHhzE1z4YBBRiTY5OyRVU0b90WzVFq6mkQA
74WuR8+5GyCVm/pqVdjuh9VInx7YFrHhhQuWcngRcppUgMEZ272qrqvxpMgx/bZcs9u0dXRq/08x
5fi07bQqInb5qWXg983MYijk6yHDZ68Tc6KcLcBpBKfx5yCWXfm6WPFIHAMJWhWsqZQvUXfLmLSk
7Oif6jRK9k8zA27aUyueM1ESrXBWp0szsK8plPMecjogpaumzqQ8Ka7iytl2WZkOP/tLj376BoVz
+zVZ+2Oe5GdIl2Fp+O4ujeGIMQhyPxQF2BnnFOpBj71j6OonRvzPCIEOgWhDxkg/SL8qSWgiQfNd
KJYUDkzdfQ3mSmtY2IlFiz7sulMS5jK4eicrfJc2X0sTjaa0s8Y9MA+b2e2xGI7zNQIVsuHABgsT
UMizUVI+ehh2Arae9plvdnVGv24Rg3T4VFQluaf+91QYmJVfGtSAbM4uWMJX9TMTWe8RLlgGTvbE
6Ah/KZs32MGMdZeR+AhY+F4JbNFQd6bHGQnJrjBN2ycqmf5mrHHEvb+7SBkVF9Hm0NqaeJjiHMbH
06jyegzWIqwAOXHgxNkYn5M9xPumza0a+XUAgYkm/RzhSgUsusOoDNNLXUqS71LGUln5ZwlQgswY
/MJ/qaWTy62TCklXqeoJCFiiRA+c4Ps7EAvZ4L1U+HUi4x9cipJ5AEhv2mrEkVhZ9wU1+uIwVk52
L1JB2wZsoHxKEaTXYAi+NokUcIoi0RUNgLNCLhq8BLSxhZG+Fru5gIuzaWfcyd16bY11zaQo+FOx
6LzLdSU2H1+as478FDlemgVi3U2stAfelMPG4Wd2XqLq5YXpgozpkqpTJBSkRaJpuy5dEi0cPOUW
70hahezqOGjToLDiycB5GpR9cJuFRhuCSZOoD/ZRE2+pgtU1ZNZPyuwfaEJH5go2LH7esqkV9VZZ
2sttd+wKXsHJF1ALS/6pfPAxgQYOTZ3FivQyk0nrdD7Jacu5Ma80zCZn1jK04AgopgZsmq+gr/8b
sF1NRLHQ0mE/teJ3xRaCFwKmwjGNiAp5ME+OwDvsfJSeKFli80hHAGPligwmfIABoil747EdGZrH
2WFeir3m3VuqwrHUUm9yc/xt/0GCzU04nfNzwOtuCkUBsrkQlqgNNe5s9K6z6390J85Nt67bMTUe
hTcRZpSjYXYZhmA5eaOaa+VZfjCt5IDpx39CHN4qdgqbyB718Y4VVpRskRl6e+9xIxdyJGzjSaCI
HEbaxpRiPP0bCC0h9YQFnur5sm4YKUVtO3P1qW+rXwej5FivHKqwauN7MVOInUrBAr99qWpocDME
naLw8t4zyjPJRp4gpiSJGL8XYXYm6u7cneimL9HDqkOvZsFotHUCAjPWjPDmshOUbAnpuZSKFJ5J
/suFa7vAzmgx0w9Xwo6zMV7F5RwyOi3sz+56e4qdNF7U7JBrvNjef2irU4CeAVXG+/4Z/5NP5U0l
72xO7HOGQnzPCv38iFrqBsWyF+zMBih0VmvW4wTjSUst+xf2OcMAPpkT0dGZFcvhnONPhTUgKusA
2efEHq5v97gZ0HMnpJ99jG9/D6/sBVMdGL6eICZO9agBo3+7RKP2MujNBn5n0cZnM3khII6bAa5H
I9QAEq2WnCPLbRpPxq5i8UuUHY+RDSBnWcKIk8Bc/yDAnaS3/ZYFyoMJH04Cant5G4lDl/el+Tee
nbqGC4I6MNS9jhQw1XCcd2EnOWSqMrsPh9p8s8nFFDP3SW3/VAUl94Uqxkeqmt1pcEwevfO8BM7z
BB7GtdxVUEyGIrJNDc3UBWwiaF5C/wPjTcck69BkO97pMCWxex7SE0sn63p/K3lyu8oYJZY70Zty
NHopIPkRYrLAKVnZA2ET18dJXBuQ5bUevfCEPY1FxZaamVFPOvmiXuKSL+jygMzHMZU2QNH1dBNI
CffTVGZJMplCPfiZUP2XhaDyr1s1ke9t4kM1PzSI94tW+pc+XIvaieMNUBavDfvaKXcWCIoO8hNJ
535CF1aheIFNfB9XgC2pn3YyL6n6hOoA2+xSRKtfPcufuFKDx1KU1Tf2SQRkRuMcYL85PxjPKldQ
79clPbrNjP1wLDyaxQK7EKKrs7lxwERvx8SL38pxpfbZIGzKrXIiKIDYTV1FcObn0uvqR0DLyu7M
zyy/n96JfJJA7CJUMbhylCu/TEL3aUsSE+NogABF186jssxGZYtfdX923P9fNkpYyTIrRhPWX4IY
C+AJQWt5aIc7bjYPjBnMJUdchc6uYRw2zBfS9aEBd2Nsm45mIbgd43peBTBBHmgy7qAT2vArzvNt
seT5HpU2VeTNHx0JaXxIW88/z9T4gXGKKtl6KlWtojWaP/oPaxLsG811B3e+KTBx2nhEuD41c0ka
vI6rNVPohPGtwQPW/CCCvEAiSel8UDqLXqFz77wYe2WU/mwbZjO8ITOBerJiIyoqFaIRB57cnyOW
QZDt534kIj56w58ureRIPHyYvC1jn+ES80LBbLoUVSqmp1n2N7/30DyttR9w171iVh6AbCibTm17
J+OkJ4EVMFYCDr+5gpaYpJunMUhKfCBvtj9u3bmT4pO7K6XXOGTKUXrvy13lTbKVVpBVhg0nLXaP
V7Iu1dA0ocyJ2UmNbeBT9sYDoVFChDOc0NqoLRhKZi6R234mucocPX0rYz3DkBH2KlUhcmmc71Ak
8yyTexxYxcY36iOhVsTfFqKx1sRQa6wg4MjcUIlQPTAz6fJbdOZzJI3SoT19BijVKBHvYuN5rIp4
yBYcwKA9PbaCn7uK3exMaQNVOdE8gdjrMAZxyo2QNQTX45GYLlk+y+5+bBExtEM2oFQXi5AItUN7
RKow3kwlfnv68+hNDSGYBNVKh0M/fA/rG3Jv9Cw1gjXW2GPtHvEjbncauN3jPNQAgzQrz0xVLyiU
31a1a+F9aLlXho6D+sg2FhZueydv954RyN/n/XBuLXTetxPBXzVIlB7ZRqJjJUbgX0vvo3foySoE
fx9E7CrOR0hvhTJzJlDsgQRoL4uZgkjejeI4ZRVmyWEN2I2QMoezCAYljY6BGACRuuqz4K+d1r7C
b0N1Zk9InebWPeh27y8IHI+3uus8bS/1jwasLUsrwxsP4blwPlyQMYeXGIYpE57l5i5CWWaTsaKN
BRhHsJF2PmIc4uT+jsoS9vuOjNvloxasZVubm9IF1C9A/4plOBlTwIEzqn93InkyltDsvtvZ+hGX
wJiGf4ySrzRwfxrFj/1jqaqdwUaa/YDLNZ+YKa+Cw7x9ZBJ5y1C3i1sz9YvCgxyC8kxSZjTE8QYf
g4hXjIKoC4RRhsiiv6jHsgL0+W+JwChzoDckXkhQj9vp9FXBRY37sW/htRr97+NDCcZVQv6D3kYD
kMfOk1Nxr80Cc9rrCE485SCCh3AJBe7gvuZQHriRXo0NJczSRn/SEDQTLw1nvfVziV8Yf7Q8iiBi
mMFdZ5iL3dXYCrMi80EJyInbWxmnZMD/z5XQDFAOFQPWTOby6y6PAbAbkqZfnmpaagY0g5MX/S+d
U1MtRKvO27wmxPMdzRrSUYAarSG7znayCEq48jSvcVBeV9g80p3jr1RoCT8m5tBumyvSf7y528Fw
s7zhaeGu03fzq7YOorqfzJFtiJFsqQIQrgRKtSFyiOG8c4RhK6t7OWyD+P+vjVo/8kPQaCLJROx6
+u+0UiezLbExQRga67L99yG+IxxECbej9FHqMeZDhqJjqF40SbWf/NQN2YiqzDiEcG3ktk6AF7jG
OF8Ce/tZomR253QpX+2er4z4ZmneFCf1okB+ZmBztneRw0o6r3OGjzNaL9ZvFetE0Ew0VgY9N6DJ
e14FsrKXe1NCjhxPsOPJu7gEstyPVyysLFCXDWoLfm3tjjA4YmsnYx+ufyXw5q5px2DPZc4cch88
qqqkfwziRtuZJ6w1DwaFycMNWOOeV7nQhzvnDtss/dh1u4x5O1mTmG08Fa165I44DjdXOECBmKA6
Mmc0xOAAkdEKo6VmBH62NhlwwcDjt+Ts8OInIo0K5yFJdD/tsBSK//fNiebAsyiQ9hj6u7PaItbd
EDMKDk3jDR7NhCiV1/nWymZm2amaV5k3YcRmsdqBksZfZNi4JpiXtvZmZf8U/ohFqnvFIFa/BhoA
mJFDTh9SpQjVIRN4sRMybEIgtf6Ln0B3IvchSLPUytW65QuZcvvfJC6lIEiwSr6eb/krNIG1R7KI
9WEmoYKNb0QHIp4ybUcMfFHkmKOia3rNwfwKSG3bHTaHEaE3m7GCakfd5+zASOxdwhSrk8mq/L2G
xw5RpPZwdWgWIAvOKzhP5X08zZEaqitGFbni6k/jPLQWEbkHJl5y6p2zbO9HpMEtrbGKSgx4Z8bL
D3unQpK+1GHnPR4rXHpZ1JYM5xRp2Hz0QYuPrZW+xNr0l7M5fFS7+ZO0AuexmnIToUMCmLZ2ocUE
1ICNCtDNgm/KwTREUw8sjbY3xGEZF/Tf67y4Sye1A+FryyiGf6/SU0zc5gT958XOJZwJdS/zW9h6
rfueUZ4KDQ+2rH/9/9VSACFPhatTUJTUMSkE7p28f4abhxPJP+Racsr+CA2a/8P41QQyass6+B7H
6wm9piZf/S7iC62EaC0dqD+QgfLvvyzGLw+I8SsUSFekuJUWpeyASImXE60eDZAuYCYttSx2sA+t
hkLy1keyY+sbexRCApUmCRNDlq2PG15O46Iyknacr49XWLTZwseHDfkHYx/Adlmg2h0lJhmqg9JO
Ht6YLMM4dSpqUJxoGd42IJoTjnyJ7t6N9Sc2UYP3cb0hVkhPcSvBxCeQjZmeuXSzwp1Q9nEsJL7N
7YSwaPW+K/eyytzLDtBKoOF802xiYI966Kx5M1r6u7l9xeVZFpnDokn1N8qYAglbICXUuFJnhuy4
bQTK76Aqzs5UCAQoTO8p0ok0X9y/TbnjVgYC4ezDddmhXdaw8usyYm/8QMT2t5aNvhpLRbZHvihE
0PtMTShORxKGcFB0jjN+kLqz7erI7urTTIaZSbTRh5quT8lF8CTFtEi2RrPnEnuX0DAzzikR2cqN
RA5rLDIkY9jzBAYhh2g6D0jXbcNw6QVvcPW3TNDbPBEpalDSuAQwQd/fI6mvUUAXVqNpMhUb2q6S
p5SZJ//eNpi0a3e+solAQbokKekzfmYCfPGs641OdposLmY427WFsrfni0YZ2Q9JjRGriuP5742f
AZvbQniK/lqcXGkkNDGTcxY97iGt8gufteruVBrRNId60TzOzTdE2lDp0B29GwzsNYl2tvtlL6Lh
FuG1cqsMaBd4LDDktwUWHopZZgNPSzGpFUQVSrWsRTunbxFaWKx6DcG32CbBvy1AqJdosV4Fya7Q
V+oFgwdfqsmp+gFnAwkZ1fadmLcRqrrQ6W1FTZvnGdEz6xkb6HtZdp7uGYzZ5JmUJ96cV0Fi6Xp+
E6E2BRNP03m32qCX+UYLanvAfGq49E1ZLC4zLJewWKHRWoW5O214lecP4bCSo5vRbolBnLCR7mBs
0bGpc5A4IQ/e2t2HfxJ9AGDvR9zl7bbfa6Zp30cNdiPmO2EPCx8FzdJbPlVOEIF82oaYEAoWWG62
fbAz9aeWDRgt2iKN+1J4vR6VI/oxStmvXXfsB/n3hEAty5/r/gigHCXsPOEEJChPK6PtYqdTxQXJ
cQCMe4z684GyLOSWjih/HKV03W7LjL1Qx/ukMaLz0x+hK3/hQ7HaqWtes6HDu2KzzGd4qqKPcUTQ
w3DWNlrNVj+mQhNOIZGY49CT24Tg4Kiknnmyyl97zELFoGlGxT6zOQOnbt8XwaDgIV6DuzYLs1ff
AS0NVD48ayRWBOsjg39gAwfHOrNTQ112Z/3ihFmN84Y3GpDouGkGsIXJoxf6ljbcwlYK/ae65yfO
+vrUHNWxoyHfZtX38pY9vLDNVFkZxNx8h+LNc59bJq3yjypJEUxsQRzfV7s1NR5Pw8rTORoMsClK
xv1NeIJ5uTAVSq70EUBHGu7Z7GUrb+rqnBvHutkl4VTOijMoR4tG5Y1S6qlD1WgMLUuB4mwaDZ2/
GXcA9BIUvXwly06HXg9Cx66EV686o3JYMZaHWMJxDN/jCaMXCmuih87gNYZPLxgWhYhNP24vlXL4
7AQjDiVBVH1ooJhlRPDwM541WGBKNdMoxgVIMz3BZPj/gjGS/Cni6XlumHENEL3+ZWyV/UNJRrtV
75NYrx9/+IoLom3PGfrDhq6eKDld4rCNkuLNeQJZAqnE2BLRjyCLbPdNSFXqN/Hqklapp1or/Bl1
X3HDEUT1jlnldDUkUcdPNyYI4UDU3yMtkKbEvlswBu+Ns71ncRZQgnDlAkH9Dbn2DeEScWUjWuxA
TEchqqYF2u/3gaflPTrPjUz2+vrW5jmozK9FkXhV8m/f3haHC9bY29S4SOJIQnLZneyihjI69hZe
jIuiIb2lZUpaivvAzN/etBN5t2nvl/9ST8mPLzmNOQ/ImAiN5Jg5O3wamSwsFP+L9saf7qsiuamr
iXyNhQUvqyGjWHiMN/kofU/YF5DDb7Qo5pLg44dXp9vejA54olhG/ntas4cxf5QO39vM0KJRxKw/
eKoeG1MO1BiGkAx36v399So+gy9FZdx0PXhB17/PNfYU1Rm9pjIIfXgIa2Vh1HYF/qw8tDAqjad+
zxYlgMt1L+7YRW2Ry5MWeIDiVrVvEAkHt9VQGFpNxdxsAkLfAepgBFFZ2RsMJzPW/aPYLgy1ly6Y
DvL4WJ+w537iyXRmzu94056MDoe5QgtH9e3LWHqtT1f26rMAX9XeOXc4xxopYhdCNSa4KzarCu3S
YLGcpdnNPYYrcZCD/eceRpQ6SJw+jTyDRKY5dupfvv2EbL6B4R7+Xx1Ly2Jy8kCWcmwi89oCmIgr
yR9mKekrgS7H7P5pHV6cWN1PWpnNJahrgikPrtLkFSEcg8zaq8jqWt1+udYbDN8TEHfqdeZRd1AU
H7STlxRxG8iaYLpANC9+OWR0UU0mECZIB3jAgiT1zvEk9aygVCW4Kbyuw8N3Sjw/3ZLc0mN4ywo7
lmuD3IEuiUJ/62FlySLzHaL2ubm1WhbPN63yn6jihutdIg5CTKxRCfPBaSlg3pzTeJaoVxY7C6Ke
Qb9HaFQ2QRMvf5n+sbVf3yzDt1PL0pXbJNv5Y4MMy4XTRmRChy1hbeSBl3G+K3LedSUzGsQWm0uC
/HtNZzamq72MEhprLyG3QnShH6ddb7DU5VYaYoaIGPc8Oi194VbxP0O71Itq9e+u4vguPSfuebW9
9h+Ma71Ba09cOGpoxxxYXmQVxq4XoLiN36KHYgHLlh7DgKblX1VOLa4USmGNMV3m3ef1Rff7nXKf
ZDgTX66DoWfYQCKGy41srLeU8rygf1g+xjnUWP0heZD1Zgqxq6+Pf1yFhqVCoVixZbLQ4V0VfI0y
4s0V3bbzrvqTVG/JFrbkO0FANiQcij1bVZmlVm+IoUbiE7d+BEpXdyto4Egew6UYOEdBH8Fx4wuy
RF04XnzIOJeFoEezqjjn+xaENaZ5PMKgv68rTE3MACIaZIF7ensYV/ivnSNqTJVmopux20Y1uy9I
8BUwLGI/Ne3yWNsWE7NY2uCy9SFXoVV4KSsO8Jk/yb8wJPvDssO99KGwEGNPueSAorOLE2lhZFqe
2TLVk2hekPpd1b9wwqLnLKLe8flw3A6v5FmGWfiEWQ93qNiIG9PAt3xQPqlQHn+3W+j58EU+RBqq
5IEg6weWyOvO8PExRo8YtJ0DbADEzkhigxCYMi2JuITuxyX/oz3VY/iMMXxuHuyn1ZIfjkEGQ41W
h/RYvbbVbn06+6/AmLuhTbJ/Ts0+XHMK4Q5MpHQlysVAToT0O6VlcarGii2ua0EjYELsJ7us0uot
djDLA5xqJnaZ/sLqTEQTPwWZXaZ9VHFn6GmLZXolmLD9YQOES+vzxkCtA6ng4hpKDmFq6XsRo1GU
0hw9d9lNttYkGpfde7nafYRKLal+hnKQgkfmMQForHvxEJVcpDKccpax6kQyrq6lnfI1sxjjbplC
ocDf551DhnYRfM1NiShG+dNUB1DJdEKZMoY7ar6STBe/LvRiTAgC94jtBTLES2SXGXYCzCtq3BWx
hYYU+W/7HJvhHn/jzrPhDMfsphx3BhN6FAvd6AFO5wjmlrrRaJ4YrxDGd3bXbe8dVxBKL3pCiMpp
GAKnKrN9CP6gHmYJDjLnBbWD8ZtIkLs7tSJxYSQe92FGKHmoPnL7hQqrZ+43X5RBs7PVamjxQoJg
wS/2Mvil5yiHuHl17DIqPYMxQh9m52vijqg1IVUeGemTf8U2O53s6G8zBV5Rh48AUnDdlSfliIxl
vt9KXYLy5cxnZc9MnRC+px/NCRyww7TzZ8lT4NCGckl2fS7anOvJscHk7dALueKDUiAlwDTjMOVi
01ON1v5DvPH1x9Hg6KrUaBtMJeRRavPIaDwYXmVr2bpeuXDjU3MvLZMtomFItBaL7itr16jebSPn
5WrbSALyQKIRCoMa51J/eRL569Nr1VKr7BDcaOkKd2py6Y7zVZ4DGUHFvmGVYPauo5KU9cjOfQ0T
9Ei32VMg/B11eyNGFY1ECE2bRkUIM+4pKCzee/WD/Fjh0DK2mg8AkGrCf8J+BSq/PbWkaWr6LlnX
4LQC6lISz43e03r/0rVixKxEc1rQfEitW+hqnyoZ2qsHTOpefpfDvt3W+XMvhdlFZAVMe30bEd3d
jVA+8MvP7iMx+ACfTKjkI/mc22DLikfnWkYwB1CydY5ha9N6/qFd+7mDXzZGP33bPI4tF+7u8DwY
Ot0OLkdd9qLlJtb2+tBd6QKaH6CMoStH/gnTxOd1+KqrvQHerXOVvHVCNI2cAXsTTAQth0N/n/yi
vCQDq6jxCFdaf8lU6fl2aBm35uXkYaLMigqNbAET0eiJXCtyFRiEXpfdIVPur3YoHzj7jACrBpTo
HEoGmoIqs95PbHQGAJYGr58DPFU6mi+kwrAaHyQ471TULLNGADMcgHfI+0f6ure7zbcbi+spgXmj
abw8Qn++fqtie/LRy4WEBDPdMwoEfsqT3TpZ9FdmFkN1N9F6D3szfNUZWF1nhFS0+b8iWX8m8sGJ
DEVpuBqpz5Ek90gnvxg3ozMaj+TgelKGgYvTztXHRkrMfwa+5ogbzYqXcKC4sfvtf+z7B0jBMuXs
815rCR+MJCZK2tL+N5mtODXJw6M1/I/MsoFGmqmieQUYsMNEKokEsrgsAM38Qfls7MwTP3ztgqKL
g+0AM0IfAK1IgmSvmqY7XTE+d0vlKC3dbxXaHe/wGJcTmEkkPKWl+5L9l4t+SWHx3aSMSsR7Z76B
obHt+KYqKv7lnKU6kLGDqLA/mwzCfBqQquL8Un2vWFyrGJg3V4zWD0aM+aymAMQZr+oK+4jkTYxj
U/PYiX/VEkYWihGXI1gHGSxuBsPmo/bo1tlHGV2T+jY/+Abckmn/ctBQaxf+sJThkK4nLUHE47v/
apOb8ebbbBRI5LsXWlermXbu0urm2RarsvTvMBRJNSPaU+YksIlDu4WL1RvnHi2bDbbDcsCdYBnh
3Vm1kLR7UHNrwPg/Momv5zrWGxEVUkVCK9xIEyd+PjrshVn5THCvj1ebZudRSRUMxF10bbe4f2nO
LWnXypti1TFcvAu1Eg91TyQANjwo2Qcxju1Oj2whW5VA17Lzd+wn7DrBp3gdxslUARWXDmRCu84H
2N5F/h3nU/YytjWmHNhv7aFcaIpCtXA8LEhzeKbvdNy2OydsKXM6UhPXw6rGHfxrPfx0OwANlGma
1l7o0dpBPu7iYhpfrqs8MhRQjASmvayTVCwfc75e6EwvkzhgCvAOY2Xchu9DRFAyihDvQgZvkvm0
vEn14VFQjB7ebx3hybGQxlTSTKhZR4+KSGxE0Qzh5blVHUj5VtKM+GJYmhN1LLj/akPrkcYVlmwM
CQJpd1W14++fh7hWKqc5wCcjCgiSqhEIBOPDvvi2cSYutVB1yIqXomUkZ2cIQQDHAycvAxgzEs6w
Ur/7EwSKDyESbIii1QiabZUmpJ6Utu4luDj7VHElFjpQ55i0C/UK8hh/N6kWL1XskNQsb3401fgQ
HWVtbZdUFILmcGi0qXzSsExZYkQMHzlHTxGkdmipWQzKLE9Wit6GH69H1VP5NmV5sw68sJVVFZBr
9eTh970OopKV5u7dUsOktJqKnHlGTRLaXA/7kdUqhwvz4FO1a1Xs6SUuOMY5E2+qch7IgACJ22V1
RBVD8qVxybSwzmgGFlP4FyDebe2aWZaq0zBi9o4l0bxlqPmZycRa5PSaK6MljAU3nXa6BdSx+9sJ
k28kJBmP7i8Q2TvESTMhY/3DOapLGkzQboSCyOYOdhQU2rFuhFC+X87IJvd1iECwfOP9WjDR0KYU
b1Ahxo+kNdf43fBPtTyNlaG2V8RUNgJ/gbhvt3LfW+iBCi6CcVcKalD6nvgn4XoNyiwNuGSC6G/q
TqJtBxzFy/lVQOQybLWuioEz/Eq8mYNNZlRqetz7IFoWXt3fDDffkf96WFRT99Em3H0ZKlgjTA2j
dIGeNQoaiPcphlgQnKZqZlswsvUt/atzRYcNyBLhqB+zI+qeathOfpG1bMpWziyqLpLBVHiALtHI
XO8Lts7esV3qCO7f0liUCmyGGORyWa6WXQgv9N7OnuHOLqAmkTkwMYheUD4d/k6r9xtz74BsoIUi
t0OBBqEMLjpvKKe/NGDGsWRzEtHx2qLgrL8ZM7D501GrrpiTuEdHUUSVHCZUNK/3FdfGdRTnC8yw
lpEAlXu6TJUDbmTSAFCDchdsUP5u9C7Hlzg7uFnFMVG+pefbiBliSLM64P4/DiuMKLQMyP+zwI0Q
RP8TADTx1OVYzbCif6FQpAucGkBecv2xpVSXciWRA4s6MdTjjpza9RJqE4s+aSlLKOOegob/5Nes
WN9jWmZdpIH5hyXYSWJkTnOf4vAc+qGqTTC4X0Jcjjxolh2Gz/+tHG0RxUfMO0G2VV72qmY5nsvF
Doq7vxWFrQNwTJHhlkIOn+WysWguFd3TGfutoUlkVxy5/P9j0YTw8A227Uk3limV7AX4y86srfUJ
4kjOqnAyuBsd6RN2H0aRHlmCfiIeKM0YwBOsT6+l//V8FzuX1Ug9TVnSWrkiZb6TLTvld7KE+nJ0
d7vmpbVJ/kkhNd1xMTeUQ3eloCDnyEI/8H0hxCsyOWonvf2vUHJGFOFSMsYyZbYto0HPMXFsj2EX
cvTpEn7Vi4Viqh+cntHgPG1iXVqAn+ZeDnYXsoKZpBLBae7zgnZwdzswh5I/yKdUit9KaJvwBoOC
BpiCZV6eztH5vk3fsRPk7djE6PelNnmHwErHSP9OEAZNzaKEJRo6WkQJ+qY98J/CNShNSy+SG5NG
1Ywo7wISEadeXLiOd/JKIQjoyJNURSjbyiTfhjomTpZQkgElppQ9klQPnG9JYsIO1p17TJ+SXFWf
WqFWp4pXfDo4hl+2AaDoObRYb+L6oWvclQqOzNOs7/XFpa3b4Wi1Tftlp4DZyHi7xCMYGiFmzWJ1
71UJl35DoWpjM6CjvFteoLNChQrPA0tgGufCb+fMDYFMTwsOGsVOUF7g6IN+r0N077SCju9hypxt
noBTNgdbl+bMbWKxFxyvWASGRfF6u/4fMjVuOQMNEjVmyYEcVpz3ujoH/rTvxYdGafG1Z1amSwBG
mn43zwt7EFd+dnZD47Y2yCbIczCODSkWkQe+VNsXc4dX1fPqaAVVwlgPxvukwH3p0KB6prVxhl2g
FsNl+hRxE2qmgqUEV7lXm9nZcVU6jvcqnKj7hMz3QyOyob9Geq//dQ26sAy3recRtYrEtdNG3ti0
BYFOtsmikNbcBqGug8SxXFMl0eDTovwO72266JqAESVnaGE61v5zk1tSZs9efzOTflnLExlg/Kfd
Ks6Qi/KQtURIpz6wcFCWs02g13CfjLknok+aqOTcllxWZKeTzK5m/Aw5c/A6LOd3bLt6VQMHeQPd
Yle0D7Ls0fn9o9xglnGjc59aOqqVUdlyV49D6xrcABU8gQaRBiAneVUu6hiETzjJiHf6XXf3qhLq
mSqbg0jkay7M0fM3WNXIulj1c+6KbPvpC7e5qv2UtOJ895tQWm/ybh0uVTs2ylHj2p3gx/HVnecK
jbnsSJuMN4N+jVEyfe1YEOOoH401Ya4Lr/w5OjJnH+NFaNTNfuUSkSLwM6e7XWEoibBYtx3mRQ7Y
xAjFZM2xXv+wPnMi96BPUp4YP8f6vQY30Wjuwq76x/AjXvlQBOIHOHtFh69gKmq0e8JWMk59ba1V
qZ7IP1fuR9O2opuljoB+hW3XQOZ05hQvfz/WMTS3SfuLuBHmRHA0YpvNmf75/Fu75pMnfdU+Hy9y
aLFQU2rzcv6Ff9ewp5MKLolP5UihopGe8h3wuNRzxR/tHx+Bfeqrd5W9rQZ6S8cBgqvSUBHkYSZd
oge4JNCBMhWOCqyQlwIJS+mmIjgGPtA9AyM8ICxRXmfZrsMl5TO+JfpBRI/agH1ogRFO9fTZsl3x
xld7ujzIS1mU9gAScY6M7wz01A5JGxcPdnzuJMUJ/3frDNX+hu1CNH9RfEW006bNlwuWXg5iWLTq
vxIS2sPIMZgKcuOU97I9DkekHNZr0HwCex8L34cQAJEyxsux2VxHm+ULl/vU9hpK7PQ/w+owPpja
VdxtXvc6j42ZjwAaLLOnby6js+zTtgjtATlRs3PPWgnwh7f6HuYilPwXMMFM4VWAHTEeAb7UQD+k
mGx0ZkLSNKNE9X3WShe2gZZ27iBqLkeZZRXBk9UWEeb/+XSSwkrq1u/XavLDV101OX/LAKOxXkZw
IBeq8/FlgpBZofvKgouvSh9F9M6t7g+v14qMDcNDIowoAsHvlCKweRRK8r542WPQGyMTrMWzre1Y
wTlmGZD0SfokEj+5oho6VjlDKGPm9ZP02B0pKWIInlBKWY+MVcd/6QjFDmiaXErppmBNpYCXNgGO
ztJSNqJkR4vAYSb0AWp1ciRU7BfaeU4h+ckn413lvduJBpWDoSsb/bwADaT6MYd39KPXcoBxa9lU
GeccGatXeQXOI9uWV3y+eHF1i+eQpvi6XvpE+Z2zNgBb+Lvy9ntJhxZYONCuLwd7dXnRJpo/aJPp
2THuWD9wfCfvKOFkZ7pi/Fz9Uu7KflqTZ+DUJUgsv0g3M+vHeTEqKCXNlZZ9cIb/3C1fiWA+N3Og
3VwbfpyjZtcAm2viFMigHem6/+/kCN9C3kHMV4+NnqPWkzrgWoeKMyV14Q3enPefN12T6n4iFUgY
nJ/Sh1PSsIyda4/vES0YFwF9EwW5ZzBlFHtgfUeoWErKA4xYkfbfgQca7Krhkk2oRy1blRq64iCw
QO9Saqk/llMcpx5hNs4LpH1GuKf2EF27c6SDdrRBdBMxQf/R/qpp5QUDa3bHfadPQm3HK84olHdg
Kk87U4jUqBNb8wRD9mHma1b2SPhbzk9aZZDmGyXl3TLlcGqosiXDFXIdO0m6+msNB8gKKIhL6Vv9
JIuMd+o+iwMLqaNgIBRJ0nNtJWV6M8KtQXKHthWBzUOnELHSLOgzZghTkWolQ8d/AGQRON4OGv9M
3IQK2i208Or2+Gp5zfkNx65mZILucWfBfChzYH+ifFusyIlengUKCCaF19ZJAm3E35oAvmgbRKSM
oQHEDVBNxjl4UAsQAKcECjYbria45rC4zRcmtiiBBLBhOnin9nlAyY2Ol7qEttAs9CzINjBBKNX7
PYMXYhEb/0tjuJvqji05h+ioTlltvfz1QklAlNTqNH1OqY3yDxzU8+DXAgO4Us70hSdQuqB0bcj9
Cw2T4x8MstvNkc3ccr2aboqTS58Qgma52mcikzndjhjgjCk1NulJZPrUl6j5pjhgMxZlfS4iNRA2
RaWivJTip7etjcRToDt4doaKGb2LoMYLfngs2CC5HLLU0EQUfAwc4LfTZsPJpbGIPaPc3NAvXlBv
VZ6remBpF9eI8TFYh80s93M3X+vbutovHvGldiLK9EHYJDTe48qkcXy+TcES/QjrUrTlp/3xmvjd
C8e2nREmypayRHTBNr1gWCIBtEbNWv188CVrtgWCptiYLBMdBioqAC33qJyiEHYbLx5OErM+CkWH
Ef6/QuHzQwJDR5Oli/V5NLpDMT69/g9ojJtMIkfQVrYJZxMiXzkwlpEJk4HNv1PnTMbwMnV6AdGN
EkOx2wc2/Xv4IFT7lIFo5MfnoHP6vo1r3IyaXw82Xzg2aUG2Sjv7ONyuePxHErCyLmTNgb6XSPat
tgZRPyUHoKKMaMKLzUWAb9eO/a/hYlf1FQCLpAnYEYy6m5qW0IVviP22MVSqEgWWq6fE1Ash8Q+H
yg66ubRakDOwJK886Un/0yyKFzT6HwVHzF1nP+Az5QT3zMoDeYpQAYiassEFB3e+El6ORwenaapW
cR+k7SUmGlKkm9UTBjkLGtdof61e1+5JEoKmhXV1W2gIshMCMmB/MVveHGJOrCErcYtTO0bYVj1Q
a7ATTDLMyNjvXsPQ3Na0rBMf2W1x0SUvGkuZP8U+mPoGMnYH/iyKMWwBMend3L+59DSCIlG/3aY8
GjJY4mWETpDbs9z5olWvoY5m2JXVkA7pz2CZ1k4b/sQ+Mve5hYgpNrHCiFUVZf/bNq+np7UYMRpJ
ZewmsDa/J1yfz/8wBzYeXNxzqw38qn+5kZHaloKYKKoNCznVSmugtTnjv+3yRIBvFyXURJG4Nnx/
W8A/RKxMLxEj80cujge1yS+WfCH13M4FV+6umbSQ5XnJjbbWy6DmkvnisoAibZahjT6Dg22XMdG3
/fUjDU5ALH8EpCDAerEo3/0HERzR5N8qwHykRMMdVEMP/RLR6hT9wOtvFiNNS6eN43+ld2sP0na+
56Fk5qdaTnwxO9IlhOPlS9g+5OE0qLLPoVlb8YRVtPlbXtwqQO2cyESN5fzOXQgshS4hqa8kEybq
HMc3M3N6DRY1CAt6gvPU54VOD52x4mAi4ffwSWeH9r9x83qSepNnQLsdXVNhageDN6lXBZLsaXqY
de5JErajE6DC672mimDkUDF3yuLCH8y+ZCw5qFdCCcabMJLicW+zm1QhHCDbsmZYuca2RCeNZiY4
boST+jg/2ZjPLle1/v2+uvTNBZENePvHX2OJwP4wDIH5YEjkj6FjZugFam9JQKAIuffo5+MWx6a4
Y4b4QabWrS75IVQRShY0KvqVzgSqKsTzqIBeiBYaTZuIRfgqxQxl/0p3hGMKDG0kKwvNK9Z2p4rs
QFoDaTXQhEg5HnxzXqUxKO3kXmaI4eBtZIv4d6A/byNK/NNUGYn8kxKXFsDrWotC3MHxuHcdjhMt
FOLEk+oAUa+UAyEUnIvphL51iGWIlWWqDk3++LKY7cXie3MWqbmYknjMpDrncm/30cJclmNW6oeI
o/vNa5R4o5GtQJhHqx7gCQ7kWgd/ds4JHiFxC4MB0NN9HpsXzBpuzP9o97aEkJdUlNLg8geDHY+b
P83z7kJVbeK0btPwQTsSy2xoVHkoF8WzO/pMKjvptQmFXtRO9ZXp05bJ2DDUGKCCHwbdOgDMlV21
RnDl1d9i9cqWbXPf1otG3KsY9VL+ao1g/PPnlCWAjfbE3SS39Rebb6C4c6eJlA+PAgQkPfrQ11Sw
R/EV1KiqjPh/f0Tw/RstqJzLLE86Fh/h42BZjjfkPcJnEZ6YTNToDnTkIwhnpV3vQZXlGEEwCp98
mmr4yaLkgHp+XZ0wraNIVNEoY/iJ9CEU/zOyc8hwb9yRuqE/o8G4oqomZh+8+yjLY4hYGFszvtMh
YJhK+QELU61MNc3JBoQDp47SzZ/2/P/0OK8HA1IVjPTwERzl74VkqJIgb5bpDJILNBvPT8Oghy+k
dOvOmFfCARaASJyR276mih+V6BO1BkT6zLbv4K7zPeDjoD+O4ujLAjOrtMuBnTfN5DEl6OSz73AU
0/CNN6Q6IJHAujUDEP7Wg4ubZXaa/WQAOUnONCfCbjCdMWAIf+OTnB3/Rycz/xzliLp+aRrgMnLd
ObSnn/YpaIq5V6V1XEyewp4SonPMd41VqZv8seffKQsRymrT/zxTrTrh7y/8AiNcYVDB+V6HRuES
pttPaKEdYU9KkAMHwCXb66I9o2wHHvTEoLY2JUJXLgXZfhH9QJuH2cpPW04I7VnJzBE8aGnccN5U
m3klOL0eDe6ZANOSwDh94VxVH3CE6+fpPq6RXi/EXw0GcMRCxuFvQIFiwe3FlsU+1T6S7zO5VDlw
7vo5BtereuaIzNzLQ+RhPIMnr1OZkdx5uXFqvZmvgZD9Ofu/eGFxLNJ9qmHGPpBcQRmY+HN6/iCl
7LvHUpLItGBK1820trWMX+0aMi7JMMEybe/LK5DvX2gpQU9Q7pDSyhAThZpl6aG5W/7wvnNnWFFb
471ryV27qeBjNu+dwUrax/tNy+Z/Yj71Rq0ERM0NDTEp6o+adt3JBRA1+J6zAZ9So6273bIkn22L
yZVBWugcGVmn1YE6dodNiR4t9NHEnP5chxH6mZfts+IZBWib42vhDH5fe47+TBfX9opspuhoV+1s
jfJHl/68Oar6AcQyHHfQIo37B06MBYse4TFCeTBx0YflJeBU8nzPg7Q00Ky+CnpkBeearnJETgSK
Sp3eZgXG71tD8Qe47j9DzQrfEgCCrUBez7XKFAnE3ygHexIavH3aRwlH6FL09xYBTYjGvPbH26jV
I9b/LAdHXUUnnjWPTdH3vmzaWPNIZzCr76I0DJf6mJ7cWjSs3oHZ764ouL8+hNcdQ9f7gray/3v8
/cKokizhpkqUjKmL9sRGOm3bqRhxXjkfy8TEjUppF5JeNXRmo+AkeW2AV497vvkfLcgzBT4KbXpF
NR3msPBhq4yang1TQ1dVQ0N0TTXJCshnlId/Z/m57zX8KgByvQ6XUdCpDoUBQR4Rkl068JMFvqmx
rFh5f8a5rL491hSdP11rh6sUdQy+Pb7eW5XSJHWzhcl2lsDACsYUTwlfOLUO2alIr5+lzdikxbjY
CnhLIN+rECEXgyyj+tmIZeF7VV407pNA/eOKFg0wZ4PtUJ+oIIPn1oLHg/3DvWvJl37aqVnr6wxU
aephbLOi27pLky/8tJfPVhQeHGm0smsMZN/mXniLdawhvb6M/8T4jTUqeATq5xKZhx0vQA1Sc+J4
/+NoFbVpCcI0kX+w2N2yzh/7fBPgod9ntmk+H4u74kK6MRquFfvru9069dSqBDOV4RxBg4Lp3Hlr
CSS4tz+iMxhoynMni+h6IMcrlE07g+cp66NIuezHJhK6DJ2t9DXL/q0/8Ks5Iebf3vTB4HT//VNC
phn6ZW6N8QjuTcsEZ0qAw6yUScSo8qAtIlf51pJ7D71Q3yK23B/0tZipg/mdn8U/emMMk2MDnEWS
H93jlysNZjjXmFdDG2lAinQGPrpV/zPmKCKhUJhxdUF73Ff8zrM0tru52fm7RRh7yfEj60M1AEHH
s7+N7hLE9UvDMGVsLM/Ul3aEjEaqwOq5jev34OGw+mgUZhD56zWKfXgVCtXD0esiyBokFdH9O7hA
rlhO+awTnRMg+sgmwzHllcXe41XyK+R42Ac2nt9VKAwHGxwyCJT2l47oc+HpJNS46ica5n262gR5
4awo3/kFFjI9zY8YtQidoarbUI99MhSsviSg7Btf29qfnfYSCt5RsZsxhev3jhPQ4W89UXByAXFL
DBZooskGboMnwFiFaKN/FWgowEQZrp5C00Z7+Yfr90FmhpBiETdBG8wn7NzwdHdpue0iO4+U4Xpu
zof/J0WAQ+Nx48XnsIO3z1x6yE+3+CnI3Y49qbPEjdrR4CMjVjdCaJdU2EYwpDvovCzMrsm6Iv1N
qaHB5IX4NucYZVHZH80t7siWjsdYlpAeQ8/Rm1xYanpwDv8lqhZ8wfXdIOrnrOJh7tAhM8EGeuWa
3EH44odIzcXHSnSQnaEgQmt/4aU76FMFO9gJ9OU80lSYk6O3Kx9QQ/wmVftYOTevOFjhLoCujx/u
VU983NxdeZ9x8zn5GUOZcY6iSF8BdNHaT0xmjRDdnRAZV4fSsZ5kh+J/Y5MZvBcSi9pt9HvP5BhC
eNNheFiLRJ/t1YctvnoPZ0n7P2qN8+eJjjd9KvUT8mC6PXhm+02S3vjLK+Olf7EQFtYU5jGuXAgo
U9CnPxKIxei9tBCBhruw4Ii/5a9x1VhGlJBYM8b3nXmc7Ym8nwuGaRApqJfWNbWO8A/BBzijf79T
6gmick6S4yq9XsXUT5tYTiKhnQPP/dHiHZOScPC9QuMqI610TAURHcqNCJRqLTJG7h+2b4wdC/ws
mOC8O26Au5X7AR6CosHCr6qci1gpMz/H9zr/87z0lQ4A27ghYm0GdOSFQi0Tz85YGsmhUlZgGpcW
DCWf8gbbWVNo3221JZlW5tSWGhbHnkIK3TOBKfxe1qc4W+QpuC0t2wWaAinazj//EiHOR75RuZ3h
xUKdixq19DwpFajmH7O3+AswCyQremovdYNwax92o0/vmnGw/SNGNFeeczNAfX0Ua5gbDp06rhqz
VbwnaMgOivNF6OsUKTcMK3yeoIglPwNruPk95s7H5yasY68pgTBkD8IBXBr/xUceQBdaA8bwK/wI
IY1OwCWmQPmtIVBHI5KayHuXFi4JIhl0vXLI8y0OJ5CebpDRKVitffi83HCEwsMXJWrh1t5lGe1e
ZzHKSXXvs3+aGzz9lDEqDpW4Qt4H5P4HST6nl01C8u4Q7/1perfO/784mS9pjUPocFpq/hCSr1CV
TUaSw8PlQKv1hkYvJejlL7uhkxS+WHgL4/ZBqSx7RRYZtBImPgpUStweDPw+vf7x/nbFC0MSv3CX
Ep9XOfe6OgUKGsBrzhGJbLL1OasZwThsI5qGsAUmexzCjU3pJSLi302rZiU9yoOMBZoyoqjtk9wh
kHtj2+NOrwbGEviW+8dtYqQzaIHLODJ5qRYqz4hwiAYG0D3oPG0lRgz4/2B1q5S318UhbRBY0TOQ
T0BraNDPYWwAw9Br2P+2I6YunODVE5do2IToT9mqaYO1lzY1iCIg7PkzewCI0Tt8vE5diiThhwQ7
qNkqup9QkwL2/KjXybgTpWSSGvz3Br4aJUW3J2PzED/mDMq90kN7+2iZe1UIkESfTGbTaxgJi4Xe
Qj6mTU+6sDosmDw2MSMN9fh7EUCjoF2DQvSM3oe9HB0bw/FYgcleuR2M5rrFyFbQEl/C0Ki2AVHn
W3WZVGbIcK20aiaJLnWNEFzbzXZh4pmGRIlSwUEpfSBAA6vU/IbtVPzlPalVLVmMkpbsGFCHOQ85
inxRU072ciJg321FyJguBC7FO8uF+GzQj3SC12ZeMpW73PuPl1Z5bbZktWq4vpcvcWDfiAkTJZwG
Lcdn+RGdpCgeWwSv2atyjHlugJ7vbbGVWT4p2TENeK68dlO6ZoUI9GwIdvvQqhVM6fmT4PXfYqW3
mjWIlu3IPjnspPVCVdiCsIvrxzR7tmJ0KqXGsvUAFobuiZuLet/SN2+6qkrUNX9PveXm84G0CaB9
aA2u7uxzSXceyoy5tsJlleqgX5KN9Eq+UHx/aIs+fFrUrzobihRd9OmtxgnEr5KdTwhF2/2M5QXN
K1fwET1vg+7aosAOOMlfS1QNC5tiI9LOoSMGHMSP3DsiSHN9ZGWQ/rO1f8T54U5RVxa4nWnJcvbs
OnqM1cCxaDgq7S/JPE3hVhYLHiUL/XZ6XurFNyCN4vWZwVJw8H3Udk3GDMRvWhvSQtDvuWLyb09b
2TsFCljpRAGgdNoB8SkVPJzExuIIW7w9ZKVpWxhG/6uz7W15g06Y1ZIpU+v0Kef9WEeqIMYuSLK5
Qx/Y6Lysjm3GEWwIztblyY1IuYAE3n1sy8tGCFEdAy9tGJS9BRBNVyxJ/lJ6FKQtT8XINp1BkMYr
wKZJ0SC4Yd31vKs1+aTd/PRCZOeTbxPuOBTOdywp4c8l9s1/qXu4DmDr7Vmi6xpdnXD/ekT2HtgZ
mUTCs+9LxwCc+RYUR8skdVHlDsoq+frICfQ9Sv7RL3B2NDgM1uw2siWkpJ9G21qFeyJEi4Ea5g4S
TfKSAeo9P2By6Opc968G8F9M5v1fCqXT4Y1/cUu3FmEMKJtNFBXyPU+gV67mT59DtJAveuaBEKcY
E6IWL35jPdhwPWHmiO146n8PM1dYb2qZ/AeeZH+22z5zNvbVMsdOwLN+5cuWGyiPmIgvtnXy7xi3
eBdub2S1iLMH6O8mcFprgFfW5WZy78Av+TbBRq9VU7hJTpZ+8DkWKwI3IaqOUJv9af29HJrYWn+w
zZvAjs4vg5I0lY1mvVNqqVoV32ZERFdVyaadBkRLDB0OjHBAxDHhZlLWNcGKwpxISGU+RX4F7Z5J
S1djL+PvSCVrSOqAX+Hrd0V2mHhHg6IhdJK7iRxaS6aD0P1vytZCgNTBv+9NEnBZRPh+OBPwaQuk
18gil2fC8eGEHDKakWDarlMTeGcbhnW4bYn42mmH7bQM9IXxN8CloV9CmWBY9utsUSnuNcC+XJyC
1HDgXZImUEyGZR/PpPGbBj2J3R30szl3tiaBepsytoHM1sdYGEl9QcZiNaoTH6uUSCNOveqXOVDw
n8B/gxf97VHZTichEfYajqCtK9qrphB+DXgzPX6BlHrqLqieY12KCqzeiu73CrvuYLgu0umtr1yw
fR3/9uLsrFvdhnIsiHr6rj3OIoUqQrow7nIAe+pAHqdR5ZowxFCzGRtBy0My8OWmZfmNnN5n18Hr
OsHzEc/n8m7DGFjgfkoUoZ/fuH9Qt3c2SYeAQ36Y9T/gagbsTATHRwrQp41Pefqxh6gH4a0fr9az
3kYA/ilFfmKhAFCi6Uy5ThQ4aL+jaQ/7V6QtRM+a8Pw2w5aMddin1AzlqTopGWWTeNoeTymUY/xA
aR9RHnr+kebRP1LJove1v5M8m2KSDgE8tONGVbe3nBvYyqMxmmAGoGLGfHxq2ZPDKSnL65JXc3XB
OYgS0IjkFFyL9wvKHde9oFico/Tj4xIMfiZkghbYj0YyJB0FBRLn6Axt3o3BRgFwgejD5cb5in9s
mObnd42R8oC4a3smwdULJLoXxzvHLqWjsVqaBRseWp7wbTWkHAXSfUmM65C28vpWS6FeOUpd7pC8
PfUQ/RuO/VywuK+0TewtHsMBf96ab5nKsV3rXAvYyDy4Uv5eWylmZsOGsEYXD5V6MW90l+ozZ7tH
UfWXPxciRLXBWbzf7Wgi5m4yIb6S+xBKjKblBZlnZPEx5WMZoPr2OQkUkdhE5RUgtBk+mpaeL8et
FBvpoQAyXEoexlXsU0z1Zc4hd/YRMdS/3/ctzvZ3jIU5P4aU19xcnNft7XMxKWZqkZlO+8e/VHNP
DQKsStMTFocdz/hkc6ZHOZMnxHyML0MnF/AXcQUXY21K6RR2aMDq2eqHurQvuIJ7uKm/a38uVnXo
lcOT92DxYG5K+QT8DBSIdCNJHRUfS2uUB8OjPoxyLcre+GJk6xhHLYQlAidJDJ35RYauuLTLybkW
tJIsueqTV90qwRa6w8yuHK1agbCyoVsoj6HTYeqmSj9L/JAY0NLSnNLg08wszgras0gf8GrNCjNw
usvPbiXOJYUGME218AnhcZgjKcg14FVcPjlS52GNuY3elcaTAE5PJKY1Evt3OHxz3VNuRcijzsxZ
6I5r53hwFy/oldQVfIvDg6lHL91LUDbv55duZX94m+YYURB7aAxP3YPv/f0ejZiOH/NPI06g4Pyl
i3yp1Qbk6VFrT0VMNrMaAvrQs0Zt7z3d5xOrsv8EzWDbIfem6tIPfd6+kfr9VmNyuz5qcNJ/cGY6
WLhFglv5/Rg5m8XP8gl/O9Al+fJQmFD+voBJVnNBJ8D9CyPsn64YG8gEyVCTCnNTXCfpO3L29By/
p8kNlFXuwTQPoyObq2Rf15bTM/iymeycvbticK8g8LQ7jCyGJJUDvk0J84eBf0UNrp/8KfDOtqBx
PCaXSyQA2JKkkzagTIveV4M1JKIYu+futugf5GMCSuQxOUlLZUfFbj9C69SLDsKnp7YuYgpJoL0O
eRrHMu0zqlufkUf5BdfHdoYuw93580DLLio0efZJqBOicRe1GsMiP5h2P40K+Ji+ZiMRy8o5JVkL
RStJiztK1pQ1INqvDzipYVRr6CB8fklGB+eCaAvsUGnaGY45WSulMN4E2L9EdDzv/Az/xapKprcK
1gSEbWNlvEQXIh2UG955fjYt3FRM9ruSBLRTOAQ0J2U5wz3nwEAw6dUxTCq65xRuOUKfhsAvvPez
hq3wtyHWIXs8462pQbGULrgV+RFhmQQayqLc/KzJ14Umnj5ts1XYaCuRZcMYb6fsmD4EZa0vYGvO
eO59wd2faVcbAWcWJ+MV2dhx0wAOCuFedcCJ5cNGrLwGQ0glw2QVS7Wp7glBN6GU0IsPYLcBwqVU
8O/uQbAPxfEtS87YKTAF31Ie/+UL1NqhbcKQMwWUve+oGi//4oO0Bkpe5obpLH8R9m8UNBBjnKmA
j/tISn/zTMg4ovrPmPcmAFRtg+4WzANRgqlKjODAR07wbAfKxAREO4chiIi1s3JtePm1jS3OPzFE
bi3sZKQQCZsVTwkL6eCsqa0wKT3AEwQHaYe+bSQdwONc/WfDN4uhScRraXp6Zyze845OlUAX6ZuT
wcSvGyOlLKC3wEU5QXspaJ8i1AfC21xvF9LjWbpFzjrw+fgwzSEpYUa08GGjJYUccFY19oYP87tl
M2z/mbHBx3Mbcpr4x38ERRU14voBTWm8080+xgdas4PRn0SoZVOdxF+ptBjHFDw/+KXkfU5M5+NF
2abypkroMQYTNnJGdsHtoyEX2LVE1AE4nVEEu7Z6fQI4SlVgjNQ/T/4yx7K+xpntD/KlVG5fcuzQ
kQl16hniT710EFMXEuhNmKQsoxbmyJB4o5A4YSh8ImmODKgaXBnV5hQ3DK/qL9a1EcgeZbez2Sty
Abd2TfBCdw3epdFiF8aKBV8VhKCIE0yIZ+pLqrQlbZNxQoGkXasXDSxzFUmW1jsnPv8oUB4lFTlb
i2NlKgRLsO9IEAeIEoYa7eHq8SCzsocsQc3qCAwYSTeqdEPwcKpCgWB/IMmbyKWl9WCxJoLlSUoN
mmn/ZCW8bamdNcO1hMwAuvAqlodFGnpJLVRGgyWvumpeqKVt+T/ZR3nfiFCG3L7Qjwo3Naxajkw1
9XUAJxtWLOyJRtgnCGmOI1bXAVucEH7Zr8x5ogfBGIFC4xjKlkiG1KU3kN4tcg2vke+pKgUPEfqm
z3nOoR0uI3CN3FjsrN0XhUUD1EgEyoQ8fiRS5HTOE2ZSrJIhzz3NLkwmgc1GKufAhHVdYOsym4/g
SBbE340avpxBxuxU3YHpQpDUO2SRG2HkgjRub9qfsLaMnQrYbMPEN3E6fyy4qMyr10BWZpgK62nL
g52hHeSVp/y+f5desoeWZ38H29FzBJ8XafW5FGVGsEFr/idxrbom+CypqG3LyTIVzwi6NmLQzT7I
l3cDGGE19kbz084y/DNqHqX4vA0T4gLhA8xnn1gQA+XKbMt6yphC2wudVegEhk0fedn+z4XFPmU0
9mDzw7VcG50WHejV9TcdiJBtf9G51+SFLyUPaSfkUFSY16jqa1X1loryhLELwVqktMPSsX3e1Tj+
i6urB6B4iQvbEuqhvjhI8QPtgvd2fy+xbchmNMm5tlK+g8nXuK1gYv9dQX1wiYLhxRdb5CRBswSr
7jPVOsgA5uXoATyKnWWbmj92gUhBOwMjlvNleckY6o13PM3L4fn3oBpoNUMfLLS0ZKvrg3RsZByh
+Nqmj1/7Tk+x2VynqhPF/Qa6aJbR/ZzeyOllIwfb/ocmf8+UxCarfHE08u7CixOFFjE2P6w0eSrb
3IldeHh1zLRvhvCA8CYFxk7UAxw5MK0Rx6afkGFQJPsVOxuO/UFdFmXpCJ+bXfI7K/AHnu7TGYX7
oa+BdLM8XDlNiFn7/6PDt9iu+7wPVswlzOvJzTuhfN6s/wKEoaEM5360MI12Tw48uanMt6Q/01jb
fjC6zXrJaUoDosz2u4nlGGFRjMcOWqbzTilWKdEPkTE2h3ABZaYJUFj15pVkQKLh/BXGEZqqN7P/
JqO63LOysXZ+RPSSL363uN6iS66OUnC9ebl0cAMVgFTCQJYvydGIdOhxPIoU2jsvfbQJTXuDXk43
HbzE0HPc8DPMH3KZ8EjLr/MqdXzriJ9L0SzHKlqKWP9agcq2szVWr5yLIJ/d1BC1nAcLWI25/vf1
hc+7CEdOzT59pszW9zmrmeBtO4l+APSgh90mamqDvnB6mxBKxp2VJ+q1EEujnqVBxRyIeVKMqv+D
50i30oVKsrP3axCwf3IdIx3ZBAu6gwIBE4W1090Pvt3dl0XSdeXeBCmngDXj1FOKkSh0ENgBTJgO
YUdaK3qmD29bKessnuX84PSQ0fWWnEtuVLWL+hZQYSXxatjTZdw2nSuw9u++2LfksJSvukCU6aD3
aDUJ03bX8nQYZbovw+m5SZkhLsJtc+XgRqm7p+8RYG5WvrmO7GrvNqSD4TOFOIW6rmhhb0YYeHmw
iWMJT5W408hfBn+oqfmPgcUitoDuS+OXJUmNZQIORPt1URqbePrDXKLpsvZF3yYzNoFII6TSsQXj
CNoYYaXtdJxiG0lOSxYVOraH6H1v98BifmCA+SMu1R2Cppx8pc5Qyq/viTqE4StciQEcMgfA7aB1
TOYylHLcJBKNM3wAsstJxIe0cMC8wp1fqocEGJtnAl6qi+7qxFaGGpOzT81r4RehjwA65OlnRlhK
TYbRXHpFmV+4q5r7siprawA1jLS0EnjGnXh0fR1upYi2NcGkQQMxcDlQvZriFM0SK7dzRnveMziH
ShGU84qwFvXnxtjxiry4tkTKmKGD6YEMlqSpvuBHqKfgx1NmB+SvYT9fWqocGKx/yIN+Wwu4FPdp
I2DlX/ljODPwKIIGO+QdMFTxpxhPgmsK8i0a7ZnY996xFcyJc249wtTLMF/x29Bbs0QEP22lye+h
trwy5D7dFACren1CBFCJDkzzfbyFNA6t/x6aNkwR3ImXYhsXqJzfCRlN0NwQcgJGLuqLHEeidG1H
uLFeh4JbzWu3ch/xL7tpMyTI7oe4ZhSbjF/6Nii7gYRXaUIZ+EhydFk0R5U1LCKaeS5oMJr9UEOx
K1fg/7UKDypPLLFlONtuoTZJ/GywJhkUrdx4IixZsTwNKV+kx8axNZqNtWk1cEbRpbklbIPpqKSZ
d73p77bsP9wPQwNXAL+Mw5AR4njKoApNdIGJR076BOj4f7zo77VyOhU1PJfIRMatWeOWlKQofXMk
CVffm/zXJpo2B7FcYc4ygqKRMn+/+hFMND48FlUMMMASaJvHlO0Y2QYGesxhvuOEVPC9aYibP++r
6rNYDjbKmQlgWH+5+gFjzfN7gsKIUzPt9NF2eM/kMKe+YaCIJdBJfMTQ1YNUMiTYZNcl5Jb3natW
eZvuqHoK9rr4WF1i3dqThCSsoXuue2T7OniIB+avZV9PgDj49RmVVpnetjTqCdccyJjfLm0q9zNw
liz8+G3TFPAvFyVUc5obOdsyWUyoJeCPjNbf3pHFi2hKYKd0sqae3gy5V7JgY7VXs6vuCQklEHTp
8JRDTLtJhMHpCXebJbqKlP+ID15VeKuhqdyMMSmt1UA0pvA2oaUCgspjiKN34Lc+d1su3AeI8bi3
WgNcGcIRJJrezuf8/Hi4dXonx+6Qgi9wnaHo7s2PNQHga+wu18sueIk6C6X/bD4fdyS+UF2o4rG7
kY5EzeJznFnzod/JT2wlEI3Rh3yECt0d26iv4l3xkuv7nlPNz1ZCrz5JjHF6QzgcJi7Ley2o88nN
Z+8YtFNsqNhtqRbJqnbrXTBITjBzayQSmbLgje0L5YWy7YbsrLD3fNv6C1K1NF3QmFDv6n6yeTwU
fKe3Caxs7lLz8C9EB8oqBTKG5ezi/+zXI2XADvosHiweCv29k3ASzCqQWSyQFlerEWVRHPQMlhxF
8Hu+EusW8rcL3Gh9yycoB9VjPSQyFpxrvfQ1hPhUH40nXXt2M23zktlzYdGdgHI5BsJ6DPXwGRY5
vpXyR1tUsGYZehzIcmQD0wedrS/q/TIyzn0c5k1LdsaGphg1ZK/z+v+4GJtaJtOkDllpQ/0G7ONf
fL9Vzj442ySrG91XDSVX5Rps0/D2FfCnHAmRIlsW0UsrC/zmr0fJY2kb1hoOqr70v/Sn002E7VFO
D//kHOCrjnBAdVSX5olzJPaVodusuO2nHguoAtz9x8jhT3Z6XrXecnOMmhMzcO9Cmz8oeD/b5lMJ
DxVs0p9JHcCVHhLJDSxQ7+OBPt5FsY0wXgJVazI44n0th7YmZCZWp4RPi7XJOyozwOMWjqpCfxYP
+7KmZLESkXPPh7SFisADBplGDfMf1aEusRawt8hZZh+DxFmSsm0V6u3RyWrtYxcCFKWHuyI66E9C
88fmRMYoO9ajSvWDhyUsYmCDsS83kj/fyA6LApkGGtsCrxCwSroqx7wKHwChrC8h6gy+adyEr2AC
GLUjwdcjQpfmSBCccH8j2xeIIh6LNXbcjZ7D/ewH/rCD9YJuRqhAJIt4eNWm3IE+7uopvqbKLmJl
w53StSjcxmifOu91jbcR0/j9oXXtpbczacJ5O8biRBWGcPMmOSUvH8xiX6llTXMyaaE34WJAnuyM
oNlP6EYInMGLt/vwYtrL6ZDQ6XwLO4Qn39gCfWXqtEFxblV9anPj5KriYZJpxb4OsEMZ+B25Uxr9
RKISflNzfoEEQYl7dhwkPEvFcEBOjULy9HVwBvxYZjXMShdYjlCQ+lkNw206QG+FbEckywcKCnjM
Ou3sA1DNzayI8Fmi7HzzB8hnxhw5HoBNUKEBSqxeP7UAZICB5TMKhsG9Z65HDnl0gGYB7l7vNa3O
g99pQL59biWWVA7h90MD1rnycnqKTz4N6z46n3+em3RM4s6dUj9R+CqWdy2OblsK/kRyEi8H6Jnl
JNVOHq7R0G8XBv0wMdqBWbVnIDcfshFFN8CPqRlUTBzFIgIvtQ2AwmvMtxMskEo7OkElRTHdiYcM
DasA/gEggEoMK1oAMv76bZjIBdVycHZEJEhJmQKXXNnmpXkMKv19HWrmHCpddmlzFO/1WMdCNyPm
6TZm70GTMZ0/gESsxipVpd/EcL7eWkl+gDZGskhoFtmVmHH7tJ5TGN2rnYTIXg8p1twK08tjhdaH
RxtznEvWRIb0q8bXiWTQusrb4lIaWL/wH/JqXcCpzKuLrsIdDTJzGoAeTYdDt4xUFbhWorf4EYiJ
KGgnutLYfm2xtS2rJ/7CC9M9cWgiHHyCTYV2TYuaHhgbYft/JiMrIvF/TyRNPhokSvnciE8Xr3yD
1GaTytkq+WmliaJ/eTQtvbaxBGmTqim6sYsHMhfua2DlWFHKZ8H77VA+2+1rIPKYSb4QdR7KjPho
U70NE/BIxwV6Ux/mjMA352EuR7JFvgggJMdE65vCzj+83kkzrO+oFLsVUpoahUodyhynPgUIQf/C
/WjaaY2xRloYJ89vpVkezpUN44iAZiU6KvA4hneesYYTI6I+sWVqcFap1IVu87W3oc2AbQHvIidU
Fa+nwHlabFxGRS18LqtPLM285C+SqXAGA4snWTpgEdPZitK8Ql7u+AZGsCiKEd6MoxpirojEXEPd
Dyhf8vIxroJ206hcEQpYW70VG1LWxYiPHK11fjpUH+siyMZaPdTli4G9me6lFMglS/1a/lbAYemB
BE7qGuB1ANI3VX4FLDYM3mm5sJlbzgLqsROFnEb8lURaWkIADHJJjipcAvi9rDHKwimIpMDnmTXT
+B54Gser5xbKQ7pbBRYc//BEHVP85YAUEI0NIhyewAwOcksX4+PHBW1btqkU9Sqi1Js5CRLyJjju
ZmGYMaY655YjYLiI6Wq6RGJsn7T7lXIQM6f9wpQzzhHYnsbeZZREUjt4FWa4xYKFPLFgpU3j/eFN
+juwB+8qCKh+XwmoDf1wQ0nsc7WMTNH/e+MndrFHuAhJ6CvYsSrpsAKe3AGd7A77+nekwETol+UJ
BuJtCiPoxgyTQXxQPRM5rwjQJNR9BpI9CS7TRZFL3aqK5K92kWFJNZ0jLwtOVJI6+cDxWYk3SL9Y
5dFxnCR9Qt5LsfkNcgl73trFnP4GdCns/bOIaSLJ2VMqJWoxuRQmk1nZ42eOR1acL7M0jpkFaQVi
2Vb1LdF/D2vr81M6vAnGCvbuODrFoGHe9HpLA9m2IETU0LH7ZlfQD4RvPK/BG/qQ1QyeAo6cP48K
WEcOYDSLRmv3DbjjjHW76D0GtWQGt53MOWoGH21vbiMC5tOi+OL3pBVlZjV6c+VRq150pdf1LQtn
5SR7hTd/hFqZgE17ZMWn7sPy16Bhril/AzB52vcSoqq4UQkXvqUsBJwdhcDkwxKmVzD8fG/Tt8mZ
6P6i0/TlTn84PlR+yxJIpz7Jme9RK5YaROY0xuChmrswk/x0WwyJiKGQdqQH9LjtJXOYg6G+1fcV
CTKzW4l1NdzfWrqGIvPQUaXNT+MZ3kdNxvqYmA13E0gmGgMkwZzyTIqF/63Ghd0vvNKp3PKwSPoG
op29DHRR+vA1kwa+8s7JUn/8HXhCcirz8ene9VyO6ZquIF/lzA1GEMUg6vNiem9On/5PZ4AThyRy
ZHGVKJBkQ3kFYCiM1x8LL5NqVqFGaBjyGZbB+kCU4dxSDizcmBV7qbKtlBCyFfvLhBuaW4qGbAgf
TepziTsEQyezMhAv1wawfBRorE36+hC3ntw+Dmq+aCxXFmw26DxJGHrQVlTUeI7KfsMwN+ZmzFF4
28wXxsYjzX7aYN3hHnLq6RvqWVTRET7W7j1ljScmXey0e90xpRn5AZctwBnHYH+dCcdvS2YymmHE
hNPLe/F/qOasI+YX7Dm/J4ZpZQqwFh4JL1A5kZ3LwukReiCat9+WFfQmUXfOI+SSnB44in6q2432
a6JRkmFhnmO/EbJMQbSK4hW/HffDy/2J9Emwm6dlLsy3PYKaBFDAeD9i+txtwz9AcThSFuW1VNBY
5Hm7BYUhbY/z3iSaNvEMAitS6SYfTfDxPI+gjypgdiRjcZEDBMzQEgp7HTxV68NFjh5r+QqjRER8
pZ6NkuB78wbU0SX2vQs0mm536/SQayExuk8yr5DAj9aszv+IlgRyOe7OA2W7/XPdbNAtplkrHV3y
NwQSQmuuPb3CAeqmmg/ItXptdcYwR1xywiezlnMFv5jy0tFYbZlFioUTLD1aBZn40hqi1xr/Wbr6
ff+U4dl2gISbQy07ztR/l3ldlpcxEZK9dOvu0c92WYn6rqWFRKTbvg/GB+GOfVlDaDFOe3KasbMq
HEtb+kqAgS4pELiGx1c6fQr99hVG/ua4rqEurZn8UFyPUwVLMdLRUiVlLYV0qpfx1SAINs+yvRpQ
wJi+mlzQkS4oCmJFLlb+UTAj7/omb2lvk5jrNw9aOymiNvV622trC2RM0jTBFNm7M50UVAz+t+rW
IpUcftYBdQ99T8KNAHM41LJdYn6jsBXURjoJEziqiJLUyZ8e8ylnnZxSLskqo+N8bEJXn8whx92D
WhlmqWDoy+g9607Xk2LXKZTWNgZIyD9bdGplqFogZ8GC6JhBS8EXX12Gq4UrVd6plpCi8Mn0TW+V
zqc/SHJsjeHj6muvF1aY961TyWCxm8aTPn9RtnDlCAPw+oCpSL2B8fcZobaJwREylrTmfo4obmzo
AwRFntpwnrv8hOTyIotjDjq/KULz9PhQWqCCWkkaS3ehujmzW2erv+pRMXJ7CQt3ZJfXA9it/YV1
jT8wmdo2PhiK9EQVYEYyNoD44Nl6QiUaOHzW95cpYDAu7zLbKOiONixvb1pQojUcqNX3ElcE8B1F
VDnIOUzYeHJEMkdBl/PWJwvW5O2GgQVZgQwyRPuYeXj8+dNdFzUXgxvFroOfJRiY16ehERBt74sa
ibKb90qEkQaOKDwA1wj6EErWiKMY3AaMONe5bhTr/wWiAY4g4NrFIhZIXcBNr6qlf6hu5JS0WKPm
CxVPr7skHfsDqzZqHE/igE5LEWsqBlpfB3mfmL0ZdWggfG6BsYNYc5Bchn/qOxm0pCNc0CFAZ4L1
ZPwrhLjQSVlz7uHOWYUL+BDxvSUni1cj94KdZffeJISF3jZHL+r8f8itTvljHADdfaRf/M5u3NE6
xrLWPwjmscdq+LpSrhoCAlQwN/cU9F16XyueNURKr7LpUycuhFdLRViOrEjTq42n8uDKYFG2cl4c
H7oIvJmdnn+bMF1tf9LzbhIoSywYTk3fHLuQCNgwhQjqKVVMcY+xST3eNWosxgkI1Q4D0rtqan/V
4eADeVwPD5puz2FCu4ncy51N4vfkNolu9eFT6PNMIiEMELRtU3JymM18ONumyOKgSCgzhYUwCdKH
FwKqtNPZDDioFW7QpfcBcraw23klAu+iFpZ6DQPgjwkjd9wHPgc9UWJyeteg48EKUqOzqedlCS9z
TCD7uTedYaxI9LaB9s/Fk+KFhuFP3QY5XYEViBOL1QXlBv1RGEeIGDQpCEpqi7j8ZKYAN826KvVT
QJ9YTg5RzzL/GiV3gpdt+zXGNuIVQTtPX22LZuP11QaQb37fd+j2iYge/HxgFK5EIa5maONbYjFy
J54ntyYSI0OH6qcH/Dr/kQUFrRB3RfEVAsueIcCeDjTYHDfo3UvczAIF8b2kp+cAxeI4uj/73wpT
DNi2NEWZvL8Tr7FogR0EneopJFXLp2yQzRoaIaj+eNgBjQ3xDMwwsqqKQkCT2E9JzrWM7K3YyDcB
1SS9TrDiqGZK6bf7MW4s7tvwBZ7TmUN91ZF9fWO4EaHUZaI1v2GuLZHNrQaQP9axghYq4A0f7f52
DE2cG9Imm1fALXQVD8CuFYDbVIMVrjVJpFQuuMsa+2Z1z1ZolIBLqWc0RyFGPYKbEKuYWIq7DX5s
2Xz62b28OxqjVs3BzMUBJEgFZWccsbJ2m94sWUOztDUc3B3mEYc4M1QCDuZkxnE/5/HiWufUwjFk
TWFCZM3fa4kGCS49ShW71KnVGFuyhX8xcYJYuFtLx87SA2f5+0a1LlIhwxP+qx/1djBPbgnThDt0
fVS19QASoZU414C99O3q/UCrQkSQKLx6LiwyQCK/4pzvKIMqH/PCSiYSZoqns7DuzhFsraioalwM
UtZUlCepOY36/QDtuE+LPR2svhLOZ8mSJ8gmdo5oNZFTl7gFrHdItiY9Fi7sAhYiMd51pjcf5QHi
C3G6QCsB0ERK15YU9/JczZG1VN8ELppggwhqjgU9xilkWYeF/fD2UUXbDCRV16B6Ke7zGi7734iG
fkT46trRisyx9f2CuK+iXLwwPZDvNQaBiH+1QA7YYGkDa1Q0ARWX5JzMDXGHlMgvyFdiR97+2G/w
41GxqCmYlDfVd1SOH1Bu0Y+PBy4sAqfplIhKj/OSagVJYIYR9WYDdx9+uXkLgJCUZTcgOMVWcheC
RaYRxihAIRiP04nD6G9lewFzyXZJD0d/FIjclQqpxl9yMVkRWHp1D3Jod5kGmo9RJuY+oCbiuWVY
IaDfmA5moqKLRIlEV8EqQ+HmSWq8Th7AJ/t+LFhaS3N2Ybpo5eP5nvXV/NSkCRjOcHn2dDFxDNTy
NtQ+P5+sgUnwM5L1nOk7olrhl1fAC1bbKDx2Dpr+GbCDeq/jeJUyvarcN0M4rnKCoGgGe3thx2WN
3pATqhQhsLFh3gYrph0ntE2WNsncEFtHM8tRqZHD/wEFWzTA6vkJOU8kcqUDbRBQP6/95369rtL4
YIuFflPY8LmyxWJXEoZk7Z3kujYSnTHZEHFzZBS79zMXiRMII5oF1DVZ54NmjDpp9AKL+F8duBCq
klR9YwxGDFne31O/b4/L9TC6iDMWPfXA24rCtRySdxRZFcmnG0T8GQc5v9lWhQwYOB9F0zbKNcYm
FGjLDO7xKOFoIUulPnqVWMwHtT3JvYI68JfZhVoNpL/XDnfjapbbFsx10NQG9Hf83sATafOGHhfg
anZ7/AAXShl+2YV/DpAHW7O1bkEWkXX5r/UaeqsYzpbvhJAcJZIy2tn7TpHr/fwjH3ZEkaGu+M2t
EK0kzHbayI/EoeoDwY3ofFTxLPsqN7kKdT/4eeECD0T0FizCw2VqKYqFaO7pnupw79euRXS2AvFH
T0GK0wcBUEbCXGq39RJajKlQgp3b+3VlaS3ube/m6W86YtldIennasOm4eQPth83MvvOzzO0fK11
pMoMksfZ492F9qmDx93sB6dBTPUsBkWEBIK19vqKNfy/a9kc7hnmcQd3AH6M7CcAvu3e+plNxZ4H
DiqIvk6r1/81Zc2Tc0Q6hFia1CgYwU768GMm8hx3zWR35yt/0PCI55RsnFsEX8hpfUr+DZzi0DW4
/ItITG2/+f8XKXtYpnpImiTvEAU6qbKJPMI0nu4dE8m9GZFIpR+xdDaKtSaBBppH9nE1gPQc4gV8
b1Ou6Rikv+tg/YZtKKVHUngRur3nA5E3hjr9brJITm4QyUp7xz5c/BVNg0lfrEG5TNA+uS8EzSGG
+69KJvTyywZ/lZw2AkmdMgtA8ALMklJ2Xp59uWjFW/vw2SYiZpI5JvYYBYB7mZNAO88BH51XgNvs
dqjqm1szfPAKlSk+gBcJgUkXGRtyBEzXWGknKla9xV7NQp9XVBLbn6MYrCPyWk/PWAeSCS5vSSty
FSk/UyRO0MIlbP74SF+7fEZX0DjB8CBq6as24nKJOcvk5e7LrQd4FQLr/hS5gVyWZrh/VB/1m96d
1eAi7eB9lIBXsIx+GpqnOHT5WmV1CznNXVhzlQfRQWNuddGRSBDR/gHRruPKdgxGBlFfGf30qjDO
tMWUCO0K/0aojY57J+hm+LcUqnGldQay+SBy++WOfTJUsmZiCE2BAXhIe3m77XgWv4zztNX99BvP
yWWnul4t+CUUEDQb/cWc4SnJ45BzWiPeGpsIoVUh9QCnzWYG8l0C0C8dADJHsTRlTRX6acZC7A2/
A0FiauHyc3arLbVxT7Z4ytSq4UXMo909mZimT2DkpJtwW3g+hKkmUoNOjtwzBiJCUoR4YBFenVJ2
UJDFD5wRgsLeFC1Zy70AdXuudd97Vj21VB7OiE48zjrMUk8OHYeS+cjNisk5jV15Sk1dCwDk40c1
tFYBCTuu61ejEdR97+Kv9SH+CdH5IAFlx2/G+Wb3IGFUeOk1NAVXG3aXQ87W29SQhuLUL0O19vvj
M7u2CLQszjGc4Kdx2l3RRVfkI7hHDtF2VsxpnkojqHIEX5BA7xGf9idRxRpQHIccdjs2TI+2IBVH
KXUZj6E7uac09sZzEih+stjyl61vi+HxL5VEmWKa5a0SCIHr8mZkPRM+NWqIqplMPGrA31OeuO27
qpXHFM9UzyMjz/95kKcbEVxC2H86ffPCtpavO4v0Zmge26LqFOE0hGRTZGdm43cOtE5w4pq8PWSj
6qCsTctLlrKVQuxT3AIRUKJ9qDHV7g6eif93HMrUC/BVzDrKuHVx0C3mJPub/6Y2FnjKky6kQJok
hH5Rrlpw4V8DtHETLtfIeaKYi2gunyv2cea8E3mCgVoeNek3yJLxpnwIKEU9Egs9YAN1Z91287hm
U3McNFttk7moqBAbOEipFwt0aYVF/SU7Noy3zAocmBvMCb3sqffkf4jVavBnWleBMc9Ntt2ASXbC
mucGVjZRtRh3WlmwwxElNWcJXjpSHu9z9XngrnxrYhKP0DvxylGOURfqnC2tGT1kSroAZJGPEIhy
ac+g0JeSJOFIdgTC4XqrvURQZrjChP+21aiPcvpDQ+2XZVJ7CyIe7BdSjtgKfA+neZUcN4dZbKbL
QVM94EgnFFcS3W8pgYPTgxQBa/a+scUrhgML3mCpRsUtUjHXkVdhPuNqeDDGwkSWy5mF+Oh+xj1P
pMbofAGlPgl19rtkouAYANsHJk9dKuzs58P/zmDdhdUTuA4nBZ1WXjIgYiH3hTlE/TkUXqrpFZgV
mRdaceAwI4zW6gG1GSMEzj1M1BmBYCdN6LZ33Jijyt6zxCTQgzl7l219vzbiPpF/4Tdv6yRZqQ3p
ehpzwQ1iiRfpP14D5PfEOIAK6aZc7FFVabblhg64QrzkNQ1CABxbib31MQ5ZoYcc11/Us7uJ9qD6
ptxD3ccsECNOlsodCWJslzRuVkfOVYOdnS5l0krBSvKi12RFg+iUWQEIJsG+eG5IHE8SYj+qW/fe
OGQp7cUuGh3aqyzFA6QlgYADhanANQkhtCfwsqJFnBS6c9VHsqzexoEkAsTqvjpinWNNEFJbaY9M
qNm2pvfVlpjmLBKukw8GE9tQP8oyNAjUqDjK23fK8yWA6V2o/Cl16IRNkJTkm5TtL7TUrvpMn6WV
arhuRo/NB75QUYWuEH3sVNZSKT5utMyZBEAcwZK91eYRNjuU1/w0dOtlGzwbFTK1JkmgWtFZi99X
jTnykY7nNgFAHSttFQ5Z80IdmU6w0K6naoSqMhmAZ0/weQfCU2xviVdiRJpmQJQAqv8gwF2yZ8vP
5pCjoNzL5VhUc/jtCYzc1mUn0kRYrBdOxMy7C7YmTZ6gj7uL11cCSr6LmqTiqMplqMxlJgNl5Fhu
FdODcH4F3JZeaxfgJzQa76oQInxfMnq9y0yFHv/MCwEE295mV3jXLRZpIwZw1kAGyHkdStbWX7Wk
FXNSo5ZFj+IhQ8m/0T2Kqbu9Y5XGFBK4iBEl25aX2m6qbcp3Ke1sRv9Vujz9BrGIj5Qx8gDH4msg
PQjyR9RuoyFS3aqrnQKzScFGN518L1NMt6G1nvtgjMWi1Q7w1zQYV+wjxJHm5BcIc4OKYmLNg/5P
sH6eSIsnecM8RE8KAQNB5EX68nVXREkIGDvtaBP3sNCkg8Jbtq0lpTUzFwFK0XlxPqTq8KjiDKlj
AU1XPHAA34EfZU2gAM02l80esEQs3kMMrtWyjlgF7D71UdzbN6tf9f+JSIjJptIZqIdlv+/KEiQs
+V1j+wFBjlcebZDmz72a57OkZgqzzd88rw60H7t6zgAC8HRsMwykIcDaUwFTtD8IEWExNUvKSiks
4MdZvuITaKmkvZT4HXsaxP/C0EU+LBrG7e9iyjbilfJtJTR5Ige55FWTSD09EKmtMqxrRYCZDTO+
TZE8+uJhNtxEhvW9dYA8NtOU6B9g9QuPXRR7EAl3dOPnY9s/5Wq7fmO4pw9NtFl8ehF8nTAa8qKx
Gffd9icvXZc7lji7sHlmQyqoRk9uNqIK81Z2F8LIFuX9VI5NcJUBjO8Od89qZ46nthSvB17hQ/3T
HMWDu6K/o9j6Cc/VKqNe05fP47nzKjquiHKGNlUpR6lCAscovaoH+7Aam28k/6YHAnGnG7aF4CfT
l6ao4I1pqIfCTlUrP78Y/glMQonBy+eCPAvvKiu+bBWTbEm6mCS5Ok4iBxBwqLYQQiKjqtPobeGd
bbaOzx7F0Y/b1i5xhB1WE2GOdCXtpsATAKDtwxgL2T8vPoTOKg8jE1ivvkt2jTNlvIrxeaX32uHo
5XOdGzsNxdcwyrhTvJdu6fVqvExRC9B++jqHnTI184bL2gBL5aKucwcu8+J1Zm58fTg5Gfa+m17o
tjagQrUIBqJoIhhJLx6cqzXIa3ZPvIXiP5Qnevp9Xdq2Zmckg73ccUd4z6s40OpDCtWmihs8z30P
ZI1gd0Gl2YI+TYP0w74to/yaCOhBpNAFGC8VilCEzjSWbQka07QLwVnL8y/jImR9H5Hy7LngbMW8
ChFlY4AJkNEQuv6RzkAq0MYDgPSZtvj0hWVX2m5bVRk4cuukjikJhF+5gWAdeOoJ80lNxxuCdV3A
fFl+cA7PINMQFnA/yGMwhH+6Y//4Ff0GAik1ECGHyoyiXvBBhduArcKE7aIwm/b/ez+otGXo8cAH
5rUR4F5cKzI48hsCIlXet9euYsR27Ryctd0SsFeOLQCLUuF8hS5GRz/cCcUtndm0DVDJ5hR6bdZw
jkXmTbtoYQrTolnDrz1OFuAj0DMuXog6TnFUpEgUZTtAMzWSkzRxzHCXtGC3oTuaTNIa+KxFmup5
+W9C0i171Hlk8Mn39kuILx20Sb4Umw2N9rGsIXUvCOZxpOVG/etrrQdTeC88Qx/dVLb7pWqVAFUK
ovfUqi5wN4+20zOQs44KROoExWccKyxtO7nNLlcI8lG/yz/gWSlduNQQZ2QY2WHGHZmfLGZP5eCB
O1NMqLNGhKrEaTF3R7rvaTwDlVng5NuIXEN7tI9tE/1Z2PM6bDtcOATuG/Lm0mwYs7qGFw9zyqEo
OjfYDZj35aOODjfYlGvntTpHB30LRNO/qEJLRbfs/rOK2ndgMQMwLxvKxoLqYRI6M4KVX7Ypdm8i
JaHsWpAXnrIaRC7Aj4qwDJHyWL7Rt/1mCw0A0E2SmW7ad649VdU1hAYErAueakaixLnCC9pm3hZO
6OV9d5TQpuY0mLTr/bxUxhzRon8yvnR2b3+2t3wvOXo75IfLqq9XaicIQGJUky+5QehcBxys++ck
7t04bVehllK6Ixb35b0AaX2Wpn4DDzemTo43ZWaFs36+0XUW76ZhEm/AGwWZ/UJabzi5IBrHD4gD
XdaefrX/3hu2MHBMCGFJBa4w15cH4eMrAjx+p/v+wkdmW1gf9wC/O2n8RrPIHw7WWPUMCgGsk5N4
umupvmOhbgcdTedKO3Y4hE0FQ74uGESlSY7DktJl72HNJjGH25ObnwVVp1F59wjKOubfn+DcaFtl
LqDWb694yeE2Ivz3ZydBQuNDkef9iXsLQ+ysHaU0e+Q9Pwru+W1xur+LeqVAGlwgeoJhiLvoHCBc
8mvf+XPvV7NBn7EA6HA+IzZ3mDU12/GZbiP2wQyhYcbMjaPTkB7Tmt28db3ig7zU0wqU+oe3xpx5
ePy2T0vNLXWpeKnX1O799NpD6QkUJBIOCFnP6yH3/WUaZO7JkgYtW0DRFMr1NNWPg7hnwXHeANZz
NkG7m3CUmWZ5dE/+3xKBvAn9A+Dfa4NkSNnTgs7UVikNezQ9u7jD3gZe/evYEl89gVnVIa+T7Fs4
IxPzmXIZA03/LnfVdb/0R7LNwEO+U6f45dVX48mpcXK7SNyGCeqEfOsDTSojz363G2EMoWhKPcwb
tw/yvbd5vN//zHcLYtYaeH2kcPhfcKtrL3FHNj/6/XE7Tkq7zi+WZ6B7xXu8H7NI1iV0wugXRfgL
roWi3Ak8De3cZIetS/2MlCy7LGhEcnPcWSXApK6NFe0Jd5BjLcKXS+WoImjxZN+OCMerw0Qb8zO7
M3O9dfvmEY48UmTcCDWRjR+YSRDNM38WC/ywQsP2FGRxxkt3m46LExLLr2OA95E7+rigmGr4TBLf
yOfCsvmeeRwmJks1b+cgPlCQs9XlfNKc6GZ6Zw0GfPObRw46BstbUqfv904v6T8sjmdJ/3mvaVSH
EJ5vyeHAncfPOjFCUOGbSy2CA2GTiAdPqySHzTHbZOVRFBEgESk0tV6OtO1IEhvIlN3HarfWdiVL
GQsnvxZoVlYRh6BCo62a3vVbrH7/cH2v7F/Sfp+63OYt1e+xy1Y4mlr/Zt3QAzoBVLdYxslKqfGS
IR9Rz82bdQoNauUNNIwFZyqGbGFprYGBgmMRiLsfe4fOtRdK6d7QpjKab3g+cvfco+u+rWxj/ugw
o1/pD1RNW9kmeuBwI7XhsBI3QtM0DMcBaIUKfUKw/t8UXkU0EcPCV41SqNwTo7A8ZSJH1zy7puBu
yzTsTN3FbCIeoplHCJWaz8TKGxsL6DECS8w3qal5Wv70INYq6OVRgjq1lmaiyrBGCaRlkLqoJt03
f51h8qoLSVm/sVeUjLS30cIRjdhPRcPwBEP2wUhx1QFGLNJsmEi3gR1k0kQKqNz9O0jBZQdJzWka
Ra2Td0L76osQO21alHi2QjrSvZvjtkSVgXe3GX8CZHG6JNI8L8Iz+7IEuebbs/YdGiavgX1Ftndu
W/czrlIgAuv6Lrn2ynP0Rsl0+XXN781Gz6thhxSbJJEH9Mx0O/9Knrp88rFr6Y5fXulfZkJptGhF
YhE29U6KWCSWNbJZPg1kBOTJqazTO8VgUDZ8Fu75JxR0eKTPPsVCLlDtNwEMYrvU8L7uKy6JQe/K
mL8l8y6KyjkNJpEnhAGWO6cEOHw+g+G9XpflN+A+4glzcj2HQyOlyPutlXlYPmnSOfO+D4/LTfQf
I7itx+cXrN6pY+HPvjhGhkltipASDu8l5pB/6kb21JRmP0C+JZE3o2LE+UcXqbw2OyRHSyBmHtWJ
hfTfMWe+Tb+/lNHHMWYKGFgpSHCrVtVP1BljK5Hd58rg3q0/DseRpkqomS26s9JmFdQr+I3IhOKR
RrxuKYnunsb89DQXFsb5ITiXMWj+98tscW8mb/HGfw35IcCqIzbLxsHfMYwxZL8W10WOheDqT3S8
UEaAer+2/VpRkenVgHkOm/FCg93EIpP/uQskhBHK7hQHlSrrEdS0ldAiEt5y8/G/2BWzowmip4XP
icHhpfEkvFEF6jc3SYRTu4MGIhxUvxUGB3I+IusjTQ+XMa4gnWDxZEAt2EWyPLatuTp6VVkpoGqw
ckrdsFgXk858pc/G+PGARBBVH7+DYGm3Q8c6wdLlI9KUQAbUBKxJlWGyVo1OKo5fOHeGB5TGxj2Z
QIptB2YOUUS8z1+guopMHwtVVKxAFxMzZjXq65rW/RLhg1crUtwZKEphOe7nh3n2P/rAZcyQ1Fx0
MgctfrRk/5jIRMS8Yp6JFq5z+bhmTHHjgu6Sx06hDLpE71iSbkEbsrTcCIw79XtpCwXPy3f2jvwZ
6VieUvWDUFNvTDw0pGSiN92pmOaQxXJDZzKAUX5ohHI9v04Q6qelATLw+FnYMrchgmGJQ4F7Mtm3
RP2HePTG3QUn6xPN7mzrK6A+yfeeNU0cvgj4c730MgMBIUrTM3g0FRw8xP4mIT5R8JGWWE4aUJ9x
Ap7AQvvd9BA797E0cuGdCtwX+FqMXJjm/NW+0YWpFka7eYwuOcGej46ifso6+PafmVA2l3mKlmK7
fPLNcwd1ezSU4YJDxbWZgWU26j9qpecjN/tRP18F3UkLVFi+rNjzBrKVdi8ybVaNcSGu+2HcUP2+
UNmJ5qQtMjbsuYc7jijtZwB5GQvOAPxkNxEZYCmvfjLSsgK+G5bB9D4g2pb7cljKdmg/XaxRlzZS
r2aFu6OTyUlJSOkpPJrGqJvHxBtTq9uUSYB5Cp60TOXmU+wQrF7vdaCWJF+i0kdKAFcs53RqZd5f
lEQweAFd88+kaWVLnzRC35F2kL15YAXTtDUDom6tfwRTkHVKC8aekEWnI9a196eV0n/zoM/h2yV7
smFN8T/peDq+z3Sxo0AoB6wX57Ms2ryjLr3Cbw4OxpZhTBu9SmtjZmEASGRe0CGC/puVZJ/zeHg1
8/5cxIECawdNkIrX58bgZWwE+bWi3s8Zipv89i/nlduDb+yeVGkX69fW6JJ3SizFZWcPAG3BBTkB
iBUbQON7O0ewRSSnAJPrutjl6xPKIZaKJGAxHVBobNzayGh76rK6uF2RQv67H7O8W4izjlwnIYu+
HcX6y0UnzKccdm/VrHADktDCgTM8uuqPUNhLLJnna4YihVpgfm5XZaAl66SGgpZ1UskbokUXuEk0
qdbXcGV0mJswtj7i29RQpiKY8F5RYTin4vjPwnnCrhqayuqYceKdG77OV3q0NFfCScyoDTWBj75y
XgQSzYcyMB4eW7gh1wvtChK9KpW1yeONr6iXSvPAtLsyFrW5EmoF69r5A/1Kz7Po+cta60JAyrux
obM0QyH8RbvwMobfE6xNXoXU3leHbnZ+I66tBFXYYzMJNQkxViROOxHOHnbFsDNU5SvMyx/9NGDF
rwAVAnSYZA3pnrl3WikE2CLOuBEpYyxsl5uMC8YWMQf1WbGxS8rhTM6zfqgo/mThujEQeEhQa21X
Kl2StUAwlB/TMVLsazl01bgHVpvs3rpenyXpLeas9FIlbkPimSxrdr7Tsf2KxBuX6QYrQ5ufE/ya
Ulfu1wFLLLgXlpSkggXyqdWSf/fiPMuuY78oSX5yaRYuLVd7VEGVCg3/LGf25MOc1uhrtQ031Yqa
krXpxGZ6SLWi+t+ookDXrfbm7HL7CtMu4p3H5qQLJMiiRakgQX8o/BPwkfQbUVeIWSIpYAzWid6g
1o9/1b+d8IzcKIGlm0N/e72qY5qOq1Tg/jYEed3VMrPpesm0TNs1UnTI7QQiC2b3KIp+N5LanDbR
7HM4JJbI4qgpVzBjMhJCyRHIVbLqVPyJmIIqLobA4KFyb9QyfGh+IKmb/hyWwvdWcdHTzZK1x4Op
mNXW3zqB8enhiBXyglrcpXFlNEPInMo9sDi7YfwnfS+2VVwHizdH4HCpTC05zNDg2+xtgEkabQW9
QlXeL0CA7NFMgo1O/rEg89sNoVjQUbaSzaGR149YKmHoux5AzNqa3zxPj8/J/KLaLdjOebaMj1AI
iR3gteJjxWf7/vyLsF2N01fLlCE1aWo+9RfOAE83+GDwEHm7rVhUKmQRpQwOTiIoix++WIht+8Wa
Dt8gsFrqqrLIBqv4FwpCVEX5TNYJuIj+BJbPHePIErDUc85R4D8SFHjB/I0axPi0pDegaI+6lBC3
mLrW87PKYUOQczqGiDx4iZ5dgFZaQXM+QoCTVIfa02aYaR4IvxY2w/u4KLYlV9YSeFfPN3LWZWi9
20TlsUuZQNk3WG8+wUdCWU0fvreEmLoBR/zkx8jIQjJsQNrciFooOVhKJfnQk/8+eq1nyow+xXTr
7LIwV29NBjLflnlGS+aMOei13Xy8/watN6LJ52SeJczMuarDaNCfwzJSsP91meqBGnmICSp+MtZs
5zYDIasWGLINxYt9MT5vADBnlel7LAdi1NL+AKvxD9Xv3mWcGpW+FbHer7JboN0/p9rDN1F3sjUW
V/Sjr6u5YNbb0zaZuYLVppKvuE0XRoYPs7d/Y1PE8PRWcfbYSuD/O1paaPj2dP3l6THHoxz73AIO
9nywH35ilGUGZF9zb0gqBy9asjNFvelbnOS5TOSNq3DGeJq9N9FjlXxsDwqPm2S38iGtz5vwjFLx
ySCagdewOknxC1KoZZkhOpWHJWGwTR3n64hCx4ssolYjOZrzKTDpzd39esEW284ttnZb17BX83dN
3hOb7J+MKqTflDhxBfVux2gjPI+TeoG5Am9DFhtOus4tMql4HCDy3kagF6Z2d0tYDduMtsqHLE++
W2EqX8tGxu2QfIQWTuvvmO833OYpSvm8hItvoB/2sAPnA+t4S7Kaww2JzEPpl+0/pMt62naFTxZo
161q2z9JLv2a7Q1ZFXgEjPuqPcClLoHMmAdOa0YsxBcyzXgbq9LJI6WOaVfNehB3jxtZuIkei+Mv
da1ya3LndvFo9AHI9ywR6NDwFXJ13G4sQpYusPmpKk6ZVipet2myb3TdVrW7lxJDAARBSe4AOIDo
kFYqfB2Xe8dp3aWY3AGs5LzmAYEkY/5FN1I1J5fPF1bb5SWA1Ibl3n+/0gR2PzcPWzu7xxHq6BOK
Vjo4ycVB3hveXmQ3wht4GsE0B49jlGpT6en/8pPRdQDuoQFGcNxI72waSf/MdjTNPktFvWQq6zaG
6/iW3K6lL5eqImylOYDWcMJSGWjaKkVWfbKny4Sd9hgM4L9E+dqBCSvL//mnVJLcs6+gad4TgUn7
SU6vM0KmYI188CBeiex9gSU5ENYZEbLNz3pc/KzKajLT5Mg/NnSVCrEDHhH5NAQvYvnecOZl3pAG
69OxMr2FI+U502yuL0VsXhtAOVkvIMxeW+CQTaLRwA0psxMPdUZypQDbFqi0FVTz/OTB3N8KvIvq
VoIEAoc56gRkuJ6kyeTRc7tJ97nakXtkSnonOYPRfBsVOfDItuaWcKGmBiFNxrYOmKb9mE+rzLF4
24W8JTWhU34G+LagMZJsLrOC64THtce/BdvLP8VlttMjxd0Yqe8EZEjry/CWry3FED2FXSSCzDPp
svk3xI0PRC3Ok/c+8c7VdrfLw0YgFws+0Vu/DYPn+zWU78Je723Sm+AixjGUEKNMuwfg27mM3lGt
BeaNKc+doM5bE9lLNRwz17Sx3NoxNPn4SzYaVsQKtNMDX3AmWGJts3/ezWNEpd4Bti3KatrRFOkK
8xeMugv0V0JA9bjUgFXNUV4dwBqi52UljsA55p+IvwDgK+ilZbNeD//3IBfplpt+3/cEUZHBwwpR
gA2Gg0Hhq+/m8HSsLtmgMTtD3UJ/gOH0vyuAFHzCg/aivrPvPLnL2KAmodNLNkJzzXZkKITFvhGs
X86An/F/X1+IuWkgG2DsPWSixURdR0Q+3iHJ6kDaklB2tOFVQ/i7rYxiy6sq1CUQYGe8kprCRv48
7rCE2WUe9EhlJOBQLrW2/Tcn9jwFCNjFjKD7PDiql247bFUGRQMTC2IAAf/MDXiqxxV2ustAwDuP
FKEpkrsmU6cmTJtgQJWT3l8y4UYB1VgSaJ+yHasPjUxeD0QZODqm1Zv+AFJGPvsQyExlT2xQBEHv
aPPWRIIVnIqmpGqpmxnec0HrLIzvjHNboWGhNXwMPoUTrkld4GFYKJ8kXVr95TpFbQcVgBvkpKzD
PEiTbKd/Y8mR8zH88nKxed+PaMNOrL8gPtgVH7H5u3oH+KizRQdFMwfkomrg8KpDJGhY6OBZCcpz
JnrnKGxUiyxHgRVJCJjMjZfgTdT53/kpGrtN8Ka3hlA4wQLW4A/kzzai/9zcQc6hYJdhQCUsgwSy
ZkWyyZOAw7sT5YU0ugpmzRZRAfgYhLJcEOUW05BG080YS0+iElLwgvkHyLCCSrFXXYrIYmxpmywe
JLnrXfOtlaJWj4INnzTbGGCMv1fH4Jv80OaPSoyMdyxowCIosyw/gsdJ5mrsQRDPrGNHSgzpcSzX
wq4MpHNC14sPYzORrSmyHFvohoJ/TLFb+G4nUGJeHIqT+P8vqS47SR4QqctuZFWfmeo10IJeEieL
ywQSKoUPfbeEzjTYyW0aRnmn07ntx/x2Xt4hQTeqU4XP+gD1wWEGZ7LC0ltVtBxFIFQWtW1JxJZ2
fuMKP41WH+CnlT0CTWvEAKjjEE/a2GTc9GkKx/TeReQgc8spVu54an/LdNAJCSv25pjtfmyOc/tV
LFq7nn2Fktxr9PraSS8WGQICdcs8w4CL/0S+vINYPoK35MiEZa2wGqcQ6klXVvO0/+dPlgT9DFcG
ZFrmc2Z+MX9O9uhg64kwZiJE+yMf121NQKQ3s2rhFK8j7UiQKofJoeqcQ1K0Bj6f5Y/FbZciFMNI
ZCua3xmRDkAplQsCODvK4a1bOqNb5W8TQtB2lvclphuQH1tmO/2tt+a048/4ZamTZ/t6pUgzg+pQ
ak9154VaSsi8fkZKu5VGzqzE7SGzIsp74XtVw4yZ/hlbdI1L+3rgdnEe86XGXaAjVx75VrpFE3+6
hp+4W0yi38Y4nRhA/Lr7aGgoQMMi/qDMmr30WvGp4WqM/EAXxnG0gew+YjYUJjQLRsO1uP3Ckvcr
vifCjcSbdB3IShvEq0TINwkCZzfIDx3ZmrEr0rWsqnXOjw5s3ypFus3IYzXDuPRTyOXf/NyUQbOt
royzzoXBxNiX4RWNJv2Oz6nUHLNH35IrFWrnw+GueaxpKiRtnxBJmZ3LfxlHdxy6w6cp+HAZvJTF
2kxOZBHItSXSAsCtbb+gziFF98DR/9eP0CqlnApxlaUWjkzPU1foR6M19uZRaoVdz9Nl+ZOwZGEB
lLkWBsifvWfUkKoakyfsc75de4IrT5ukja6sN2GVnJRx3b7e7QnbUdDlBOkuCGnoEP9T3DPXLGgR
FiEYBIlxEsHFI8b6TlUre6DukALtXhd6v3gtr8fCdiwNbaTeZve2/aHgXHR7YrLZmrZgUuZCBdZp
81aOfTehypZt7X5Uq3uMfFxZEhJEsson8q5NGesnmDYxbnFcL8tFQjoIesHQax2/RnC113NApYfX
trtTcCMDpyRwE7E+Uxe2M8jrBgVHKs4glVimVqE9WHxdFMRMtDrLnZR6hxQ8ZOxRZoCyMYwvlfaB
bwdsfYjFnO3Gnz0042n6TQ2YvKH/CAzCnoVeSiyL+RlYMN7wTTbEzsxzhdntmiTIXaZfW+VDaGrX
BmOkugjqbs/G+rw7JHjlQZLlmtE/Jpvb8dVnpb9lLru9Q58VE165nPUQ8t7iqlaV+6jqCtPjAjaR
4K8/8RMYueCZebjYoEYsxEPqNfwhZSkYd9Hby1dyeR+8nvfbcJFV48/Wu7U6bzbBdmiwoKzCs8P2
kxZp3pgZKpMaWKmmx0ruyRW8b6rbi+HWxLAOvrfHGV+9e56yQPfwarkLa/nvKZMkCG2jdXZ2S7g2
uf2RU44oRCZOmzUo7CanCFGMbVq9DSUqBR0gTbXhuCSiJbk5eZcAYx+LLSkedxJCwEnD9fqQCjtQ
CFpJpMKxiWg0U2nsU465yPNMuOW0c7qZ1zUAlX+Dy6gGpp4Q8BOqEjmPrLH5DISKwT8IYnp7Z+3x
sdCdhGjMcPmpr1XjsJXaPoFgZbNC+h4VHaZZ96frhB572zHjsgwAKPk43Aw46iFARti3EC6WxR6k
ZK+6LO2Dx4QbzyjfXy+a6xe66dsaNhYuUuW7bpjl37mCRWFXil+lBEx0g2jL5+JMKkAAGON7mcK4
JtAbTlToBNeJ96YHutgwOQPz5CMQ6dochWNm0w7kPKnp++Nhg+g/0p72Oh9Z7SzwBprY3eFcN+a1
YWwqG4/lxAXzmLazau0x0orHfFyb4LLlru0jmelg6ij6oDK/vGjqV81stb+tk9nPA8GLbPooBOg+
dioP9ciWv7Q0dqGVbtIN40IiwEHML5fp9O62NP9kUGwNeaHj3SohaWIBRHikXirAnBZGhX7asByS
j7maD+usNzdFJdOfG1gqHlWUSaGQ1HjDvGQMS75QK1mjav4S2qY/5Zjo5dlqgVa53d6nM7DxjSnx
Nq/urLl5D12Iyhf33EG7VaSQmbc2u0h8x91io0WYe2Cs2UHv3UJZiWoL+2tcuXevUblZ2WhPL9Zd
LCSFRLPHYDuiG5A5DtSqoNpN7Cs0HJTc45lZv27wLyl2whsfti4CuGbnuYwQRY0bqTbR9Qj28Txy
OmZMv05p9XmkGPfRCtViF9ue+vdXQXcVtypEPrFjB1VwDcCv76aBossnp4ZnbnEwFkiC9zk+O1kf
01ZoiokGk0mRD/snonEV04dQtCsrRd4CjJlO30Fc8RJTV1ys02h6Zo5nr6Bn5KQYCLQdLphpqTlZ
tbJga43aCGaQJDBfzO3LGQ1Qel+2tJJPktAus7a9HzIxXeubEj7/47vvnzN/6uXDcVry2JfXWO3Q
BTlQq5yQG1YtKmSUE4/M+SdRZvYOoeYFtnPigDR2LTGCxE664x7Ob7XIclasvQ2UsjiWyuaYrj+q
zCEoqhKx4OAhMkywtpiTDVIbYv1tP53N8Z/Rt0rBFFsa4IGOmF54V5SrExqVoM0kSSDhk+eSMuIl
Bb2G9QGpe2Lx9yseLAOnya+owuf2oFhSE5O9ptGNMefhgu7xmGuL+TTcyMziQziM4k5pI3dUXd3F
u4+L2CLR6ASkdX+e31KCOswp54y78VgBlIrzM3C0l/Rw4hHIbcT7FC1uHhNQEy7/NcWjroi6KqJh
s3c8EPjILo5bhXQh7OaBO5k9MRK5f7vTON+4PwsIL3nNsqVz63ms8nBdWa2LkkhRrOXLL5R6qHyV
w2qWv/asqBjM6F5p+t80umvHeSA+RibTcLrLomBmifa6O3GReLJZVFrP5+GsoRVg/N3hwqI5cLcp
6ERfPUMVpSXx7J4ikvqvTytsF16BduE6S8cFnEMzv9mOzIAmySC4wYnVkUcKFNoNFpp+Fl+WAKAJ
2aOvKT+itpMOy8zT1O/aGQz6mrMsHDsJ8teLYHxNrrCQV1hupmJ5UCKH+O4fHkjPa5cc/VMzvwhM
/Kb61zdR26YUGOfHH2VPhXa/q09yj87DNlEk3u+jRvfteXL3MWrYVlJKg7rw2dOReE8lqE1/jiKi
nH5takoIhHeCyKF5mODQeWMlBUZ++SV9RKZ7A9GIOi7l/bvFKrlVkY/yEgbLRscvS/XQmKO69W2c
8TBU1uJhQ8d/n3aUU760IJ9gUNzBH1mOlqUwQa4q07S3Brkhhz3SYFtUZb1JrkMLGHC6gtd/msOl
6DL9Vmj36Ue4j28e01tkpTpioJwOXH0PyjneYtr9aQZ1bYlwr5aTCcvzcwOwHyMAoyMNJsjOm9Kk
uUOxqtAMwgS74ILo+OZ2vcGVZlUicfjEzNQYLgGG7mCYb4yXw3vFVw1Ytnri10uIW5RAC0v6V2Jv
OEqJghGgmzS7TSLfvqLiKcWLsZIaet3Gl3h9jJ9LjEm6vQNJCPd3ontPZAsyHNV6CjGmliyUn9oQ
V5lm5cfY2nvbSYPk8cNGLRtP+kvV4YyrZrPcsRoHjf2fN+zsqaZP0XX0aL9kM+Q++52elpKI9uXa
uOtKhFWtLripnBD8eYnS30Nfv6LvGYO7u8JPgkpQYDMRn8PiNF6CJOyXGcnXhtEGHhE4XZST/xdk
hS7+TzbB7Ix2cPLoPPJ9tap2yMutWTugXj/mkU7ttJU4VzdVmj32OL7fpSadPp+64dFGfkEcHw9O
uNCcvbFE5XSrIKboS1kedglAD1LGyI2gzxrjTxhlFqOuvYPtmTsdq2+oPVcbCQhpDQo9xiGzS/xu
1pDTtOtKXxMu+thXXwNUiNn7SYIowZHLRbHNu9H+w9pYuM5Wjy3unM4c43AKdkWthFW33ouJcJhd
Tgy0HNLJoUpG+gr2LmPQKzKv/+ScQKj3SfqJLs0p50AmjFASMT5D1IVNg7B4rvguBf2EhmIp+0aT
FDGWHVdAVBb1It0ff8OeDQNziQ3HCynGkVbsh5J1Hzl8GbHYOFZiUAput88jGhPnD9CUQiindNHp
GTkAp/C7mR3yuXeweOcSgsmYBP5BDPHYLr06zS1bLNniocVRO1n+1DyPSFfrCQJ4MpmI366chjOr
9fvdF0UzcHFQPiFZBOI5e5fY3Adu5tHu8d7tATmXgujuTG0Lishy2T0k9B0mCaU+fIFd8OjgfIaK
4CD1lwAYkLdiTl6uZ1oQdkZZ7V6OB1KwER4gVzOiwbdRvly+//Q/aU8MYfNkKhth12htyB1YYuKp
RmiptqiweSf/oxG6fKwRyf5oY+QRAG0A+ICnpgGQrSUhY4b0zgfdv3TziYTAXc1vOS6Adi3B8xwE
th9BaoyBTUNNk8Mf4u21EoM6nic9OpL4cZLTG9aVMS/xlcy0EvM4y7P8Q8edQhq1aFs19eB2S3Kt
jsPdCvl1HxMJ9BZHkXFXyH7UN93z+U4j/yjDNNY59AgfHizFbmXKihfRUMVDw6fwnhzRK7p3z4ug
mALgIVrusmxJtokrt+hOV6WMMdH1rg4+dEfQyEeO66WAYr8vL2UgOAyYp6jFroIlCkjMDr+P6yBL
K61Sy2+VBgR5EFf0HKKSDy1NZiIgj7v0WptBJerUSrXSGR2F5sudfbSgRuGgx5fvfHlZ50vDTvj1
m9gqSEEDzkC/chZ+iLYNiktt/yJixhPvtEM6r1wnfAYEHg0AbHirsZ+qcEYQhMKIGmNNF3oSk9Bf
K21+0O06AZvlPE1ZcKiLQPTB0dx3hqpYuuJLfm5fvBPqpAw/t9KehJOMXBtNHU3YbXyw5y7nF+0r
nZD3B/IGdGXEZfINWMbCbRsXjj2xDS6OJ1MYxN3am9myPSmKbRxodYJq+s62nLvAOXjwsKCWjmPa
MFdGwgGkP1Hke0vCYYakS9LuNKY2Bkb6qXRQwFt23lj+vC55PQg0KhA7XOAHn0Pk9dw7oj2J1tSz
BbqUlmAgkcOwCOiHNCiyAjGz3qIM4usvipdrp324eXsGCXB0lyADTaskGje5JwvrBMfZV3/y1E0o
+qpdA0kPTFE1GHJJ6d6wyjsa9mCxem/clkkTvxmVF14KQOy7vbYUv6++GEmmIMBrs7AB2EMipl3q
fJCtu5DeqsikvQ/Xe13+1hfXzkJxfQV99EtjEdfDsBwS31YRQAfTnH1D60XcvoT/4WJ8LKBsBLtF
JNvdBkI01KzRNWoQzBKWL0s3WsHo3H2lsqFzyw1VfBW1xb6boOGIhtJV4JOqKObNUj8UHi4pv9Ua
c8up0kJ5hqjznoesyujtTYXJNCpJ/Bw9AqLRAApsHS1cmw07jcCQeu+zU04MeMReYnFK5G5PwePj
SlIOBIcSnyRrP3vqaCx72rAYMhvXq55wTOUu8W0cJaezo+XgiVE2C63qwaSzSa8YK5gso5B9d2zM
5xnxIjIcEd87q/hJkRJy5UOTimorCExqLQVgoPgWja3ygEcvqCYwSXg+iXU3h8AN2z6P1+JFEY5d
cxw+XpeMNeXQYf1B82Te64CgAjGIILDKsPlg+2KtXaoGQQ65ZvXSCWS+q9uqzzbLG+hvhpJ0TBk5
Ofxtdn0ZOjl81FLIJOgRgsRoAUXAHekMQx9/ddk1Gj1my6KkdNfBn4f0AdTUwbvaiGokEsRMDF5s
I2JRoNkhQ8zZo1ltH3LluC/DdMuqDTEph3OOorDNWoptLBql0e2SAT88IwGd2vpq2l2qbCGmlTw3
BQyLoAjQ9FWRa0Q+RmiflL1tjWfeRMxdK7qfvmKx1c4RuqQqVKId2F3xKTHFHUdpyBmYEJdQuA1y
u6QSuazACHc8TRkGWYZeGA4HRYycWapgwWMfmd1L52irSl4goUpi/2pQ0NrmIryDeXvJIc51rAKE
EQRVjXuwWT973YHUxbqLNE2iddfrOEnyQ+3vPjhkaBRPHrjMgDr9jDBVkZGtT5J3XuIhPHt63WUb
DtyyRQxeSgQnxoklMwln0d0FJqjM/C0eHwDYWPKXcSXm6nIHgdkZzqG2tml5Gkf359UODcp75zwC
MlQTmc8cQ3kJ1MmE6JARal9BurfCGCTWpIGEab1xgc7C8rWGPFjP8Menw8o0NZZ2qBEGS1t+Z3lr
ichbzrsEuI9ATllB8ihhNoO9YzJYLsKieMftZSIU5U402GGwVCB73/Dpj31UVz83dLnAshG90vai
QEcjjHaPImOdo1aAVITPKsec8ynXylolSaR42WaOzKQCLuVevfwOTThGaajjptlKm3bRmysH1LMf
eqduGG8vHERP5mq+v+ohJubIf9T90nak6NA0ceyh0KnoqonMfP+3h4OPHcdDLNWrmiLq5fMado6r
jGgSG9X9BUe+/pwCbHdE4fkW5SbMpGf+HsFbNHdjBhznSBt/kvg1XfGEXNwqlpibNbd53wEGkoli
p8jekRpptcHGPH/LwuT9ySWZ/92eojBRSekvw6cmraN+xjsOJchBAAViG85xxgQq5SCfAPGdeYmr
GrMSDJyqbnb6NrsOrmpZi6S6PZKtV1lW/WPpgQJsg70afZH+C7pztRNvKlym6YTtBfF4VuPu6O9U
xWZ3CivtDcjfDQpn/L75H6AP5oULQP5eErW7oMJM54/cMjzkxNK+agTN5ykb35Wjhl1MnFDXJ6hr
NNinydTw108/TrtvsMwcqAucj5lIWkvun69QM3IBAjhpyIVjnX3XA1JBVONY7p+oZX8dKUG2SRVa
MF7h9nOdiRqxfvuKnuDVRzqr9hl2m/bPtS8ekRTvjKSmH9vLTNqMX6NSr+RD8qKFdMfVE32H2a1e
8yToukvzwJ3074YL6ocsh1VxHuLVcAqVvq5wAq1HDfDsGAJx6KPPNHtI+I438FEk6pw0Iq7d0T+b
/1XmequIOLgK9XmZU+yxYQHkTTDhpZjfR12JOi+j9GzTD0gM+iUBbrB9iN6s5UrosVosbQAZ4sQj
eLJpgnQloCACtZGacwVaqU1DcjjyG+CBpokMeh295YoZG49zTIpAp8Y3qfqerfRL5d0hkQSCiC2O
nZhytY8gUCAdm9v3VOfTDqG5IxsfuEK8dcEFRbgYcAwOpqYlozJuxTQuxZdEtgtbGyj4Luyg8Pqf
MyHxwpE07ecBxlyDvm8TDTlo+H95mjq9wk0MQhLEAMdHgTyfzOwO7w6YjUx2aY09qJuwZAZ0Yuu6
tpWz+o6lrow0xnEsY5P4S6p518Cbe6J+NUObSLhi3cG73vUNMUJzA+C8nEnJimyXzJ4bnNxIs3hR
ns+WJsK0a8NZ1uld9mxNU+/UzhCFUblMGRY/hHVAEK88eQLqlPy+NONpnznKdhsudE1nkoP2H8i6
ykyPsnoZW8v3inuxBt2SQOfXS88/TQfsPS5P46TCT3LXWhmFKKjlMdcQp+swtrIvQOQaQOXe0QRV
tVZVsou9m+Do2SFc7Bn4P0UIKlFUYSaEJttKCrNWht0yTX9OZ7rJ+nysQ3qg9QNlaEvChVngMHsA
RAHW6WiVVxdnBgCUiL7/+PpBbbmSomNqjqDpQoBjr1JfFLgQ3JH2AntzjiE496fimbqBHjglMgFz
LNOqQL9oWSDGA0JqVar2hkRvjqm9USz5KfK4u2D1rRWevrcy4fbMcljFX7n33/HmcGZIm89X4ku8
Cq9uH5FyUP+zWLyRMSYWA5k5IXayCxgy7s1uKjvO2fksxPLAuvG7bdJueZ4ctqbmLq6meebpwSEy
O2KsMmAwab/f4wlUmLKMvi1viD8TD9lOVXGfs2ZsLvG1aQRcel0WVS12B1PLFdjBNGgZ4Cs4azih
nMFlLwCQwV9dpyW5vT5pewfHNq49aZ3qsuK9ySU0qwuVuaxncdWO82QMdvIOqQP1Q7DGN/bfmCHs
+xDXdBEr7cj741ZIats/uKI2U3dDl8opjs+jYOqVhEUvGCimOrb0w0qCrDHT2UKfDnO1/OIsNSM6
QYdtrJ6KcHrU28QM+8ymQXPXvjhnnu+zweMd64VO1y/Yo3L/iY0xX6iyD3IG5/DRcE2/bzZ1ilid
fjmzXI8w+3z4QO/H7uJll68IZUtRr4iX4K9pQXXHP26bWlF6XqTCzkmab+yB9YBUAh3K30C+ElYo
J9PGOQujUL58Uo+X+aEkcZ8MOU8lLUzsDcvGMx87OohrCoPXTYrtZf8IMdktZ9wbw9lEBgL+9lZD
e//pRNA7FW3rE5P11nbpM4F1MJZ6TormfAON9xjq0Jit28mIVigI/TunzOogdb2Bw4AGS2bk1ow6
jAjwzWNgFYhxNXQ51cr7qVdimWGP9usspJJB7UbDkv7UL5+M5Uym8DXNfMWh/bUUSCojnc10eIix
b8jHAs57uPGVrLB6FhqfLOWfVsWygGdkaqs/UBi0joY3DqWVtg71n8+Xe9SOXw8jrdhX3XCfAVd7
MzTRAJmgb6byzgbWXHAzSt7qRPKqDZfJ4qhe1CUjlY3Rn+pWePoipGcijrpvatEVjx8qQ+mtng3h
3uhrhfJRo64LmBDr+jEqEi3jrm6Jjii0vgDlCSqBFqqOPKNylLdumQbwVzE+lLvjVjnMYDIGVdfx
GnFILCR7jsfgvNbVd98xZc1MEPRx/OIvgWvn9Ufl3uEm19JMU6CMqopuwrslKUZVrsz2dqIhhva/
pYoSzDlNaske573mHmeodYoOIprsZ62M49Kw8hjPF9b2E75ZrQASubvL/7wMU01qjQugK7Bynemi
u6pVicxbCLWLhVmDfEcy4WfbJW7mb/kB3UBE3q70tnG0sskTz1JS4Giybm3E8sczycWOZ4Tk+/F5
YvkkiU3oOk4iC+54iIUTLkN4CjG2+fcvpYCp39WEJEAo30vj2yolkxgzUd4GxO2s+EHA3Wf5ubWG
Xa4iFJ+PTZrbzPtuUaH/tlHdhgusIxtIN0J+CXcV5Sd/IDN82WC+z7LSZS+ujG0Nc61AtRn4aqNj
ESv1iGSWVELedIKGWdf8aFHMFlB8KtgdqWwu49qGLY8B6yXYo8jK6vxb2VwVu26fQD/ddbbJaCG+
sGyPBcbECHGiIyFMFbZxgnDbkYz4BvRQUeJyBzu/DeS3M9xTEN/LqVSQpD++miz5tMCx8JPghbIF
ito/ys4oBDmZH4UEYG6E6swhds5Dx0IffjJjRky/BmZwnElArV+rpIdvg21oOD/MJm3aft/n3zDx
ZvSdYKOIN/QJxv7y/F9tX+sfOr8pP2B9mgYcj5X145uj+LS4J9m1CjW0yoNgBHSIsq8zNQjLWi00
IyE0mCVz6m603yb4KExBnkVnOk5BlDi5YHH9/6iBm2Q6Zx0IZXjgV+Tmc90C0FEAVVlFTj81giCm
KolxRW/ZlHiW6vqfiG/YwE8dm2GjbMxsuIPw6qNg1SdJ8oJKo4AiRdhZc0WD6xBKva3Ng0pyJLVT
XsyYM7tSKhYsklplYygP8ob4Jf+aOCqdnldCGgIBrBS7Z3USVqkvcFDX9EerCMy+d+Zhb0WcG9Gk
KthvTuRPJyYa1m4RT2WYiI5ewfiK4aADa925EDMfVd57+Zr+1vZg+BMDRQaMrjMf3R8Zfg4NH4Dj
NBas8Z7ZVFWiFIECle92BZeOeCNa8N7MezMcf6PADm2r7d829x2QA1ZGpUF3qKKaWCNnrloipFxg
TAKhuB12ehwK4TqMsGPG7diPly9xjn2dPzEB1OmqvUqLLBZZ94F+sSxZtiR4j/HGVTUenFvsNO4+
i6KyvMY0IKwroITe7LOEHYYjONouqdzlRzN5EzrgJybIvhNlYcpX67fOFC8oCP6DH6A001wzX7Dn
/AurvJiZnfUYFIxKZ8QOtABh5tnMAsGrwBJhyT2NcWJ3f9vkIuu2TGn48Y3bMuZjcmz0eTY5m/qT
vew5H8DIGzGx6mtPEd2lpx5qhe0ADa+upBM7etEAetuhsQCiUE0Ga4vUUzh1No/rXwAwjzXvNyAB
YZgmw4/a/6MCR3lA2WzSGWRuCjaD+GalSBHNBDeu9G7EgY4t/Y/wspk+UW+ivXqsruM5sMpklOsr
W00fOqx8oQ/TOpQJKT6OmAyxiQ62c6Yshd9BOTzE6V1A+IHP7QfcWYTa8DktcdZsRxezyUOJkPlt
HpMIV/IvPSAa8i8N+B79AFbQPNWWlZK4AEleaxjQJPnEyItvluEmpGAES3V/5QtplWemwdGV5U9X
6AZB71tfAlLtqK8UfWjg8Pj2cwEgbUreDKu8b+HyD6T1KSTJHZO6CzY4NdJszRwcubBiQbYpK7oJ
8fA6m/wlVHccC9sU6kqKHSVbX00K7RfUrZlPvEVC5Zr0fABlTCk00hujufcfcamJB1prssLb6O5h
hwX5HPGkhwqKAhHyLz2zYS7rIimbW1d1ZlcTs+p829jm10DCjQZIX3fxjQfR2WjApsxdgKf0qOJY
pgO5Hfc8T6tQWMtfjoC4hFqfW7wJuSHpXHY5i3qJbUrZFnM8P2qQkjvRARjzhDKahuCxQgaZBTd9
ZFRgH3uEHHSqayFYW+f4yXlhuXXz5p3AF2hDTWHyB7ef0GzdCmsqO3KJkXMw6PqZoq2OG8/fCuap
SbqK1HEVxi74PN8zmmwuG+fDsEc+8gYQd2xbKsM2zFDe5XTIOk3p6sUjmL9+s1VAjHFxyTwsQ9bC
JQyfzDyn1Pfjn1mvBISpxSlDAT8DV5eAKQ/OmcV9p75l0A6K4YdUw6HMEHdI/HpLdGzidLSep+t8
NF7U1hY/6XLZecIf6uxf8iBEPMY92R3K2Fw35JxPxJRlBtm//yuKy2tWrJ4XuJkmPu0+ptTz8gku
vobTIaWE1h2i3Uqr75in1ANZDVlS8bfaY5BjasZ0d7BDqkj53CJ7Qfg7Wmox4adF+H+PM64JkcZD
UGkBOge5aILCMzLVatwFlNiiEJQh6jCODWa4asvSbGlzqzOgBKbHPye7rnyAWYPnba02tizNmhbg
OCCOG5YtNX1EIUxEM1Dn65mFrphq5UKXJrBMchs+bMz+HdwEA89CenEGLqgyfWTaVKYPb51sqGWc
U5ljQDCaoA0BG/E2hHWwjXb0sQMqwWJHRvCP+IAYWAfoKSd++EeEYH6bCpkWzgDslpWbIlbWr2W5
5x4YCR9do/El0U5fDkhnjMjvzY7damcTAs1pg/R73UwR4naLb3TAJlhUJESjP3Sfpeooln39FsGr
2u2cBN2408ocx6kQVpUGafTNC8VY55NpoEXasjUiorwAwXDmKD58m9WcH0fPIXybz+FC/toNwj2d
g9iDm/BYrmEWhH0FlItL9kmRwvOQasDqNZv9BVr5pbSl+bmg1mqneC4xBfGZkuViVhyMe72E/XXX
GO/js84gUiPkykuKd6mZBkBOv/74hwE034NYbE8KzWKCzb7dsPAURoYGXF5vZJbw87pc2wKgPiw/
r92joIDwUHC0/rQTaxKfoQayeZwzmNJ+LZCJR0QPVXXARk2Kf25ODH8pCd6zBje/BTGFqx92kwEM
RBiD6Ck4S0DK3rXpaGvv23kTBOuCEIVHd+9AlJegMkaFi9FEJJY/YQ5oIp4AEzabVRdrXJSd0DXy
dShtY72U8GA+tcDkUmjHJlBNuHGM3VWnbSNW97hr6aV5sCdtkQJ4pDMeXjIXLj83dPhXl4W26uH+
rpxIQwYWmLQcSN3sEMg6Ug2FvYvHsUPwmwqEpdj7JXBtDjsol6sr/pwcAsM3AJKI8i3yD/GDJNtw
UJqi14BxqpH33DWzGhdQCXGis6mfov/QEgIeea19pZWWD9ItfjCtt3+dhkuGd4DSwCTeB8760hK5
XiCwEcerYwMrYC2bNeefbwR+YGVcPIsItHcoJutd35yBSj8elH4gdjOZtlp10tCZjPFa2rsYQBY2
+SBvNXsNdH2CJCyXECOtLmG6EJ+XQn7b4aOElqs/XI4Z7Q189QngcRIKoN2ON9v6FbsFTLA9e7xQ
ItMa5Idnol33rv6kQBveUxrz/go9Yod4zHdnYpQgHbnOrr8lya/E6OM8+ciDn29JnOkCou4nCBRu
PHH7Wg/rBRGB/PaMT1sDY2BTybJN8PbR6vdE4FxF9JkrFPDqlieZ86+A/c/7StWUidVXiAvyw0oa
j5qhHdPQvT5l/RjEGcyIDEOzc69umPiZogYfpEmAjxyS+hAup05wAOfhecwDCfnEmncnAhzeRLPG
sDFBJ7rZCkN+4DSYtaKCmvccF3NJe1WnsH4rQh8QuSenwTceXcFWVEFGauYKN7mMkg2/JoltXIWI
N6LOJSV9zxugLOOLx07QPs4dXSpaOce/wvxkHRvfcu7o0XeVxyzfqJzv6enrcRAB5uNqz/6Jmvx2
8e0ALAVbGIsvlmPHS5Gt48robWgQdWJrkvwvu5vKEbJw/04/72cwxLoiiB7wzC7YG5gJFgVwejUA
oaBm393jCIRv+vPIQO0uieNKYubWElViL3AMJa0GlfveDJKF6wp3dT+V8VNJVH1LhX/XjlUFDHgG
H17EaADZaKejGYWfQuSygePTeWDfXIsrh1sfnRqH+3dths/Sv+Hq4cBCpTygxPt/MwOAXOvpu+De
Lx4RJ9mNtA1YU7xyJwoDsl35uEgfpRaRk1uhSWIqbOk0g2gv7aYZahqKJFnUs4eOQkBgwIZtlqsH
CXAtl5HrRv60g2b9qKluct20oF3cjbxJZQdyuTSsGSkuLmo3y7jsGrJrPbFEYgbVgIDEAlGigYHr
+5nRlgfkB9IFjGNHcPm2pXHBePC0K6brVgH8ReRHBkBlZ3lPaGu7EiM6FNF0RnYBmdhroKG3TWHJ
YuF+Pc/PK0TGhjzoHj+qnydlarnn6j5QFr7OiROip+eFeaeNyuR5MKWeH9vY8UuKYa7vaogoCHnQ
0zr2vkDMdOeWHEriHWF+fH8rQc8drDAYcpAfVslWYXsE8Hn2G8BvuCAxr0pElFudD2cmxDz0Okls
Dz/2mXL1RQ9/6h72fhDTTp3FkkJDc3o6mJiXffFwBUua5BCStfCf3Q/uavCwVYgcm0aoJdLVkklX
pXKRtOQbHj4N1rzIsd/YLEM617mNX6UfAmXFvy6wigQHGQboST+H8Uq8l4K4cEz+k5ohrhItuoBB
TgOPbWeuZ+0OPVD/sw5ChO/G+0mPKf617Fn5GW8PpNQJ7tdfx700ZwV3dc/dfnrxVVjJ1818PR5L
Nu01fd5Ut82Fc3guvIet/iEtpui7RGrFeHxF2eOzpQkCfWo4I+hkYv4HSEKdNkVnqzO4NRG3gcjt
5OiCcs2QhRQVJnIfnaA4mTHnHOXUsod2tDlCEteEfQB9pAy1pXJ46lb8iLtuO6zTPYlR1nWc4ymF
OgPJvd/fMWxGQxJA+ZVRJ6q4SOpqCu/TR0CbvRdA2bUPLgu3W4o1y9d03B6f/AhZO5U0NNyvOmUt
kl8qrP3HMC68l1j8gCSXvaevLa9corBT+eJk75kkEHXRad6VIOqxFNUlB2CVE0C44If9H9tsdxKo
tAAoWN6UHYVQfmrZArvZ/L3ouUYsrqOqfFXZaAo4zgLHP4Dn90lNnQGhrxRftw86QLGguEfV5kdJ
y80bfwsBLC1zF7aywFYR2jadlSsU4LN37NhuXj6Gi0/DcPCSDrGuA8MqjpNJDPDXN6DE1izYaWoU
ziapNqDxIBbQulykewy7jykxibsO/pmjLG2VMe8J1ofI61fLWixAuWyolXqkSBI2eJnQPo7dSDaE
mC0xwVZ7A8Vq0g07zPXih81eSyZrWh6hFH2ZEYESZNhpQzJucK2OTWa8FKx67bXAD+HBCI/rgXIz
5vjFqDc6DOnX62eByRNdyijRr06WYWCKV960QQzLe/6KrJZQPEppzO5jht7fJ1S99fGF0Kg0VZ0E
vbSIa+etrCx4hWmZmk5M3LQYN3m4yAo+1NibKM3oohJkQjE229utXELlPU5M5PdyaWCxrQGjAk56
ktTpY3lCpW9uVgiUQS86h9v3nLTPA756rRDUzfIHz1ogr4un5SQJIIOan7cX4S1DhxqFmZhiwGfO
Jj6Gs6ACTFoEaXr1yL//RbR0dw11nlbVwxnZ90T+u6HpIOCNIhQUqkqhjjI9SL2t0YrnDRj3CSpW
TY8ia8Xe0KsqnwpzQwfgpMAogPrGeYR4Jh7lYY9NmJhdgA4YasiChkhY/dT1R+71xiQh0EUEIfAi
NEtkPCnmdDYfiJo28IpTksD1iCyExUT9K3+Ep0D8NX1gz6npfabkObCTPdeiosj9cJiuMTythGdk
B5np5tcQj6UUQU0hwcYxdcWU4zjcBHY690Igg+CnCxYuokddG7cPk0vME9jj+ydnqbpX8Az37u8G
2um1G7IeYyGCU3May0FVyktXenT02fgboIBGkYCVwv8NvtfacV+maqSHmZUO08u6JDihfmz0aDw0
CaXqNTfTBwGWOlmmzOVTGlb+Nt5xi0pUka6EdE6hlHC8PBF0JiBDHdKVx56O6BpQ2Ric3Mxtfqy6
3u7DyofG0XfVwnBHK5JkqCad2LNcK7QrNfhQM+L3fzs7KgYDg98SfuRuVIGBtDDvC/fazv7u0uca
/bJ3QB1SvK0P8shcoTGN3FD8zF0mBHTXa3+RqB7fT1YtLRmn45sDCVmaM3eRDIQNeWdhXQcuCXrM
FSz6xKeyJbvBxMdOFqOlZm9KaZQqYylbJPTyNsbki9XX/JUfVfosLm7RIZZZfi+YwMfNoctyYvi1
TB0qCZG6WO+FMDCDwFlqgiaRlXo63RNfpNJYZHzVqC3C8sqj57HfHFzWZMZbSNeKdnvd+8Lt6+SC
trbnPOFQOdV36GmBuV1Byorc2qhjQWu6Nu9PErpg1b2lVDHJPhFZxLXAVHdvMyNWtvpgoaZZLUay
daDKfdElB6/GQJTtpKaPl6rN1zZ7DjsBU5sYB8RYR4TYX/hjGSYRtazfQtfr3KZDEL7A8KwXAZ7m
YmQZRX1q4eg9GDqE5Lv9ZqqbC0bCWPeBN+H40HuvltGKUxEIUzg6XufWzt/j1x6XUTaZQJVaoK/O
Uhu1aXdLWdaIE+vaC79FGFiEAVrVU2t5PYIUMeOoL2/mYlxCD6ECVfj8f1F5RkHGftLNlSa5KMRF
3dwko63shTmyYzXWCU2ANpxzQjVlv44/+widYkTHbp8wHGJe/87S5/RDkuUF6YnYSkSm49RcDVcc
5HH2PT2VR+BszbZlvPVGCJx1NNHnG7fJdwAPMgltrvvqdH8jgaVNNWb87WRjj1CegHLZafCi8Eh7
juTvACYVYxM2KuJDdZRk/7T/O5t7Bdqh41/TY65+aScDq2I/CkcaoXChkIFj5TGXm8BEW+XKdwBs
pfW1moT6mS7mhygJh5quYI0at54z3AZFNYtOxXbuAKR3pHDBlTgTZzVsVKT8pK5C3ZPPz30VzoeW
zLp+jySw9rdVfYu3LCb7wF3g8N0LXaS15i1WED46occUtCoqG9I1AOZ3gRKrMJMhdhG6WuQj6y5A
WayAzko3T+kmcoiFpz130G+82L6h9gpkumbjcPDxlKRLI5SqarSzFi2HUCueEVUL+BDnfcuAz+eN
yF/0aSPdwKeImcmTyywdAmgocn/McDZ8QaEyN9oewpg8iRafem4iH/TXS3lXNNEtGSzd4JcujTBS
EDubAOR2oWClBTe0aHnUN442WaGDI3WPG6bfYnC2Kc7tNbinE3Lv8e6x/XxG9zYxVfo3DuidHeJM
tVcDXOi89CO+dVOIpuGrDCHRccmrXtdcub85ANADGfEctIoh/URt7yQaEm7ATwveZLo19WKXECew
A9bO4tkF8b2Ro5UsqlnjrOfGArlidu3CnGFYXbtixNkjkyvyiDGcTm8PWZL9Lu8/ri6dG3B/FbJY
NH+pJyHsjrYjlot6e6VmN2ZS6wkHbaqjDfrv/FaTAWQ6ehwLigEPjzGJ8J9WbbXvZ8yv/tcksHau
TZMRs1bYiazubeSToH+HKVzpcFCxgkNf3gfAkrV9oidHffPexsNjsiT/l/askZE3PDyVaLHlZ+aX
Ipqhss5TkfmHP898861/ygXx7wIPwl/m9DTtyz91hjQcx5N6jm5Skca/jMy3SgJm8lqJsKxeMPz+
EzItdyi9vkXdch6Qw5MtO6Hbm4brJ4pmVNo/nOWC3JKYSRZYxYFMDBo5CKpmEKtDqweMFeXh5q8F
kJ1cX6n9Jfwb5E4Ir/HznzVO2gKNRRk+wv/iodRbFijAxCLHUqQ24JeowLk5Quscgeci8dGJHQmk
RdaKzNGrxih6NlZbhVbUU8A0In/XsvRIYNAZrQp4XCzi8UL1+flm//sqkdfKVLBJXwil8/3jRa7L
jpW7iN9lm9ufOSCcxMduOR7r7izm4e8BfPNwQ1xTv+cx4H4LZc782ZNj6kpW3JzaGj/Imch+GWoV
QwjMTiF0HCwIM/jtvr9/SEAbr0u2ppch58gP3SATN4UIoD7ifR9IFVKSVvWljS+mRfMc1s/pryd5
RbqVKMuFb7HXlOOERJi3EQYgv5wBo1hAUOrF6M93NcK0xUrRBY4lLVtC/YJmSsbyaJ5fNheo3cgB
trra0fBKBq3egeYbJrmZiPa29AumS2Jf7LoKc4xr0nnyQubpRp9q349fwkSDIgIggIFpMXkFpGUY
t2/Wi+EuuuaYU5yv0ciiBZyYi9+UuBvPSKb94MMjQzR88sMUya6DXQAID/WihhIT2xx/QWxdDDzD
Eq1LmlpNqGzhCGqwvsii+p9xO97OzBZdemDttdK0tBuisoJ/AFyStOMeQE/lnl8VC+HxouX0Hzb0
B1WWlEqVCfFO12VyfN3CM+O3rT6YgZn7HRYOdbBKkUU+pO+0t/663HN6yWDy7DZVDWr/iN5gjtq+
nc0aVL4/hWxtWKc0tnk/vh+sS1Xeqvpv3ExnyjGbVdOowKo/AJYJN9ls1+3gXgGepjc777dgAsNt
6cthGs3eWxpP2jr2UXbdQBQdTTWWIvOU0eX+/WoKBUsbYov/HkAWTRuYekVRFIXGzy3lnSYiPAKz
urky5wvZjdDf6vmQa+fttpazxybs/cE+w9cLJbwKOeodIcxp305GZb4mLJffScwdDsn5GFVoGid4
CRLkjCRRf36ZRecddMENGrJyN37Y1YmWADXs7I18UXhN3U1YNo+g6GuPUAeuiLLplVXrerW7RNBP
OTMaqb0Ft3qrrhvjXBXco4yilKfy7S3DI3seO8COFkxM+DDnaXhlVcHD3Dxnt7BdkK4DH1rNz6p2
OI8YYagiHe08F0YBQqQyVPMSVtGMW+/pQeqyisXfzdWUSDszUqG/F5vDgYbL8vhOrfn/Fwqg6DCP
MzT0d8xrRf69SxtyWbz0cx90DTMKXozzGzRcGbyt2Zk9cFj4e2cMLy3IIIn4Zv5Mmx3XrQxeFQ84
/qo2Dci+8hoyqm/Y7SvFGIJ9urCxUZ/e9W6IqXxOx0NWdHvVEVM5ZtK9BxdedWo3ug/HyQxWmUX6
Lha6BeVqfluUrs2kKcQdvj7fNfemYBtmntCqyjgNJ16LpJWrTsknT9oJ1/5i5sctVwcxQNyTsonV
QCruAVJoLBEoi3Qzv/cluQVaaLTBAzJH4mJ09icRxNuxr4mCqKWnaeBCcsJ4Jc+SWAFGgakk0yZj
F58TyD6cSv7Et34392viMTtag8nTWPyU9+Kfj4B2WhfLD0HnNcV8z85AfRZRwea3NlSNBpC1CFkR
Xn4ZzaCxPsOLq9pLf7tz3NZ5j0+aQAKcvg+4qCGL2fdgUuPZvJ6UK0TVx5PKR4Dn0Br/Ua5zJA7+
n7dz2lVECPvq6GiEtcMjgZ0jsTMwA40mjU+0J5L42Yw0U0JsJHfewwe7y2Cdi3TKL9O5dBY0SGko
SN7I58Y68oUwCP16dM65T7N5WqH64HZvXvo9QmaH10glx3xyp0qABsoUCB1yVEKQCGX5eg5TZ8+E
HeBvbkq0mQ7XFK7bLa9U7VXx7FakGEeFOAgNA7nZjpIjTX+bWvU5oRpzsBbUCmaIzjKjjgEtC03K
z14OxTaIyFpYc6uib+Q5pAjnyTigpd6YawGj3yaACL7oddU0zL8CNad6ivbdFe8Bwc0RLUl/mAxD
PsPUAsTwF2okNpp6XPRYDwy564fKn6+kCVqVroEoi5cTsS5PwPW2AdRk3nL+pzw4Ne7qmPn9DHk1
GBdhBWRnMcIgRUWKvYmB6UHLeRJoiiFvJnvYXIbk96xpQuJw/kTbqrafcTDP8MmfyiF/otZ9lksd
8+igPDOXnrmRKOly/ZAPNg+WVsK66BNBJi3AbLvNzNUmLSoIIWX2mZNaVuj6lc+ipznXPYaVZo8Y
oz+8ahUq1s/b8TAMbkgqJsjKsh7E8bvaWvLcMPnorMV5PSCWJtyfydKD05F/32jlyXxV7B0emw8H
hRn5YN6YhmVkevRMM4YyM18AxspD5OlkQ3ai2LPKj2+PlKFt+dkANtyBouELcro0l+Etb381GezR
FUoxQ8ZoYSoHGnohDai3bQ0zO4m+h8RK+TrUHO1ojPq3mKfbFVHRuKPRlWcrMjz/s8Qb91FYzhgc
EntbaZCCWuaN3zX+WqSR6IVNnMMh80jLNnzX8u+2qvV5cnSGiRRgLDux0hF9NtIv+YGcKLwAv+bd
pFllBwVIClpQHzeGtp/7sBmxNn7WhLIDONigb73rUteifIZ6iQSe3WxQrZkuC3AAsrla5N9r9qYv
TuoA8ah+CdUN8tehlbm+GqBuPtAlbUBARxfH3dR9VruZKAF3JdcWXAxXqtKSdY8vtuvwO5RSuTv5
qam2RoODohlN5jQWSOksW4mTcYbDdsh8c8rlQVZ1PKQPA/4fiVN2m0t5hsOUfKQfUwuCGjMnKqca
5ej8d/ulbZF4l1x22siYabL/gsUt9+A0YiJ81O0G5W8e9OW5+xi9PWPSZYZnAB2AMLh79FXbBEJZ
b7EgY4lmxjNQX/sPSo4l2tci3ylPdgjA0tOPFNie5aoOiocreeUgJZmQuEsaNHH6lpUx+DOt+elj
cOyFLhzbn9CzyE4G7QwbswThBB2bpHj8Tk9h8sy1tMIO/tTm/7K9i8bwaVPM13pzVnB2lrtMZDd3
7J5eMKVeMm9T+pk8EnLri3a344o0xLlylkeKWSxzpU1YferSHXQODei1oVN02vqExtTObDf7I3CY
U/ZIe+jtvNA9lJkklpQ4mNvxvXxxu/LZ14QSCjMg0EbOyUxsEafLyXuubFQJzrOmYik29MqmlYLS
oQL1c6zHgml4gk0twfEzEp4s5IcfUSC+qUZ4mmlWUj24/YOLhIW9palgY7TgInHfCjPbVeQ07gY3
8wvejUGVMe88fLc1zVOOTMywGnKwwFA9/zUpxXLOihwaziaEVLzaBQjWXe0ic76IWzHOhDnexRDf
iYqVfjTN7+ovy01HbtLJ+5lqherNS4nFqiIzUUYFI+FH/OHmWM2bKc7t/cV8gL2d+EBKkntHMQ/M
t0vV3GXUzzV5mkIvQXqquLu6Dn7IRcyyUAcWYifywqLtq7JthI61gE9BVtrBGhsnXiQGdDD9T0ax
1GIIKj0sb9ZsuXbVDsQPbhv+s6W2H4dRIAW2hLGcwNs98trdfyjCNeE99e9feek7ahGJYb6Z4QxA
9EO1Llbi2usPGDrYDQ0ledEo5vbcDX68qj3KM7SPzkONEcG5TEty/siPKMKQWUcZLjAtsWrDBYsH
GZhB58OWRxbllF21YjURa/s5YehwSI8aKex//EB5IuLmFjC5LS5dWnUN8Cc36VaWdzBb11rKnBqL
jZEuozly7ol0WwXbL4AlGLHQ20V3zxOdNTvlqsN8nEfaPIBMbIJ/pVmX+sWqWOpI+qzHQiJkbpVg
6meMdBf0OnSVqow1YdexhEQ2mvl4XCYTyHb/+fcn7E7xdg/i6o2KgYEokBzv28bnCnMVw6xFoX3n
eVz7FIQKh2QaP4JNEJkRJwhRwxahu/fhlYFhflTmwAK6fujtrBI55PIOZ/vFkgNdEzjlBKEHSBLX
oQ4a8/1FmDDQ9img3biQPveGMo3bHAptQte4hw9KADK8fWbShPFdp0/cl/vUdVklv2mCY9J1JfXT
vssA7SST20V2iLJMETA4d4n0o9gQmMi2ftamyJFEutmJqipJyZG3W83q/DKeU3L7+BEz1p7HeDn3
3N+AGOCH3wYm7n71hDIFKQlil8V7O4yPVLWxjB6FvBDtnMxS5FLi6uxS/FQqTngYOZ6VeBAx+qA9
y/jfE7NNcL/gM684F05DB32Q2vzKzM94x7NdQc0NQt27z+9CFVHySm8N4eGFBHnq+5/J0tDs4AWk
hHXCTWe0pIOFhuyPJs7z1oBWYceYHohwdyTAuXEGgcZtV7xdo7z09O/8Y69ZjJoujsgnyu6MxJAy
JaQpAg0Ht5FmgnfBOmxCKoFWYFag/WRnN8uYjJDph586sg4/8O1u2gFlPNm5In8hcN4cA5TFwFv9
xHOWjq2YBXK/vbX33sdOSRqHhQGJfT5k+HOARH7vt/6zit2W4t+9JvScFr31vHmMdpix7NULAuYI
KQK0uv8BjY5rxwgU/P+cszFi0w5cNxMkQi2qzKewUmrD4vj/Q1ETSXX1nsHRwaqsZwJey8d6uhPm
hrXLeOlcXTAv2BVaJ5Ikmc+asv1M1OMWjK7Cd8ZV7RcuH4gBfbz515qnfXcrkTVRHnlhyFG4tvcQ
603lZe/Q2KQz1raw5G60oFy+ztyQofFwbxEE4IFWlmIyCD6VqdoWtk1xRbGuX0QBzljRx3iGWUGb
6B3emMlwwesViy+BNKVrdXzdEChPtw0ncjuagReBM2NrwjeUuTdR3u4ybqLW8TFchIStM+BiJ63B
KzMqbZQzkUF1syYlXLkEAKM90ZvfcqbnmqD7GQlN7DyCWh2vWyKdrAxB9tyLFeMu68/r1w/66pKK
rMJs1MfTgUxl5tb27mMs3iok/ZCNaBfSJtkfb/frg0UjMHZvScUxBfM+Urf4OJ62CvXt6EXySqTI
a8M55O9ATmTc2ZZJ6PehfRv5FUxeKrK6SaI1o7JN7CC/zlXXbdIanygYlYIzNjHHg+QgMXzNJ0CR
AgcF+K25RvXFfEHbpe0SJdyJCVFvEHaEgV+e8qwi346X4txDoJY5Uhz6iHn4HYtv96pEcD1mi4PZ
1YzSe0zd7zCZnGE1S4rCplcb3hMoW/eft0f7FbldOhcqWLoYSJgk2MKsSEkkEp3WyGeKjeiLw4WG
7JNJts2ZY7WFdP9o7lHSizPGJshr7KJQ0bREIl6sVBeWbcYflMqk9ej9HHu1BOG7K+6TC/O8Oyhd
caegwm3stzhd/AnAxTmjQzZnEXT22HPCUAn8fTb4yKyIv0UAatkuyhARIZoqTbA+CuMOG3YlL5Fz
xLnpFQ5LYNdgi0FocNwd+Ux8j0qCViW+mfQZdgaCEMsLwo/CJ+M84ApYQSI7+IJw+4vR9Qly7xt2
Lj7g9MBJlCkbzRLHCNMuJEZnwui+ewkGuI4OMIp3AgXzTZJDOD9ppLmvq3kgQXdYvpaavaHWUQtD
4nE70/U3rRhntzYgj1MRcfG/xlUROc8WBUzYiWfcpjXw6r2A9/vcYSRKvgrOnZvxarXc3fT5elJ3
nEUyK8ntU5QDPCd9Wz4e0QXncDQDNUizTbDPJFXKLpii48Qtf3jDDdOTUBKBmEAVD+794jAUi7FF
pMPZqjetCfSAaLIfi3lQUIGdXOS04NLTF1pUUW5cZ/Fw8xQEq3lfJz3ODbnA1pgNBSE6hpKaNVgn
YHSUNNiHKJpQGwOSVh0raKKW1QIwPQhd9Aky3HMLA1LqCA2s6A7vIBCH74IN6AQwNnoNyxG32yAp
0Cfg2HevORDF27VamOEmkZApWfNewjXeWph6PSgU6tCYvNNpVR6b5H4lGqJXyWzjU6+CLk3SmMi+
Z1k80WgNwdzg+isqmPX07OBtp4yAWVSbN11j/XTg03ClJOt4tXehH2u9MaZVj4cy4KTRhReRkdYf
2YKQPnv0uxN6YpGNCs4Kc53JYzGY5+7FykpK6BmEHImzm01d9OZDxoKmLUfZG/k9ZLCQLF8svAJf
1SPH02RrKaI72G2UAzPH4epjn4ygoaadV5qsmIcseisw8icGkUDmbVoGwZfy+crrQlAzgmn2+mrM
pU7K2sKt3tk73FSaPrvKY3Th8OKFiCLPoFbz+ZuDrGwFqCGEdO7hQgPAQxPkmqDStmgn2VB040Gd
Y95E7jfCWbHJoLqtodSfDsIr5JR5au+7Zy+FEutA/w4WQLcIlb3ThEDyU04Vnoll+wzvv8jLJ60j
lbjPRtEQTypy2J10ADLYvGX5jE7TsLwz7EsDaWTm6/up9dzm+J6CT+g58PEAj+RzPKyvqwN39SKE
5eybt8pS7G9wNmhGdZMvdHylmqYU69EA6I6YMZajhlCgcfcI8deX6WN++SKDRpEkNMK4nf3FEhGF
B6c+YxbdKrh0TQWqT9ERwe1npQC/fazvlMbWW0w15iqex4W0lYknge7Gx2SEDvLKGnfjsF4D55YY
R9gTRhDRL0DUSPjPP/d90POPHNrg6WxffSb6a2fClPjiPsx6OTf4triemwhepW9RxbWsI0fpYNd0
60a9PBZmK/j5P8gj1z3za3p6ObJjRBiiz8iSde4SqwSCavk4a3wCTkc22MFdDFJE1ebf846F2A7M
+A/hvrzWLaR7V0cWTBd5vyyUDyEMvHQYjT30eYKg7eTA4kPu+rSPIo2T11GU07gnmFMEHMVN7A30
gQ95tRiIcpqX4lquvRvob7TvAMQfBT5PdnEciUEszLPj5M5TPa1fyMf/OzMlrn5GVL+z6IP7QpR6
3GgMdWbz0+HacOg6YSPfbkybMXA87svzA1HFoeo8vfjIOvdB9OAxzN7HPkHPl+XuyTe8D74x9MoN
WRDKuzcjlg0Z5UT1W7xVVpq8s4VD7u6r5XkYDIvgneXHUGnCs6TKjEuAcy7Y3g7/UYdCKtK+mFT3
lrycoDsROHgFxOPvAUx7t8yr7jpBkrX/w7UyCCgUiGPD2lADCvq7s/U+iJmENDblLg5PrHXHQdMl
XtoOBSpQpXi7rFeg+YJMYMUjfdzBcuZtmE7sjdGHIjVBs/Jgl+NqnUWTEJdJWdCT4bXLamgc+mgx
PaUoqyGJsNyfN1oF9g8tFHj17ZpJlTDd02dzV6vSWXxB/t+V/w0N3fizWnzovf729zTKZd+/1yna
LmEKQn8vRnGg6pStSSv80JWmobtYtFk2hHGngcb0aOAhMXDrDzb3d0JTeBHowyf5zZbErUsgEwui
94Fks3AWbpK3nGWYXRp8SeGBXmXrP3OlGMDISn2vpmGJ2X5GhOc4PyCphOlZFdwPI3rE5OjQzVKz
feKUgrcZH+Gv9L7s6RfxZxrg1PdUp/QEMhEmXlB86vKDU8JPyPnC+XMDxuKQ0cMyYKgTwHl3bq52
xys+1tq+5QA+BsQFboo5OhQmwIEt+lAVr8fARBxvbCqL+eq3CxEJn1utv4gjnXNv9SuEIq43BsAD
rKSZcaYimhMTYBgWTTJXgp2A5Mc0VR62dk+42+W/rFCykOP+2sPKAYi4HIJxKnLmd4Q1dBYII3ZA
t+VUua+eig9zEHj84ycO3ZQZw643R1Sd0J1pKzXi9MOvDiAO/szVSLlZDauZi79AfFijdk9ER08n
WbGV0MI88j990qkwEig1N/90vXOydpDC8txFu1dQhyEKDufeBz+EcGUvSsv5fUMXIdHlEn9gyCjX
7VaJpb3fhhKPRsTL8Evhp2eLKi89G2BXQYxHuiPXEGvAasCOf4qp5CcG8Du8ANtFX7zDmAkxiexQ
gZKCTnXfbHpmE4gWB3DEdyLQUyWc9xowLBxiuufDJ/juYjIgjbjZoN327A15+rJEs9Q1usqJW9Ay
R/Ie6oW4/iY1/+0JJDzr6fVONo71y5Dj25hnnVhlNmFXbfO4uExHaxrk4nD6DzCqimThCIScyrxN
G10f4jendrx2HYPuK3MU5T/YRy5ATgzHRisUk5c+Lvd1sv0C7o6M9ShTw6GWu7i1ntXwpf5sNFH5
5xn6wSX1NWp2pfjHEszkUILQraT0z9vj9z82cyTLyiWsWzPYXZLkN61xyRUxdL8jK4L9RWbG3cps
q42ae7iJ3jVH47/ht1Gv4j3Tj3T3jGpvevhYNcdyn2kRbzOthGkiHBaQBBB61LtcEHfz8Z9xpcb7
qZwA0YU4+jVZCvtpUC1BQqvV0PQ/D4q8tv9FIiEjpDsbn3WXpUp/8vIOmz7/kFVbKQNkzHxWKcWC
PO/PEnTOAQs20X1YrJnpE/2qZy0TcALP8cEWcZzr46G0Ri0zBvTM2ORx2u/G3R/vfsiYMzP5RvPh
BRWisqMuV+zQV1/S4Jdvm3xDuFFV1MtfaM/FmnCxy1CZme7qTLcPoM/ZSzJxdHOZk7lPuXlvrRCE
z0iLBkgnqffI7x1rhaoP9g29E1YRRUhv/jcDTkB9VgJSNfaVyqgPB1R3kkXQm2k0qWKs0zf7N2pD
wpbPyWWeqY5wMagyCsRbKqJDOzLXbhuuCQ8dttdnaRb3npg9e7r5P5wN3HdgoyCPZms2aotXtRGo
fegrAw3IMRh8fP5BxWvyMQpWWHV1nmSYm9+tLpIhvdYzTJtUFVo5qoMna/Rye3HiUp082Me5dBEd
bzIJqvoDHthZC8a33sIYMxnKo/U8AzfHLrvExWpuIMFYF7V2MjEnr8v7YCEgoUH5Kt3lbn0XkXuH
adDl/pyD42L+6A8Ns+JbN3va4M2RjSiOwhnaCCCSe60Eg26RzmNF0HvkeRn4rm1EHWkhaoEIQchs
TyD4OT14o5Ui3t53jkbMxprUneqIHw/alf/Eq391kU830BY9vNK8YTBRCLe+J9nbNrf4li36MRWN
GX+6e7dJOWsokGmLdxYxoO4AliaWgMGX3KuwqH4gNeDDMLxrxYztZr5BiviTGgNVQoQwx/K56heO
1Z+I9bf3ALxH1fUo+Gc+TnrCHjKNAGO8kxXNS/8miRITVhqMela+EXrFkYwXgotzY6HOJaMktM2q
384oCXtndh/lh1rdfm15Blt+KIi2dsecq5aC2Qyk2YOL+xWnXQ0iJpbY6xuoc4EPE9vf/Gm7Lx4Q
89YLaWSzyeHV2UWcSNK/YpKNyaKhGViI2pjuwQUba6Dl9PtflrW27P+zJNqbzecctll0v471fvdU
Dy1J864hUReo59SM12R24vSJ4d9sNunuZQMQ+PtiUzHmTF+C+bvEs9/ChGe3De63lbQS/Ol6RIXp
WRwlEOT6MlIgshTCfstCNm9ie/xtf/4yxgEsCh/+4+aFwo0VGczY7GygDc7AGLe2WlUwJ8ePOS7r
JNASb9AVQynGn6SxCYPdniMxUnWaMA8BXY+eo+ewyQOkvD9ppt9SggzNbLVuvdJKPlYH0kjH25L3
hZC+BtkA+iP6waUkoaVIYaLD6O0yQwWnqJ9JUMIq9vCm4k9z8wRVTKlZ7JgL23XOwc0zRYGUp4Q0
v3OqbAITqIRZxnQshwMslJZOxQbVZB3z3eWwrLhqdOKM7LOl1gYYSyEM+zedEiHQO9rfGCixu5R/
M1ou4Q/GDWOx7ZaugRfYoEf6G1TE6sfKTVpJuX/iazywcDZWXuQisCvdhNyjN6m/ejATlS5FHKvu
uADaNY2FaEHM4VmTz3oiSUHf9TWugO0Nm05UdWZlZV6k9bl2sRSpYID/m48arYJdT/MPE35xOB64
jQ8/yuLD2JYkISRRPas6BOdkYvJkEzRd0dYOEBir1VRGlPTh4Xufxl5hnQeVhBQm4DQpv0vf6lcX
r2inKo0V8FBtdYfeiql/VacNYYnZmFEcGAwKulGy2QoB9sB1DFMNkPVffJ1e68pJtl7PEg7bxmHD
J+Jw34HuAMCSckyKNVhdOmTnR+AqGcFExuANIPg4o5wE6X7KnFaNxOFBOlG+FA6wyofnR4ZNVHMe
jptiFrrwYJ1dh8bXRPkCvjNW8NY0+Nc7f0RB14ltAE+WJF3tvaXgv9KCqJf2y9sAv+hNC9kYR5FM
/dQjBu0KZqgAtB0ByzTeqU/Yf4VRl+RoC7QVmCsvQUp4vOtxBveJNU5GwzJJd1g4zrR4xXkqJ4J/
Gz3H8hVDuM1d39New+/WPSN/NBX3U1jzvWFC48gpapXJeVxIHpXFCc3/d8/x7nPFWxzpqMHjz8Qj
1LuISGY7X4lBH8S5W8Wq0VCO78yLAeAmr+tDWj25kEbTtdmCEx0qbLK0AJMddZofvbPX2HEAYfAH
SVsIm1vdpi0UJdnBEPtE7EKZgJjiNrsNWeY4y0oa/cgwKP7tNiN6vje96LK7SOGiBaamclzu62Ss
IAaWczZICn0hxijApH7DrT2dp8g/alBZZGu8XdvOp1YksqytRpjpP/zGV9jqjB64oIqs4b8zlEZG
EO1Jb4Lk3sflB4vPV0snno9rbfhBalVfvjqYLorRv4Cag3+OW54X2WOmD+28Y4s1+xGaPv2Ipmjl
c14W31X+/bDB9+yx6bu3Uu0Ov0aPkvpQnRYt+ymctWlSU/0yvHXkH2dsMdzwFPebQY1rV3r5x6qK
HrGHFgBSxukSgvq66TE/lIkbIFEAnFJdL3KQa/WXP/bcfNaGaXep1gXvYYg+cft3a2aRtr0uc8Oo
kJ7l1Feo/RoyLmlAB4GRCuCC14gRX+G+KEdCxJsLKQI2rC3+NUB0r84fkRVU38Jr2r9Thh1V4+Ky
K+txtolC+T0nnlAVuz4SqYCyAqvo15VWmk43FZaNGTq+Upw5+kpzsUwObdSbaHHqZZWr8StZKWSn
+1P1WqFBiWJ/LEpdoiCACAcdaK0imPYA+gIJyvleBcpnR6+jtEYcoos0eZamsCBfYOiU7/qPDP79
mh3wAznU29iJXn7KhxLept8bXjY5mkBns1XW6DSLM7qS3UEcxx14qAmRNpgozTahiaEhqXEgy7JQ
5YYpXvJF2+Z1wtWoRoRKxp0RgbuiLsFuNVCrJhgSHAai88ZIOtr7twgDv1ZjKHDWbPmevDyJEtwb
w3gqCMexm1lAMFcR2eK7i/U6Ffks8gOoiJx8ZJJA1d6Padg2tGpwtHFfA5gj61eT+05W9+C7XVu9
Y6ahwcPqp/CXE+2bJPukS8dgg3TeWUXkT5WyIHiIIt6P7jtWPXdYRgoWAyuOvK/afsfTerN9LWlQ
9Cm93IvODTzgVvsnPfVu9BzERJeqnG3wMXKQNoGJB0jdIAH17arLLHpF3gJEqU/zu0tFL8oot/i6
ie6ZuurwMxi/I/4VznBcfcWXc8TiHEOu8zb47GoRcOsujnCnHpwy9X7YJ795qpY9XwrUnl1bSeM7
1/Uh8SNJWwihr4CbeQ6PIqhXkGQFMbfzUi6yimG/nkYY3LnjpVDSgjghuazxZngMERl6OcA34H8J
KCQ7iyEt87FNArfYzLSUbp87oe+9iqH0DotHjfW5B0QDbZhthitQDR3em99GfO6e5Gl5Ly18Dxrf
4XQgtJ8rVMchpwpSWEpHikbYRy36FhQHVZEfBhz7GJbLNbd4Ytez8FfL+mHdpaaBjDug3MlEZ4Qy
mQ9fT+tU519DzQ238ZR17522C//jZzBWSlJpAwBu4C9KywHPP85LR7z6fjoG4kWg7zm6lIOm15Tu
FAFNSRmvgwViYiGBOpXLQa0o2E9bV0/Df4RkYatF6nyCoswBjgW6PaGVRIRC3VtKl22oxddS/HDV
ZrY2KQCgWdmZGL6/nQ/oRyfQ3h6ErO4KzKnoI79gTQiwc5BQHE15qg3wGiWnP6oCa0rTs9oc7H77
GA7YzN3ZBleHrMs5o1U+6taRHQzV5mnB/nglRu4jhBO5SDDt0S53vpmqZJJOyEF8aE+YHFEoB7HC
HBie6Zzq2Ac9VypmR7YjdIxXBpgbwMn9j++3t92r2dv9Hgtsg+WOK4lvC+eQ0FnEkC04dGEktMrY
E9srP0Otqr5Z7Dh0peB9lDGu1zMn+LOAqUF55llRuyMbHqSULqhzCusJyWl1XDrbbRJ66zcGcdqI
T3kozwIe2tgE180/ZzwxaNtXWvPF5I1fZYywqPjYFdXP8/rBIVC4WbvMKpS5Q1Fzeva20MvSCF1P
wpuCLR/dWd50wOgQNJ37jeW3eDAP8tiEJ3BK/0bI7a3hgQ85/cY2S+seb4fcd2gZlv+ZIOpQgpth
EoEbdkyTESlAwWYtHz7ixAESUryPDg+Imq39d1nkWF2utWvpyhvqZR0YlbNQFLYtJ1t6Eci54vak
MAxD+1QUQIzVLhbnnL7VAO+L3E5NbHVsYPIzPE/AxUUqia6nLQO47mJjMOgoUAo4GuDW2Da9VSpp
k5e6bshTH8cbZPMA/2pu2lEr52FqYZbc1gYLiWDRKT8+EeIl9X3+F74bbRBcBTDL2PM3i5wtdE+y
fiKpbUPWGQ+XhxCwNwc6VpWTnbTlcl9ewDA/w/pxFe3uHKs8eaTSiopjFGI1UfZ/wR3173pmQKxv
QNbrHuY3RnTWbOuBuwzSzu8Yv9L+dVjk9iBw4j+z9BfFmOqQO2/NOlF73Oa9OsoZOrS3NQtVgJIe
4ipHwXkjwEYV9owOwaBlhVjYQBEiIvpVTVAvLgnc3ReCTqRfWvXFdfDAVIac6LGd5Jh6RsZtlol7
Dk1gbDjRLDzGjHUttJo/vDpJY6H9aIRXM6951PQ6fCSHKo1K+BuBaLk/switmMvEaH5hnJhZrcqS
B7lrhdTXuCqv5oKf3kqLZQxI+X5XPAmP2hieoFCl/aTYNQ5lBfi2r/ifllmD50+nOTC4GyDbxMZK
Hu+COkb5EKJLnTZ6E4vqrr3bHIBBp4OciujcYKiQU5/vU6nYSxuAr1XTDG45OKwlZOiilVn8v8oD
Fom1xoOLuLmcUaiscZ5OptyfDvvyp7CrYXqdZy8sQo4ZBu+Tj725e15TyprXca/TL6oYF2f7oWfz
MsHa6JTvY14VpvWDmQZALSEzfD2TifE/hhbqshHxIosd9HA0v81ZvRJ47Hjeew6xEkzWYopqm/W8
oWiq5fQCE8lSb8ffDLaLWQcdElouVBwPmnseodVuTbsj58+oxMCdhgx2fpnbup5BGniIL2gHTpx9
6RO2qPkhYA612Z4SCauRHf/nqHWr1N47OUZmcRLl2lrxCkMOYorRop2jDXhEh0nrAxiz5OSs+JvX
W5YLUDK3XXTtVJgezR9lSjoY76ac3K/pRI0Fuczu2SUafXB6I988FzWIc6WEDv91fqeVMcKRhSML
BpN/XUKzCd7sPkBMWG8KD/dG2WAOGFG/htraTjrPwkhwikO6Rurq8fi0kzF7HdYUHMjKHv6ybVL+
zDWm3LL0lIDDLqQZOEgXIi2bGWqWYMPlGpXLYiszafyjCHi6kCO8Na6v7IMTQzS2v4twtmfKigDC
x8XD5Lb9YwqdiBo6JB5Q8nLsy2zMsPb1I/SsUG+ouXwXauMydU1LQOmHO6ZrJ1aSeVJ5EYlL2+KB
xtUNixX87++Jo18/yBty1/d3tXUnItQJqxf3g6AovqS8o6RyhxvqdGeTk6L2YAf18EfZasYcilS4
K8qQH6RLSu5Dvnmjcl/fQzpMcrfQWBiTieJUMpgkQq1KAquOSW/DG4bT8Q5iayoioDFdBJ0/Ewgr
B/gA7CjC80ramQNRX4f+4vOrz1ZBgbQitnatYHugovIUdmHzYEHo+I+xPiRcWaMQnZvyBDRQbYs0
jDHPRE/j2s6eCgZ9t7DFj34yFH6a06U7joOOHZ//b81X1zddfCEfDHC3YuRlV8vphwI7Zdk1BVCB
wjcq1U502XH5Ayn3BXAzsobgkoyzRZbxcXq8H2Q/69+yhU7HCgPk41eL2YiMcdlcRa5WURNrvit/
g5XKAK5dhlwe7cORm7y1nW5ABj5UkLz9jn6o2/h4zYnlHWfAN2V5nBm6ZinmdWTN6O/Iv61sPDuo
Xy25vr0SAoh5txpGlL/JGZOUcmnIJtAc11mAMkbAOh0vGPvyOy51VS8jgPK6amE/BCpFO/5cY5d5
33N7YmOYP8CXEkIF4uCkPIhAys/0MeQL7hp6x2mwPzbXxNz9IlT77Ls5MJSCVOdMXDMeA4g4R0HP
yrQuDdf3b6nr1ryAs+Vw+lhTfKb+4CpbrW5r4NI4IL7xLavsR7pFBiVMHk7QrmKPKVfDhpfmzd3T
ThhEkO2bqrSn7bD4wcOhFr6A+niM9pP70AgtK4hcsonwy/1MtyNnXXTLr0JOITWw7KI31pC0Ov/w
vdlxkOZufvvPWYnu/YQigBBkD60Bd+tClhfyEsslBKUMfI37D5rl3AeGuIs2zqC+Rx7Od10oveZI
02qYiHW/hvsLdAtcIzVJHwFLtTbH1NqMbfJhxueO+zI1COhB5Dx97Lq2SVDyb1rtJ3tXVT3eZclR
HeQwmxQkOlub/ihPtHk8/SJtYAb2noI3euf5keAgkIl7Y6lDKcp+ObA0XnyYOlcAeUvWnXSIq7Le
c0rZ9mc7TtXLNfxpiPSe0redbtbe/9TvQWCSSceNkZZ09ckbR4P7Rvqh6UEO1tEArZ5ntK5Qrwdj
ssG048NvGbHWPuKgrOrfv/T4pI4/7FL29zk9HMDzrJCgH1vHDz5rg/ZRtfwkiobn994uD4C9vYCu
OGlKCvK6pgNTfqwwrYDr1pwjeHzsmmokYa3XYzGJovm5c0H4XYnqdk9KhtKeI1W1wwpmO/TxoXj9
Jf7dqOb1cnC+5RbMVgJi5w0XS0bkK50oxJalGyJMI0zLf9iEJSBdCR43dHzN01i5BhIoZgE2m/P4
NDW6J5Bi0adsxYFObTPeEVB9QUm4K+dTfNMQlKlcDSaQrAXOOv8bm8UHcv6HO2PycQAxz3E1hLbT
aS9Zkc8+Fmo4Q9X0iOOQt9nB7kVMrCErGArGnhcO7e9WZLzizmXasNZsjdcjAonbbGiLLkRpWv3R
WV9qJtbcI/TjV6zLY2HO8JaU0KpLSs3dpNxm42r72g1kS8LjWxTxq5nXJR1sHCLeHZqeTayzoBcn
RJWxSUDsAuIzyCjk2QSid4jUA0hJ0pJIPBoyXpmLvvqWW7vQjBz7cg5xB08vsLsWUmF8gDOF0UaX
VZyWZERq5tLdSZzMrSqaX8OwgJViQRbVlLlMZEU/qc7JjfKwYnz3pX5M3DYcxMOtW4PN/5EZFosQ
z/UxM9y1W0cTWPjKzeFUk2rzOTokFvR3loHusdYnWHgoQwFYFoM8FhWrjx9rwR1jls55aR7G3AMA
zQwpjNO5Cj4XA8TgGXcr+a+7cu6n00e3spFdQhXC7L7FjKL/GToACug+mQoDrXhQN4EyeACxwTlb
5I+3JzSv9nrPfC+csjoyND3PvIZ6Cd6HKlZxrPj9bA3ZdbGzoPQOpIN2eS23WxPT73+tTdpzhUyF
2rtNoIbwcjH4uXn/BvIjySHz3vQt3h8pffVLsAZagWrFLRFga2HEmq1QQbG6uXpVmB5hoMailm7p
Wuetrq5GXDyP34WwARuVxkhec9S1sxwJKUPJQG8L63NNWB8s1J03uFIridAcl6MqaRVZgEkVsZAg
DXX9zH8fhb4/US5iAqrfjANp/2n8uwPhtigulOthm6+Q182TXksqD0+dlZovHUTSmnDUcj5MMR8l
Pm8lsIhakcca71p4VhYX3DG0hfNdKvbQTKn1EyttqU/6871pTvLO/30myzPB1ee39ZxAgLL0rFwP
Byv9KI2gLX1Fljot1UX8w3YD6q06TCmoioPE53hHhO6MnVHb9LbywEMWpDgYva/evDH07aINsU7K
QKRjt19+UsPXriTstFvwOpJqNSGjyTpnFgaNLEgykDvmw0eiGE1hNzLJWG8V6/WyOCb4mkIuezm4
DyJ/nm/Af4hUUgqRjd/+pJNu98zXyXhDrTfms+II7xVWixbHdXZVTcSEQBylcg50sueulgaChbOe
bGiiszIgzw04K9sJeST6IdMkx+0FG8ioy9PwNYdA/mjh0XS7s81J8BtpFxpD7SiIswtm5pMP5zK6
jvCfDxK0Xro48hkP2ccFHlN8BwxwX9X1MADJq4oQYniBSfXwWLecC9xmfe4un77lyTMAzDlIeSys
651l7XNVni2IkMY0DLx5jY0PxJRF1btvzFil5U+rw6UFYapy6phwm+CtxqtrwT8zmWDy8ClqjyWi
JW+ZVg/NQVhk4emaVe6I6TB6bZYMuGXZLl9TJq6mdV0xgfEjnE7hrRDZOScIhcT2qzZ9Bp08CccY
dl1yDn/bLm2ppqM5snDUjjnzzWd0UQcger5oh/0JS7/MH+dC6U3keIkgbPiD5WksB5CczglGV8sY
Iyi0FmAd/jPRL6evEFaTQFxC8gdIQKWlwI4+SOEM9KRxuw4BwggWw9QFcFlVQ9sG0vAJjVIwm8Tw
QMNL+3wUANPRln2Sh74CdT7i6K++NccJ5MWDeeJIUFliMLuvErUq2n7Mz8oisHw4bl7ty8L8eqAG
AtkObDJF9HEmT4ONYhY4drjFGQcowlXry1ugNEfe9ajmpCbRlKQ1FLmpr+C3av48m+9UphaOjMuT
6Eenf3ur/sgWEZ2MWmxOSZ69AJK7ck9Ojhr3soXAUCSK+KmJ2dL4iI5lDmNOxh4OlFxA6ITJi5Pl
xTDd22vrzwcOcvIN3WcUv7jC2TjVNqIgBbcHKyAXQ/EwTmsrnfloZSh1Cr91tRHdlNdwDHq8woKh
6mam7+CBQ2z6fpjiYXdsfrzVnz+pp7zlHaPNQvOEf0JP4MI0RWyyULGe7KHfAA4Zo5SN1m/epG/s
yyyENJ8giDaWGlj+lKUW6AgAOlkyqqic70fmXAKQdvVB825NfxzCmSE9462KANXa7U4oEwOTV/en
B4CudhWgXD2VYJfRw6WAmumQpkI7iujhbyFP3A30P8gNwY9rKvrT/uK/o8meKA59GvVQSfGUB9ES
5Yb+QOFGEGIyyplc8KFa3xy4wJO6ECVBGrnsq/81VobvMrwryo7d7vlHqDjyJMtr3tRB9fuXLh2M
CbP6RmubL5kYkP0Aj+d3Ntcpapj2GwrOt4JRiFiPJ/2zqgeuB3irqiiuPbvtOPasFVzMRZ7FW8dC
rZeqcq/rQg1/LaL7wRpVnZ1HpfGB/hvYHPLXeKQX+Ggx4afMW+ubs1FzhegDMmDnl6jwouKKOMRH
1goi+sj2QJ19b0L6CCZOyymqx/eeIXJxqS/jDY7jujjHomOYZeryCk+kLdsnd2iNK5xz7S86hpl0
9ombdNnKR2w/6OvxFadBJKmUmh5nEsWDCBTJTeGrj1qUZ19swsLO72gfFW4BnrATf5fpkYbs8APY
aGdKzscuL3dQhTkXDoJZXPfqfgdmL4DGOrGbyB+02tp1Cc9QVTdXHeL7tXblmHBgwIVppW/W4mQ9
eGEKW36qit/BD+gym9X4e+CRt0dgo5E1SzGAEWJb6fAb2N0Qc6q4+AVXsrZNEjaujhnmy9sVO3sK
5sTis9YgFSPcTdJjgdObk6m8JsF+E0iRsS6aJ7BnyQMsTqebfw0chqFbE81AGVA6T3CXHAGtElwF
iP6XycR45wUSt49pqU906r7Mb2NfYMVWpZTX7kJYc/RZPfKn8fZli1C8K/fNz+06MWfYyfkEsyDm
bGV6IarrQ+ipkmh0ExwhfAiiL4121UkWRx6AbNPKZCBoc2SohtBUjFsr8Ihy/7WbW4PhVbaqlvX3
VVjoZ5x+3DVO0BMfYY0Sd31bfRCiZKpgf6ThUTwvjwB9khvFOiQ+TsSeVej6eYrIlAAu470sPbmA
ceq44fOowrn5b/T4e5MRFhfsbBlrigOtTxlFJKfIzGWt3ScSgG4jBxJELIKbckU6gx6B/jV0IW8e
nRkVJkV5PXapwiAkJauXzH5NPjZYnXC+Tj4Of1wkJopYAbKOJUrZRaKCvP+btK8auc2yiuBkWw8U
ThFe0HfR6emzV8KlqO2DGI0Hk/kjOfIrBvcwdyE9pHP0R+Br8e8Eh3YyXLrEXIvdj9EDoAqWWwec
VaqhEQCght6ZjeTO4K1P7rvYMRbGow0KU/wxufKARYHMv2fgzVAj1c8GJcgMImitEGa6oV+2N9Mo
/hLA1Tk7L+9vJeL+8mZrwbOfouJzx0NKH54SkWCxN4xfZI0tylDbx6VwhJsJWM9D5TbJaq6vwmku
Yg7k9HvUwRq+GxKt+VU4qb7obegs1Ivx+JuT3a3s6i6/fVUXFie+7ocqPSxPFgmZqHt+8utw+xeN
nzqqWhCK05hNB9GZinorRyOytkvx248imeeUqjY9T80m7BBMCMYhdb6DC1r3c2+cqSpFTM09v9HT
1Thfg4m+99i13drzSK3xcXpQ4KLj3JBNnmYIpDIBoVywi6v9ZRAx2Yyeql9IIZtWirJLDt6G3kuh
JGzWT1D6dSpYTzeZC7rhEfCyaeyEb8GmNcbmwd2LVLxAZa9kiCu7UvLOebjjnYO0c1cZ6oySKHH4
mnDQrLkkroF/sXyHDKOWz76lcycTYHO8vrc6Ed1xHT4NbDGG/OvlTLf61p6+TO5vhG9xOqO87iv1
fimRUNRGt1gQDYe5/0i5/SmxCF+py2AkvOtgjDv65w87jVgxaXP3/LbJrXPFs84QvLTUBdY3brsE
V7uadhyDdew+ygNdTTVccK4wJxUpMLpO88Uo+332M6BpaIlcQEwaIzldusMn1Z6pjhmqBHhuQjCY
PQI+Hrl0PBPV+Hln41QCUUIK0XONWKhTYndUg0XpPmYXsRKCvRPjirxEKxFJEF6FCqvT1/PSceL2
JaSIaQd4meSZvbWG226Adh6WRvZJV9UAYLs69+3XwPVxen9ZyPJPHY4o/0XPRgMOnZTmIJ3zu3dR
k8sSPitQsId6+XThh5ES13U615qbWFdWwYWlwCOIn7RuK9mEn6yLkkProfqf0UaFh+tuFIlo9DUw
MYoidI7/PIPPI4NgBCUiOf6DqeXEdfmMDqu29exkHXR5UvET3CK2TFcq349Zex3WCd28SDo2/Wxc
51gjduNwhhH2m+GRGaSNp7NXk9KyGHrDpcX/P7fSYmaO8gzHlENpz6gb+BnVDn18/GlmuQCInY+Y
t8nuNwBAt358MF1/0VjhfyEzlkjzZ7AaPq34VywFU/g92bkKPvUxsyLWNyGmz3JepDPYMuQIYdcf
vsOIWzBLE2A63RpDECEYDnNkwJ4EclWqXB7f8IAtfj5K29dP1gobVfHcTAbIADLCUFdMR2z5L9WD
hw1u5gXvzZKvWf/ug6B987UjQSkw7BakXM4yGtCk2IN2XxfbF99ANurFUh4xAUhdkB/K42XaN6xi
APud+ulirQBszPvTvuNSGrWyxoerNC4Bqao3NduqQtotbukM+xyNQyx2CvKphlYXaA+EqTDaFCS/
inXTBfs7bvTRKZ8aoJ0Ny8rTwrtMOzryzSjf3+NQw8Uz0neR5h2sifx8TP6z3e7YeA2pCl4hwE+Y
ymM0AFKoC8wpZEFQGuCQchZGTRy6T0YiT7NnrslBxyZyxyqE13gLf3dlPORDmJCwyJl3M6Z7wptY
H3d8TFHzFMkuxoPAN7oj6Y6dBdlqiKyxrB4zKdvyqoevitxbNP7LQ5gp4lBon4E2uV0wqzI3WUlw
znV8XsvNFTn35dsWjGJgjSyw2DeS9olQfrCsBkr4oK6gAmz6SskzdLUpjY0whQw2qdbvhcAUlKAp
dDWNaCi0uAUDsYGyWQWVzXK1qZ3qNJXhrQmL0QKC7sL2jjIPayXmkpyAAebNYolniO1lbc3V2V+d
U4yIr+55O/TwqNV/i2QlnxksJbETD4yuMjIfyRQQururPy4AMvlkfC1mBfk/UAQfLohpZrSUY15e
8iibTaaWAwuu3iQqSGMld5nuQFA+JnUleXn1mepMK7rqWIJ2sAN+Stwb74nGJcAu3aQBQ0RmF+Yj
gDRyeGEsHMmt+JF+uL+WJOvFgTFRHcEB1EFT+7Y/upUUhbTkyQYjOCk6mWiX/QiiV+ei6ZJJZaiS
b2k9FEEZuHf/rzBirHwoPPcD/DCcCXDq2j0Lf8jCmhWfveNn7MobybSoYjLZaW0tHKz4Lo98ZoZS
JDXMDN3lB6WsRfEMKO9uluDYRF2pMzXGa44nAH6MfGS8i5OCawRlYW1SxldgrGoFJf0bzYHcVrRb
mtnfh2SjKNbLO5gAUYlwBy0tVre0DsE6sbfC2BbYRWFBunv5VWpxENEo4upG4bsqxxgbCW7laPlc
kllq8A+tz7IEMZsP0STCLg8O7caG8ES6MZxIEFZotP7HS+C/N6Ha3N4OGsBXNRsGKd4kRX3flOTZ
oiE4Tbjh3hEBfmRIaOMEbgn4ZjrgC/fxtw9YnYLijo+sJJzB+0Th5mcLcfgX83G9sykiicQvt0ur
sTYfocOp/75D/67GwZcfAOhE791GvFVy64616VTmce1NT2vuymTanxAhbyKwmWYk5UjFAmUKrivA
/bd4pCePdXjaJnzVh8SCrVxi5NUdvX5ROOounkchGXTHpm99HxZVmTni1ZELerUuUGNXW3zaRQYf
vzQCdutH2ERT7jcs1uTUwFzGcrkTm62toUFZJzNKaeC3zhUdHa1BDnHy3rjNmwueuqg0RN8/kSuX
flzRr2Uqrkud4HQIqsWWQUoRGOCdD+dvsS5KCN3oA2/XpqMJ9xLkmu1eHQTedQfslgKY5/OMN1or
gVpw5ajYkt/ePid9R0yYPmaSLBGsrwFeIC72cJsqSXzF8bTBc4/ptf3nes+rrnvepFK5Prz0kI5V
ts2vZEiM7Cyop30ZCp+GpOgDYtmddy2XiQ1/Ps9Iz5SSAl/eOPMbUHL5Dh9E0qNbLyvjYLV4FliE
mpDQSMj4tRn7HM6muXSaqVCx6njUTfr6hWYftWa6wQyDPfFIpot7QOlSAVb3F4+yhxeUo0HIGvbo
jT/9bqDY3yQxA2Q5cvs40K/zYMxZpK0MUK58giVIjezi7uG5Ix+hRDayXNlR4Gqa7k4GQlWnVEu+
Q+GvZk35iYJULAE+54Uc+eyQ/HKvH+5cHSA2bOiSMtOJ4Pb6tfmLxgcDDrK6gNGgKdlMpEbIWZlY
0MciC83BuUW9OzqLYIVMIZj161XmTGsXGZhpHlvx8oao0l5Y0WdD3lgr8t6KPQlbpg10ByEBKvpZ
WqiU5dk73wFhjc2s5dsFrVoBJG4/lZx0O92VDdehhit1Ijy8oo41FnzRniGVGXRu8HxaSW3o1h4+
uSGPagdmPP4fgH8dPkD8mTlVVUhCzXNeigPH14JiFzb9YrVmFbiEADhtfw6/buOCBA9n507HD4/C
ww4wlXnLmrTrUwA5hnbM6vwnrfdKF5S/iuKSjX2Kz7ABLnTlnJ76W6jEH6kw92gr+H3TfGWvBdzE
yc8/3Y0ck+pq2rq+Px5XS896WvSch9BlUU5voGMeVvOnWzpcimhFpCkcwOzrL1tcDcibMG3pd+Si
NLHC6MmqY2uTjAhjP1o3HUQzpCupKpsSQGpYhM8T3w9wSE3FCnWu/HQPMnjFfpdlFblaGv7vFwKc
i/321MFf2RDWAcKaj3qJIDtqhv1Iw999n4DL6sVVgunvezn56Y4PzLdDl45oMIKATb9cXqG/XE/1
0PsOOj6EhqnNB8Tf/XLtmKRNZ0fkh1X6QPDqGWefUS08mDlFhpP+PWd9hniliA4ERgsCppeLJZHL
ZmRiKaDpb9zJn9x4TZ1pDUtqIrkJ7sdjXokQEwnWMpIRvurSg7+2+scKm/OWvXtfR9JRHm0gSSdo
zqGb6WUioIWbRnUdQudgA6syRiijDxFBZtmji+3wObf1LWxCYWS7qMGmnCpZpu+Z1B65EULB0QrO
Kny0bVZljvjvpdgAHlEHB9MtJkFYTneMQc+L/EP7PoEmkwEaGb4LKNW9E1GyU2xH9S0uBZ3M4viT
JzkiOB3drH3D3BprfxH0OIGVpHN/Dvr2P/mqSA5telL3OePlZQ/p9cb5ggJZFaJP4TXkX0jMnQwQ
XBBGRqyWGndPMz+fZf0IpC/Su4hzjG4yBZe/fPwENZ7VkbE02H5t3NGhmbPbBFPeJtW4zBedv8DI
Vn3wbsTnhD+eK96HKvL0MOZ32iBft/QiiM4oaX2wR7WUTTm3RTIkhyroWis/KzqcQEHot78Wpw+K
nCGhTC7mFc6izt/xmm0SjyyIjEB/IrK1glRIpje8N8q/IcBmvzsz46rV4JDGSJTkx/23nPg75Z+1
H1GThv3bAw7cvYnM4ryu+gUrSAJpWCXgXKIFjuPpbmHec0cW8ROUk0ia6sUbX35AkD4HrEh6aR+Y
b4184Y8LQYuMLzL2WXNBLQeElNVKfN4ncp6ya8NLJWk8lByjt77A416rUsYZ2I8lRNG887pisNrS
IJoqNIKJUtacDq1eTwhSaf3QRTzksKYcAiGLEnsgHYlBQmDhpJYSYC/qIqRuW6snKI8DHIG60HHS
z2CBcpnseTkNO5/+CRRVnVVuAgOdKGK3+FQwAh7xMcpWPKPgOWh2z1BrS6jOONbxJ94mk3mEE11e
Oc+yPgtsa6BFBTBJUVzoK9vTMIF/tJ2G83n2R3nbdQT211EBWXODSMh9ycYOxhXeDMXbrT5XgWN5
SIYEQGUDFIkp2ue9phkVl4lmnEKYGyOW6sxG7oMLFtHjTIR3LXQh+WqZkmMdtiStioX3IiOiwQpL
zON00P+3qGzZCHqdFzjB6bkGsT58dzRO4Aw2rbiUoXxNX4sSNX2ZR14NdHLHJyMZBqeY0xOujjY6
KS5YNNgyjD44lc639jrzqMdjzZwcorXCFUBUYNFsaY0V06Pruc9J6eyJZRZRGH4Y5ooectKF2NxM
2UMczWZazIKjJpC4v10XDhRZsHR1isbkH9PA3WXYQp8ps73gaRZCSAHkjEqwCgPXzpP8X9MdevwT
L4s3pdB1kQa40UHlJW0gm1gmNnwamGEvRRl8gJflMf+xr555t3hZqn52cktlGlJtV74dSFktp4b+
QMebczuv5VUiogz6U0pP2OcVIlNzIltRSd9rD+O/k2ix2HTUnPK+8zKIgNSv1O+KHmd4lvcu9+6k
piXl+oyRP9ogK6msZvIvjMoTPfrIgS0C4hVbtAZeg0aQ1+GvYIRcWNHn8qqStpzvFBU9IQiMn3Ne
XrJLvK2/ycZWUMtLKAm7NhqxmGe8Xx3x646mlbMgMsZ/DL5Qw/CzHYqNPsJROne/K1DEswQ3lVY/
Mx6rWaWRU49ciTWSeb586PEiyuybpYICEPmo+sRZZ9rgwDku8gsGomD5B+t/t4ZvqJTiEN5a+gRe
p9OZH3eeW4uyLlc209eGRL0kPmnj3a77fwtB6gQ5FlphwpDKQUxrg4AvZedaVL+OOGdEmv3/5NcZ
Yc1RJ0JZVzMFUqRycKk+mxE413PPl4AFpGIZa6RDvxxl/+quXoHGPiTb8v6xjDYczXwfVf+jBCJc
ZDEmcV8FeH9j9zHg9Z4vliqjekiOmIb5+EINN6oADw3UlYUBThyFGNwaL1kF92O2RRv+mRMDbeHi
/6Yif1bxpioyroUzIpLOBUFPED3roJPmVH3OhhJr82sGtNI2wVDzT2NACakMToo2FZuNvBRf1S8e
w/gIHdLNNbout+RLZSVbbUGp9xNnYuRIH7jzOhHA/tKKlkxy5ipXPp3+MMViNOb68VLFsHXBm6OX
jtI8muVnjiPP2TgSA4i0RvkgG70g1HqeeXsOPQWRAaLjSCXCS53F76uUzzEMGOc4SSSf6klTpmzN
IVVR9cn2gSVLzsCCyDAcX391mv6owvHhwFgtW7+2bVzp7Qw/iBKvzO3hBe0m5F+oPjl7Ux+NR5rO
/VSMzcyxD/GH5bjhDJJFSoSNGicAM/UpgO7/rInjqM3kPm/uCpfrdfHgUIR/Eq2GiWst/az32ZU+
2ACu248Rd1P+dlcdUVD4ojQLyGqP1SioCqnVOlRAWuvGRzkr03mXvjgbryMkbmaTymGJuzQ5T+kY
04mnqGvz9JcNK82OPMt/pT6U/pSHHU2wPJ0gWl2pdNqFpCAs0biRRt4iLECuyW2Blrcx/8bXlIES
5HC9S7zYR+t6I26/kM2Npk0NGOfsO2Vq/Q+lmNSFjakEOfjKwvxJ5zFtHkBMuB8V5ehs1OLrGCWC
wvPR6JoU3zX8HWuv4V2HPJhdkVRt3Keh4WuJgESqqMwF/ZGkmneOvGm6WIPIFZDYalQctB0Sxjwz
fN9pNzmyADzjIKTqY7/Qww4zVI9iwWBzH12uNQZH6YzWVkeDKaqnn+25RHdIiyDpZhdddZkS9A6H
5e/Z7d2aJaFECWg/1FM4ezwDmFp8a/yurNkrM9tsgkwkoHOSjtTLi28zb0F6s/3pTPwDpNeKMKHA
wCoNewdNaalaRAsMGGxOnXTPtU1Zi4ggRtm3fXTH5j5ovXGOQZT/ze72eLIuuyTJExLbHl0GDW3o
7Qp1VVSSqgdaTAnV0rxc3BK9LCIbj/9E2CtckBMvGZAz0Ona1GKiAx/mfUTZmzVmFY6WqX7cBnTc
8f/SizD912ywTv8nfXj449mIlG5rGGd+0LPVo7ptoCrIa5eUJXyNN2PTmOPuGxkPX51gHZuMeDBm
ADQeU8zIAV76Mt4tACDDIZC+NjY5BrULMPg2xMaweW0qCStShDKZOv84BZXOqXqnOuWG0gpl8MNo
BqunVy+U5dnYvDDXyrobYDxEH/WQ+7qGjC7ocm+pRqhp5L8gTzzAAsVMDb3roARVbVbPqVuyQ7Rh
dw26E7krqPxTTl19EssM6331f5d8UgtoAMpo3Pose8j90kRdM0k3GDtE6ZrVZIgg4sf0/pbSNleI
z1LUcB0iXBCFLOtWdkd3aqok6FMi+by+nwEDSM8OOEvJKpMVvb1nwjxptZ1EPzzGcohIIOATRYul
PXIxd3JImp+hg3E5v6FUdlNh2aJrFlH+ov2BFwfaEbw4wBp+MP8/R3sPKJJKJulWooWyaEL9D3O0
MOLtfzVrcGN2rkfauFnPokfz6U+XiakQ3j00BoNmq/zBtOFAc1qsTndHdUsjpPvfC8IfXAbz5zcV
YYbFXCptzSjS8srTMS0MdiN3yaZZkMhclIBkfNGLMjAwwPPoRk36/CYTM6gqYk0dKU4r9dgMC2R6
1qqNAZJ2C4DqhyzPeGk5ji+xiXN/rAXXB2Pykd8nvCcmqq8bI7jzc+iztsfWIXrcH+hBKV7N1zY0
krylzZ995K++7XsKEfuj5Emr9lO1aNOIe6jBfHcO0NI1M03NyMy85eYQg5qiQt5+/afj7CWKBcdQ
eIHTVgEK+8M6IxsF5JJ6m10x8cUBHZQGpSj6+RS4K4Jrtmx7zk4FCe2aoeAAndI7iMAivCc3fIJT
qeCPXJMoNr7WbiQyvHg2u8B8zFXOggliKuhkwZ2V9cTOWYu0j3JNWv0ZROT6z2m56K00Yo69uuIZ
4tp7+Suata9/TxkAuRWBeeByeT/4KZ9FCK7TnDtvirEZp3hC7/Uv1bUAzZh079c+6YQvaQo2gCnU
6zh9nBHQvLzaPT6T6cS8M0mST6A7nXjZjQ10boIqsn0AkJ573gLeIUsQxnoUtZC8p7OLSs/apSbZ
4L8oTL5h4NGn6epkkS3+4SokDEv91sGUpRKLcFLTVTMI5J8ILZA4YqqsDAyt+cdjak8ZIn9f5pHu
esJpNESzWMdxHHyTFVRI68RBVo5d49mWyly6xcRNkamgHPNGp41uWZoSu7PzEsWdmiaVxn3cxHH+
wWl7DyO2jC4PGcO8MxYL+9w6uO79JzGnfDwxejiHawdBGU5GCDJere2xMk3+2QX3Bl+LKzexUdrV
5mN2WaIIh6c8gawr4ldSAlSoiW7c3glOAuVHwYkD1ZKQeGSeiEti0hGfRHaqpDBbJqsSMhoWsjQO
TtVQ2vv2TecMv60oxohTGIj1lVysVWmYnisyy4gK9MrED5Pm48p6AoEFwLDd3zx9hHHTIk1MfkUQ
lwtoA0sId2dEMpEMABjr64Y9LggCB1tyDE80fMGI1ODZdAWYCPTkbRCiGX3nr3VF7wBq/RZfOigI
EQGIu4pT6s2csFUNgL5ZkAdagDyAVsy/Sp4L3MRzja1Odn5XRhisEY1ACWevVuxkexF7chFVKFXH
RLeCGEJ305BMF56mgePGu5qQq9HoADmtPGlBiYhrDzEnEgOLcT5N/M93pN8+lR9cqU5ZwyIRW1qx
ec4rRuhVW8VmHCnM/+ODNwnQcM0zYNW6RWGf5C+zo1krpNrgScDi7b1x5zW0jQEZ7tQIJdyYAcsA
tU0eTQR8zOn5ayGF4p28ruVADHWLkhPtpbr3Q5iyBaWHLgFkqLkU2hNsuWARHEeyiOoOIO2h/ODQ
bxq9oAOX7Wc2K5Y1DON6Y/ah8od2BMSRNl2KkLZ89KQK0nwKN/iCzHzXWVXf4p6wo+RD/z2IxjVp
z77XdLSqZP9BOw1nqDaBusybNoyATS9XOmON7ZipsnLlW19pr6AvfaLO4moIjE5YGK49N9pmL8Xb
4rO0kUrYFoaIWvQHfMV1+2XeRohl/flkcTJHXyLuOKx16QyBgYWSILOOxUvB344ZKvajip7aBj7C
OsZWFwFzYHprmhKjKfls6soYDGspHvIxC5dWvERZ/bPmXWywR1wDfaJYMZrdHaP3LdC/iTuTA1HF
oiKvoF5BVt75Bwx3AQjQQzedE9MfCQPV0xebVbzLO7pNrcr3+0/51Hbd+P8QeWOnaYap14SITVAC
uNqf0x3QNymac2e7tjqJtcwe1MrLgVOVcbUayuVMQhiyk9nHwHFcOp+BHF6THHUFpJWiuWy7JEg4
wD1BHdSISfLwULijAMKYtmNt0Cmr6mqshiq5UVuhnUa4VOGCyov0IeLnrta2znETeFz6/Pu+UC3e
u7CGbIfY+5cQb48VaSZ1RePgwFImHEwmKzmJyKuvcWsm3eIYRK7XvQIX4gt4yVKqX8493ekmUjfY
XoCptbJOyW9sVOFeET6XW5wNeDIhvpfyZ+9zYPHKmyTm08vE0tmUwd3JJmCPp5WU4XGEoyXPCgrn
FmzMfB3QZirI2e08KdaCgAkrkwK8hx/I1e5dAnzpOOI1DlZGdYhj2EWPLJt7yldUN0ZAZ/JwxgKO
tzQ7bE1LaD/+bLFT4Hb40VEklcc21mLTjK+r+0zj/yAWwpaT/fhLR50B3FrbZLje0Tjw54dFjsJ6
mvQIoMxjnOmXwelGnY9myC/2vLMet/OmzOQB0uLlPrePrOUGnwPt8IL2wqbDFX2vkfh/T9mqHlF2
f3BFzg7Lev7RwkOzMqjBdK0KimQEDpyQGzUn7KHkvu9ALTaFxmA+G4N08GmKtJiRk5SHlJ2SKWPE
JusFn79UtiYTq5NHnX4elrrG/9j7rEDYKUhKWFnWwg3wH9iCfgOL9o7xm9GZTUAcJYIw8Kj4/O/b
V1WOaMThBYICMU++o4CxYvr+bm1GxDJrvx8e8MMxsRMZH22v9hVKssQXAbs448rVup0pcDQT/hB7
1VOwjvrgYV02YSg9kERy+noTF68Pgd95+m6HHRurasKQHVwg5eOkMwV+YnYBfQeAle9F2bUfrkwM
ecFpU3MkK59pZHBwSEs8CAAltR7h6OTFI28ieJMFPorNVRc+y962Fi50ranCrBViU+qa+N6S7kTZ
ZOBf7h28XREwTmsnIMYlY7XY+Crc6oy5UnBMI8ZJ86ml5TZJM8pBK287HoLUw5V/BeyGprDGTYio
VjIvsb3iVSeRcRiEqexkU8d+6PZVFvNX6aSng5bQtATdYtkU60oVRDLgp/Sqs8GWmf4lRMFDg6pc
hv72xRHQKAKZ2F7//FpAejYC9ilfB09U+YtexddeJYNGEU3p5fHoThhTwwSPugHGkfab79A1qLPh
GLikuejBYEpsidBBuYudibmbD7F1jb6D9aAQzrQSPiZa0vA+J/IIqvRloChEjnWVm1KPOmnAeVqm
cpEDlwlknS8oD4S5jOUFD9DRV4R/5U5w/cGpKrs4RhF/QkZs4aapL+AqKmYoJMepVmd/LaGPPgBN
NFWT87gdvIkO2fIZU+9U8bQjtDeoUVEEGyJ2HrVbeTgI0ARwdfpYH9WvQXG+WZ1S7nOsezbrEAHW
7aOTmWJ52gQ88GGWkU2jOqyDNyXvrX8D2WISWZKEHFI4LQslxtV14DvhE8HtnNxXf2bFAX6sXFJO
323lSn9oVne+z2hcwO+5Dq7iu3yhTE63Quoz++uReHxeGH0dvMo0Lww+0cqd5RZItFphvbtF5ud1
JV0XFVpGjb0+ji0r9HxAYqfr55ScY68MzLhzQFuLHpp8zHe7tks7uEu5Bd0gwGKSKUd4n6d2c5Xv
ub6YUEjU/L+n1RcVZXev1ADMTXOuPShsWQyLGOGEp8Z2xDechBl0uJ67nYdNkH14VdYeCEY48MCJ
fViDOtFhpFkYpX7JKze3DJ8nYkp7fdmSmxvr7MPTXGJ32+kL7rL1NxXGxZIy9EtBu0U8wv5Nvhwb
eYNo0Q3FQUQuCHSl0vIZ+ZdxTy6Kdis1mcJ7dLczoNOH/1YrOBfVtrLdjT5HRkNIpyg6odJ7cQK1
NUwcYt8D6Hq27uv3hm3T1NTTtY8uAwdzT63QxcbmGlq8bsPbwEVo54W2r5B7hMwXds/aLHxEXbBq
wWD6fDa1REnd+rdmcgjikgtJagGb5rUVZzCJIYJ9ffYBGxCvJJdUQDUNCKpIcvai5HTnkbzcohs0
18evxfFUVm29tT85zbvOlGd809DhmXxR0DgRQMSndIIcIQF++Ymd7vmzAwYRUSOdB+ylCurgYbo5
sJcfo0P8uOu5G/1DFjdWexz2ly+29fxrd6fWEJSr5rwrjghCq+LQIXNZ56fhihtEn6blNL7ZeuNj
kcL0CxFEk5NZKb2sbE3oF9tscQKvZcasfCh8PUQeGnJVVOlUOvJgRa06Pfydh6X9iTqHh4wN4whJ
HIDZ3ZaGkQln5GcEK4WeEgIZpkO93SKcApbSA43+uO5LWTMQNN3B2Uv+3Km0fivWvZyFgkwwwAti
nGiv6glUV735WaHy8MTme3lc8pLbH0IO85GoMNA6Ib2M5gjB0RZZdkWi7Pu4xw3pD/h73ZVpHEGa
XuohWNpO+lsRsnjH9BlWr7u2rVoqg7YR9+Gd35gXy3kcYPeybDrI+PC0sYcGLYL2qC7EBT6r/cWj
83ZA7eIlDBNEeQmkAQeqmKRq8QR7Ce8VodYRcIoTzvmFtpp3En8Rtk6B6GEwE1YL4yaojW0je56E
0fN5QT8h6wMtUaDG+Lj1NhQZBLq5WG252kYBFvyOnbmSOn67LjzivAfr1WD0mC8e2f2L1eHTxCxl
XOX2yTqmW8Qm05b7Anu7VtWe2FrYQLxggI+7X5AqfrNDuUcW2wDA4bJE0khzj+rmJYX8/piJry88
HFH/mGTB6562XmVT9jh/vsGbUcmtBqWBMGaezUxeV06ZtCrDgW6HwFheCrxbvS6hegk8ZPShW+8B
5pd06pS5ACN1kTqIRS0k6hvOSjvDnOQCC+ABXw27ixu1BUaIW4eloCnfLk2ZjXjA1nWs4X17Fr/q
mM0MD+qEJNWzrMsMPNNZs3OnT3DsopfiHYXq6RujE4zLGEbQMhuVUsqzVaouRCv1+FzqucZ7BZJ+
vfQ5EDV0j/oO4QrJlC91dn1Z926JiwpJaXgqTnLi+lpfr9+QLjdvBMrkdmLcqR20CRPF9TgwWODF
rXlwi2vYAVZVdB9mjUMfbcnv4zukW/nuhTE1ASRaCxmNB90ETE4AFaEdO0FFx+XS2jq+xdMKRbx1
Ss2GtmOsxRXq34YkyLJNsZhanIfaJuFKAuRT5bUCWeGlhc3luqdkRq5Yezbg3LaPt5PsAMLKNubD
don6QUkpWfoE7mrZeGBkhyGZ5/03OcNHoAdrbzanwIgZmWsyqcli1hWOb67DLS4f6y/IIXJ8IU/q
FTGUQgF6WkYL7+aTBBSOGhlgigt2WK518BnHlKNJUDj5f8JUD+70Urj2cR5hv1CAhZ9KN0OsCkw0
H+ZE3Pc3DPXj2mPWwjc++V4I3HLPNxORg5Dd3Dr2aNL/8P5ibQIeTh15vgGn83P+/8KatUb9TZTY
fZtmxki1Xhu2AhQWGgExLxa8UvrxxwaJrXti5mVOLzVhSvZEMbk+PC2on200QBmNy+lj3/Jh1oZg
vJHMZEGGU8nT4/2QNPkkDrNVZPWF/Sg77wf+Asnp5DN3jBfZw+jWiXLp720s5BpIByMBGs+BD4eI
YFJOlSpZk4rqw+C/QRV9dZSF119PA64kWWNXiGEaldgWg2/6K7xmKo5WBOGFhOBBOtdRZvGJh0qc
JInKE9Vg8Ynu5/BonKs7LiIORvGqlgxzTWLCnuyFkVpoPb9KAZocIMAY7+OpvqMWLNogsLqr8HmR
xHYHzvNfu/xrEIlbgRKJM4qRpskNUdLoZF0f3M9aQ9gknUb3YARnZPm2i8scFsAP4awLkF5T8xiE
HMNiEotI7CqnmSRIBLVCIKpdV3oCsa8jG75VPPXzWEjaED/bfPUZ5oCSNNDeFlDYfBLD/S2UQaEF
z+ImDQINM3JVFyqwjTFLEZTFJuCpoztrd15yOW/NAyZjSpNbSiiY06WTdCseG8FgE9EMuXYJ2NC3
05jkh/SGu0ZHL+b352ZDFbyt5pw2oAz0TzaNSm3if78e2O2j77wEg0r8vNlUhXgRldgmItnvfJ3K
01GsPoNq26zjUcqhYfHpPCcjJj+09E2fPips9NotVkMv0T5Bi9MNDLYTg2JMtQ3oZNxjkIuDCZhS
kdTP75RjsGxfKnptIxz0iX0tPG2A+eeLYDqQw8GliHs2oFNnNdlobIfwYqYO03yAvJzz9FTDUN5+
BhKmkdIPQL5NYK7IIZAqy65BPnREjIbIM5AWbNV58D+LtQidpvcSyn1eGT0ENPLV680/5PNLcMcD
W3cBstCDX/TTlc1dcAMvead6XXlS1SuelPYVnNhPl8WhLoX/h8i5PnxC/bmJCeqo6/fpZb77bgNW
IHNvlvu+lFIfocy785kS5Y5oBkn2ZtTQ0Rbl8M7BTkC0N+t6axZzs0VHBm22WrYJtWW/12QAHuiK
5UIiqpjTQcVoBKlAab6GAjePpDnDj9MbmaEZpuWbNUu6PJ5FgvS+8X3leNRX6x/Pp1HHK8lksjeQ
dlme6e2EYsAAQ1gGUuxh8o2kd274CrMBWOIBnbZyINfal896SPK0naUdmI2sHPlv/jzbkmVI24RK
A3C9WmEoGO1V04LzwkGHdu3VBnmMFkFoRGdFqXN2ZKaqkl7q7jNZ5JjkdHP6U1R8YAoduE/r6fLW
HI3eXYxL5x3A2r0pTZpYzcTWeYY0BlmXwVu4i+BIpCDKNEVfKdWxI8sMZRR6T7+Jeyu2hHKjuhRs
vsgdn/JTqo00w9dJQbCiBh7EHuqt7G5GwzPqpT4TgPag0Wr6D2OGgDKlOBfRhxXUlvNV6EdEjPfJ
zGY0kbHOgYYGX7dUBvB2Sc82l6TK1aBRao7uOKIuW6BxyVC32ms7O8dg+d9SDJK3VJLomOBt+BXm
gBYkJOt9F8ASIrWNh0suhcFA5PEZSA3FqiKw2BF4EAhGkhaCaFc/CY2fZDHwzHOSytIZpGhZko3h
jQhS0cLfV4hS8kxb6xuIMo0irp1OXQ6Nz0OfcWszDxgkuYvHfGM4rEX0jmFcl2BOcrdtMAn0EQlh
IrmV7Si0PlvucakCVKuKAtdjTFFkIYBobL2RByK/RXaUyiD4OSNQjuELHItoS2xHV4ZpsFrUbhtq
88eqx9WPPXRi2u/I0k9yYvLwRiDQqfUK6ebWz/0ihWa4mLjC1x+OGfwBIlWvEcWiP/qMU8lTUI4P
p0/6tguJa3sM779mr1D+hH3sJaRb0Dn/d/gBx5cT2cheIiojap1kJZseYI/cQWJh3+8PI+dH3Ve6
7VzR6Pqc/XzyhYxxUzJmz2zs+J/4Nghjyqy3WQRbtWcXVjkmYNFjwX1S0TAvmY3Qp2xypYd9sx75
MRPQ0VvZbYtV3Ns/Xxs0MBMcIbJWABSBnkM11FJubxXcG7XyHlQOszqI7lYtVevjXEZXdHvHu/pe
rIByVxK6XTHWVqIeJWLA4NlYwPceFd0AeOSGKm2JR7BminR+uvrL2jrAPIhzyP6Jr4rx4ReKV9Fo
kOP3SUD5wviXp1dzZRXfAGFyfy54JX6almE4n6CCmUKacID1O6n7XqgFwizvbtqVCRu2V9AjC4tV
v1ukNrj8S8H4FVjUZN6kdqkCRO7FV2F9vZhx421VtpaVdJowYyZl9KlFXe1CKZNKYbiUiwJmXhMm
+9uAJ8BqBL3H9EedC1Gf5SdUNA6m93VIr6glsumsRPSkLDX1PjvLVWnJarlLvyL3di3UilnPUoql
s2l2kRPr0y1f7tTK/FpkhZ3nYxspHth54gpOrn4MVRvwpLHTbBjs44vN6bXdghxE8F1qxRIa7wZn
eZlHh5hT9KAlYgDmB0P1PiTSCUVlYiwRtm4goRjt3s8BVGap+/XCjLcReAiWaJggzZoc8a0sr6Hh
s3o1MTa66zDBY9OPiTffJpNeQPU0l/ZAFe1rRxydo4jl8cXOnXd5FuYPjQKaipy9oY4eWmoqMr0h
n7DNt1dK5bUHyq3wPvM1sw3k32v1K9Tj1ySlkJXUPYiBvDfDfwheOK8j4J37++vyAinAanBfOd8U
6159b5zr1Lx/Vf0pLYMJcb8CklI3zOKR5rJ1hbq0d1Z1VXjQY8ZiY/wBX3by4o0PEYvaFrOTK9n/
nTYil69GXkgp3CbjNouDZ+hCUGandl3dzeegpSAOj+Dxm+dRy+gJZsFb7TBWXbZ3Q7iOf7eevrih
p8q9fBoEyMM0ZSqGFxH4y+4Q1BQlTkeK/UgAMXN1YXqeZ2AcO4CRAegU0yA1w8dq3t8zj5QZZH3b
43dWDJ3hcj/qs3MmAP8VrUMKPamlyF2xX2Gjbp8rdlAsSf1EOtb+Gwp6Qla5tp0fHd/0ag1JKyub
Soxu/oSaqrbgnAhzmRPD13I7afEdMhQv4n6E4yxpPWnlwugxoYDmRWgcZhc+nYhP8lxSicOJP6QU
UsCP8wXMqHXzKTQvuotHScU/ceY3Ct0izDYH4fclpAXv1y0JAtbKWUTMd9PQLctD/171iRXx3V/i
kwsyHRo/R07841BOqs7YWyH6xGKxH2Vr59xtEvW9tKNRO3QFWVO6bW9VsMDVAOkKAPr8QJbz9D9t
EInVA50U1puQninmi8bkhl9wO4OSSP47smK2W410y1taYdDSqDy6QyQQWjQDGsWJsrnGOgofZfvU
bs/Eg4/nmphMERQ9n+6t9+RZ9Y5j+lpA9n4hyaQPy9TLZXcbRjV5OM4yfdS8wzelxvr9iqI1BcUa
dK2/QpDDBi+cZrtnXL4jJ++ABMHyYodhtglQ91Stjy//WZMlGvFpUuBYs1TytDR2y5ZmVeH/0r9/
Bk5juQM+z7sLz+fpI/0ztFxEZXPJGbhxCdaNlPqBatngcBU0AeuV813L7l8ULZpU1bAqrPG1U1LX
Rlvj6lfnJFtB/YvzS9pT02Hi20eASp8dXLIMNEw73hPo9XcA2U4zjw/rrIbB0Jt5SmPjN6PO7rrT
EQiVQi5PwfX2729HYbsothExGyQvj6ovniy05h8o+1G+3x62pQu+ET3HM/QPxPAcJ7ZkQ2moZTAJ
Gqdc40BLThNVGOmpa78N0pFLbgchBf+gj8Pz8Ze9lQ63UMun0sTyf4Cg6ALjnqqQ/vYAmVindg5J
BtcWAzQsrAyTktel6hLXxodvtvNgPFrGH0JY3MmwgFuq5KPffn/4ksKFP/rtYMmV+KUQx2IcZc6J
VdP0VBHbVGeI93AplR+T4Dg8k3qY0jsgL8GFCTRYFHhX+ZiOiLrBdO2BaxFKAA5bmYn68y14P/32
nW0qRvYF1bFx+94aspzRx2MvIEUYhSn1MDLhXKjWQabzIi4iqoGLrmCrfvdajU5MOSIaQ/64mcN8
WONxF+4ITXJXUulG/ILQM/W16IcN1laPB2qaynWVrsIAT3DX8Tl1DK3gNfVAS+pmB1q+SFxgXh9u
MkduwsMraY+ddV4+sPmXSADPj/ptHecTryevB81FG4H7Nzo7BiD2daSRYmLofuqa2ElFxUj74xv2
pUjvA4pY4qxi3CqeZsfbiCXWODmPwzxpWrIx/KOEQKbWFcB2ENdzA1JQiNwfHvGre51LnkDJOtx9
FuRlTS3/3gNIvuN/HFtAJ/cGoT1HfrKnxgLi1jrYpRU1i8d58WUAv+9U2eQZjQe8ZeG8M0ZC6ISH
XqEJoFfzu/MMkvMvB9dYGrHScPp+POIgEgR+Jx8amDqcMam7vpEibxuM8QnTwI4XC29DZfCFyZx8
gdZlpJXOeKTECwMmZ5kI4QRZGkuC6EWZA0yya2/pAnBPsQMEM6FFhCCXRYKpOt7riyj3Gnbsv0my
Lm53JxzUOi5H2Mb32JowpuSc4rS7asJZHbayksrhii8ynXpBhKOnHnNcSTntQwgZfFtZuTtLlUQN
sHc079U0qkebz+K1LJauHMaU+S3KQNIyGN71GB0nsMoSyZz6WVjOwEMziF61klNXCI0JjMMpaS3F
JkztMgfD1SrD7WbZYk948xnmUiZk0w91DXEvT1JtKgR1YJrLn6x4z99hBIyp+QlB+qJIC78f8alA
yjoRhYL5Puka2oHeTrqSNBtpooLALazmcGYIMW/ovA6Wni3riDRiLIxuOpO+o9/QbizJT+GvkcbG
RV6g3+dAMgxcbFE0I+A7GXWKlLi2lh/BwNy/BMBl/mmHav95uwgT6Sl8vLi8jYHA28045K+5Uniu
kQm9LOhmQX1dXmXsAOD0VNgRPA8BKb5Sy09sSciXmX1+uyVMJ3tkMdBYQo1CNchp5umPOW8b/XkE
x+tmtlHM/TBIr78BSw7/8HFTpZ0Ab0EroeDRChkzczRmdkEpZFaVHJRKW3az+rV+akTzpelD2Wn0
4ZipXhZbK2GS4p6bUMfwJced61ZrAtBr25F1P8tci6liLc4SaFlL5Xvt1jIu0Kivo9D6/pGGplup
SNYHcd0ENwjBbMMcEkGPf99I2gxtGo/gtcgVKWKGn3q1/tOISfwFawKFLzbdYfYlxgEt2gUKQHx3
ddbcsbkYnYkToC85g43Ou4njh2JdbmknRv91hjb9BLSvScwSDL9iG8hUDwc6gFmUJNIqInJaZBiJ
jr+9QaOoHa/SlURpcMqrCU5kgMvSPY/mRLPWfWDMKlz/7pGYa9wE2mABUo76Fs4krQMBjk0pasOj
X2NbBSgnzZFttcGBO8uJy5CRwYOhc4r5991bcm/bovl4ZbtTdFlfgtNn+7XmOJYAkWHwwLUNxvTU
B7chRc3V6NlaCmu7ca207cxBzB6WKlvzVpPgC2ZDIsKWV4nKHbykHhMSysV7UZpECmUOdRuLd+o2
5NI7nUktKySSLJbHX+Dz2tLMW106ONadpVWqs8NCNPJ5ZFAqbiGaeeJpdGJNOmirn5Oi7KLrsRf+
LP7hglpKqsygObEA+s1hX/TnSaFGEIKqjx4q65UFEWszwHkCSMZ5CBV5oHA/Qb5sDJ5INtXG0C2L
ehoTEHjI/W4ZbmmP7UWHCRApqai34K8n+hEY3CkTZe3tCwLhN2ERPH/rw3dZwljLFebq7/ZDwyV8
zxwVb1/HWuw3apcv+PB5TivjaA/XPH9wIPIzVKyiKioNXzx0Dd+Tk1q/ursDS21vw3OitcZoRCe2
boAUAAERLrCtOx3ZnhdxWEc8HbqjxSmZbnFlziC36H15XfXBWWiLNIX7spquO1JLMQMlBSEqiFBp
Ni7JnN5bPPA3uMfOCGsyC5Oj8Qelzi3YA+Kt60nE4IAU70bSALcsmVZ8jcevzWEIDVK+91kzXSPo
hJl0eF+ulYKyKGnvOn5agWoN8352029xjM8bXHqFm9b6cBTc3lV0/MoAtuCFoaHNwHRs8tOHnYDG
89VqEd8NeOFmq7TBrR4UEhX1yw9agIWZfdIsesQQ6h62KorNrHP8vSeJe3TUEBR+eM6QP9SMjU1J
CR+orUSV3Y3oG2DonP64oRgsMM6BzkxGjXw0x9TityijxOh5G+NNQBxPQiSWJuLLiiZfMID0kIds
o8+8ObKjAChES8d8jKDC6LfNWxrhs4nGyZkjlSbjgF6McWeeQ59eL5arA5F4+DnrPeuzrRTVDNs3
bcvGO4se+R0sn1AUzZDW/6nj92zFpqZNlYvIunNyarT8TndG+4gg3LpNRhEP6gNEgBn13Ls6GVZI
PwWeYBJp8y13/1gykmOHrgZsT8EFNc2xEjro+VRUAipQO2kkDtTfGFqZ3fer7q0VlTSiwC/uhAp6
JhnWzTCNFCGhSVkVJrm4xW6A00rXhY9LFnew1xWoaulur5reLOWwoN2P1xExkGjS606urDBvPUAt
yHE9RldiUbJjk+vNEwSBdyyQc41B+JLr8HcY7Foy77HRLYX0kwdjjmxQ4fZxWgJzDJo9wuLfI15U
+/tHodzclH3MFIje0Dq78Fq892RlKJ7heONszuLmbhxuJ0leNvLx5EjcRo+UmlMVIhx5FHTaN7kF
p00bqcxzCRW5JvqsoNkIfOaXKJXk4dJoCQvburj19hgiZ9X4JUYmxRxrvsYxyDOyjm0rhVgG/6wc
R6tzWUW6yfSaNU0vkGFtIQO2VopT/HLJ8P6CSYfjN51E+bwU9TLIBNKJ5rfBMRr9JhtelDTfmEwy
MlgAJRu8qTNmb9X57w3ry0PEG1LnlBcBU0ttY+wac8SJlFcq9Up0tiFtlbB4DslVqZHVi3Kt97m+
fv62qtmoiLC72HJzis6laXPea/qXW9SFa1tHlI9W+gidXJtNEyO3Q3KG8liGFjNJkwMgl07FsGXs
3IYyFDqgWAHeK46teY8VzRdUo++un+X0hHKDl2kseDttJQhNm3Y2BJ4duh+5MSlX9yxci+NCtlzO
xQN5xDwayLmzdncXMVrTR7CEDSwpZa3+bDZc6Y193yKZf5l7EPVmm5TBtRvZaKR8q5L8s5x2ySED
L46+JLcG9kakJJ+aHtujnx6w1mxxS5gCVDvivvqOu7c4ty9hwkPn0aV9DltfGa/dHUf0cOIhxSFd
la+jgJYYdmXzjcI0PnHZQHrHIe4quqNKkWBw7U9q3/CVEXh0w0Q+VTji6ssvh4uv8duMaHwnSp7G
cWKJiOSo65ygNkTz2bKKjmNO5ALDFivQUGe73h00hcLQNXQ2jVtF2ewtf27Uf63uUMmwUCWQuwdO
6oCeADxFniwe3LKgIgDWpYSGCBYaDmw+WLJJxra7Ims7SB3+YWNUlu0t0Ze/e31su5B2W0GpS2A4
PThpt9ps7+iy8nODmYgi/DvfZscWt7e/IsRw9qfPoso2p51a/uoseTFn0TR4T8mZJIBxproQsM1P
rwcPFYibmhRpD419XDN9P0gRGBG/sadyTVgxWxniRUPFe9ReVvrhZiRVZ2Ss/3X3tteJ1ZpJX7i6
BtP0yiaZsPcPBachwE+Yd2ekp3hP/5w4kfs3q9N+F9mQNr2ZgD2ui1jJDNUlFc2hH4ZczbVIEdJ5
/mcFBLNkBDHCmlV/VCDLNTMVGVTHipw3t4pMd+NmwRYqunR47EGpWP+sF2mFpJzO+x8ARnrTdKL/
G7TfvWA4m8eGYmtwdJUeAl7jup0bv4qVQWnL1jCLgqTTYLQXKba2jOHEmi3A35yrRTt7/6aUwsy7
zWZkYXOhHETM7XOSKoE+FxH6DLPKVQHVJXZ/f7UeGIhjctaMYLDq9SM7dRTX+IDiFAvRmQf0YsBb
og9GxYylPDrexpP+w8L8MgFEL1APBE6PgiFdPKKf2RDG//8VsJCVmDh3vo714gD1cW6vX88aBWDh
Q/rfNi7sT+kYL6kBfZXzYvl7IkLnLjypDUFR1ZyrG9WFsUPomQPqA7HtNp+MBXhjVRTKYmgE7cId
rT0xU0zRpiL0QYmLdDg8021Fen49Ro4M+uBoIb+HGYOBe0Q5EjqKaUmGHyT8F2a2dzoS45KY7U6w
pHxUCkVuhUSLWsOJBpwpnyk6VYjavY31aOTQsKpfkAvBOx47SV3+Q35rpWit81aKBfXY4eI0+JnV
spI2GP0d/dDXSh0o9uYq0fU63gXydv9KS59PMUola5SzvQaL2dpYaOs6suYjUrlDT6FroqjO2Fpc
Nhc8Yi9LrRtucx3obrg+TmaJAPqcq3GMMZmoKC3Kblj5gHX8Zmjaxzi4g/xGc9ef0XszSF+knzNd
ICEF5v2N487GoViL17KQ+Wy0e3prm9oDJWnQsbt9xhvpsgPpiwj0cdKdCjvpJY1lMtqbKhSSA/gd
WklT4g/V+4TDtlLCHOazUF+e32jubf3lE3GRLb8w0aZ2A6HoEcE7v+C7q0RNEMhIDFDyOIz9ewJY
eWWIw5AQelv0RLcpCfDXROtU/F3QwhOGBwjod70XtdeZeSSbFsiDCAPlNeHe+AkTrJErdbn1hwdh
0bcVVLvR45NPA0U8irEqdkSftL/ZObYHWsMnmsOn1VYS7ECQd+glnFvOPXA5EyoD92wZ02QOAMNP
8U+WN+bHQzyGfJbS6Pw/QLY7fGizW+KeIu5VXIfoRmZrvmebAbfGL516EDyPMf+VEZZlv2X2n6HN
CUj4LLCTaODJ8a+kn5PR119muNykECtw3BykbpOfTYlqF5WII/kZlGREoEqGQ00ABD5xkX4yEuEL
9RJRJiVnjfOl6Ri60zb+NVY54LKPGKmsN6xgVQGK+7b1V1kOz3D8Uoe5deKru8XDrLtETrSi1CMh
GOBpd9fOJUCzus2X0qp4vKYwE99ZwKeJpsmRBjbs6Fr2VifNBtS6GCNxi+m+gsxLhMgodAebkWme
2ERU2mB+83HNGBpfY+qb0R/9agUDCo0+J7dU+wndo5Y1SqTNf+M/76d/twXNY3bxwQIhrQS7VtUA
4ICXBn+E+n458Br4altaTyelFb/ikXn8dU12uBO+RggMS53pueIxeQvX0xvEVaeyOwkXPjS9Fmq4
t6QpoZrm+szgNcIp22boMhpjQgyCc/srPdEkKQUH/Izubvow6cBWE9S35hoWXKX/03L7c3m16ZiG
DWj7wbGjJlszD8mbocLFfhbaOjbFaAfPUVSdOWY0WAVgH72DQjpQv3GB7w5SgKDg75Za+Qlvl+V/
ALrI/9qIPbueb+mgMduDcYnN0svykpANCcdjUFsN0Mp34ewEuW/QMNYoAopAkdvmbIAx1OhAyT4s
7PG3dE7yTyNorQd+eG5CcDyqy7BtoHG8oZkGZBLyFH1rr7nK4vVYDpjadyHP/3nKzDlcV9Msp8hU
IX/NBLvNTnmCrvFG47Czx4mrJTH6TxGFGX5upTFfLLbsdarguoNW78xO1ZNhSY4tUInDkejBvg0+
FH5TabQWJ4tpxqrgsspMG32a7JlT5WCSgC+htkSxHlMOB3O9OSaMFPDUnGPMMRbGAyO7AZ/ghIMo
gGMbWCDZQKcNnNTuYKebmtNznWc2YvtD/M+mZomHbedNUWa48Ni0XHjbqXbzzeG64FAFqVK/b80w
WrVmBuFDpfyUVUIbsW4gIczy1u1uf/vAEsc3hIxb9ovOdH1veSoFnHamKM/RwkJqya+MtJeZ/5wW
tD6sRl5CKzHEYp+SGgisO9HoMbkOukBkpSuurWQa/rvXEjWs1RRAVopwqI3ks8bRwnAW1B6EwOUB
P30pUTJGg+78O30RMBPEcKGuNtYbXbS/hk6FeDtudMo77Ofg5c+e90PDyrg9dVAK2E9QEyj0ifSf
3u/4puWl4Y2TujBPfpV5I1msZ57JXihPWrJQEGy7IjynXSgaLBDOjtJpjZrWcP+Mz1Bq3Wk9aT/j
uqHl/itRS0J7JdBfb/KoIvUW2YDh2r8I+x5u8lzf1GA2v3EieqEdzh0z0ELSB46E4MS2xdZB6UK6
04/XMDDLq8aYLWcrK1OrrEJEI6SlGJuyfxly4yLFobxfQtzcnwvefyGa/EVWDyGdtOqPq6MI/Yzb
vzmsS9R4N77fwZv3wbd6aszMg8gACTBGNoi47OqchYQUGY/44ocr/o7aBfxKTpNzSwh+Cyjmhi/4
xhhBY7bMAbHqXT0h0qBblWFa+/MqYCNGZSPU9HF+gm5BBHFcgSXPT36e8e0ngmygqmR8ricMXRm9
v+ISZy5UidERxzuNQtgm01koPmoJiIoe1w6Mwky/v8NzNSca2PqlzEm+dxWpH9fPo+WFD3oFWAvR
rSL9frwicuBrY9q6Y9fmh4WyakdNKHnvDIs1cdP8d07Tpv8IeIbQXDN4V0Kor5DL0U8s01fPEkHR
A2QVIQ0nYYYsMkElZwa3MdV+3c4163KOZ1PIjMVAvG1Bu0u4rKZsvkL2AXwW+e0tVcpECinQ08gQ
iQ/6MBfOa60u2spT5kRFybyn1+ed64eejGTAlNJzpk4jGkDLOLd8GijbT39Fp6ZXVQyxtFHGSyUh
tVw6PDWOI2LAQz3C+f+iNRNdU1YCXLZHce9t+0n83+XBJN1dLQWWVZum3tCmk7cNMM1Gv7Qrl988
QAkKNf6rjqtL4mHEBInOHs6bv0uwZatjKwXApiuaT9hKrz45F1P1a2iXJSrq4nNEg6oa1f0X3nWE
wglI7O/SKx/PWNzskyhAMydpsiLVWT6MXUg842K3A4AcVxhliEawj3miw1t5nujkdMJPVSda0H1f
bblCpAi99DTYN1oirHn7ZunvORr89eG6PuKxgCt5sC7EgynPxuxJjMiKjGRTNq9qHBsDvLIoD4Nq
2yEmwGjAgUZAtzK3pmZN1awIWrYylz2DTwDDiVde/NoYj/dSTO5Qp1ZeeHW79ahxxiAHX5oAAWjF
mW1jmE9JXktmmW4twV7lLyKr4vkfuLXoAKcVP7ki+9P4OktndMIhCneFUFnbGfPbin0eMZtTKlpB
WBuLNXKgWr6F6zjufkPJeUUTTbziL97/BEu4sQMRiD3qWbZ6K8igvFHgMaT3jg6tjCL3jIeHce25
+V4E/fS1cylGYscsu8/kFv/loMd+vjTj7sctu4BIcQcb+gcaLmdyIaDpYjEOzrm92UBoMVQI6ISP
6FnLtDK6X9O5V5SiP8itciFtv+HQ93DUrfe3vdSbZXuZEwlreyjmScawnY5oOxkXizGcR/PqwcKE
jCD0NGg608dNug02r8qkn2b5Zh2pVN5jMaAdVh95KH/6gnxORMUugfPN93eogUYW0+jUBjv/dtYM
JbVHFjRSzyfoVWf36m8OC55L1pixkDePD5TI2pYDBcAZupf56J6xNiqa+GYMxQtb1c7CbgVITz0K
88NcDBdDO6NEoF1l3zO7YnecYfasOXPHL/r9EPMK2yjZTaFZufjtQwGW38GXfQmq0wWoJ9QBxt61
I4dbm83OnZ5T3xZ2DPqVxvBxrT4P6DxtROs3zg+1tNewl5G+wBBKzWvwWa7inEX06gTuo6HxsVco
xkH5L1bXwpSJjBCXwLDksP47Keu+sdJJdxqZbi1lpqRlIRxHrBztZ+bvn8R0RxvMIW6olhlrRU4a
3eo8xUu9m3UP8vSNyGyZ3dyzjw0pszOid0KuDElW9vDxPoiECcMFQsTjGWOtEdz0OgicomFl22Bq
Kc7BF0jhcBGYq5NadHIJWbrfxPwvMUEeiYjTsx5PNmvHu33rtiRUthLAIyxePAlBsCY8zrQiTN8w
6KkODbcdlMr5Ks7zUxL0CvGNhuWw/bUGxfBBdq8ma3B/im6jWo2+4btg+QJCO3H3IT02LVky3kTP
HCLvT699FjSko+DVxKt9u/HlFhrK9GVNUWd0j1Q1DBqyvv6e8SWu25+1+2AFP/IflSwgmnAXHio7
cqbRiHs3xjCVO5UIhXdAUl2C7jqp9gst/phGUlQAuTGkYucsf1+2YcrQtceyboB6aw4+7Wi1+Iz1
bNblp1yLQxbvQkW+lhnMcN0SWlMU3/1NI1TYghcn6VoJoCvifKDfNX/EXCEcktUqvPz3KzQOpaIi
sVOp6x3mWEy86zRSeINMRgaNKK1Ng6YyDXy+m14vo2faWm/HBgTgKV9iRBaxtdjpv+mrwNOqLR/t
TocAkZHQLg9wKzSAcDKmgGKT62UgmfUydUtSzEfWov/u2VC8SdcZcM7D47FvykMicxjytjU5RsYB
X1hKYzjHtlHAMgCNZuFNAt2cKxVRdol/kagEZVAyIPUj7G4wATjoKnSzeBUj9fico+cxZ0lq2u87
vQpLVqks3/IuQ/938tAyHX4SCRg8bXIV3fSS9Zf/tRYhAEiolpWDH5wCS1Yx1mR+V0gt5BmWcc7i
UNuF4TlZ1TN38wtdNIx/CnkUkmtDSklaemTszJYnxEvvWBBjIkiOHsJMZ8TRjdnz4Cvpy/Gu4IB/
jKmzfPV+1jKu5j6KXlofteJNvzkJEkE+9yzpIJPnOf8mi5TqL4j1oo71keprY2lFKqrlLssq15AQ
gGwchUfynjwsM4fi2OfiJ/9ugNv6fV0QToQOTVVwXleACtOazpQyRlD+yYxlCCyzWp/0CbTcbyGS
rP3nF0gLDqEx1Ycg3dlN5aVcSyUDBbyODFgcq8XfW+QaTIU3Bz4qkaLf/evC4w92AqWmnlbmIX+r
FzSQmewmbdVqjyriiKJpwsNvQnBXgnSg/uKHrMehFzBDZdBJCHIUDWbizTBtGE9ydmBFeaadVKlS
qhKn+X73B9o67ByTCVP5kmKY25Vn3FdQi4oYPtLuMsSOc6/B1o+m5KGIIMTpAcjxSZW/oAd4paaw
4TBaE05TukulFPHnOb0OtIHvGvUoJSJLpTAQDlCjoLWWISKww+3wJ8axdKjraN+e+A9sQlhv0P2m
nyPCw2o11rZMdGQBPnkQ8QlC498oqVhNcCnCCYkkLdHEvU86hP75r+zKbpZXeyXOotlBQkav7ZVD
Oqlmt+nF8InuETPMdUtp9nvI5Gc5qusMyYm7uNxzqHo0Sux8tEf/uXE0i39atI9y2pnE5phGDZWr
QG/uAnK53vT8kOOXIdeBoTH4Z6N76uibC1v2Y7BLNIYPZ2lXkdxevgV9Qe80B+59JOaqraRj1JYu
YM+UFkLb91Yf93bZNLC2Bs9Iqb06dCn46/DZYKuw0KBinLSQWMlT+ra3Zmjw4r8jBETD7/Y/Hr87
b2NTeJTXS/xXxscIdQ28HJmIR/MP4JirjOLEF+4Xe9rktmYh+/NGvzotPlaR9MkOzgQNdyjosnky
CUiD2Yz1jmdvYqXPdVLc3nGUmUb4bIBe8lnG3/88M95QMCNhDwvzZ7PWskkHsBb8IUqvnvd3DnGX
MSsyaCoSP3eMnx9z8cADqM3wzL01Ahe0bbiWFosyEuiJN8lvXZ3z6oHHOOhdmmpqTxsFSJ7qpyca
aHo6zgBNzRCP9rijPorKchHqt9j+BdFIqNEGe3zwXEpDbdN3SsOV2P7esd24fzUq2agHn+A8MnXO
n6gmRElZJQwIjCQLPPWFwA+UVRTnOcQEe+yPbl8bq9Fcv1PFW8uEAw90Z5NgSxbM88KLIU4zBn+f
CUnco2HuzE+L152oPmYQkMXi7LUuEE5NiS8BWsW4T+XW+c5g5saFPSWWGqq/u5i2eFOLppINSW4b
2R/UCNalI56KRnzpW05EOPt/ic4YvLaOO9vTWpcxsRPJA8mbu5d5J57bUZxL8TXqWxArypcvX3px
CHV/nAcEpzNqga5CTrwa9OafsVovi2h5QG38t4pyWz/8564/p1auWqFaO89NJMPw3Tr/1Xr27M8E
+2K2IxcRAw3a9EEQOkBUUh9wzHm90f/fiBTLjh0c2u1hMB7JM7uCIQRD79/sbHDl6MRJy/7PxvM6
eQcmnfodefkr35BYj9RQseFGlYB/hiQ79WSQuy1+Pwf9mAqWtk9ks/b4W/PRXX1Pqa0pJGgc+fnU
n2TIY9K7wu0QT7kgXgQxAin7U/lvzkxnZkhKI4pUFVF1SzdsS6rke35SZeaSfcih2wTwxaV9L5PS
OXozL/mDLX2BO/W/ny1rCqIbwyUl49sSTnxhpug7Codh/ucZIVOUuYjVvM8NIRyK0/UFBkbBTUCo
wr/UbhDPdCvluxALzQ3m4m7pHgPUycaIPMjgfJt2o8peSkYfDu1uYx9AxVsAx90pg0s93yL/zTkr
fNL3I4U6KfuAB7Zn73Ag40AWt2bzRjWJVsuPX1xJ/Olf+o9YKmEqMTS0M/cPvE5eaIGHdDeY7F0g
6Jk38Bia0LloN30RGzZqyvznEsejqWyFLmzULEofTpF9WA7JL5ACDsTWnjkJ+w11JnaTNxxo9rry
GIOJM//rMKacM/mICCd8jO/1lXsZZUisZxmuo48PuRBajZJUeaXtB4z29kErf4duslehBNViTQQS
iDJwzq4MzuGAOxfU72EbZtHkeSS55/V2vm/C65rk/I3senuN69r3nFP8wXbMAMLF/T169XAIP3pe
gFAJkfXiJ71ugyqKYQxplVi5C92ascUeeLaXg7pr1SBUp1licy2y7geghygChPgWDCw7/TbLL9SR
EsR0I8aQJNPuLUZiwZqPqkMDNUAzrkDSq364B2C6se5Oxc1uhmA8dEvDV/0lmh0NIAq9u3kOC5XP
eac5RIdSW47oB5tgNK8NI3Me1d8htITWPnXLTqNJHgv8R1nrCzKLXnySFKPOERxgKGLXwGQy283k
7O6kCOVTUndjXI/zDoIXUAtDRi47Gr4c5PfPqzjUWPkpN7ZyxtIi4/OFt3RCE2gTHD49vQ5opIJa
cg14XPBI+otWN9U6qY/R2tsIbOPeXWxyiio8TR+ErULEaiRyKiLBzZEz5pRN+SODNQqQUaObIVYH
mEhao5BTeqDltFRnEZqLofNmsbfG0LyGt9zhyA4kwp5x1osEEoSK3Znp9es9x5hT+1qD7TeVR6Df
Bg8cTYkPB26bmZ2gtyWeVKFhWiCHVP4ARdLuRXJAMHjwr2XCzm3AQelAz9aDGuaIQIFsM0yKUW8s
EFe7vWXwq6kP4fhih1PuuHMH1U4EaderHGf8Ecd5fGKX8+2dIPpCzTdFF3xKAIesQwkYGfLRZh92
d6ZCjzKfZ+HsoOLItbbeNV6CLbxh6/pTMR6r3fpU4HfUP0opaW/TWcb0aTr+mYVRaDFkMgavVWha
Ql4EC3MFZTqtGXN1C1LuFWOA9NbbBqIiRlKfeP8qGQSy53E5LOvs3K2a1+PBKrJz4U2B5QCXBIrA
M1ORSm452DkyJxiiKbGQO8O7ix2/EepjFONBmZgpSGpQ8RwwmM19RQ/1LPBkGPNh+1vdU3AepyaH
AhrU93pAHpNlZltcXO3DFMpEKt/LB7EhrRqjKfs/jj6BJa2+ZmRsEH0D79vHYHEvvoD8N9G8M1pT
SBHsrcYk62r7UMk5fzKIoMuIQX8Fe4+CZUHmGIm8ngXBjWlxDpC+SPzuRqncXpv4gvVS18FwoHkX
tFueuorUrrjXxPqa7FrYWG4bAWTebFIdUvhCoekhob4yh00dO4Y4zw4ppp7VIIoCDOOCeuZloE39
8oaS0pJECtEKMLOVnmD4mPu2ZcgMB4GvDh/H7snZM9kc/YTtv23rhTGmxQ4IKYrD2itLyxtN4jJ9
Z5X13uwBfcZFXJD1RxQEk5Xo35FHxAqP0tXlI7qPhULZBblYJek5d7mRSd/zSw6n8sHdZ/5i2JkU
Xi1+NB8te3C9OnLKU7CrSSkD+cC8xDh2bk17A37gsOZtsLaEbaetAMV15leWFoqzNMgVPlb6ey0M
xq21RW921dUchMQfl1QPuhNnKEUKOhDgBOR1cMom3c9NogN2g3Ky5TJKAEnlESa45ScPcdfjcb6H
f9z5IYKs2OjwnFfrNWnbtUs4VCH1k+CxtOaL7rVdfkutJeIqlh5FkMp8H2eSoKhpk+X0Ag3ue9r9
llR5eBpSCQbHrrk28pU+39zMAxEiiElj4DbZQcDCRm09UlKm12bVWI0yf+f6LVnfwVgfdc4uVxBS
sjo71X6NS1u2zTjIhP8gYevI38g7Ad53sE+t+Oc9xHacqQtYwzNVQPsidXqgZGsWzodTzFdZFQ3f
sU5EbyY9aKZ7SPkKAvOcr88achUF31OPEmjag7DEiDLHP2ze2YnWAgClvK8YzDn/zL5HOlKHJXqy
P1+gtQ6ypyug0mhCXzO7QIV3bTrZH9oEFx0KiH7kvOF8e6fpu9pUH91pbbNW2T1uZ6CyduO7gs7i
PWzgBXV+N2BjNrrD48CC+CIkEfIShstlrH+Ev3FNG2eQ+bGUqExMfu1iJfxmv8nBdL11+fh5auBk
xP22okkeZrjUYIMzw+eHpgCqJoOMpbGLNhZ7RufyKOAfcA34T+icQv38UBsYd8gw3MOer+k0pfhE
OlRdPuvh562qasNcK/VTbdPSh5++kNWGhmtut4QGbLLfPRYLGqxCEj7AR/FROI5/FPmKGjjrICm0
mrhtjZY56Lh1uhP7MeiwIucZ9JxJ21s+juVfKKExTs0FmhL8oLXwUnDsC8nTtReaIGqsMUoXwY7s
PnwaSJHE+UjlKIcTzGKtPVdmzDBj++Y7+PxSDjoi1tJTfAbg1bODvrfTG9HXsZYgx+s/mn4DnGsQ
amWdGzzgMKeWWqsHe5XdSSxD4A/ni84qd0eF8N9CamFmegDjt5b2B00O+AY0gcJnyHfHd5am5gYN
zgf1smy/eWhc5yzHsNiq66bm8x+UyksLyKx6kPSMs49grIRj2wgUvGZt5kHAntki0LoBGumEL5ai
aXlmjfKmVjDLflAefmd7IqZIN48jrb1hyWTBlk2AMb1vSh0A/KlRZAJOyICX56wm7+5Eo3Qx/krd
IH9539Wgca3lfGTVQaUTqNSUhxeEA8YvSbUwNtz5MfeVDKY1gJ8RSjoEqpdNBcmmGJLT+hvgZcPE
XhwH/XN/7OBiA2wAvB6PI481ZPIujYO5rww1WtuRYNXZUxcqiwkPxkJhACajOktinxtqean53n5Y
CPjA/wHxoH5Zmpu+D5Zrw8NXfNlMlr8zC3odp6Rqzle9MhMYfPHT/vGA+M2EOpwnuznCtuPvRCvp
PME7yXcN1Els+ohiR2SlKk2NCs16n46W59IunesPgArGdvDddGB1i1uCytIYqoXA3OaNVVptZ5w6
2sOkEaKlbYctmnjkq8lON5vpKhCJ3OFMFeVwuR2bvIx6iPtwdZ2wX4r0Q1rV1Sdw2IXwHw715cuQ
+L0CCjxZ+Ac5xMMaYdMxj1hQ2qilbKdjiAbYAlC7m4GmaoraZ4uX4HKlj+mXlJPrGg0hN7SUhIJI
6PqjXFDG0j7Bk49mFEVkyxOgbXT1E+/rPGI9/YItehLNudMoFE1RqwS+9aEeKJyEDDu0cZpWzSSv
QRq82+56LopI21uzEsdcnYTJ2fdV1Ajq9ctoB6m8ntP6e/iCzZwaOxPgPhM1yCOgB6kyk/DJX/OM
bT1lSoGEyCqXhnlV9LPwkdpSR/4rQLbQgPns2BbAvlvNkTUZhaEpDzw/gk+MfqYtse1weuWphXDZ
mop8Dp9K6ZpquqJdfqwx0qNQhx2DBrC49/otEjspr3TlYJthgCoouEHkt99lmx2fGaNi0GZbvIE3
D4i3IzCmfyMwCa9Oheyd/0Q242YRIilkuBhCT3j8RGI4qB/ryRwnIb9S0V5eSOfZTjbohmsd3WmT
6ADfnmdqWi69CWBH2jJ4e+EFQipawuQan5oFBPFa2QdLjTYdpfn0Zu0si5LHRNGuwXVuHBUc2nhV
zDkT3Sxfg+ugwgBvGTlqHip2i9mfgR+F8g92yJsW9AWPz5Psoj5CuyJdwupjpsFZOZfVQQYlRsER
LflZoYTqIj87//vkxDe7zEMMpRDW+DiRgCg1xkzT3mADY+8zASNGovKCJXigZkEX4+v8Q7DkAUJv
ox6NrMJjeSUTvn7BMEsYrjNF2n+m/z+Gl3pskOxi9E3SZBekDOkbinWCXTFQKtRc6p/iTCsxvlUe
dO4uEdTo3qx7NIUc9hIodpsKE6ibdWJ7SbF9y+LfROfkYv9LEVhtkmiB5ZEow2GhwgsW5e+JGcC2
A5L128ApsA0+8/DL7beAUhPTYGdBIjFilrZtfZeWRRrYHEUyKXn44I+o6wLkdFANjlVZygRI3rZ0
IRIty19C6gLNbHwc9dp/z/Kczockfk5W7JYwKPKIP8qwsa97sLoxhxxBNulajf6ZNjd4ZNlEqfqr
cX+uwa521B0DahRNirK12u+6J5hI/YTxJFIMEWxUWmwCmEma4zhoX7gi+D/ZcaITvqoq+SrMECaC
YXReqVuesxUYPIBmx4nQcsqpYMF+Tah5YyLzNeWLJJYpQ93YGNJz5J9zGsM9k/jDWU25G74OuN2H
ilr2bNEQXvL+6ogowkB7q8TaNU7ytsJJJizeaJ++z6tUk2iEbQDxyq/o/k/6T8ntTnyTUjZyiXTj
CIiW0rswGjR5ugnxM6hMEAq0c+ISow6HtNplRJS+cYHAYFgp1x5tm9uMm0sKBck4qZj6gWALuY94
EIpzCIX8GW+EuVGin2G/hP0mVcPBhxNV40gIulYXvVuPvGpjiYLeBIYUZge88IDUTZut+LunStjL
gVY1+NgMrdQH68v8UBtLUTW0sjTZBw1lhA5qYprFrqnR470fBqPBMt7GGH0F2QX62N4VGb19jqPG
Qtz3vvnDxLvAJxtRIPGL7dxuJHDHi9TSwM766Yhbby1droGfjRcqosv8mZ22Gkm+YfBSiKUTi7pF
F/NXKHW54UbAQf0uazkusI+oGdAQAFEd6vEjzoyfv06ZJJVoXOQsOo3JnIiki34y3mS0bslb0B7g
2ZOw8xgV4Ax/7wRfwN+ZNV1Sn0/8BQloQvfrOx92JG8bNahN3d3cgLnYXmLhwj7LGR/8ZlHaGXTQ
VcAwpXouRug5nN0zsnNsq14dSxNB9suymwctVvrppI10Nzehn3IWa/gjkNKnJ3DEjUTPlOotCacm
EEs8VmCRbvXg9yGrQ275JYhNHpzgGn+vlYeazut01LZrPIdr4n4sef89351fdZcV6yV2rVhjSEo4
4Xqh4tCL3qK3s0s+E5Nefy0Yt/1JG9ukZmECLUx8PCMyo5nDLA6K8wNX1z7cpGNAeU/isJyYS+I0
lD8YdJ9RFHcU5xISU7AChkWRW9/9D38gqKE+y0KTVCBJHYsuq18/W/D6vjoWJm4Uh87f1s5dRWP3
fND864TjJXCn/Sd+p5/jfGy+wjlNeRfiSLGdUfL/FX5Hgc0NXAlxtchKbbtqk+crFI2FMKpqs1cn
2Pvj1g470QRIm5ON1LwrrCI9+N7vm9YNOgYc73Mzv2cS5BHXkzdtYepLVb7oNS83KWuGYH57Os4F
5tn0t/kgz4CJSIEqRLAVtSOWi9SYhzdljwVTpVmNoctC9KdXRa/r2uhWRcK0jLPAY6ZveXkwyCyu
5g8W4zEbDW8yj04+3aOybxNUoI9/ES7sAqcrj9K0CItR6bG9iiy1jecFaI+YTMZ3rJr8ZZwinoyO
p9tYf82bAceRwbvSpZsvGEZP9JuHO9SEuLFPUbme4yThSqP2DmMoEcJ25CbfotgpQLqkptl6i31r
47W0YOf81jCd+HECtWqjQ8eVJmkv5HJQdwHG5r7gLYP/K0CxOQpTbBkexmrAvW3nDf+xyImjrn1h
TpjRYCn2UNHX9cqrYjXRFplwm7AmlYb1KPoX6The8gdc//XmEFe5upuM3Cc2qDHDvEKq+n2MeCok
knxMSijR6d79Xl5Svt6EaPtO8LhJkMS2WetMQVBzSVa9uTAqWYGDpGSGtADam0ICd5tIfBV09isK
ANV/XdsD51IE/JTE3LZLFX0RWHG51zOzSsF4RJLepK1px3uVJ8GkdwjG0l5Qid1Yq+fCUcdOUjaP
rl9W7zaLA8x5TVPYK4V5k6qzORLPf3hG+wiOMBbvUS7J7uMn5luyv2M5fDpIBCeuaiy5ZDZyoWHR
9vIfe+hI64NXl91zsgJMGphMd+HszLrgIj4y2kqNfwUDBPvp0FS5ADa5XYf0BLBNJ8qSz4MmORkA
7jlHNkFRI/TBBJ5vd6ja7CigcN9FIgWXaBoRbFy0MG4HeqSADhzatgYyKItAOzgbHC4OcoagMJJ9
ZSdGbQ9VLBBT143NBPBn/Pd3wiSdVpIvd9p26L8PLP+N11wMK2Y46yAdE225GWQfM+vq4bTQ/gUA
FUmkxrb48zCzjD+7tsuEee6UpT5zEw72wRS2+eD5cmEiZS1+D0MZED1FX+hAxJ5BeLU6GbTbKLIw
dwowNhessOPnCC7VQFlEldD8OyUSx7oBcYML4cCYc8CrMUF8iqJ9u/6aazOWxojTzWnZlwzunirw
7TcFr69sh+5sZfbDKTpczquN9ye/AABd4IgsnoldLK2u8qbgw9JWM1N4k3m3sGaGu0jFlGBv8SK6
jmRrOX2WuiGZ4hEagSfwqpXgkS8Y2IWBu+XoPAqBavuNuZqEPrIqgdfzucSALS4VWp8mMhmDzqiz
93xpMi1/pfSAzQiOgIelfkFnDwj80yype85JyKmCyHnoKSoqVyLCph1NXsDHBm+QdGCfqYQp2A5a
OCGIFT/VzyrBwkt2ePI/ZIPWauaGMAwYuCcBo/wgLGKc0uKkjLoUFUcLr6bT+kuHj0ncD7l6LGdv
M2OWslA2+wFUAm0xusV/TS+pQABhpig9UZb+rmFuiuuXbdPJfvUs7zLRXgiGbuS9FvYPo8MRIO+b
YjaM3j99qUsg5AS1zZR+eGnXk03hx/gF+76xV3lB1V874/nBQqT9JTx9/R6r3oawtyjusdATDiWU
Ls6u6TunYmSI1TbyQXVtPvK8PpX1EN3bhlhbtU3xPiP9+B5/fVWDPJmZBOO/ZMrWZP0UMFb14TZj
oyoYfoa9LdgrA5hAKEeLbmr1t6ICLUF/5xZbcpXiMYhplTEU2aIqOBqfU00DvQZhzeEemE1/RdXL
EtSRH/7TiqJ4MD1NQvLnVt9uOArCgvN0V/VovsS2/zILxinVs1ziA6X46u4kiNV6QnHo77c8E9GQ
iawPgadQrkHBquAQ4/4KtO4Xfig67hgxVoDtNJTCSImaVptoPox4EbLw+H5wDOjom71nQTrpEFX5
c5JOQWYluhyE8NiABvChATZKfFB8P5lkND18zicR4zXYPcgi1LEnUEMCYe79O1FYl6OWbXI9TVE3
Js3+blrTPAm5hzsMbdxxcfBaMW/f3QmFlrH/yuDMHUYPN1qZQnFgF45Fd5vqxj9UjyoLRCdj65cs
VARupjOjbnmSaZKykre5+i2t48NNjxuf+WGj79CGj2cSdUas+HlnqNPHDLp1JLXsK0i080IXF3dy
vVwW/ZhI+RSb/yu1DgAv/gumHAfU+B6YXBlR6/lHtdIL7WgIVmCv7R3zguIaOf5VvlUlfrhCfzbu
L0TM9qzp0bHbcL3UHLjAVJJntOLACb/COtPeIDIFEU29HzDavqrJF5OvzefRGzhfS/GnkXxzDgNB
tjgV6X+0h0V8gFIG6zWDYq+9CRuPOtAoaHb0mdldSnJK2SARnduFAbmDcPVCE0w+C00sMpsXdLwc
d+jbOLvwcc6KG3e1jWCfD+tZrJwxmWMCYCBxN+GwmVoTXtccorhp6AWhU2tg7Pwh47BZ5IWpX+Zb
9K8Vt8zZamBda/sFyV2cSVl8uegejDlPQgO33PcKy2RH6nAJSxDA+oJ6kd/g2nF87L2Y01ArQ7nM
K6g4GgGho3AOsl54MN0JToyi0ppL85fQXdVadybTA9/MHHMRmvpwp0awYc3oRwnaG8y2P5/rtn5X
axBXFcTI22HtTsCRUF91sd+OVdXai+SIJP88zxSnzolJyE2bIVGEo96/MobIdo6x+503OAMzltha
sCgqwGoEZPwKWM19+nWDYuAvY9nLBPtr51ORVD8ThI/xzvrE2ZE1BhX27rUDVBLsySU2F4V5VS/n
syd6bHhFdkd34b1vR9+m7/9SUrOLY/V/cQJtZEuVZQWt90RDF47bOKfTNn1TNa5g3JwU+ylrHXgq
ju79rsZdXzMWIrNnlwghQNV5c+hE8EV2Na8JUSOOWlusr5ucx2NM240NJDHAYkI31LkvHFeNd2rG
BhtgvzmA2NRHfWxAFLEHcepQzm92YbrElZFGF2rxVIJTmSXbw6T9IL6vbihnUqt1VInQFdQ6TCOG
fqXNKCd+TzxgRiIdrEigMZh4JJ6nNzu0S3EWD0tVAxAcDrEZfbjjOuxVUiviZ+BqskwWc9LNOri+
nW09XDivTjWNzv5tDllDd7TaeMvqoSJNtePav18konbnjAbTxIjA/XF82RLvFGVh0UBfVhpQIBH8
l0dm3Jh5O3eOCbBrQPRk2Y81rF3+dv34ayzDbn+g+5SN4DAY5CiVVYoxzeuNrdHPpOkv4JTQN0jw
Vp40y2BWWUuCm9N12rvfa46Vg7CWNTtQK82TF9MmaIJFvJTMY6KwNdcIemCA2vgHCzPsF3UwvmdA
uELqLkxjeNs2EsvC4cXX04HQPIQRi3ARz5iLJK5dQOxmIyvFLYxr98kROm+ali9QiJGOAcPvKnVo
BbN+REVQFNkCjj9vpGeFga/vQjse3zmSWblMb86k8UvNjxdwUC4R9DkBZKJ9mP/ZS8O2UkvReznZ
dDntC7ecREIg3tmfo6TThkq/QrqmCIpCWt5yLJDPxiSd9ov0htHoM7kKB9h3iK7rfsiFNfKgU3i6
LjpJiG3+uum6RveKkbaK1TcoScxwiVYIz9hXeMCFH4ji4QpjZh3go/4FqSktDXn+E87giCZs9VSU
cHmbesd13Uxm/W+xSw+4Ir+mohvqy5F9n1ioB5w6t03RtzljnB5UtBoNoZ/VMjnfcAgNn9SZhHXj
dHCwTLN9E6PK+MwpXFc30LnUL1MottxCW4xsFLCm6tPJwwqrayNARFRv3xxLeFV24kWoEyHuAcZ1
bLaDOwAoa+X/E6xM3VSyS1xilBlvc9dvxNVmlqqdydekev6Uv6RlBOiPpN84Yi7TTtibgd0vXBoo
A9SHfFZ3g5gmaoXY19qT4PovsSkMmWOW8RdQUtG1O4oskycg/j9gM3jUTQkTTI+TKGyNS/UbzMa6
J8+GDA1nhes8qrWWrHI6z2O52AXGnzjihd7VfF2//fUfIJEc6KzGKYiziLxYf9xPHArfdv/KaoZq
daTZpIHlPK9z640v/QuJw4dxURgvSOV1S+1hUgcbObEFWLkujuzfevVi8h/BYASzUxYp7uAh/0Zp
WHZ78FwpOjb6O22HOORp7mv0PKzMlCERp4ukObJe+dFmT65snin/Dt15EZ7ptSWmlNlDM3Cg3avG
4K8y6EVIpEZo7boNFGjbXXalP6x2SMS44XeWEpDpIXqRnTo5+IMS3v8Kbqhl6WR+ZJmv+CT+NnEZ
2VyP4Ev5iktkziElcS1ebjvTPxOxmoh+Aa4l7NyTCOygYUsM83wVHWiDDrFvFmdfQku9ULqynL7K
yJb12iN2OBirm/ucU7mot1ZmYpJ3EKhZwLikIaJQHyPKfvU2EmOpFjDGehyHolhrL01HozyVjXDZ
JsWAm852mXG3uh8KxOt2/YP1fbZHqz91IUq6BwmccIJgjvXz3iurCe/hHaK3XPr5ivzwYk9cA7jg
KorwJnR/R2YWhurM3IydIkFf95KN5OzNmfK0X+loAj0bU/hZRDCq9F6ktiTNoxPoGi2g8y6Moqkt
3l7dcjXdty1wJmu5gERre1QEHbb9D5BSMafATOuywELd3uPbkfuMBXsBirxqFJ642UN3Xy14oCca
jhVjhGry/ev3qm5nVCECeTYwhFJ6lCh8L2CtP4pjk2VNdB6umlg7WlrZgSo95hOlXqqqEJn6fSZR
uiQCzyFY8039741ozopmo8ePLiAaT4ztaCz9xxfPxSwFLNgOiCfE+mvgQXOwytHJcJQ2eFTpqcSc
42JZ3rudsmwCb4HoFSC+N95khOBfSR3NK/Jc7a9edIgu2ifDFn3ymw48InDcrI6R5H01yS7TF/KI
jkWQNgkG+32MtWwYgl/SueQRHCMWjVHfmD7ZnwOV6umiHRrVVNDdgo8Oe1mLYun00S49rqIM1e5h
ca+JaH8EK53tAIBeLSFNbmMP5SE9IAnVp6ZUVwkGRjzBpTKTUxTvwX4I2I0MoRyD4BHmphkWzUrX
1dUH38ojWsl9KnhbS7b1cTkfLiIgO0szbZXVeh1AsWtVVcpE9IJp9SmdbkxB21MPiMukaL9oxPCl
ju+crdUmPEP+VYDemdqgLPaYoXbe65qFWphpu4FhHSfPxIAjxYhFq24dUD1gG4GsmMgrn/sSbptb
EAQMT17bynZEv0klkI6JauhLgCg0KU3gULoN1BmcHCKP8MuArDA7YswWquDW7zl+NfLHRpmH7mAA
Bv0TUVlmwaKLdSeWBNdJuNKgIiyKEkr+WCK2u06K/sSYDBWXMFWkHizQToL3u02R0Qb/tV5HBauC
6KDTiWB9LlXFr2VSHy2vsgIU9ooVFOJTe3ogrRS+Zk5jj/6PTvkAFzh2MdPvzeaK5mPwx8xdlHN1
S9Gd02n+g56+/QNjYiovx2LJ2w5mZzr/2SQ2SFyuGPwQb/7VYVM3jgf/0hFhW+zeZKSVHA1qkkhW
LFJmTwtoveDykO6ym9OjA15pDPUbu2L7vcFyTKOa0gEPFAvfoimMhzUTdeVwWP4mUseTqk5ubXGm
kPYBcghiIvxrQ/YILRZ9xGtJSJ5BaY4BjnPb5OvZeoYAYKeY71UiPtUN7Pbo4t01Kydf3uQGDphj
b4fDJjkTXW3CV9fH3VlrgBe8GUel+xq7Lr4sZmsiu1YgHQFVZ2kf7eVwcmOJf0CxyzO6Y/nPQEIO
vNLqCi1/gqBdP6z6/7b74AXy/a3/KtI71F1FDxiyYs8mdQh/Pi2wrQLB2KTmEvmX4QddJjLanxHp
o8PM/pG/yAkjBQBu6pVMYhWRCdH54wAUCz2nhCTEejg9Fgs652fpFRvaU23zc0pYruKTk9CsMg6A
YOY8t4WBXQsDfMRtevzeuDb2QXHhfN4DEYlmIEKcpIJ5eKswjBlHcZWwR2P4nc8gVKWeD4Pv5mem
u2NY/p64pGvemju53htFgykKODYUAOT3UBYwMECVw/aklJdGki46MlpTHrOLJe6HvYWvLJ9PIztf
btyZSn9iRFtI6W3FakqocsRUvN1zD7sPNL5b6gefZEu6r8eS+H6t+R1KNJQAKD315MVL11OnK0Fq
bWNvuUO8NlXXMrGg89okB7sPJDCM/NrHPALLiIrqcT11EQZAF7xsDx8KwKRtB5hqQeSYSKkwlLkm
VYdlrmdlK6gVgcK0Q9Ep6xaJrioEAq+L/T9wr1Lcj6prQ/9ZzoBcCS3aihYr+pKeB7uQ58eyg9xU
HUTpMRIXhCJJnHaXDeoHkRWljJwDE3bl9JY8xQJzsZuDi9KOOf7mvASPtH+LFQnNSI3wSmthY16j
fVIp2J3nbxV3f9zyCebK43F1wgbyFHzJLEGohpqHyeOyjlBLAaJ/4MMZT6yp/Y6MG7eFvTCBixJT
S3YonT9XZsg6qRzanp1zQRnu11HqDEKi3aLAkLPEVcrIV22j3jbTKk/AnVPm/hLyvJOF2nVOspZT
ZNKE5EHK5WcPO3YpiTZPqHYa77QmEnXXg1M8DnQwnQpgsZ48BYZ/fhBn6C0cThxDr39CpoOjkWtR
irfz4RYO6fNxB23xuIf1NHVkbWUKb0DnF85Qhl2wsQPb0teFR+9ug3FoHWTqJYb43yCoxzMcqDDQ
h3z00fYv9KyJOEHjLH2s6jK2KoQgKUxLzmU3llWEDwPytE3VIMdACglwsTpp7xdOWMlw3g5PJuxm
8fuMadsH7nMB9cM84kyY1BqRPdm0TFgs2Gc/NIjmHa/Y8GU0Qib3W6ss2DRet55VCPE7gJW0qEK2
SYjfUKC0mcqNBxt/wz6Gy2VTVy6UTTa2UZLaIM0fX75fZynvHx9mf6Rn+SEHZD8tpigQmpHOAX0C
xBXWI8qAbpI1uM0rITlS7rdKodxXnFlufDspAHP/ppCRqon4IGO1FvZ3l3h00dBofgErwh7q+QI6
EE3tW8a3BssOBmm3Dd1CXhvcNcy0/m4mZDy+WzTA4hB1Z1UtPQmmaYB7vcDT+GShAfIPkBg+/1dF
aIbRmFgGCpRVQtRY7yjw9zqRH6hIJLgIR91a30tHgXrwbkSx8LjoIDqbfME2zcmB3ZVRi10zx5wc
6MQPo+9z1pp+c5xwOx382gvYGoYIFz+IyAa5Vg6789i6Rm7w40cd7JXU64SKYP896ko+kjr1k7Kc
oHp9CKuj6CGdi0kRcMaFN6NdwPOPLRNnynOZorWtjSN/dhfuU09utlOYUgNSCdrT2LWf2cLenLz0
Ftmce6bSEOJYmgeiehLc32ms8mRNY99GxLGwAwJmNFsw7mdxVZrnHG6RSeXtzn+d0WAfWdFVjC6V
LttxvGbNhEq5NzLrUvzg/mzNnwiST3E7HvUk7okvOoIIKzfQKMKnbXnSvjUCXSZsy1AriVT+ZC/G
oWnQRrKOeJsozF6Ujc2BDjJSwbVOKKOb3rdHikgDyN7JvIVUznAzXVf13XB5VIPK+qxJa1ht+MVj
QMrm1lMhbROjinzGmGs0AllJ6WvOdip2bO0+A5zfeJ8uPVoOcu6v1OIqJrKIE0Dh+VJZZBGrA02z
RlIpLLwsB+nZpcqWJ3sIjS7O+/PQVM25vE7QZ6sSb4diZg4dKBaomIdHp1+3taeUdIuoUxsV39ni
zqTc2b8TIjeNmiLWM4dWuwa/qVsEc0/DbE6zfrLRhE9LjnaBirAzTYZmpm8hA1NIGlrwRKzSOGas
IwliGZcMkA/HtcTX0aOPDc0drsAL/bieegSxjbj5QssbIKJe7FLRVV+IZywhamnxyXWh3/GUlvTh
fqf11J9yS7xEMDJpQJYLZ6HuPTJyQDardiF8tkMfv4X0ZMrkFn6Ll/FhNmC3ZZdbNKbDG0N12iEP
BxBqCx01O6E6a6MWsPtWwjTXWr9e7wnkPhnsugUDJkY3sPAjhbGw19E6whphqDd0mJI3oMzyqCFB
+yE0Ol68AKZkyQy61xFQB6mFyZ2Fpuq905URUQSp62nfnEPDtcfyGCN21zyhZdirjrVf17WScVWs
K+Mlgps5Mw3SCHjWyfrpiHBV+4jcpv0dUMP/pTZ0FPXvAUqaOzsN+x4ZfgUk5e0J0CgrT6xTgIwp
Eg1DxGJInHp471hrS+XCqOJfDx0TujOtPpOBFmS5Lg30ctkE4k1GtrFYk2LuidftrToKxTFPg4ry
a/eQhJRFkrUKuvomYdJHH6LjELIFAdTUAQH7KvFDQ49/FQRZo3k6XWwPmRcFE5lGQJncjuUZzcBf
WX+uXAqyRVDwn7TDwCTAmdfr1AWdRxDmYp2Uxw8LZMwupJVWknJp81PxP2iceOsJF+TS9ExOUFKm
zKNSLn6Drv5mGOaToWP7JQgcyR1b8o50629vtPR+J119neUwWj6LD8rDvHfZMO617P68Ro86RfZm
aGYf58upgbd3/83YkABlM6MpoZisjUamrkaMWfA0n1hTm0/9NinVhCL934+pXxNLJGCzwzoibYIb
QntjXpzN3CW3K1XIDgHWZHBtSg1xIGgReiovKzjHMNjXsdvm6qPUxoIkJ8Su0fUN64Q8bA+oTBrT
XcKACC2ZX3aoIK481Ank3MP8+8FXAe17LOd20+L0jOOABqFgmEzj7FYjWH/Du8n6rAaNce81U9EQ
l3Vd+6Yc/IBDjExdTPlSCMnFbfjeqwZcdN4TgxRuiGUfoF+73eYIRoDzwViBLeU81bQzqYZvyrCp
IdirGTb5pl4AXM7K0APMD1xw/v0ZnGanCz5DEfNZ+sdtCMGe449RGmPuxKD4VGIjGi8x28Iy+3SG
ptYnYGrYZDtwQ4ZAlke9Z8BkBghqL1j3V/TCTTruNFrcN/N7aUlm/o0W2p0wv5Mn1W3xQQwI4wC9
tneCt71IiPjlN5CQ6xSC/KWthop1Q5nAwOPmOega7ReolKk3f5vrStH3duUgYpSGi/PoX2jz/mE0
vv56kgYX8pB/aBnjrW8GJdCc8OppBGBGWlzR6R7bsGr/bbszNhDkKqkanuwF/zybgCwTOQiTbtHU
2CyaNxZxkelvHpWNUkLMzB2PfoRhxOsrPmn2zE6p6tXskLhIlS3rE526qziukcAexztzLZHl5/os
QvJ47ophf2CjK29PVteoD4eXpigkrDVd7ZbJh3EFxH+ofnG6UnFltekawTPWjTmE7BhoWEx6oKZE
3AyXh/A7BABJ4c4AITdR9sRnllSXYQ5YVNa+xmHPsdHLu31kanvDMOrslZ4uW84bMN35v2zvjobJ
23ZoPtwUXoMH3KHkGQgvXQ5qIc32P2iMKuvfrc8uKyuPxoyVN7BzOWbfSnSsgIb9qU9ouy0lnWkb
3FmeMG8F+0T/MpQT5aVcbnOGvPI2JK+K3uQcx6QNub3oeplM8NyKMtmJVRoXAyIDPtqxIEKsfgao
W99eYuDU2VMPM1f+Q/wHCKo0Z04u0MvcL4faZS5xtSW/dDrApUFe6mMkzxPRiQGaewUXfm+WS3Pr
oEHeUaTbDU1lFnxJTB2P3mkJxOLF9jnRjRAKl47naLMoMhyy4xmLZyW2B1AabORlre9qe48+gd6D
vJl2WVMNIin//9RNtWePtkpszafChJoOAD7HMf+JmoEindnKMQzkT3qymeQh6iHXV53M3bUe1RHL
NuY7ABSSXq6i4aay6CeS73yN6h6RXYop65vv1KbUcO/xoYw023xLFf4XpsLwdZAoaywSaK+6ysU7
Xe5s5aV4/2g9fjnp6sHe2PWwYeW/Y8gCNm8sOCKNVtboiFgHgjbExhPqTb+FZPgzuKGXgJSUHvEW
dtDHrIESsXceY1SOXHuop90stAuSPkmT0ZIPRONk1iQEbqSdn/0wcGYm5TzUZ70y+gY8LXw1zSal
xj87Tk4LCIspl8RV6Fi4R91UGx5R2AVm9LlTuyIK0RKLMcqRuEGnduJS3lsjqxlD1AA+LOvTOBaQ
/jr2I9pYfQXWSR5qkuuYjqfH99wSuUjn0F+nrY2LQeH3pB9G/YdgGei+iK+2L6eA9TNIfpdIxKpo
4Vw68uyXCfjdEZnYEWYW3oATp2iu+nCXhLcryMPxYugl0ZRaLbYOYkjAGq0buDmFq3fc4ElCQ6ik
0GO8J73+Gj6rosN343paoYxW5+BaUXb1jS8cH+bXZLbDnx6jK4BQpg+nHohcvpVIabDOumP4BfJO
7Fk2A7w0wrsGqHucwQ9tcEvKmP6jTQkUion8ljCrFLpo6V1Pq7NQdgDJ5GBgIvDoq7ASNGU1fzeS
Zm1lwzfOSjmaV/h33j7ejj7Fl3wm4JaVmaoFcFJCPYgDhKaJokqsEV1roAobAK5tVtfaNeUvpkQZ
Xv0POUZ0VbwgVNf1CuVe3dm8vWRveOXSOoIuEYqE2pDefaGi/5CCIHd7H7DU8bFL6qiSokzznXOw
nTnN7QfN6devuScY6ye6qJq5NckjMFujYVh11+xvH4Sh6Pw1yYfZ8csWj8AGc2RtPwtuZh0ak14Q
Xo8yOMTWbTLAFb508vnLQkLIjLVXwDQikhMpmNfTt2lKELqqFFVCBgvPGxlNlGh2yh//TIFcBgEz
JxT24Q3OSQGN54LDhi7ti3BfjWpOCgz9JOFUsZ+iyq5VEZbu4RbS81vjpteI7uZtBg1dVtvPYPv5
OmgXtzrusxVsrOuBbehE4zXc3s0KbA5Swxs0Bll8o6uTg2Qjk4ejxA77dqXbIZiqZWRmXsv+xOF1
eTcHYiH/xEGSVm64lXLIsMR4IrRIU12BNwmxURxLxNwgr5ETQ3gdaMqHssgPM6oz4uaFy2UHa3TM
vHRPVbFlsCrN8la/1cYWTZ4LCTs79DsliY8a9E5bETGSX+eO1vYBW9nD3rJbmpBMd/eRuJa+9ZEe
8CjMzzeyM9MKpa/HMa9tcKlbkreHiu9+4sxGo0yTNHOJVDRt3IVKYmiRyN9LKfF9tBbjhspfbwX6
ceYNyAFHXWQ/cNHClUQdItvkW9BiMiRlG2oo7QJJPq7cJocYvJ7B0qTHUqmoklKYTXh5OYViO/8B
CMtEAcOLrXshqtkCqJ6ntev8IRtMzGKA3NdJ2spEU+hOefzruDaaOP2IeQymPZ9pmdnwtGKo9PBx
Xz662+Bl+Rl9DjKBtItjfRGGXYBTMbRrkdM3U3FqI21rprI8H1LI17XAtQGWTS8kq1296wHsLT9k
GKZRG9qpWqdCWdNYm0JzYtL1igt1SQtT8GF4T/Oqj9DEOJtOmovM2wity+2sVHncAiPp5K6GcKh0
2ejh9+1ghnkQ6F6ynfUzkxhnXdEI+F+x0u9dS6WuK7MgOffSc58QzgiRaKNi5dN/+VuVwR8n35nf
6vuTjz9F7WExR5Sdw2hUYA9/4yhABWU/sAMvaM1XX6SsB3RdJV+A2Lh1Rwth7elFyLxuqVieQMaa
iqhkH+kWx5MdFzDKK7gMgzbTrN+vYMxNvMp2Xq4uWTJr8spQGxHC+NM5cVA5jruRX64fb7VHQMG0
lXGtXIYk1HXfLpkjFMZ/JYa71068yECxLodjsp4KfWq1R1vPdPLJZl9f7h9TRIraAZD65yRADm8C
q+Y2owJAuJwUY19E+nTQHTlsh7CLCd/jjFA41IhQE35ZgnjuYp4IMD4mzH370OCSVUDnFQYVIsqz
gp8o3KPTiyHDviBQ7ROG8yT4jM1MQOO/Gz3aNNDOEBZkHg8IR4Kj1Oy6aVaP5lmbzhYLJ+uzYGQd
jssow9WxUMxfc+5YuKnvPxl6LT1jO8qCIpelf2kh0nUsIiAhWdxR9GQTdoo7T8rXctKqrlZf1CxR
nSQKbLTTnKEX1XmKXV/5Bs0lonrGRpI+WzxLU8OT5FZa7PaesoG4847ArPDvx1XKi8NR/Bm3k56H
XdT/MTowXLdR724VWkwQutL67lZU8cY8smaCVK7aC9hABUyh+TbOPZ07WsF9eXHLWU88syyVC8Hp
u3CpO7mGNTTYVdFYBPoB0Hsr6qG73oL1uZ1+oq9sbwh2DEHrVbOe+wzonRXtCebavxCQkq5UECfY
nUdEN71KERmZuR8Gxj5huBf8YM2zTDNqUyPk9TWM1PGp8xB4JwQBAguk1bjAPAmc5l88uGoF4orI
SzwaFA6UCIugwn0KxASCt5JlNPhqxDXbSccaOGJti7LFRHHU4BeNv9qBqI2taK6jMzFuTPUF38tZ
Jx+0AecBTnbC/se38lxvOYMOLlTbUt8RK+oUcGwAwqZHsRKTc4FxiMRolODBV+X9ClQtFc8kGB0s
W+zl/FfJjZ8wlg3cPj6ZiS+AGLUsCx9+RPdEl+0ivJrqmukBPwEqnj/CkPuSdoMoCQq+01ePDWvR
Vj1G53D5Nv7OeYckY5CYFt1t/ncmsBi7UM3PTYwix6vGsOZpeJKXIVNJ4mD1T5PrpMFuUAEgDyu8
AuwXtKZ0cEoExwUeZ5/v4o4lO08/T/YV+XQbmTyT2dlCYqMAu0uvgUql5FsI1MIS9BLctkOOC0at
zhBtEAP6+ECO43baIrwVLANeQiTAPJrraiE2P+j2kbFULfnLLvfbaVR2zLCnN3mSXiRLEQCiN4F/
jmg4tmjNzSFtjo6OJvhFHNSOm7igIIsXDnz+Du6QK2xIYf+LAhS9frV+kpyrMQhgLzw9lvcW4ZeW
QnfOV0T2SrkaRVmeu4uXyH1Z3LVryZyonDWibaZVz7AgUTc7IdbiIPQ1fA5hi7IH2WGpIDoqtiHf
gU3yJpNmfO0xYH9w6g8ws9HpDfUu8HZrmMa1paHV4W+gjRYNXXu2M3OpQ5dakPPgICMewk7WlVVf
RVVn+ngJHn8g/9MnJLlER45b6hAKInvrtljcvli0DSg694FUuFSXewRDUbeP87S+H51sJoq/aile
TovqRezl/86XU1kNuvjevU9JrfXtcRaimk2/EB+7HLDOmpLsK2Rsz3WaGn9bbBKxhWoVwGDq7Dj+
XlI+2n2VoeELNAf5Il+MA0TBKqr8Av0MPWfmdeZnpJADd48FoJjNaNfchJmrNHfIN9O9lPp2ebLe
ktW6BQ2siiUBGK6uJnggAp8oNnEIhwai5ph5w3sDq+SuVAPruvtecOZyBjj4awuDsJGhPzzXibfb
PIni7GVVuUIeYb2wwFEQDhU5IO0bHHMC12ui7O2ha4LlnCFDx0GdKrbQJCo4n0LQKE28gcpA3GNv
KqJ9I83oyNsWshwlyxe7WaM/jawzKFkDXoYvtYdaNGajHFAdz3SfFbkEbCSkNyBKpJKY7Cm2RQNs
XKuPwgnsn1c38WyX5ou9uL2DekdcIAW/1Vxebq4v383Vv8/qMljkyaR6IMNs44C+kZjVTBu7zjNa
T1+r7EZxwBCllavM0aCyI0oPDcR4bvIG1gMVx5LHtKGmICFaeIYuBbYhMqufnvByWhgVe4fKWiO9
ZA2xKUap2g+FWPLsCE7td2V5r43gsYlWbjvmzMxIJptLRAbUIGDNZkYQGQ28j0iwW354zQjB3lb1
kPugBbfe37IaLQaNZKZEq1HZ2seOpYj0/VSoAxRroP2oxglFrnvdFrnFfIWKSm9CfojB+UFtKxz9
QZ+B+p2FRFVVZ3wdJkWi5pSQqGmG2X7n1snvwW4Qm3gFsHWc1FCStgn10JXS+sw7Wt72/5J01nFE
e39iin7rcrdvJC6IYJGT1/rB/nJpwglzsOTuA0RHuTxaIxbAwn7OI56N9+ZKUIjtSsHHjuMhhBD8
lBo9E2mdonZd9vKegMN0OzctcSkQmv1TfQ0fv88pvI5N1wJwdMdRjSwe5Y2lVe/BkdlQP4KKuGC9
Gsje32zlz9Dy4y/UOQoehcQK1/7LtcbEKshWjrPM5rCkBS2MmSgmzcz5hurt7W8R0Cnb4mqYjYBM
KljNC4YFJVoJ+/F9r6N39zG903nDPSOdfsp67GX/nOhskPCoLocVmULzkL/JARHrei8IKjtGXHvC
lSXvASAQd/xaHEsS5I17xZMNqs+m9p0024KgPEVJoMXMRgmsgD0ipzhb+qkYgJzvHCzQL/l+eMCX
bNk1q2hyCd7/iRgWRhZH0yafNqdJOTgnjV2IgrDp6J16qcjdKcgp+YgPM0H3OmjBfNSbJRZfm2XP
7vWKbRWkrxjBYiSrX8CPwriPiPL+j3LGBhQY5LLZ5lJ1KpPg9oXwqNYPP4vmntOZHsi8WGcb0jJM
ryTEVQXNbLUNEf0uGezz9JxSkxi+fLS5h86WmwUvsiEjUfGSicZC2CzQ4RTOWRl9KmaD3oHcg7be
w8pnyU7qBedZPu4chxoU38OEfx/gmhdLIxanganqGU7bsQyvTYTETNdnSYqTuJAzIrAOLHzS1YHU
eBJZH66ee6JX80w4cviUzY5QphQCx8hMlso/1cwvbFxKaKmaXArmS4y5MRSistLGNEjYOwgYcBSW
e6pT1P2RHHtB6d7Om0tfMFvURYNy+fXNhqOJFl9fQ1bSiJMxFMfpVnncswOFXnLjf9CGgu0+hgJW
FJhuaK46HxSGxdXhYlABFqG393NDhEbS0GjGwngDxjegWflpS+1PIwkjCEiyERjvkXE4DztuXTpV
6V6X7UanU3yXDvS+d/EokCpJ0bTVXTenlx5C5IIWbsngMIcVoOnTwV7KCD6mxBHzzWgIR+oxRD9D
UcqlFXdbAhoDmDTn+12Kvve/wWEvhpJ8oUiTHnlAsioghYX84DaXoEBfywyGPyrQHwqRs8vKY1r3
NUKBYQc8uFX0kxU9rkyGKWGe4Ysp+zGDEeypyBxj/K7FzRPT9mO5q02qBFItiMTsSniYgZ8UazK+
jFrWGJbcUBfj8anIJ6g4pc367WDPf56jLG+mrtzoqpQJ9UdOXzudWbhKnBcG1Oiipd1KttIs18Ub
+u+gsn5qKGM3doRrCl5wVSrcKrfEn2xxqVmMmXYj3brKlhFTeGkQLQHTIpro0589yXiTKLqExFcg
Z5tur7huie1v+8LZW059zfE6DZIpGkGBaRRVbPxZkp7KG0vVioCVfKGdUfAueJJE0QDhvBDjshpZ
k1TfJJIj4RKBdvESY/1gaQr6OfEuUBPKXRx3dOOUXtvvdGiIQ6NoytdtbzvpuxZgXWMovBejEZP8
CUZGSZSke4woNWXY0B+hQS4iR9d3s5eAi+3hycc6+nK4gyXecFjnXfFOv9VrfIjEEsjrAm69D9HW
ZnCw1XcQn2s7eRejlLODn6vgEyrEWy1F52wZ+31TQZNMU8r+QP4apbxGXtN2PMpKjrmb2m2rmsW5
ICCnRAcIhkx60tHCRkvGVHkBmA/9+h4nwMJo2ojoI6ae9+P/Ts1yBQP89F83jTge90IZF0t0K+t2
n4Saty50YHZeGPRBOiIWZB02aFj9fHSktby+ksam1ofJMgj8kBwhMFzgqqBdkF5JKytSVAQsCAiF
KGdUtd/O1gonPKT8omcKCfcD/umGepYSD0uDJqUvG2J09tacJyLugNolIYJh/GRAsq6cD8rHAs6X
y0iIbwNU/pfgkvmR+yBJ4eyOLgL56vlGGuBaNHUXypR0DArUxhIDIyTl/ygF3UwYo/eQrLIHBS/E
zmRZHmOoq8PvhddiI4Y/eVT2J2dGoEA5jj3CLvZmYC6SoHYXpAQCWuO06Va0yNrojP+Uyqqol3TW
NnMWNYq+3qM3IRYUz2kgknmBrCHFomCLuUuY/BMab8G4mI14WrjD0wBu+3BDjZI2LVt5Jvjqcm/8
awgtyHIQPLhgqJK5Zl4myt28nxyH7bHjA2ioy+x5exafUqqQkIuVvrglcnkQPvSEwNOKvAQ1yGgp
MJLOpFnVtl2aZzgk4EDHj2DieZ7gFSayQ/wQe1Pu2M7XzTPKYaZ5/MxGqkWhD0ucNt5AGZAOVhED
ghHCUVRzIXcrGpnjU5RAUVsyXU/Qxxm7L8U1I+YON5uvUICHfd/xcGMFWAC0QELDyO0lEOQOzl5m
ob7nul8yxl+qGiYVHUf/YMpjTscwq0snBzBEoA8t7ly15N03dzHzeW1CJ0+aFetZmZJb4yOcWCl9
VPL4/5FLrt18ErAx+Cx5u49raulJlXV98HM+6wSp1RZNU/3eBlg8eu6T3GCNWFB2irK1LNEzsrmS
6vnxYOaf3YwFkPf5CzPRLpuLA9gquOebzJ64m9XYYtpbEBuu9u2O54bCp5KM2EZs90kmkrXXgm8/
f/vlhR55ekK2S7tvqy+b5tBlBrY18pBq8fhxc55KPp1wfDd5fcUY8Dw34kG0EUuP9PXTt+SlV9sc
gpVs464xYVKeu184HMTwsuLBSMS5tjd8kQvLDzZfsRNZSNhgy3b/7/xBGnhFZXPt16AUKl7lr0ZO
1AHdJNl2aVUmTCxeDDt1XVrwKxKl5mwb3Gus0JmhdQbZQp9c6VwKyLjmO59+6lxwlIzBIQ0U0WOc
Bkl4P4/ckekpup/d8OSFlF6xvMfpN7m24o2IVKTg3c8gWSVEwPxuJvbk2GeISc9gPqlc/VdxSrGb
ShK5Miuq5d7vvmyACxlvcx62tsBmmEboXMZqXRocdGXJBDWomwI7o7WPwPc7kmR1KuCqXq0bRMTb
WqD2QIzCEqmvXYq37nkDf8ZMsxEXGmAwecds2Ketb+MoLbvlZ++XkviPuPwE6Pn08LDcMLMohUf0
JjOEKkNkQ37yuGAbKKVVc4+30xz21QRkCDvcTy6KhI6CFZb3J7ZsS90podw8mPN7Aew1tP+8VDzn
4Q8JHmy1TUkaDpmhKSoNYX2tb7tfpUH1R83JrtauaPdDcyiUPQ3pguBVl1DtI1B3klHynWYXC42u
cmCKId5mLg0pN+6hOLO5HphjaF62E3YJtCer74v0RUsSTfxKQ/Uak/kzEszyi/aGpP+kQrqSOHL6
2fBUTF0T9bYq0OxZiyFQjfl/ApYs0S/v7RXVRlk5829rfjLRicjfm73drq7e+oDaQ3ksFZd37zME
fVubP7jfD26PecNj3w2TwHrIUXMqV9CItWl/sHDkPkVe01RfHCCAoxpijOb30sKwhIbQaBAONBM3
V2cHNq3j07mTm5lErik5y3o+UEqrh9TAUxhKXY9Odxjw7hFFbLUtmgKneABvizOKtpwFOAVWX+8g
AlUMqAEwJh4hzJ04jgRbjkAjsTzdX2KVhgI55lw9RS43CzKLjZHLvHpw8oQog2+N94fOiNmrunNO
7i/n1RGMEtWkI6cPJYut1OPyhKF620WA7Cz9bL6fHZEGS9rJPFgJnXl2EiqCzJNPUS+heBKmwxj2
E2MBVfq0EUMJ4vB2f1Xms20rRN1yzjM07wSOmCUW61iSXVYXhan6THSWD5Sa1Vz9uhRl2aKzvEZq
fsp04PovOa/pwDnQqwQDf0mSb2QdUd4o2w5+Ga/c0KiPdFp8z7ySdpaMroCImcRGZ3TYICxNVViU
yqlNwiEFnBaYbe+Fv8iMyH7mwMd2uJkALhsDKMIeitorOosj/M+lqWDxgNcIeumeZRW1bQSDnzBU
JpQNdk6i2tCwg5x+xjaEjPNvcG0SMwHva490HqFRRD49Ae3hs/mKEO/YI3Bti5lEoL5jogCTe+Z5
U0BqNzFcUkNXzasI7wTUBVZ9Eo5FwYirC9eFC583zSuVPgQtY9IXH8pSxuTyvtqgyE52qzu8lvFX
R+4T9y8hIhEP6Dy7AG57LrfLaOLbUrxFmVDbrtmu5br9/IonPavYcsXu7scd+xeDtfN89y+dmiu9
S0Zdgda8Y9HKaV0tYrJx7Jiefx2RWPiw9DCWxL6iWABe/oEGgg1kJ8YDDgPPbyy7rh8g7bUakeFC
dY196jkdOhpzVzGRjo207+4Mpn1HB2sWMnEpVbP3KvEaYnsZOV9120Qmgj+s29PAGnmiFu9QegL5
Nr/Cf1HfMkeZBXZUdWPyTTw37n7kD5edtorWYon1tPLqLRpEL9TRJAf4jSo6r4zVzkZYt2OHX4HS
JpyO5tmfzUcbPE1XmJ4Yvkf3TaM1hVrGMyBszWGpEvOCZP1nAk9WTMchDOORBQKW6yXbvWlA+3mC
WA6MrffTKKqjYMJEy2LCME6q0biK0zudymiqMkBqsBpPVMB87iH0wHZAFVqp5quFJzkrtRT9/6do
c8YqKI4VDmvaIYql5f0tzixDPEU9k2vEvTt4xRk3WzBq5stoTokmQdrAEK3mMZwicGB8mnU9vqsR
DeMA69v/fhX7sKIcucLufA1Nb/brMYmlOslObqOTICthTu8pVDwFVeu56XOktFobRTxnArCCeVWc
ItECUtIMZlvFNYHULSBOzgYQBio4fvfAjffNEDfniQfMNmSod54R36oIcPszZzd8AWQaxJcjESoZ
KbR3KX206fJTr/ZPF8hcTBtaBKcOlLKG1L2WBftgqmHKXzVlZ5lgK7SjT8W3WeQc2vuF6m7gJuo8
GphbdH2Y8GryCB5bQq8nfh95gjv63ICpf7njIfqaCHswYC2Xsihu6sEFgZJKiTyvP9ggg8Dcjbkx
2Y3OIFPP6Xedl2+sh+O5Jcxvl9CnJIXXCfbdiUjdxMLuBz7YB0D1i5trC59kFoFavavZv00sV+1y
lpvkmzDp4Kf7s3BArglj+AoPP2CSzpENEXr5xFj+u5c4D0wLIo3Wo8GIqPgmzAjWcQLNH/c83kKh
QeLjVB81voFcYst9Fv9Kg7r+ljBXEA1Ar5jENf5fu1HQk7Ctamci0/WC8DpP3f3tb6YOV/ESB3qk
GzksqNXgFWtKNaHO4nuKEVFfqegIK5YC0GWULPKxUEIW+s6PF377VB24nNY5pDYAiIPHEHdeFGan
N88RMVQpmACdOV0bGIHIQLWAUFj5tXaJWtF5yt1I9bQHKbJHOGcxjC7SHBRVYiryfLnEqE9CQlvx
DT5LGHqxp6bgNvl+bI/wkf0Pw03nW9W4/KAW2vr9YlRr/QouUnjgWg67JqSnwu4sMY8s5gUEQLT3
qC9DSEQopdW9NdhwuXSf0fZBtFNfm0pyMQ9WehLQuNHdi4jIktUHVRbcX2pq/EUjqXZVshHSVbAM
mdGY85KqixhxCru0COMS/Fcc64MGV1eTdx3IaVoj2NYUPIL8UgrpKWPlIxZJd/Bv0spcA+hhGdNC
pHAgOP4HzvZPoe7eFhbT8BXht5o0l83OuxnJGJBGk+Ea4NbvN0gwCIYfk+uZr8Q6jwd4GpLSwj/r
0kyVoS8iqb8gLYFGh2ogSIW2C+idaUI+vVzlsbOwrhA0s+watAw0E1cSbcSXkT1UiBAIHwH9ezAo
sCgNVVJRki8osbvN9XUfzlcY566jY3db8shjHoiN5aEnPJePuDNpyDhYZ4pFjtVNtQu9edJU719A
1+ZG3dnO7nLGOhdAmzttvU5kTvcaTQeYN8qQLA/kla/dHLLR6L31x711IkWdEIUsr+foL1fbUXsb
6blREP0WuG9n/U9e0ygwfaHmoA4CCkq5h8x9/aYEfl/FLmfy8/mRncY5zIchtzIsnyJy8K06RuK7
xEXPUS9rGW0hokQzG1F7b9GaBr5WjUItUzTcEGnJIFKd9JWCbbMp7f07pxME1AckSbnc64J4pn05
1dlNQ47rrp5X8eKjNKSwL7a/7ejHmZV+OkgdQhMT31X/dWfSkauncX1+BK6tDaphVq9T81R0lxGw
uE293FMbwLWr6e/fmbWETQ8qiuURHfU0vOZjlVNlRG+FHcpZSnwJifK6aHwFiZ0nVh1X+jZdSjbn
2B3eXg8+IBSTzuSwy+nUQjLgU/imeLQETHZ1QkD83R2SYtqFSAqJWn74vOVJG9OWtqOKRaYQ8iBq
RBEwg0yKys/HB38cTKQTqqSU6qjfZUcx+bdHQ7jPMUbm44P/tc98WcCOfEWeAK3g8D5BLACrXA3l
xG4XyO1wkyMFijGE+K8RAYJkwnIOWMJFCXEHl79VEUmvpRRorXYOM/DvbljD4UNwRI0VLF8AvjjR
SQMP6lAIHQt4JAQ2dzASEMWLEZDt6v0oJyGCATkBAoX99yIIv3FTJbcEzgq0YwLZ+5mOv7/OSCJ2
TySmJU5fDcAS//CF63xlzesRmmV17jWHzsCOjagi6T/rE0Jrnz/D6NMbG6ZqT3adLmjFIRyb+xQ1
p9dKGixFcPpu5xTfVdtc3cuwtyS4GqjkPAbKgwv3UapPcBmGfD56KrpofXMhUqR01sBe9QnW+A/P
jBYJ54vtayh5Od6F9/xjYmRL5/kQ1Y35gY0RWvM9oFLq3vE4LgGqQiWz21mXjGTYAKKJGg+7Eg9w
OcNYxgYewScEuRI4uuAS8x2fKX5tFw02mhGNzEt3Yfwc1kq51SoaYXI+dTXF9AMOyW+9dxyPP6RG
95hnGliv6QwabT9iqI89AydL/DBnCgfMCT0omA2JMpa8tmPl3thj2rTrZORuwuJ93GMA4VbzgkOR
QrbUO6dr+4RjWzDfdzAlTCbek6aL7/VQ6Lm9tPUy6PL7MVplgGFEffnNCxvv+DfcBNiOrZZPVSsi
eM1nlObe2+gmKdWX8xFoe9QQ2FJpcvLbqfogW+c4hBpTDk+jzMzAoRGCRMtbONhXhSWG7z6ELqWi
7mPKeEeQDaVHIqDyfcgD9TsSlMfSdVKE1QoMt/Fhdn+1sLjbv9FCVh+ZfrvaTVTC5CV4z2y+7ThP
U3hooqNl5xvgTkQgMrdtQWYBq0fVGGGfRf73ozkvEIYYYRcD8+1TVWlPvLGfy0xzfqCAPc8Yhmuv
47XDMxgHFPRGKlpRAZss66fMXmEsTywfkT0aQZk8hd0hv6Ph7y1QA+A/1FdyF3PAZVCaE31Fm0Pt
OOuT7Cr5OLWqEamG+Ds/6MQVyA5wI8ZBtaiYZyUpHsbh02ISXOBVDBgtQZH+NZyIRu7LL6YVIXrB
Cg4WKeYDySTihNO8HajiOTSEsUXE9RrYArsN/lAS/NVxmejQILTOJz11xL4P1WggE/KQY6MpLxuo
h5mXMOszjHI38UdO6X3hfmUWmzrOG638fsjjjCjdLzylsR3OuIAI0vJES0jikVD/K+jZ8uWMEI7t
L+x/nmi1u7R6EhJ3xBZFlIyd3rWExJyhkFV2+/7pCewn+Jx1tPEtApdhFnhbKApMIqxrawvx/cXo
oG0a4cDlVKSgLgA4WLG7TX7YzNFZd7lx9uqEPB1oo3kb+blwAWu48VfAhS8n7+TcqlIHNbmId00F
AF+35t9cjD5YxL4c89EXvUqYM0daKUBLWzVz73C0yKJQQUP+Z1IRkTMyCRwckvm3oQRDTQDnZwYp
pTZPhvvUp3VcVxjsXz5eWNsDzggMtIoGNriReUAq8hCxfew61xi3+BZnEHjSg64ng70vT09hB/yS
pYxccVjP3y6KnSD2RzcipVvnktOjAlsDG1tVyD4Oeh8zgzCDdM2NpVXLVqXl+u39eluI2nm/4N0q
7Q9VeV88vlB8I8brtjQnl8LvhyiS/yTpOmG4ZCJLGwFnIWt63PJxDHMi437E3tkDmHUvqYVQQNS7
sv7UMtrvtgfqP/u6mkAgIzS/0jmgDNyp9eZw9Pdty3VaqtB3ZjmhD5FAJ6lAWFLPzsPC2X/ulA+9
4mvSVsPITuOQiqo5Lg7hs3WaUfUyMNl2n9nDNocBAhSDinqjAj43qp7RJ/kevTYHtyE7mgeFaoZO
y5U+I3OY30fuoQrwAtsAJ/ACa82Okr+nQ2NYrqlBJOwmghNA0ZFlVcIPXgyv+tyNP69eJ6SdL3J/
i2fZxGswPvj7n11HyG6CnbaRK1XDPTIWzg8SrTn+z1n2H2UkMnwcvHvH1OAhaGvkTYIoPBqNDJkY
sM8F6QiZQbOIM5rWenXTcRoe+n6R6t8cSu0DcE1fYfYsfwyEy3fYmWAL1BniNZyd1gMHKSzvmLij
Cr+4X6/FFVBqWDpXy7PYS9iJ2fUMzOq2YSZxjRKm76oeE7ogfYzAi5OURaKBs+49BjbXr1ICGhjn
dsVpphfqgYxDD+h9827YeFNhSr5nGanAjy730ap12ELrgWDxeNRpqsbgYQXR5D/AQFO3o6sYxfon
I2B/K0QyIhNczUUSh4D/lnW2xalw4fvjhkY4etBUNhP9xTW1gT1LFPAFJ3YwcoBZFT5WbbYxPOvW
dhGUTkuEPnk8r82dALdS81accDIBZERKsi39ja55o1+YDKLECaWNeEOCq98d2//BIDPyJ29qobF2
RfTNp1vqKcTo5fj2JqG7tSvU8U8ywinBQsFyLwsCbbayD7WltxrlnUouhVNHbjP2oteCGD+aSSt2
rZ/JYCEYQuNSmcQwFGetSo2CSo0I5EiRDTd75xfzdADdhrOtXELQQj/5AHRIeA2fmOSNoXY+45xm
9rzY0w4Pc1CT98c4rHBzg8a4BFhHGsejvw2tftG5B8odG6h9jGsCpjkLDUw7v12HNdjG0+lG6hK/
l5231cQdIEYwNnwA03B/5CBII6HzUBytl/6/53qfi4LowWS1J7ww7U9VxYksM8Tx9+ty2eWPAY9w
YMKijOXjp6NsW0ad+igqQrVmqvDzzTm0sil3kyKRtc7H+gJo/JVRCKuc4+bUTop+0zciy0lEHNW2
gkIEpx1ny8duCS94Og2o1h4qkpgLYrNcEyclWqzDYj2KvG9jMumgeE3Dj38LFQySexUh9jDX+A7W
gMIRp6tybcT2sw4LP08U2SWzG6twoVB/tf/PE7qvG/ClpXKEvjX/z+Y3ma1XIqW4BHUuWbQHciVa
oMIaFqJRc1bd0pSfmPqj6zOdCAK1sJQ4x7l/gzzoyx4JxZ1umo+GGCe2MnUX/LQVa5QZTLM4Ui/o
Hi+Qc76U5PAfsYcEr6OHYT3cblNeKfOwiWstGDqrEKI6EcjFxwG8dwc6ZnFuZJZZiNUcPXsC8x5c
CFr7zw8RrqW2OGmTheHOjs+7CmI5eIxVc9EiqCQnpUwPkOHobVd9hF2RByFgUiodWYBB37JsJEwn
+pDIEfVKRzfnceXLzAUoXGIl7cvgiKzlyG0xzEPEbaadmtD4shajaxqCDfBRo8dF6IiM8nRAHnSa
Qharz7P/oFeiBuhQ3nDBbDANcddUOaWiOUeUbzmQgXRJtguV1emKxkG50Gx4xg5qhNf+i5jpzKZ7
pKTqRsVPDrudfmvlvrtyiUpECJcB1m+brYm/GJSEH+BwWRV4Iplgdg/luhc+Nrk6kxnfQib5d/g4
OFH9d8GqpK/hzLc3jiex4ArmbuR2fOt2wSgjMz7BRW594W1Pe7nyPdtZT+gS/Am2mGpnAWzbK+4j
UoCnYrZahFm4EhgnTA5LXXlNLtWavvn+ZUo4Avx8vYwmMeeHCDJtMxAu1HTRX5c87RKfJmYoqbI9
LcVgqSwgfoGJbjoAHQCp8syjSQgXcC4lOA2Vk4R9B6zZyv1M9S5DgdGWVoL2qsAbHBtecVGf7LCu
I+KYI2Ce8Eq9/wzr4oBKMM+VYPFvBJKjYaIeZkkv8gQng1xB+kglXeQ90kku2wfdSx7GzZ4h/Y3e
pV09HO2jrNGYzcZO68ERlK1/tldgWIq4P8xGhQCKli/eHYIjJAU9+PdvY3sKSZmO2CY4p/pNNKTS
GhoDffBHD+4oBLiqJD375998r6Am1SSEIbN3dz5RS+5R42omozNcgwJoaMQaqF49VB5lfOA46i1S
GRXYXmgDfqxFXKlCcRA0QvXU13wsbvgADNpnCtAUMqa9uXBSvE7mZIi+APSpnGkDxegL6M60V4L5
Nvwn+aU+dwhL+K5T8esNeDshjaTbEImWdTGy55snd24PtFa1h3RMQb9slARrpwRzQ7OOnXL5IjKp
z1WkHUpPMUa49Y9sH6FPS10cIGliMW5Rn0okbr99TUX92h7UKYe+zmL3xsCw0PEJMotofysBepVS
VymRX4oktQc5A9/D8MvvOJFsJOOh0JzdxsNuZscpL51v44FnLIjrG9P1EJ0GgQVgyl78oG7ss/PD
USS7PYqhfI66k+0bh1sdeMl3QmyVGGpoGgNrxqKyV3qVH0F4WNlCEqJp61qpFXINBmVkeYTt02Uh
50eLp0uGkMNY9SfuwPIdQhNLWIS6sMt/Yjr6sV4WxRrU7K8eACO9KKRhfT2dHKWea7HtiU8MdzhZ
H/3fNYM1+4/hOyTRQ7pxaEHc+BzJc7dX8l7GpXPSFs/zt8O9T0CulWs5RMQCZDR6yXm5lbkoLe1K
Ip5H2qRmZdzOW9UjVNAwvXO8wm5PMRYr3JZtD0nra5t+TYyb0DwuDZF7lGBYdv/vvpGCT1NCuus/
CJr5IIlqYI7undEZVxnHSXvF5al1OrjUOLFz/1imMkmSS4CHukm/vy3ZlLu97mkFuIci7WEG9f2R
5uETSSEr24TJTwxfcZofaETjx2S+7I32RfuD2jYNlkfB+ppIFvhph4HXI/XaAxtZ5dakxB/TUjjP
02PeJM3Ben862BdFYDxopmXbzEwLFWglK5ElUPjdqo1JHcVhhLvo0w3i8JRSz3j3HCm4wvovhBIz
comrKk7SGLYY3e/iLlPUJw4EXTt3xRCAyAOSBb9pmF3GBBi3UDjOu+mm1LAYgyyHV2dr1E3IZYkd
99hhR+vXH1E/osmvxAuT0ZQlYjuH5K+Xq2TzPDVpMEcTqt29y0SD5bzFg/0ABduVPZbyn9AbNiGk
z3v3aC3xoxmU5A+DYRuNJ0z9LUGIjhm8zQ0JvEMBTHj9bSXNX1eD6ON9hkfMa6zl4QAVdlHeQJbb
HNAxl9GjmmXGYR40KSq4fXJXFZo3Szq3UpyHbziYn2432mzXMxrji8UST0VvcCSxDSi6X1BmKrCN
ppXuWzZR3gtgUxzQRD0+Y7rNDXExs+5QEGM3H21LiDIrKgFFigiImrxgKHlVvWwOYx+hSrlO3Ml3
y0Ar46GvzW7e4qX10fxbtVmWXkFrTwwG79MfYUTb6TFRl3iv7rux4Q5mmv8Yz+83tqxVHAcbll+7
9RFiXOzd78EhVrkUe8A6HAff8vgcHaX3f+6lIptlCRrqHcQztpbIDUywSYlt7fV55pRNTWR8qxfb
R36XPxkdDEHz4wfcdl+3QU/I4tUeNNyBUeYzIFNLrCJO1VIUCtNOS2tZn0JeA0Lb5T44xqqDIB1S
g/d3BXGcOWydZ8sTuChwMjSEjdhVbnNqRzjDJKDm083xpsl+c5wA+WoyTXQDaS7twVA9fiWNnTw9
Z7SQ9DyyQTCiyVscj64sUMM820uj1V7VVLz/DI+NaxNLPg89JgKmX8zq7noqv3AMaGSV8pQid3M5
PIConnQMBKL2nRQ5UKNr/EMeTjGrhoyjWnf7DLi/s2MxY+9PJSCQAA5TeZMbp+LQJ5OyfFkhZ6wm
Fo1P0/FhbC2KwnIme14XkOD4RqI5ZIwYnM5Tpp4hL3d4DQUvCtpwlp4/cFYGPsdUdQxXpoNg29BL
tXjLzxsomvN1XsrlovULZ58gkkZLr7F79YTVbWqpSUNolvIgraINOOUicL40aEFpX/1mo9IA0JK5
fcyWGOeXiwVxmFWlp1Z7Xd33RZCo6wuj+tDjVzenlpYt31SjbsmtwkWDMjhQq5npWL7SyzeNFtUu
GPg8jaQxzUwE8xb7yElbUf4GTE8E5EDovv7SBnHLmqY/t1qbYeFPNuPbQX5Z8ZSl7gK0hSXOiq88
vZzFXSlQ1CmDwPdLwYXbcsnJhDDDD+9EpwASZdPGcRu8JLb6EBNkV5JLD2qGzjEJuLAu0r9WWEVn
0X8TH0pwfTZl2Z+KHhTOwlxGzEZJXJeIs0FMHKJ+xzyMmftfzmZoZtUb/kTGI9pDTOhioUwmxbr4
lrpHeVpmM4djj8NOCWeuL0Dfbo+AYw1Q+GMfCgUFITUSfSS/tBXEABjNqYZ7/3YA3DSHX3FS/hV8
Z2XzK+zHfTU4owu32vMtp3afHrov8/VBdr6BKq0aQMx1qMve3k72VQCbzOqGImG34T/pYOSihJtR
UxgoN8wOKj3BuCngqIWduOPb5Eitu1VQ80jbL4aq01q9vm2aO9VOpTeHA+Az2akehOyyOhTGVJ3M
01CyrTTrZOTpdk4cjCbDATC40NKxziGzyswKpr6WChv77sJ9GSodc91Labicb1ENXU6ki2+nwAsD
AP6me4prFK9SVNCq720bxiWHPQVGywhq0pl58nzNuSjgfhGPeR/rYWTMdyKpjntkhMATUx8K+y26
HWvwjdi48PupDamXjyhNzG7Ru36aFMVTbrHO1JhqkUkRemzJKWRPbG3v/J8kvUrqBYC9YCJ+mTdF
n9GyenISJIy1wHRYvfivHKhvCtd5HLo3xYodRQHg+URCivDMSd6laCGyZPZtLDDlHwTDYV73q0vf
0sOPzp5AyDCc5pxAR7MWuDtCdn3HcmJsUiY1/KSytnbZQY+7CG+ykXR3wVJEZrtwDPxKHQPzzVWP
HEHkBbO89Rd2N0Ar4/d1gzUKPPolhYMm3PjwVdmcxrRQF7QFWfiVqHK9E6u5PbgkZJGL0BE+t9V/
Ty33p/d2n/P4AwmgoGINbM+7LnsXRt1OwQtQcmo7REPxF1OEVbYxkllXz0U4Zi9io4d+COKWRTxc
uxCDLRgtcF3C/56YEU+8LVQiVqoKj32h7HFRjRl1GoJnvJGBeU2o5ZAIKbZ6QI3TrNuqLOMcG3Sx
J56/IMpxyJWvzvIB0DSA6VaW6mYfSMhvpOmmWC3qU0s1oDm7NY9K5F+b/xSHRwh09+DTXEVlYjj6
SGOr9wmPYRUG1upjQEVy2ssWsMm3rxdRPVks26IkgXw5RQpfyodw+R5sWJPTuV8rHHi76qdSY8vJ
+OaoqgddGutMNiSBl7BPmzTN9ArSDCH6aSYMuCE7BNMZYNFQeyHNfNNywuS4xyBcGJFHByqkejrl
X1jIyM4oWY8qlrj62nwnqCjWvL1Qrabl45W+Y5Yd6IEJ+UgAxbMmNQ4YHuYIkxewrrSdrk9Js0xs
uQMR4RCeJmh94SLknKW6/5Fe/ajp86i/fnm/ssLSwM14e/ggzSqvtZ6vVfqN/w8pvzZBI9lhnKXV
L7ZieUh2qc/rlKUaRLJk6kE0g2LiLsVzTr/mOzFWpE0rcmGnn6hBs8cfZ4fr+tDm+vqczDAw6f3C
QbJ3ad8fKWArfnNBvAhta9lsGavOvoqTPr65damO2ztH1ufdCVIRA7Q858lv1F0eB7cxNJdb4RPP
w8HBM2jEvqnIE0EBblxf/uBSSG6V6P5LxLg3xyC1LWNulMqGGcXVxtXkvLEtGbjs96ts1QulesBM
pf1yzIfIouAGcwescdqHeWPATopZGJgqQ+tTAHDqe93g90R5p4bF9UBFe2tBgavGg43RhLyL4tNL
7OxLFMb7W0zemnbnW/vmFsU41xjJHQy93MaDywLqD0SkcaK7i5YDVOXr42LfAEs6dxhktC9u25ZG
do/h3CF7BuYhrg/b7tzNio0heJI+5HceHwjn7Ejvw9caN2SAU85YEUnNyKJd13A/u7Osvp7fUKM5
fM7HIYpCp+xV7Y//bdfX6qGA/73dkILqoJJQ06VsfGfoxpXzfkFJBRgklKBJROVlux0F7Dn9dcgf
GdZGQLyLwmIY4cFQhfF/cY5t9r+5aSCuDcBRB87ODJQNw/AubsgxjIrBMhCbkTUh50hNmEl16aNU
3hqEK+kZ+9BMiO1P2paGx2QBQFud6QgBV8hGryQlSc2vlpDq//P5X+cNdezFf+dkrvcXKv8Pmx3O
jcyyROahQx3GcYbk700Jk4UDqOD4o+7RSjusJrsxdOP3txD5ejLxSUNXqZg0RaZid5sotTNXviT1
extCItV56stdGPT5asm9VPWPhvzrfaKU0H2cbQu7fdxRnXulAZP2yIAXLEafXUUEnSG2oZDAK9bJ
oYYZzo8hVen9dSMUWGBZcoccrpoP0hIUp2jY8w3mKvfEHh65XjBOBr3sL/FtqquhTN2q/gYAdQ+R
DK3cVU3LxdLP+mmzeT7LK+lI4KKdbgstBuZtk7QRfdNJFT8zkogt1Uek5N/9p6zYLPGKcma6JS6h
XjSnDhADreqWNRrFZCPmLsYeGSwyY3/wcZ+HHSoTraEhhr0OKdusLCOVSWcY10FsJt4vETdhIZg+
HGaNN8VZm/dqp3FoeVGWz7VYu3/Y+vuwFe16Az12GvdCElrFuJOEf7zQrBJUSpDJzESLtacrE4/J
plUewn5zbqWRiiADt+Co14CjgC04iA2J2mVMzfpZPLrIlbdQE8eQ2S6vCvWYjvRIqbuBeev2+hdY
7DoMMl+BvShi/2A9B2YfW+BwjA2ZyRoScLCS2jpy1799kpB5vCLREz9fVU5kwIuXCF2jyzoPq2LI
Coim9f57FZ7T8wZcjEaWN+3fexjZYe3K8OaeiJzfbYsSpKfF8nPV9o9/eMc8xB9YKo+/1L3IgiIj
ulpDNFvnIw/ugXqknMTZh0Fcx97sUVFUwXl/5n3thM88qp1Dm6+JsigYcRwK5vZusY5D9fvcAOa5
/vaT2szLOhomirAV4+7EQSBuf4zQPq2MOYa2uY9VHGuwLHy96HFmbaYGa/Q9/Or2GZN4QQWl8xYL
okKjxCHdfAXxgy61Z1exLTqdt4VwuBn1Zc/2U/RipV0+5Zc8ywNbqEKsWpw1Ddw8X3jIEMNSvs2T
nBMt1/LmtlCt0BKZH1fjAhQ+C8l4Apq2m8yaW2YTvfMMLD7Su5rHjzA71lWG+nglkiVF0FS+mYer
ko+QHMzD+qBCVGfbD9Ju+oleT0edndFp8c+RXuCalKnVSL9Hec0fJO6FvDSJFnoeV4pmOKpCsnyl
BrV9XlCMO8kfrC57Kl9SPcsugrIdklJG8Jn5u+V92s9ZCu2gViabUq0OTDljsDLW+jAfUw3dR5AE
bA16n7mVXHHYoeQ43olWunHpPfCfrXP4tHUio/JtYiqTkvMCGUvnl+LcUoFcWf/L7XP5Qg0vLnsX
/5Uhh1F7N6UTp4Dl4L6N6SSQrDuKnUnqGNEX23OgdDu8Hn63axUJHqXZ0Z/ZNzmvivoiTi+ZjOk5
YbABB6pFCJZcwrqQp3ONnPTYCKGSwH9MDHtMjc8L0F90OjBIGwrdjX8wbI6Cdkjoyo/OncsuIKkT
P2nzKwdkc2fLw5u96tmyS4NiQawsJYmmyP5U/YKWnS0jeF6oTXgIFRwxC9AlMH1QU+TsFKsvLUnu
nsAsvGVsUxleNrbMY77UQ5ovTQe345BhAQsiP5+I2aK59Y8F+/Xx/vZidTTLbxJkgtUn/ONn3OcV
fqipT9MSGiweWtiaNDNqjI79/EzhAJB2FOmBmNyzNuLFZ8VjFCJ4cTr5tJwPAvmCSs7o4hrQmIAr
KqmX//Rd0G0MVdQOiPnrT/d29X5XRz+Ms3ql+mz6GPbim8Geb0wiR8Qpf7R/vgDxyPYr1cCbWpEr
BeaFhWUQECgqP3t18HDUFPnuizUyL6iEFLutNXoS6Pjpxseu6TlSM2OCQ5ccZ7fR+H2EQ1xBV980
KzgJumElvpp/RNzu+y4NJtymyIwWwiukNRTc3wgX0EAKqhPdGSiHsnwvDUOp6edM9dDqOhBlx3kx
YqBSTIZaY1cag2tqLAp/Q3YA8uHrdGVCGktF/xKcF04DlHR6VqnuHRg3q9T+WSa6+1PSERyNNNlU
v5ZbrBWgA9btCGilxTdjUi5qQzMx8xI+OS0BbXPIhV6eIKfSYaKvOl3fJREytBswUaLbH2e5c9uN
RRoFciO+hajp/xvOlOeX244x/wXVrbTyN4sPL6m3z3hIm7+5q0DkJCjd+ev8R2YTSB3psWaQEALO
cr5SAqHeEMF6XS3A0Gmk0tV/Cyohsf6QLp2Aub130Fi/WQQO7eBlkeThl5XY9MnESf9RccFVn6Xe
mb1PZK3L+v/ZdUcj4nM8UOvh79744NjOy0VKE1pFAuYdxdId216oTa+syT9QLpJcve406tXGbiLv
BNukHpO0zQHNHSQJQjL6qm9ojtoLtvrOH0/ZTmnA1Zzj0wAh70JwuN2cqPlk1zkgVVFMf0OurFvi
aFwm1y6yVYYj5nGmHepbf043c6ZWkC4KiL1NgaoZa39f9KVQjeeYXXcyG7IeRanbpw4zF0WvDg6e
pP4Fjb9Tk8DbJXBoRrpQ3oU3tXY0Zic5jkUiVbcTAIn5L+XtJPsd5xgRleCRZl5ypOZBuD7o81sP
rcd7GQcR/45fsv+yRZB7sICQq+TLLiKZdzTK1aDsUCJ/I8DqKdErM8IplOWbnh/UfV/2exnVjvSH
1z8s9gyPApn5DK5ErO3utcYAyGMQYjnWcratkX/orLHzMasV+3wlx4BR3D2Z4VTERc1PCB25oYJO
ss6dI5Dm1lEGT8/EKmOd7ey45nwYijd36VLg+89UeywV44y6HP6mcwBtSAH5NkblILNyv9AHmEOl
5yt6OX4yzUObrZmzhVdQF/MweUWmuJHWBApiO2LF2b3Zi1JcB3uy8AlI5PUP3blPRfG88D5Ys/BV
xu5BXLhEXm4zTocC45E27jpggJIFKEaSwP3BqY4IHkeMBfahdG9pzhsWCpKbbBJE8bfH5o8O9x1m
qffXMXboozU1mCOPqQuMbBYVQSH9OtP5P3/64w4cIZzG6jpfVGQPWy01fEDblZvc5slQWiy4A+xo
pezRd+DquFr6mqOffrD8bNM9kLUgLxHgq85UeevHhqikD2uwN7W8Y6FqE6We02asbVpjGaJaDi2f
ufmsW/tWEB8jlPKNVVyktanLDgJ0JSwXCn+j234xC006IJvI1EuHo+ieWDt14v5fgki3+1gI3taY
PrieNS1610sWAYgR7IbRn5LIf7w/GpfnyQ/Psebzxpf5iWK36MB6nbGYOQp56p5bEdHasiOD0DB6
i9l82r11fZ2qcRpV6SH65Gv6eyZPBTC1TEe/It2Y+Vksjj7fZ0xdJAq7D7OkkmX9MnKtM57KkzfS
p0rHfFPWj3lxu6dRc8EdtB4oi6dDyyf2fSdyOWvOSy8vjwcwrbGNlVGy53DE3kPon010KXDaoOG3
kOYBL5szWqDbrowUTE7RomQXu+jqvnYPlc0rGv2bGW5wResbkJsZQdAcb9atpDsfG5Q6jGpukFgl
bw8FKTX4HAW+J5geuHeUTiJZWXxfEe6rvBTBjPE15JuenMbCPBdVX90ikaYdRDsJu6sBxBVh+B1g
xC+qK0q3AM8y06p06NOYnjAGULSK0iafpZllv7ZjEF9cCm36XVXImgzCr3pLYTl6p4eel7vg4Z9V
K9qeCfKSpNptrZFAOKhhlxFTfvZGxCrvM0wXW77l/rr/x19EuIDUp7V/Ufn7VJHTyaeEaxdAlfuz
mheexqL3GKeij5KvvVzHDCV31peWiGEijsOr2NCERBskg1MZZxJut1eCAw1BrOlmzsJPjhqslk53
jA0K92SQDUxsdQucd1hY0vCq3qOezCVRORNzCkXGprr5/bioGN0IeGl1PrDiMM0Z/Te4zCsoX50k
eztjoq8rXDRJE5n5l4X1bUYJXA8VVm05qifnAgnM8OGTZvRA83x8aaXXQjXQFf80wPTozcwbUGyv
KQeCJHL+SjHiRSP5fpUXBtv8+6MeqI+M2AilA/xo4h35/UDxfaCx08dAcHf64kn1h9A8LeexctL4
f9ai18YscTilvbMHK/DGOPPbGTaKnc4mHqS4xXvTOI8YTwmh2wB0VTBNhsOy0BLFeCzjXyXmUke4
zK+IJ8B2rC7zSSDIG2/brV4wZf0TXixg6Rjdf+mKMfBr6fCRXwrTvS+4KtWtZErmq1FkWcUN+De2
FSpNY8x36YVGgIyp/BbMKL3Z/nfwJ1XeDACpUO3wjX7hKzf2Ok8awg8EIs0czBsEXj2J22AVI58b
gwn4vL+mFpdJFwczTDyER4ftAoT9NF40LVIxoex2Ocq5kRvudoNw6waWjwDEcxFCPV8N02bchBLV
r2x+3Fch0UuQhFSKX6k38L/XMTg7uluBiqW7KpW8+eoODuIJRZMerW0ybQqk0cuuZgaRGg1OXLWt
rrwNbMhK+Q97JmHyt65Llld33gIMHDpP8rVOdqNm6+mkjv3mXT7Z3DfzhQo6lY1Q9/9RQkkD2xzC
wJGXYt9/+5/0q22ZtGw/nEmNkyaWdgiFNEsVfyBLGvLEzZGkxtPEHjVcB7ePtRhmmOBhwdEda/B/
4y3ECeRUBHNEebUS9VOPFzPk0iM3KAGZxL+LzEUinUa7NYnGIJGXC91GD0h9Ew69EApK4BiekeZm
3ArwKjeHDQSq0qDFqyIS0aEIZCm1fg/m6ETtsSHi7ciIf5H6SNuj/OFPh8tzpLlO6EdssQs4YVph
KeHnzGUuxFso4CWWQVq+pFIb2HPXLtiq8Whz1Qcr+XQlSCWiRpSZ4QT001a5lUAhQ+2Vd5GS72Sg
HvmxWdj4Mcwlc959EEHskL0DDOp6CRgl53uC6kJ/WcAxrP32a7rpEpR38mgiXwo6MbDZAv70jYzi
0q9rSfkXauHyP4/jgw//NelElEtEDRanZJ0ohYiChjwryCJWoOhj272E2arFn1L0mRexQqm6UPFu
GzmzJ+ik3/H+8v06Udur2Kc9Yhc47yeJFgM31MqO8rsjvPKyiPC8qhQrrsNSJ1bat6WiybHGGjPT
JBV8MaEVoas3S8AjzFnbJfN9CqIwJgY82jWO7YqfmOl4nKqUbRlC6euQWrVTaHfBK/UV4JtLHid2
dt0G9JPWMc2wPPSr+ZZk4H8ygPGiW5XSjAm96HwKUgC6wyoEmimHC5ggRiWr0x2IZm7qBmYtRflO
BVGH9XZPDkiNWDauR9Y/NUJHerVutXvmbwFRma4D7KUO4kee8ogbk0MXgF7bncguTVRZnJBV1N/H
XLMqAXdqxVyjy8tPQ/lQPsU6x9iR1IQpWX9wilzdx+21q9P9TLQf6pL2kaUJlUhiXvnqKAYh9BW6
mbdl5JfoeiVUSBhfdI+CwJeNLGhrVdKr7CoLuCckK13TZhsE27r96b4HXGRq4OiahbGjRN7+oli1
dQUNg9lPSEHDTuhxFKZK0yWhgJxtvSSBLDPhprc56ON+m0tj9mhSbeCZoF6bKsKR2mWaW71LuTWQ
W1FHNeYtPSSFBWSPo7B9X8zqqzU2hufjYmuzTL1HEIHk4Vnms/FWxqmsqHn6rdW7BJmE2yNFzRZy
IydPU/zCorvMCzGjk86u2gylrLZXA7NeQ3uy91C5B4yaKoHDOVlArZVfzOLS3d6uxQQdzLP0jtME
RqLSMB06VPsKapG64PcI5Bxzuo6XJrejaCYwKNRnAfEcMj7jhwmpFifUSaB7J0mX6eyHYkifQDPh
nwO5Jxpl5mJXNqKLfzRWDTb3XtS/xXKW58pmA8TkDaxmsByEGDMk7RvgcpOVKTHrBJ03jOXW956C
euVuD2Ud2nswt2LEEicppkHuPWN8zXciZzezejdmPI6YcvtVDRJPL4tY8VOx1LWbnRVh0I1utjHB
ZIaijWCONKAxfz2Q4+gtWt/TDbqhIVMoSzR3XO7lTaB+jp2LmzpCtW+R1edRsMtT8PKd7zsBCiEG
DjiqSlAoJJAn+7Xa5N3Bhrehgr+Rk8FDyMiTUp2Vm+V8Xkb9KliX3JyXP/ebVrT3GUYCW9DcjidM
BDX8mk+PlxQaIYExEjQ7jnQP15jKHJu56NJXqg1VigR/OI9oKf4ktcQHW7UvRSQWTu6olgtmmIxs
6cH4mYiiizwh2MzGTWu63UY1Htv0XldXD7Iq2DDY/zo/DB7kp0APE4ihlPzVRmoXdSvDZhKOwn78
5e28rW0Txw3LxWadbbhn4NuL3bQ8/+0ZaEU5s/Okr9x+tt7QvwwzG5sIDPDdZL0zlaq58GoU5xkj
2VU91xG0TOKoKFt52QafzC5jzLS02vwTYWATOaN12H6k2Up9b1fqbya9sypPwJYo1mXnfB+oYaI+
F6VV8v8gHvqCczWEn84Ou8bb8opbqnyul4Cc/VsaGsBXwtq3V3DxaQsLSj2XvsRDSY3h7gW4x8ce
xsp0BEntCgvw61nBcWPD9sMRViE6q2MTY7yDgIxUgxFv7Y8g5TOMVMrRGkERDoi6mgDbmuPTIVed
4bC7bAoZbUcS7/Kle7Rk+sYhL2D/3KhOWaW01rQzSReashY9ra42rmoRG4QGueO7JnC5yTKwscgY
EvCepBJVMV9LpmMT7cnKwO8pitIY+yV/RplZyxRaBOpJ71kCUDV+3IqkJE+FUm3GDJqOFg+L/r1+
ss9qAlFPefOiifOcKmH4RXqdJdaayQB6UrhZSGSKPWN51KwXd4VbpFtBnCSR8CYizpKIGlLAzPfN
S1ta43IZPAt80Ua13nw/4246e/PkV11/9Clh8weIDifm3GrRsY6L3+15pzMIIngB/qwb/e961cjg
t51atTrvHKpZ40MPiquVjRr/ARBXqzpKV0cgqFvVW+BYNhEed4IQsmi4QgxYLkpH0EaolvQqH1nl
W2Scue6E+MxVfxUCMesX2eTlUGs69WjeHnm5nXsqR/UvjUlkl8lMGMRzn6t6b4w+UMhnQ37blIWz
p1zLLOEli1kBFjJoVpQ7qO+nlPDYC2GyOtn9M9GzVpWXoU/ns/HzquC2q3pHkqQybbsbm/N06Q3i
79q7NephzaIlUE7qxF0XDr0TT/E4i45mNlnfgP45dYQQMC60knZd7kPWkyNPAEZLGO7XPFcjoLtm
tubF0ekmiZbjwPF8LK1wKJcIdWZwmeoDZwq3TwrOAUDTpJudmFB6vkci4L+YQ4qrk2ESNH+XyV6X
Segs+Czg0SORFVojjgh1LlBAV8UEK8qb8NfXXRhSYZ0wZsi9A7vuSru5K2Amtwb08xUAAgnvrozM
wMWIP7UuuoyaD+ZlvyhpXtgD1lFrb1YH3E4NWt2JIcZMPvReGshsDaP6IzNRx/wR14oYydvz4iQe
d9bmVoW3aQMNLoAbBum1OuqpX4MwChpBzuCpIEP+zX+lAdN7eZNe5qbFra2cC/keIWu2rJWQtSol
NFtpu303/eDJcdsJFOWhUQM04DpP7pZORsn8aCJC2Q80oaZ0Vq8W1VcB3bkrNfGXIuQzbo96hc1J
SWC97flufR3OA2CAVBuWBrEnFb8uwEuBoXyy5U2+T+qIIEKo9KZD+RbMoLs+ciciwAZZmry0w6J3
HPGeJL5PWvN8fyCt4vHjZbAX39yDknxW99/4svl5MJ7qZ92oH5aGJrgF0U5DvPS+JXAnwB6k2ds6
rrkuWARVPPurvGhCfbNeViNjRWDSW/nNf5XcRjuOwohg2mANeDmXUMjymzx+XZ2MBrIXBJSoLUga
gSlblcXtSB6L06/4PZd4FQDqKhDcBWpO09WjCy3Mju38z7eqyYiYFpjTcQs4k7TKoMl4Rm94dN6j
u/VP7NY38EfZiCviX2kXxLzoFF2vpEdj/puEuCjA+BPyaGBmR1tcFWQ1vmAO0Se3CHsacs5njJ2b
+iEEm0inf8PnKoAvYM6x2scMBFJu6YujtpgR0jkJfbIM1bqYUZslPvN0edx0XINaV2pxm376NfMU
cj6ViD7o3D2FWx8p+xQdxo1DZgSs4YKbOR3NDx8M0g6RKq9n8ewHyIEKFca7WOhU1xWY/oxAMXNr
IIoGBaI2lKWpte/aJU9agHPRv4PXujwAcbX2tU4/kW/SMcu9/XoZmIENKJBU+WEHeeYRfvvwxHjq
khcjJbyGwwseQbxBQnTIKhO+d1YJwmYvh/bp8uL/mpDOvQVeyyGUyY9eq+w7dhVCbT28gEmkGjkT
yFFCb1XIclN+MsxdCyVO53QhhUT833vCSDkf2iyJtqxPcNoXB77mFtHPLiHFVWkOTfw+SLvoyeDa
SAm0bnz4lEOnNroHQKYgk/9YPD90oue/O95NSLoPLH6qoIhi2Ualxc1be6Ol3ZGnB9xUu+VZ6s3g
SYy78g6H5VhvYVcjP3MfT8qjSR73qQHCIob1iinYHcLEU350Q9QF3GHtZnhl4qFZKlhM8mfTXPs7
XGSWIMuxvfcFHq6RoVfaTgj0nFhMPfu2Jo8lBJ/9Dbb9S3N9NhdEvzWtxDewyWQK0/bZI5M66/GY
FIVsT663z+We/dteDKPJb7FqgEun4Hn2M5wsqgtmjGWeSmXQstg5z4CQViB49dD9HtbB7xRLNnS3
toR0cXWvjKuxY4UWgKzp80fxEaMKzWm4tKBNPE9pPbv5EP5+py9AFR8nqRXdFwxwzlubvKLmkPRm
E30poMW9qZRLqO8DkWc+nI/3EmyvbRYoSkfnRGIeB4W6u0b6o6YfTeL9MoLIIwR9oetNZYJvkRTx
IEfbb9tNCRpdJzp/dRHV1hXbxRNI03kRUjDlSlMU6seelvvdpYBlk6EcL/itT5/BpbFsLtVFQLnO
12ae5+zf7vYMni/cSzdlexHh2qNDhFXn85LyBAo+AepG9YKsQV5iM7TTHDX1QJiSNs0fE18GR3st
pjwEWKz8aczLHFWDkX2i2NRlDwJKeo47ov6fesPrqVOvoq8v9qVqeX7a0CT31HjNi1IbfHmRk9DI
LhSXJ5bv4BBPgLlVfrEYsmC9cxSXCUaY0G1BJPW6llb17EeGlUm55g4+fi3MbUTySleS7Rd2fhpv
cnF5ceQLCnJfqpy/Q08knlIG6JRrwExWzH/WAiwTnRdNHFS7OjSNbFmaUP42p1mEvpdQYtKXUVEr
E+pKl1A7COCuS83Qimt2922AqwD6y1VTttHV7TyxtFlZXpce+rmHLo5j2GrA5cQ3RLwEnFrDDNhj
SwqN4SgUOtaxXa8quJfESsR8j+mps+UlSaehA4wc6um4v1S1z+cWlEkIJKvU84PL9ZDP7lt7IAF8
6/Na9DhGmvwwjGLP39ve1OKirIkFj1y57eGKKMsXfm6u64p50FFOXipcJ2mMiPjEdG/MoTpYk+UA
/DgPDnx/NTN9xVIEsvM54LbWCzAd7+ICANEEwyoiF8JeRQ2iCj0IxU4VO9AxmEzEEl9enLrhpH2Z
s063Iq5HhjOKJU+LPjCO9v5ud9Ss1L1YiknXY0X8vgfzPZoiqW8oKG9aNETGKRm50XAUakeUmpIF
PTYL7TyZRuiymX9VxaSk61hZJYPfCW+PxjrC5RLo901lEPJ9bifC3lsi8zMPbyznUsuMA9VJ+JKs
O6lbzxWHYJi/cLB0ZwOLDENaIF4QYQBpv0F/lObrPuIt8t/lOe39Z5QCSQN21ehAT4MyKt1LbJie
AalWVWL0218YNMlY3IJ+dqyS79xNDop7QZjRMFN2GDGrp8GQ7oXxbFvdnQsUOQv3PlCU086ONGgG
VjMCMAUdLHOcLqocx9ppMZi9zZzuTu6nl3zQupLejcCsKu2NG9ws4moC3gVuWS5gIa9fNmzUULlZ
tLnHs0P7bsfCoBekRYbkUp0qyWLFW8ISguD2ixm65qeJo++SIT7mbrfr58z6RT5Y/E2SZEpmj2RW
vYVOlfiyPX8WX/C9oYU/VX1st6vn58SiqZ7+DfbFJeEROUilgBGlYR4M0jw/cfwoXtqRQlLlMTSi
AwfpUh3DJ6hP8G8KUujmJBrFdz+tPzL1uAdPbyk6N7NTgP7LQEhqcgrdXV9rAfdfuE13TzNFUjyX
jUcV4F34HPLWVfy7PbGbzaeXAWB6XKZ1K/Og45pwSKiqwBgAWHC5MA6JlgAtc+W6cENKF4DMYmq1
F/I9jsF6WiUOqpJspmgTGGUOWAmicQIAI/PD8nuJI5bQLviOoEtAdRgXStZQwJXFs0/Z9yMYCK4P
prVcqwPlr6k7sBZFTl8lQ+7uKWHkhUfmalOZdTOXKFhX1Xt/nJ8zat4j4vuai6BafW/iGXPf0NG3
DOtO8DL+WT5tR7qYl4fuVjD9gwbmCSS3LOYQzE5MGS86BtH5XesWKw3h5hClAahI0BAWog49fTZw
m97Ae6vDp2sjkUfyyLw53x1XP7ofM/EQ7aisAGVmvqepHMniNdVn2MzXqFGo4+kSHjWJZ0gYsJ0e
g499P+TVsLWPs95YFcUXrb9JN5GuixMx/WdNzhrzWM/8JVoT8lc5WoPxpjtdMgKXJ07QLIbYFXsR
nj2eCRQhww3giI8F654Q1zPvtCYuolZkC42oq8npswv0vWRxGjDdgVlopCxmH3uclZRs65S3SE6x
fTD5atku4TachuTdg6tGbUbcLpQ5F+jKxgzFtk6B2JHa2Oankox7kPf1MIPvbt+qnujw/J44AXc7
RedsvrPu5unYtT2BPPCd6uC6qp4P+co3MIZyQy3NQolj6PgFPGLmZzSJ4FIJdLyEmheX7iHn3Ur/
gVn65YPxgabFcdBHuGtCYFj9TzpINRFVCtUQMAWo4iRhlDCvYTZl4KNAPlzGU74iAczStdd9gnUu
2WErrIS1G981jm99Fj4fexGNQGR9/4St5ROc1fmq36/ApWZZYMTcLds88QOMkvROThU36wfoZTdu
kGdkZVPwXhgOffQ0H5Q2VM3UNEGVNabA+3ln83Tnxp7sHoAOdBi2MV4Ub/bq7tBDwCyL5Z12DJka
A5+umePKugil9d1MBQosRZhm3iyVuP4+StmNQ6Zli79y3o4KyUb0YfOJVKZUF3/T0WHroV5N2QZL
FUZVI6gydUrcJ3u2/umcVun9msUuXMRv7yEx7cB685MWRzZgYAelWiPT30T/oWsn+Y+O4fPqafcE
8jZYMZyD+rhtgNUtX5EE2mbTHsDN5mb6VD/5vZDy6yUHxtlIwJCPFbue9a7m5JxZ6xNSnTQWrhvf
02T2nk0xgRpOj2Jb57IDwk98wiRiBi4ZSNrYv8D0bfuZ00l3PdB7KhgUTdsYeSrd6yhh7/CjHnjU
5tg1XUh7lTkx5licpVcfbG0XSmmwq2zt5YE1zyvmh/d91dcemgej45aUeRobt+nUgN05dYnySVh/
A6E9NgnTmhdn11oNzzlQFJx+aZjwm88emlCFnZ1j08984+bpiX8RbbDId6O2wQbJN6IZN+S9mCJy
mf/MKn0Bc33Im3btb5dbGZ3uRl+NgHydNtOfTcONIpga7faWUhNK3aoH0oNzPgQNoVThilOnE4KX
IxvgynPN0RZHofVao5/DEPpQdvooSvKRcTqB37FD9Q6Zvr030+1zsK/b2vPEtvILp43uAaNHP5d4
7L5js9q7S5Mau1vTr2z2l68ccfhZoYbz49hEjYWA8+rM/2/KS0AqSJYNPS5qmfy5lcDfJj2Y1q+D
WE9vaEB0s+fJ5u6JhhCQ0NAAnu57AIrzzJt6SjqRcrzzlHdI/jXh1MdqMf2j4GqoPA/b2dDSzWMG
VKkwZYqd54xa6nxRnGmbE+HTCxeaSfdQ1dbzck3nC9dvfrMjLsKbWv7UWgUuf62AuWd4JEJ/Luwc
UlVxAyxDoM85k1Qadw6tgzyBT+LylkmEQgeavRY+8u7ZKEEpme240kAo9QWWBKPp5/mOP1zTtwRB
KW5/le4jKs6qR1ju6rUqSGnwwRKmKA9MTkQeDaSVrnkSMRTVPmT6E1DO/IJu542cmCJ5igPcT071
svgNMZLCbagse2VmOcpsnS1uSZ1qQoHA3DsYhrLqJ9M+5AERHT1VAQnbZC7QT7gsQj0gDOg9lGya
2Sd6znDqG4EUw6Olp9XpIM/S2nnb4WAH0uDSe52jUbPcHApC/eL0QOKnlvln2fWS6zLw/qHHP3Sa
7FAQ1sTQ0Ij0vAhF3JCVPzbH+8S+bBpwck2K3QgzQ/VWf6IlSO+5vLCatPIs3QZUeBto0fF+wWrP
84PQeyDfbUNM1D5V/Nbz7MUK4i7B1MDL9tFsWj8+Cnrhuzq4TV+c8cmogz+P4BbNh/NcJr/Dw6eR
Bm835oausvCfOhRUfbCSUHHG8l6JF66oI4yRmZ2bhtSYrrajqshQZNa3EDNEsNy2+uEAGaElxu/S
lNHhHWhXFQkx2n9I4Jf22AO5+mzO27KHvqurTGar0yBbBRe9Ikpyo5fQwFtMiajfrwaXDV5XYEyV
qFEWaPqWVcA9lP0EZ/yrevZC21r06kxI8VIpy/QhZXcFh2XeC8DhmUAAbEvtI6VyUdCdTENy/kMu
ymifjKgjX0ONd525cjeTfnrw7Sr9KFsW/uY6suIW5mQ6pzCXiy93rb16Nz1pUywSE96PHGEt60Am
I3Wx9FvzI2u6wq8NxPhRe35FKrzACQ3tiWrykQzgobEk8hTCBIUxibxjRUZbnVV+AjM81FwSrZHP
rSjh9d0cMBfcAVh00xl5c0LbxhnMrjM+ra+a5LSOnQDu98Q2A4bfBmSpShI+DkZ7bdITEEx/2ASm
Eu/5ldGUPytiLTlhz8yDXb5OhjM19i5aE2O/Z+MnLSDUz39eljMBfXeJobnGM1aI06ZTA5DFqhBV
EHRxdngGamRxo5j1DNJz0myLyO+jxm/C/oYIQWIIVQDlr4nH/bH649BDO0kY0dLfKJtZ8wX7any/
uFMsGm5dbx/IDSXpf7/Or9XSLzADe06SiTq9FunBSDi+6vZ+FD7kB+yB8hMw0ZFkQf6/O5HTG44f
nPdP2UIQjCziSzqz5lQqGg5LVADSBklnVxJgAy4V6QBV/Xnt/dWkzo2EZ592F8rIU8kKepZQHT93
LWuB6eEhN/+cRMw1PwU1i29KL1gBWTc+4s4v2brTbSoYjOLUZMBTYQ9X2xGC/f5w3nAviQhvQx2G
AKyUwIJE2ymXmbVApD8u/NhFSsSRY+hcFVBsEIB++2CV4kR1C3GRWcve9QmXxU95PhFMYhVa9pR9
b/4hL2K7qHGnAHwPh6Fc6JRrqN8pOziUoplj7cdZ2KSeg/PjTsZESVWGnY1pZfU1dwMSJ9H7uJe6
CZ4/s49OImCtawwWUF9DgnEM8oQOyd/9o26nv9rcn+0m57PgHS1Vm76FONubjmi82PG1cNKv+/tM
Oozo3d4K1U3y+fMDCESs0shz/Kuee6yeQVVIqthoEnssgZZ3/EXS+FJma+036JylyhnI3O/adbJL
P+qIYGY5m7RKfPnmKaCx2AazcWRepcmOfDX+12Gljakylj1HGR4tzKWnqlS+BMB1KrQEkElgVozR
myIlPbEHjxtWElI99rNMTeuUFO6Grof/RiEHcmcvUe8trfV9L6gK2N7ZL7wKGI+IqUQBsGCdWAmC
8xswhQ+vqdnqP77nlO/ucYb2bEsdmwdflCrckQiGbWw98/iJXJdnvhP6g5/nE6SugBJGbfZcm0IV
a11gO9+A40e4z+qOO7YGYFwQdmtKF/Pk6ZA9doxWg8rIOIyR5Nkhm4d3xdfHQxkETS/L/0Kkbbj/
UOb9swK2pYzBAI3QJ2DMdrjvPAD8qoDl5KAOy9ZrtlerKIcTW4gX2slZm1F3vNcFCR6cIJwjF2Xz
sEz9LvuR59Pm96kmB7hD49Dmh4WimH4WzJ866NFCkaqByiS2eIa+EQ7SKc7Z1Eb/fYio6riahdT9
ogxCwlDkexsLuzCQQqtnbtUJ5dkTYfEty5QVlvX9cJL/JjjprTFUyT1+PrT1ElpRUH+5oFYhqE4R
tScMhJKcDssBSMDBAdrW1PKCh5qHt6pL99x9VBKEVBBKJ+laTnu0rePxRsehyK4f/LSd17cbj6fz
NnDm9gocA/79O8yilR/b0m2kvgwA4o2vsXDlmMQ1UhWCnJx5QQRTSS+E11YDRR9t2chHGW6heB+4
zU79yglYU9XBhlik69tynUZukglAxbMfeXwNjClJigegFZ2UldeNfxlyzUj/pepx0QZQcb8DhpV2
lQ5vutx9oAacIn2NDL9cB1GgLLwDdpUP33o/t7yRsLYIZTkQcx+srHcAygM/Yik4ciGWTdgIESy6
oUDzBQxH5aWccd0oCVM5nfb+HHSzaq12apgJ38vb1MEoxJeUR7m27cAco+IqwtLCDPenfzXfHI7e
fKwrI77h5lEjGwVWYcT7wZdV2oJfAQzxsH88XBtKJKGMcGO+d5Py4iPdNsq3Kj8/1a+0iHDAonQc
Gs/pgdZAnUl1PNBa/MaIW6cP9Vm77QtgpJ0GaLAYAPWh1ANkzS/rwlf8gpzUiY0MoM0Qzo3XKXRc
pC6YLl96Sldx1saVo+UnDI9xsL/q0x8PaXUQcPNPqurYsXglxesX5EyX9UW5fbv10coi5EGcLzb0
CFWOys7J//d/O2VI/vUcL0VDHxsGabjcI/h0M91w+qEorfPNlgwj9Veyy9RHn+wnjEw6uubi7AnM
vUdiCkpmBFBGMHcJWpbvO2PN9dE7XrUW8IHcBdROwlUNc7NVtLvks6IouuSIC+7eX+HOUESk4/5C
zRBCv7441qVwqoVm3bJxoRPVY/EASfmqgHW6JziGrpVKnJUScQMDcQjq/Cu3OVeTY0qXTLgVGmS4
Co6qE6BEXE43ZqMZNEpObPv6Q92yzO9TcbptyUQVM7MzLlWYNVWkhY14vKjIpjznxAgC1xh08Yrd
hxMbtKztq7PoP2wISRkEbYmK70UZ9yrVrFoJj+EQVQHFxxu+szh+GEZ/70g2z0jnSjP4q2VWiYDq
/KhGbSMuXrlGnskYdzYqxr49GXtsJz6vMErGOe/6AOFq6N9zsT10tk6efaO+xQESvSpJr9kuIJO/
CjoBd2oeq8VOYawducmtMa9jV5Nbaj8Us7IN7YagHN/YeHhKk0d1uyll5zX/JtVhGgm5bFD1uJ9r
qoydSFpXNV+i40VYtvSXtTEGPV/0bJTnIZWhlfA0pOxjwSu2ZepzYyv9S6REbWWjddP5AvHYGOk+
OBM5FzV6neT634S3qHuwLDd+U+FMkikXN7FFql73FhCHcirUklE+HvAnuU9XmERxlzqREluS2l0J
FT8Il5LoWJcaRvA3oi9vyipQCY0e62Dj+4FNW798nJ1fAIj4iM2KXpr7AYPaBZvXDDiW0p28QK7A
+/C2+ZI8RUuTQ4D8ThhmRyFWFShGBD5zcxNelJiabMpk3jqueDh71U/kwRsoRxTX0vImkFdoRV0j
6ElTDtxB+MTpAr3jfQqzk5a4UmrrgXPpsvbNqBq0woMV/U06dHwBx10Su3By0f2/91dW8b7XQKuk
uAdCI/l44R0gM/n3qguOf/tXfjhgtmjoL3MmUzQkzjQpHytlFXOYlYVZMnxlmqAio7+RUnmLV8ih
BIujB6+Fo5H0XOJrxtWvxOFUXp8WzBwX/99SX0kbbMbcdYsB0yr7bwzZ9mYUePE9bSV8uHU688QQ
pdU+f+tqjcRQaAtT8nqhATRAoulJuonKp1JfnFlapXa3XVpcysnYUXIZcw9D1j1D2HZXRTRknPwG
xX684DCNiLA+atqueiqch7Ozhnw8VMQ6G8Yh87ZGlR/wuoP1MvdfR4w8Y5rUuu3roz8Pz07GGMyC
JkztUGmpVFZAJO7A3SGXbUuZ52YQRRDtGkRW6KqXFrZos69wpO5gmVdJcqXjAwAM5P1KdkllUA/0
NuA550QxbZAMHnBHH0NFvr8/ggSTAW11noVUyVZJvfp1TGz3HZ8IE1V0lAcwKmBS2n3JNudiByxL
4gmq0Sdh64mrcTGdZiPxv0P/tx2Sqq4AuFFePjlcbJN2XrgPGkTupFyBfe1i2a+snwp01tmnJLVZ
faq+SmxxJwNb3l6CP6mXIUV220Kg3AGmoEQ84XDVz1mMjjt6TMTtIDLnKq/7s/R7gcVtK3Hvlr7j
D+4ek7h1hZU+jnrJmTbfkst7OgjvXkkYVy2zzddV7H1rN7FuMTNb7x0UHyWJKOkE9QsWMhKcMsQW
6naC45TeHmzq7kTPeAdDi4GtBIm7HFjGL7mZIOMGbV9Ktmi0G31smbEZ5AcDqPCR6REO6bf4DynM
RhhPdUPo/qkk3qMT9dilf5AJzQQf5ZP2oryom75LAtP1xKnr1Nbv46Y4MJEnvaobJQrtFAaiVeez
CD1/hbibFc073rkSTn0DQ/5eTxH5mu5sNvpTj3x/z9+iRjUcmYwSxmw+12dwNqwxmjLmnSPoKB3S
V5HmINtiHQ10o29Lf82b1n19NqdgGyIVb91Use8ETMGhyZttPZ21gJMOi9I/sRBnSm7HrFrtalO8
kCRUFwaypxb23JhtxJbUFhb/F5+waFl+Y7u1JeKM0HFd35xNIyCya2AxW/uvThuQc8tUzC46SZIH
gisrry54ns/j6jeg+AtCg9t5t44LwpPZfVwsIGxf3d4WlZ3Z7LRbn3ERphyO1v84lzlmKC6UP4MI
IYypHHtjSSeMqZzl8WgY0qCSqZ3HfVIRKE7li4oyxETTVSmnPOAWFxrujtRKDwDdsMUpXMlTLR/2
h+f0aYENiu5NtvbaHL8XdFDwlf8vrWFQ6nim8aagUiCxSosefuxKaW4QB2ORAXGPghDEHMl5WOM3
SxL5DgT5we9X6N+1P2bFpIq65ZcWoG2U9Z9Msq3zVSb8MULsDegyDumzufhrVB/p5GQRWfkQrx+F
x+XY5I0RexQE2yLujDHmbCwNlRkWCudSs4xsJeVDOu1WJH+0VUEttSuraoK7P9BZ3SUhyNd+/cA0
IEgN8PEe4TqXZdOvJbbzzrwrfGJQ5auFhdgQ+uH7m6jZ/pYoGW6jD3BlMc3P9q/Y3kptIkvMiQZ9
AgHIeN1T0rvnxhgXqSAaFRqVzywYs4dseVwqTKuUTsLlVKoosEtVhfu6RaXzZG5yQsGz5lUTGREx
KRoo/n2M6cdKsPRdyhvoxw2n4cCWAbxG7087AoCxCRPa2aGeWweEiBSkN76yBHhEq3oEtOujcR/C
9pT/b/LVgHwhQO2pI+NwFjVTB0wmqj5kTHKrqHXsCq77Gcww1o97ALn90LCDF/QbyiwRDXrdo9Pd
2UY/rUp5RE7wMLBSidl/ZuKis3KkRV2GJue0LJbykBiz+UNKg5cjkRBgwgOZxJFM+P/1MCgafczY
syyaDHxjBRw5hlWHaN8dqGdGtJS3h7HkB4aBPe+idzDw1oe1Df0KFabMZJN1PLgL8OX46K4iC4k5
HKHoyJOvY5R4OlvUMQmCDGZqlpATh7JGNyE9jOxSdubsF7XCwjIhnhKQXTACovn76ku60poIQgEK
xRO76wgcJtM4WAKJDPHB1r8G67yxJLrb6nUmHz1Ln4S6s183XU6uq2wYx1uBs1Qmqqo7hfWG8QHr
PAFA2nwigR7xSgTMphGSy6KvvJ9WY+A7KhH41/SZYjxRQ7cJHrxlTmlwJpDkLy/lbB+g5qxM+TlB
az8+N4dY8mwmCG/q+PWJJIr/B8apt9zr/1kzU6bu6n77Lq0E65bhq5OR5BroVpqoGbTOn1k4jrrF
FKu8wPkqL8AoJNjQNcgTNgqlu7QA+zOP4bxSgFz6MLm9ZG7a78s+8+LDig4lulhngtlW863YZgsq
qQ4M4D+lo4L4s5uv/h/ZHtN5Z18NWSGF9agUoXA655pUZRdGQMrU3uuaI+bUgsvEWu7b821hZzIE
qRzi4f4RmiAGzGXhPb5zHyRNjzIC6bnWdUy6hInxNcSsJXmeJBEMH8e8xGvez7j0cMGxZfjAfvQr
TtkD4lCNVmEvOB0pZkZuiWFe7BjjSF6zoC0sNJMiGkWa93mksjrwa6BB8Zu3scG0+ZH0kNsoz5GK
nbuNdtWK0icjQhmHNhc/qGlfP3EsoOY042q4oksEWZqfTigEbbcy7F3EZIOwgQzc39FGOEPTzHgo
xqT114Yf68QYEizTmQZgfgaGCRJkq50nLv48JkGIyNZ28OVEoAKtH9CL/w25Zagrw0V6Vny8EvbV
e4ndrsL401iYTXiH4+xs1EWKBvbQ0Bvti07mHG8yD8rK+v7iI4dVSZM5euAtPVHM0FtZGiHOFnRv
yH9yxpWpQpKn3SpWaxfyQKFfK+VcmOevDhvyXrg8wHgxH7rRF8o4S04d74L9DpYzXTNLxJQdfin/
G4CPWxhOqXaS3eZCPuRjzZSnpz5f10yUaf4uWR0Y7wLIec/irynpwxLZDdzjTGO2K5cT2HbEK5TC
VI9l3N8Bv1AXJC/rivCo+23n6CNLcKwLoc49HdeTetOM3ekTeIGQKHySy6ApzNR95KImeyvEbkNF
BCCgiDWvBi39jGfKNsKlDcySNMthxXvXML6Lv290Aw1I7Cd6ofdFIUMHFvIZ80PkrWi5mTz9nXQv
b72mwlPBfsKutcRn9lx4paPKhz2B0NZryYz+3I8qYaClJWHaNjvXymw06ThwSgtSD1Ih8R7PgzDf
d1a7O+aSRx8PSDOYfbAPSyD51joei3TRkhWbeJQTOSnvkWHyVW/35h2ch0I4ZT4M96qS46I65c/O
20FCCircbFAOwVvoHNip7v8AZGAhvPYhs5qGCaXszk1EPncAn8ZMnIRR6YSBkND8pGTMSuhn4zXo
ryijJMTNoMqXpXeSGCPy6vinal8dJC57kVDA+t/lW4DDp2wZbwlql/N40HYJHB61bPt77H06anXz
7KSnN1Xdwhfa7uBM/p1LljDl+XOzOv6Bc5pnqzaNuskRfBJOXtjBEaZaipk+4i5IGVwsCHubuodi
PLthrDbeolleRD6Tm9SMD8Te0Cc3pWgwUeKNHeYjJ5C0/hqgNekryhr1YTkhqhQJdju1+cQY7Pf9
ik9JCKjY0mRXj0Fx08i9kdrxW5a0ytNgI3Mrg55KV7m0pVMn/3hT4jw02EEZPhIVuhKhzKhVKu+Q
tzcHfAEO+rUUnzxuoPeNwVGquPlCQNAcLt2n8Gm1ZzWbLDNai8+5/VYcCh3z9okJdGHzLuDAtb0q
GYl1kf0mHF4NxzcW/w69HeWw8sV+r2nTrwqOzj+reKddQw4IrOTQ7qp6aU3KkIR34BZkbQ21866b
w+tZtFZaOhes/jMYbOlPhG1fK0CLLDpNUTdWV2XhIuPq3NtrmPVKJ7QMOEoWjGzWptWg7Ie4hOLB
FVwgpVwf39HOML1eoNzdEVkBeFeOpjEdypx6Cha3B6kT7eVUHlcskFdCUcA0eRJ3+Io4uxr87Dxw
UOfJq8MCZ8xdcwHPINoScd706irA9ztNPJBrEXyunFFBUX6HTeqqIHfzQfRNfcEsBwIrGGN+B1Mi
5DM6zrb2R3zMlN+O8F+M4hM1DTeSULWotAQFUckPA6ip5B2peHhDI3guDRKiY4kTVjcA8z0GRfpZ
9slS10f2JUl7gK+FYYbDmLp6Uc3nOFbL3vi0DztIp1Bvz3EUwIOAKHg9JHOkWhlcL3b0xiX7Dj91
Zk63F2XJtsm+M8+f4tlEA1KzRyncVutNYKANKGhX2p/0yMJKjOtho+N40agRB0oFZPqJ2tPBn8Gi
sU5CHPpq/s8yX61Ip4V/snWICwGZIuImYlkxvOYxhGmb9LN1xnoFXZdPo3FIlH0QvINQYvYAGnrq
CphSJ8E3gx8dAoebBbn6Lt7JJwKW6bdtUjwGtcN/3t2SOij8uTp8RSAt9VV8zfNVJBJ0UBYRmlzq
ghTgh4jhvhxPAZl8MxIfecsLDrX+Ig/zOo7IQ4Yw3wg5nDeQYQTE+LqNwgGUZEa1PfQ6olHv1hFR
NEYJwDON3WJnJOtT0R/Gq2vvMOsQ8G0Vn8hOfR2b0qV+AJ6ImSY1svATJKFhEoMaYUoZD4t1tBAF
K8qj27MMleJW+h18p9IM7h1Av53WdL7qfvCmG4Fd8CT+xn6gnEZCku1+MytCjeBJWBZ/K7iMJqCl
DXwkiK1wPkYZnqkM2MhbRoDFWePWyPluV7J7UTpowMGIKDk7MV1nC9m1zkHuIg7VECD1Ufr+lKwy
QeoZ+qWVgxbHS6jgkT9e+/bXHC2b8wmqZpnw+oHMJY+J5ikHUaw9eKT4WN1mmjxRAibDKyVheLWs
HxD/6f46/cBVxmv0ZD9KtxaiJd0DGubuP/xOz0kqb07fnt/w3PfIIGOv2ZHXvmn+FF/8FKI0qrWV
u61ImRhpQH7urhf5Y6RgkRFZSR0fx0/RHY94jb9g6reBrskei1aBkbwW1atMRtPKfoxF5DntKMCj
N4UAT7nRKYd6WW8x01++zXL+pH56gou7D9xxvLpzE4d2PLB22BzuzYghsFnAUJHaa8Ui2kDeHE0Q
+0nuDx8eDkGHHdYiqV5aZ5yQI1VZXr4OuWyASaz3q2wZ+Pcw0j6HURQV+J+7R3SwHji+anWAFmoB
NBLG22rPQYcX1dwnvDIWOC8lL2Bt6Om7oUeQG5NP1ze4zS8xTLDy9W2Abc03KUjz8NjNkSl1oPtd
hZ0JzpcP+sfe2S36KjzNYIIhO7OSvuCtqVU+Eq+Fwhmg2yNml80hQ5cYAfC5tB1j39njkwsi0Tpc
2ewX2p5WRi9Tj04mxA56L8qamOzaHqR4RbguEc3G4EOrLDd2DaEfJj8tl53uG8VfSArU/Dm/0EPP
n8CPg42Dd4hjrOH3D/5d1np9I67ggsk0NX3WSkgNudXRakWF9ECsmNUx1Zg811fnSo3bh6iCZXqd
SYjAKB/ZWN/IfYjS0n+u7M+HNUgnRttQTqHpMVNZ57Vlv8HnQV4XHg1eMj3732sowNdI0MPbo0ol
89BA8xekIrkbYtXKmQAYpVhIAF/uRvYlFu8qz/M2nK/Q4n0dJnIfDXd8hvCwcnwNZQhH4RcGb06I
UPFV5YJlH7YbWqw+4jLpVfGm2zUqKaYzHa8JQbHruExtbkz3ILS3tU66Fx7P8gAR9A01QWIF0jg2
CfqiXn4wYwV30FCNMP9ZoFWvn3Pkt/cqlag8pwml1jq4ipsnW5ObMSKtI6k3tWKA8UOEqqw9Qm1L
wxqFKG68gtP9nvg1RBAJYWrc2g/8pqwkYGYAKCQp095YMUjSxedLB/hrFjRkDdwRrX83IPPXj+Nq
kMKjkSGSaSPIQ55uv4TE41CdBDHn5oTKcOyshR5dUv6dnQsG8PBPO194sIrKlz3uLniobwOlG4QG
oLUYhMONhjSvA1cVn8FcITuvLKIEmIj6JWIdzFYfRuYvJXtBfdhLy3Cw7VHo8byjMFH/nHpnkKap
GfvlDVf+UEBwOgjgTYuUZ9r/t8HlEqd2vWzOdwPGuxbaC0Iz8vO5wBZ1UGHTLaQJFjP+glWkZtrE
/6tRxBiUoI7DkYYm73WGR+DYfEqXblfr/IS9IkUevYSAF7kKCpNwuVu7XDRkqmSPoV+a2EEBbmDT
KGMRrF89khBvAE9z225K/xFUpPrlL/kumjIKpesZs6X3/3Sep/7lidxjN+jgYnz7e3sfQxQ3+l/F
3TBVhp0dflE064yIPtIl50U5Ityiu7FQETJXvIDySI3mkvDXx+DGVQLQgnR2rwFRv8cqg502j+gc
UV6VkFF1aS2mnfZbOLm21JEnJ035dhsCefKvOdutHESi4X+kzeKaDgdTc/iIvWsSr9G8Coao9tCn
Oifz+h2/CsspVW3KrE3XgU1yLrDw2jUQMEDqOYTvDXcd4CSctsxQAMWrBq3Y1aXDzQB90vSbXNQa
ahVX3JyC169JfBDWHUmdLDrrk/D1/BxXG4/uiAGIwbyDcgE3DmuLGJHIVThHirp+dldxiQ+GYG2s
mybt9yMOrej/+kerikiw/fQQZsTF5rK/JHNSmwuqf83yyRTiRjnXk61PauaY0lWJR+IQLMHo4m/G
qLEA23FZPwyX6EK/fBIkdEHNTekIId3dtTEFVRHUp8az/jQRqFyWPo4jkFtkniGnLn5xHCJU0Odn
48Y9UjNUIQDQXRjGm0Bl+RqqUcu3YDcppdM5lcyBwLjso3Lgtk+8oPwRLP6ScqorUA0mwl8PVvDO
8oO4m6c3DDRkUlhMWZuGPS9mYznuPYjedpLLk1rhrR9Q6ykMStGyc35FpNaW9K8sbgVehQM/r/3a
45qmmsWaUFPTKx9EIEAr1XH/gx0myJ1BeP1n2pfUXriOITvt3g2t/H69Msl/flGaHlY5GJdZUxmH
Sb6kBKtEN7WyXNXBw3pOJy2dOS46gJG1xrX+GFexh87rRuIAXBpCkFBO8rMEzMq+EqtPyU62gWqZ
V6iJTQNKFbBJoiYO2eWI3AkQ8AvWrgPN+qH7JgdlAsbyEKhnJ7im+tfsN9ZH6pQvtm2JZ85O74Ab
EpOXA0AGTfzYf+YB50KVvLuwMxBT9Rh194qrAdmEhyA1h05NSm2wtXEC0W+y/t3xbSbk6/Y7GCno
W2UgZX3shijLZGjcPPAfMUgYa/BIA+xsHv7TJZVUsvrzlUjoaZPk5mmxmnrAN8HVfgE0iZI9OSn4
2KXtfj4pLtn0nMVJx3DSWKwkBg/tiip1FnGbvg2t3IUup6ccfGi5GgKZWjfXpBARF0Wu3o/wyIUN
ROac6hyJRR2kEopUMSJy5yKmu4zqgOeAcz5VKZ5tw4W/+a+hzccDur9zVgCFniy9WybcA+ufRuF4
I7zid6wixHVYbu3WB1GqN3KOFcTPsWFETLHcEfRw1nmS7e8NaTYEBtWXmEcbPzDASh8GoRL8LKeG
tF+9msseTZvRENAONJQxEV72ta3O7zKdGkX6tH+cTs9Xlxvg/uhZftr5nym5QXw4Ywp2RPvkXzFN
FacqXSRhdEZ07xyz2xINDPUu7kntfiJ0YIsDqiRIAW1HEIjlXJ2VdLa9XElV19yPK2+/wknXaNh2
sHy5JFm0nknU+pVTWuoQ76k2lYwlOuQACO2ubSbqDyV+3N0+FeaZuCHpNglC8EvTrg2iQDx+4Y87
6zYh+moN7omCwrbUHwEYRiN3c8cgRzPs14kebA6VHHgTYbW85GdZ/YVdCoHuHQj9n7VYfMpx1NJk
PIkJ8YynOESREATyPt7PPMICiWFUwpecqoEw0aXNaCcNkR7EjKZ++PbqbWppPvgPftVrSdhITypQ
Cdd4Zf6jD38YScYbTD1L5LfM5S720pV9i2ri+ekfFKnLXZSY0WN2Z1O8PQ7NQhNcbS59XvLU7YGf
7xMmSM3zP8JfepG0A4YPb8RWc04Pn3i1YIpVC+l6+DdW3Zjmz3eegnqTkoQ+eUyWgHQ4B91H5eTh
KwWXN/UnHoCKdaGaolmXvJWiuSFrVrvumy1xI18xjbR5bjpYprMH6u75OqJ0FvnYtnwfa6x4vXOp
KUSmsgwtED/g4EfzuxrOnA2eSil5o/zRntHpDxuXBhoLn9KFKui2unuzJPMRoXaEmSuOhKOZkZoi
PWfFpzAvPBtjTRd7S0QvnHVxDtNZbGH9pQTv2mF0p0JMLSv4pkfzB2PItZKfSig/i3EH8mTmUtME
Pu2+gJj52Py98owep8tnMKr2L2iJGQoNGYl1rzD18Oy1+bPuLDlkAyYs+6rrbQJ5BCg4f391ga6Q
QsVa1nAAnFEUqSXCBYwaq4Pb0QFy+86+ywoqMXa7kGZk3qGFMr+YQGouu+m2hlv6mK5T46kuBk82
WAbQH7UG1MnjeibQIvDzG2P2aVgGklQyqNYQumXhQ9aD1odepZZmHcEcDCki0j47oHUE7Hl0LFj2
TSJNEKII/+/bAu3VhYaLThzMsPXYwBKFGxq3IZo6k/A3RiNcgVGidtwcYA2SyvqVBnfv55TSsMrw
JydhP9Q8mZy44ZKkqchO7tPibumSNvm+kKuRvcDVsQb2KYaVvKCI/A8pM1Oi42ROYB/ECMQgOD2+
GWr7hjRV+2w76KFV2x85UkHAfV823qrUuMx7m5p37A0Tvqojf/fUje7HSWcihDyd4RV/141IwTQf
JgpcG5nROVA+NvchO7GVN2lW5ZyKcGEf8ZKKhiXpxRVP0VgpHKdTpnW70VLI42K1XmsR3/z+9HFk
5X3CwU8aK9EUmIjXQaRMZIs2I2QnN0HqnA/dCOyQ8Lwig3vM3RAq1hOwn2G3a5+Vkaai0xufIUNP
6NAuhtU8Ogfi9GZle0PXuqEqZ+FMvhWCBLhQGae0Tzpe9QlHDtQYcGx/w0H/YlX1aGn5l5eyo5wa
+xQ+9/DsTHv2CgVnM9fwW9Z/NvkUktlJRMkVO0TFWmkRAXDORyDqyHAq9ucGAbj83n4gdV08ams/
XO5LnmJlER/Nk+0azfZpIkX9Kfzfp3PI7p5OY53j5Kzl1doIn/e/TFAaq5gTXBeIvajbcf9pAqgq
L3t9vXhIsbJBoYrCkHGPS5j6R5yfZL7QT4oesuAiVrrmpZGvvRXbdczNQOkC7kd5MItGYDFRUbrv
y3YQxrwln+cBNVNMxq/8z16lS4g7KNkUmUNw499sXx8YMo2tMAkitbuy8pXffqqrSgNAsoR1qEBI
W1Pyj0y2j/xR79AQaiZm0cnS4LCCzNDPhWq5or7E4JPfSQI02SiOpaDkuA9lWfGjkvlLXHLAYKdt
/BqAuGV+ApMCWFTo4d4bYX5golgUdAnpn3nsMV5iar+y3JGLMvfRW+kZuBuyA57gg0KNLdCIBjL2
kW3ghMCqIrkkBknAJYL/cICR4/qzpboi/bJh1+QlpVWGBK5ikul5I409C8AE7GVDtRJ8K9aE3YL6
p/eD91DgzG+FxLxysCEBCCi+5KI3n0jbYmc8FY/0a3dbJmeGVaMVpDEe6UrXHVbPUYzxTL0pZceD
ocpdZRnHBM7FrRdVvcBokZiL3QXzWvy/cXM9CgaZjQFMcyPDd6hNYsCCibSphD6zNqldYYhqKpH0
wh/361IYkBKFbb9n74+cOHZx/12uZKrEX1+Now1STbwlCpdoSYEbCuvtwhVYUJ3RQvsH2UVyW6DK
VFVhKbIm78Jo/UkVDOdcn18CqyGQnlkqFfrqdki7IHmddmnbFtqdx3+WE7cUX7j/zmvbe5mlmstx
SGrlzKQNUc8G6EquvIhDzCltEKeXae1MOos+ISvDioRZDpr/JUKe9IaSNPpL3sDWtvOF5mXEkHB3
oO2O46sr1cKs4WyUZDmtj3QyVRPOiL75siwHvhr+3ij0hFtiEdh4m/n56gSspdGqLyADHJOWi/QP
xwQv0v3DgjkRmFmHamofDCfyASgfU8yjtY2CmDcbS7SFcWKw/r4IIdykheRK8NCuS7A915fiQxKu
ku5s+gUbWmWjzhAEb5nlYC85Bd4Udm6CZMX6+GEqhuQ15uo5CB0zlfcFuqtrI2LNNDUSiHmBgC+S
GeF5jLj3ed02u3J7VhhSqGqR7jXYdAFRSxOIDi5VUgzJER10/kjyCJr0aGqzzhvoBB/9r9zqcZOJ
jT6UMAic87SiYehPFtknEHo76d6WSGHhuB4H0UqejwKfoNgY+rQz0wJxU9B8maC6mvMGMQVauAJ4
nadOxN7TQSTCsg5B/8sHmhjdSgO/d/g9A5jMoZjQAu2pUc5NFGj7q2w5aAjyahNu4k6aM51xJVu+
npe5lu3pWhnG+Fh1sbdslbPkNir6RuWCD9bXH8GGhTW3uJB2XScgPyK0CQEL1kaGn50MEJE0DYJD
lejfVrm1uJX724FJng+/Stxx0NX3Ge4Ou1NcjcfkHZr0iw191lf1lp4WNuUiKoWrotHFBhllSkvp
MH1YbSsK3v/TMkkGmeJ+oKq80TofEq7OGCiZeLXAMRZUNJpzystb5zOeTlCpUMKQDv+O9heyivZi
K/oUIaZMvNnNUOcZrS0Xsa8Fe7gNIhh7pKYP3Ed1RFOFPIs7/YsXOuft5+KE23RyYMUHGl+eUzsY
auHJ7H8VaPTh+kIhCorGgAw28P83zRCzRubWtsb+PnrL5YvAhOyNsWHbgwj5P3lsfJoxIyB4YMkb
WhRPSx8GpY13fqidBjG91KpbniAsieWOh2krqIGHRr7mWFv8c6Mjp1fjh2qJDFM/Hq0V8plQ9XNa
YF//9d9xATWvu2X8ABGk6SLlInZS/WylbWQ7kaQrAzQypd/4AhJZ4M6yniJ5fjbGE2Jj4FC2Uuq8
7PlFlgYzr3emAtyZN8rBF7PU3HLWwi2K/vlL1OWeX3XXKAeXaPG5D18AQvT6+BfAT/5exMZP9i64
thhpVQ7W7O+0LIXINGW9Mv0VppWuZ6TwlzH4KRj8gZx9GFatGNiJQi2uGxv7ftzPSauk3QzcaTIl
Ln7excqywFtnIVUOp+h6ZXGCvAFfEULvGSObuJiFs6jm2VyUNLn62IFJ1Z4b45IhF8/3nEKqFsh2
ZK+QCvXhHA630hvgEy/oSWVg6+Fl4enLlGUl9L4vFT3Qft9mtdG0KlEHDR6OHEfpOuYT1qR4KpSQ
hx0ChXj36HHBUEl87Vsfs/iSO4WRtIi5UV8KDOfQYefC1n1CrEkdfzXvXyTwdz2ruf4DwvKMfw/f
Skd3WZRPCoTulki7nAKyhc2TWp+/tbeiGT+gDloxd9H8HLR1wqLoKZX74K275mj6V5GYmRPe8yt4
qED/LA9In6p8Epa8ntE+OSa/l6J4irw7VMuQCGdduzn4/yU0R0UCpRZq1FSPrTVqsZkb4R2njsnc
nXC3KGaWd1xjqRt1rF7h1g3Xj5cSglqkXm26ygV6XMtFDMC3zbv4PIhKgyu6GmXsiJp7E58AGLSb
PaMDZA+beWX+g4NDKyHgcmSSqCpjb+ls3m+xVGVX/wZewCgkSqmHh+uek9biO6IHnkWBD6/HZ6UO
4aKQnBWVuex6t+5ZGEk9kLqDrrk8cqCC3Ls/vjNr5yhnGHnh9+FvkO6Dcj/XyC+PSdWJ1dyteQHY
F/43BnlNLaO3TWfWtjdHlKb4yq/2tyhyu9rR2GritoVO9dUXPfYLPa8gvL5oEIWv3UKgB61G61XW
hyDNvGoBjS55vFsNq+TDJMSw1/sTXxoQLq4pYBYYvUj87Q8SZ622xRdZLrG1wnjGo4WJkaw/rHgk
Q+l4hyQt7Qvh2uuWB5YjX1pZHS3J6bRwUetSx4+nGV4AoggWXERX0CYPVV9xglRFiwW3PpJZovRA
BJ0/0+lR6TG4xmAAzRIaB/HsE98p3j+k8HSvn/3dCiu76bgqWNiePo/TRBx5rZOM2CrCJKYpGYaN
OC5u3l3/IGJQ2a1Zq9UvfwCFF3ViXNlLZU8i+fudvqfbJwX2RqG7ffAFBURQjWzvZH5ZEErQM5Gt
WzeO2Chx31vAmLF0X3PASM8qm8ocLGdtYYVlb4PcO1TMavYndmKSYzVCOEIx0tbMSVrfcx8Rzoz0
WOfVWLE/2uNCOq1QClLZflxpM0uy1u2Tcm42D7fvb/aJH3wzh7WbkfujT8jQG3SQFem5tEW6/4w/
UUQeS0Rf5KOMmJoBcqqYz41pAhnLIx04Xso+EK/7e2pcXtgoQWMFVTd+RbkVoBeMYmhBTmiE0VsH
/tvkaqoFYtoXNklG/ZrqHGtNk+ZNmyW3S7ESf23X+0NfMEcGVimK80WsPw7jLk3b94aJFdcVjhvC
Gh6hM4UaCNm6o4FwZYLkTNXub1pD2TN5fbETprj/KEw8zIrAPn3/OFkhTSf7JwTuuj6QeITx0WSx
Kpz9lNP5fTrSyBst/sP9qusWMlpjGlfPwKENyoa/ut6ok5rHsffJS69k2vX4QfPLlGIJNFkoRXNl
99v/HbvOPxSnL1QhHsKe0I8mTa101SsZfqIc5OdcLZH7hA6EIBeq6Q8/ruBR+or6g9BmFcHIjUgZ
7hfWOIlgujFlj2rIpV2tsDXeWEoAqBueyi0uKgEd9ZuytZ9qe7ULCfCrvHHKP9WgVDozxSprGKuv
bHSbictBIsAIpmX60ArLI4/xlZxDc23QaWqJU473uYvgSxqFzj6yGCjSMtY+pe1hqXwVix2j0shT
TBbaDwR5oko9dIS0rcz3folN7ZvYo0ku7m/cFZ2dRf7vqG0peojj4fgAQ6f6dwfj6oJskBbV31L8
0L5HjksoY+raIJo1gqSe8hXkMka1g90B2ZHCG131/dQVLcaMoBpH5wYa9glOnjtQ122RTahkxFld
GzSlYSZAKYnp4F/BV0xsz2xdsv1endEMgyl5IR6wWK3Fg7X4wijzkL1CIJJzY6EnaVJfDzr/TQ0b
eSV1gYdIiiIH5yAOYqUl4VBNGG18F9wltoKRWY12vZ5PfrJw4QX4isa8fg0CynDj7ALnOaqJaCJD
6vlTjby/CLSJdKsbeNSdjg1Dm4mUVUs26mkovW8sTBciGr9mPLl8f20NfbnhTx4ZEzsH2VUMIP0l
N4uyH6mBmoxJPjjBhJixYU4/Bl4X39+XJ+/osGQidbJ8ZM3x3eorUy0cjhE8fH3wVBe3P576Q/I3
NqK3MqN4a+hYNSSjHAmcqcbnrcBNORKieLOOuzeOCqFWGDHGtsCgdAKYYgH48vrF20jVO8vmsNIk
sdKLRaBMOCUze4GD2nY7og81dO8XjKF7xqtfNcprtLWhzfQmwjQgi96+XklaYlNQ1fBU9SIq5vwA
ncRqaWcqKWYQj68IyDuqfOuN6k2/7LRLMFWEcZsImLVvJBGXL0RZG1FJDWmwHXvBfWS9A50lLbyM
TLMjE+/ms6FE8aWRBeKP7aJ/DY89RsR8MewOPQ2srFMEruzWguOqDEDaCiBZ2gIlhawjnIGxzHpR
ODnK64+b+3erwyh0fau2clioS672uYx81hpCjbQGYh/PzYN+X7ejW2d6IGbKyLSUq3yhiYxmVXTC
WBbcfk4ilUOUyk4qE6ZHZuzMzNn6B/D/nfOS6Frkuj2H0dnx8eqTgSTIuWUdNpVMX3g+cjikKQ8T
3aGrDNVjHXJp6xLfKydc+EKJVnRsoMvhef5xXzUoJPduIPljfFY5IG7EXCj+WAZOKDB1XvXgTGBf
HAioDvygo1VEpu9THwZEsz+rpLYZPoZLrIbZllp/FmCVziYXL4y8NSBgcBg8H7qIGyfT6CN6+wSx
qzx2Ww4L5pZ0czEMs3iuJQAYjd7iduqG4ZQMUKhS+J/gKxeKjIRzQ5jfl4718G5iPdp5xaRe8Bir
hDLKyXdQAQomeDPolt3c2hQrGeXRO97L+abvD8GgSpWoipzOa3L3XjmgJsaN8DESGc/n0ipLJXy8
LfQm9VBAWgE4VD8XGwmR95Cz2AfXbKf1HBgDo+UuYzY53v22g39SnF3gOYfkMYBTZVf1BkyNNGaQ
4kU4DoIL1mApdbRO5C2TX6M75zxm2O73ILhEAas5C42i/ddF9Z4LPXwGLMFV9dSClNSeqbABJKdO
yZ4Pn+sVpva4/Gwoa9jAFw0HS8xmYXC2lII/uAi3qTXfeK//qAwlS21IM1wpZZaU7VYQgglJV1fJ
WyDKYRE7pKcolMSEl7M161kDfQozLh11USrJDgAwPGM6yBxifl5ATWwVaz6om/7G/o/0PgsErMuq
vOoVIFiVwkt/lz3ajz/rdZAALaIyzkFpLPZjnyVc3zCFAOCRqn3FppK2EtHsh+g42nTH8J/Ji6fN
rZHKqSbqzFKf1M0Y7EvQbaKLV4MJadEO1ejV8Zz/f36nu6VzVao4w5x7/byOLMm09YhSHvTrn5W+
dtacdm2HkGgDlURv92BEP5EUctLnXdUL3zNB3NsRv28pBxGGgOFHIJlxTpfNY47YUicO9rBxK5Cr
6Uo6ytadW/4izh86nX1lVzyqpvKtoc8RN6i2iW/tg/vQaMRenyEasnI1YvBYkKxFwh9sWIQY5YKe
S1Y7lS3MNRcljQKC/brX2E5xTbZ4qiR2ez77D7+47yHy1XWxD/NEh+uE1SSrm3Wo++k5pfWkp52b
y/bYChv7IawoosOSgpV9BIEH2G94v/Ub3GSg8tdGCvWQqdN7zDEMo+KKGf2nWrbgAaXyIGvuKDV2
byZUgg5oZNNXT2PWC1gCdbVnMQEk6vnI4R8Ql3Sb+CgR9EexKafpcrUa+CwcCA4ZhajFVM/eFe7q
mY7ayvRvxr3PrlwE1E2xgtiD6y+PMMDiy4XYGdCyFjHTLMnq5P7UGEWhpqVs05Z1KUL2ECWk/Q5U
mXUGyANLiQ7OfE5SJ22OMov6H5cUUsrzGH4SIW8KeGFgaNQZEprnZKLptHiPmLef9IDUuoRywQK8
omzoppgsPX4PJmV184zgZ5660FhJVs9R7LKOcoEiBNhTramG/Uwi63kX1BBfJ+eFl4FDEqzoOQnr
Dk+Z0YT4Q4JPSDcTMx6Wi4SswWcay9aQaRaIbosF7TNqrIAiROrkLwG4SeW57TTfp7gAvr73HY1K
RuzTMPdxLIlMMvAltWfhUQ6ixfF+rU2jMUwkn2rQyhXlRtkxb06g08o4Bh0bJfBv7nZu3RDojTbU
733rb6/WU8FLfJzDTEgVOSeiwxi9gmhmaSGinQG9saNTy/MCutEAxvgShtlQ8x7f/PtPfbatxwPP
6SOQuTrW8DEQckRncEtD4pNNXzXrcoBF+sruGalZ2zjTgKKWvcnc/kODt0190P5jYjTfz5/Ft9qO
R71VFMbTuuk9Dz3myBr3PE2ZFODyUMMYSy99pJwWGYEDXKnZuxiTrpG67XzybRskpT+dIAfo50eh
ZXBJIcLQo/gfiH7xtw8nAml8dfd/J0yVjQ61kiDiXnukxBDuUzpCMmI4JPgwS4QawdnSzI3t54b8
xa5bTdP7tRJ+1L0YMGGBebqhg6TTNXQbXCM1fIfSdSgTKAeREIomahypjXIQtEMvnkR/180hKyh3
cCJgb1UfOaCKYYKG4Ba5e0OkeN7loQAIW9TsBy45exGicbiskGgQGqsGpqW2DRf5cqDdvIOLL7Ny
eMEkLIPs25Ugx6ynp6Sgioq1A6fyUjA5G3/rRmEMUnXxd07uAgosDqzDFKFwAOWCPSb/KGGy33pf
yEQgDkUEjcVZqfkpVV8T0NFzCBABcmgvnILeMrPHgFev9cTovG8jFWc/5exYV8Qv83mApTmxjKiC
Jf7m1atSfDyIV69sYqlbYgvlBAw0YF4wAdJCc9woso3IxVBvqoBsRuti5HrRRTR+R1AT5RIOzQtV
CSD0ve4cvehva2KQ8/PSBxR492Wtv10U4h3Kje6yRi8PQtSmAj9wRY7VJJbYzUPtkSiQCt6OyJpR
tuGw4AoRT+hLMVHBepuxc9jsv10KtuBlmwSGbm3lTQ1fUY23LLU1nDoNuRnRre9OqHcC9h1ri9Sc
iSlEW5XwbFNuozt+nIivXUfPbc7qU7V2r/1wv3Z0dJrLaS8RACOd6//lBQK8oVz1RRcxfkDIkcoR
MXwYzbYEIkYf/AivgaKg0B7Zx1Zq0roKXYJJsvtBIMzt0NUYy5srhsu7zIgyczE4nAMNaqWjCQ/3
jgHq5blJ1/0VqYBNOzrTNCE1JyJlGb6QNXDlspbTKkCoGwfGPi0VIAdv/ogG66i9mKFzrmW5LDSk
aPl1uhUfKbtgy5KGD3PZLGLPZCU8YPcRMZ7IqaQajR8K/J4HsCl5phYnQ4+BKQ0csq2n1ALWEENj
5wcKZPmIvHFUhKkzNVzuBLEKdpVJoSMP9JSZxkQNEkWU+ZafTuSMvLNYuDx0Js1XS/8cm2Jaa0r1
WJYy2lg7m22BLWtuRn/KjVQObm/yWtTawVJ9MPIMDitGQPn32O7fT8D9I3Rm0L1mzOiD40nXqP1S
M9GtLkKWm/ZLv1F7UjUBr0dHfQ4CJuU9IVXID7AcLMcGvwyWtfkIvnkmK0cbz/pvq/ZJpJcEh0QN
TDaTe0MENckFN9q6DnynniwkHVBUnfI5af6F5Ot15Sk+W6FW/WP2nsNfBf4RdxIrLTf3hNFrRm5f
m8F1U4xXwQSO356NGE1GpN8gtY8H0IfMCE3YQYoYEBtSO6tnWzarIYj8Pfb0TiY+tIDd2N2WXUZE
TJXwhSJ/auUkc2ZxbhwJ/GNy9EiyOwEZ5SgSCBgtUXwro7qkPmwnMX8iMp6MRSd7DL+mdAYU01Q5
429Ebkpfdjfr34bAkFxF+pUQtce2flqx5QETv8MX8WO1QwOu+QoILPKpjPIZ7i98UrxDInhtncaB
oYZVdh4VDGALSTy8BpLw6w0dKzccpZE6xZPhJiHgZg72Y63HEUVvmm9+PcVx7gr7rmm36UBaxxwZ
fTaUVFiQbJioxfPd4H+DOl1+nCbqFPLK/YqM8nYiLiZLmNIsPCeaWuXSKfn0xawY88FYPGa/sphW
gSsAVV5smQ1T3WMYDtldQhgzk2x6PXEC9SeL3twkzf+smZjnoiCa2u9d99cSvwJaFjbT3vPNVDyr
KiaPJt/IoLtt7zSNkmpRSxKFtfHty9CGO1BTtfp2rY+c/lGLoDcNAf4xI9S5oi5DSrh9GWCBPV6c
69j2bnqAsvN9R0Iut1r/2s2QwxbTG5nxpYsn8TBPHVZ5Joesf2icKJnwCGyVCfzhDJPLOn4exbjX
O3Wiu4je9IiHMK9rlho6tQ/y+mxFwew3CPMI2BFvbQofAlet4Vh2fiXBUTtlj286z0eggMe+SKBv
8+JJuFtxI4crclgmW/rA3LAbeD2F3636BJyyWUVgh8gk3Y62j212Dsjv8aMg8bWxcJEwxEcNdT1O
P4hpV3Jv1ro244GDIb9zq87il8TOl78GVNOCrSb1Z5Q4/aYmlACnQfVRPhI4CbcKfbbadM1u/6Jq
F+aggqw20Um0YnZv0mUCwT7afBfvkPTKQdQ+Zf8bO1NdF44+d5GxYaFeAlenu3VZImuU4PxoUNdY
UQKzJStksP4770lONedPKKxQUVcqkoBBQ63JNAfMOBuQzaK81XzaE9am6V+p79L+ClnOhEbTodfr
K/5X9jhNhCDsz1AlktWJL8k70NKdV5mlUSeuyD592QQsiWEyrTGouggWeEuB0XLrfhvv1za9IkFh
OwoaaGcc3Ut0AC1a+MIANqvMFrwGVxunLAGT6qM2zmngoVhCbG+MikOr2FI6YxCqKn72+0Aek8ST
r+/U4TxHoZghdKGNFtgGo/EtTbHAF7Kr2RbnFvbrqf4jjbmDcJPp+Xa3ED+i7b7Yn1KmuP89dtsH
nmdLtwmdLMLsW0fYfRATWHfiMtAtJ77U0akjawgroFCT6kuns+F236vG0e2vpytZSUoEwWtfxxGX
RLcLV2fzg1kMjM/z6kfkYbPfFupxC7CPZZU1eC/eidhAu418C/ERCSL3VV2WhpCy5WUo9Uz4H0RF
Gj2NZi4PgYXX2WxhgpEBdLeiEksNr/sJf1cEq834O+KuFtQVTr7Ukgx2TYZLF53Vf7fqbJDZaYUV
y0JSf2kcrouI7o96mDtdTv168nIkVDspqP5Bdl4KUyHGEBCZMzMtBwvcRHzR+WUwZSVsg+hS2o7c
eJf7aGVQnTtqP2DXq+tGWga3R0dcBbqu1NHL+k9ZHoDwH3zNi3oXOUQZu36iA1HrGze0cDzrPc4i
45xbnd32arsn2PdG5aetrSk5QXEHd99q+iGNZ/EQ1Ak7OSAdH3KWt3AV0jt5t3mM1mqGOHWJfjBm
5oVy79wH1KAxxkVkBRUY3h8qcxnbhkFBJn/upM2UM+m7E4Tg/HmxEdujAHUXOQKGdwxIt22kU01E
lpQr2Cq79tYx7FCqNMpCRe/nulhxwsOEmOEGqNtjbCsJ8RDzljDTLZvTAiRCmVMdWPtE3y8d/m7C
q2ObYb7HbYnQbnrUfL13/OVyMuC4GcdA9Zj9I9g5Wbxj76lZ9JsGs4WBF1y9bViEv0VFLbAJx2Kd
gaTJbyk3iO+yqVt3oUE5DkK00oU+azgyUYJLjhp3yDS5On+T6n03h99nwEvWxb+SrhlOsPx5yd10
QXEdZjvVLxYkhot6fMJed12ljJxU/PPIp+UfXD4o0sFbsgK1zVtBdBMwZaZpXrivi8WzO8qkj3cq
fNBO0S88UgACsteLo5l6xmaOH6uzw2VfzddB1dZofmamkqeUP5gRE2hlST3Ia0Bvhe4lX8tUF0MV
LAjhuurmzBXjFS2hdqVz10Z+IG8r1Fqh3CwV7ANA9h5IIKDYLxJfQ79OerdXcCRvRg9LDpY95hG0
yQUdHks9PZeMWZS6gIFip3ukLl304RqkCedBvBnBya5Fc6tJTJoRloTDJWj/T4cK4JGN3ArZa8Xv
E9x/3zih/O/l5nl5oObuJC4I58KClSq6stuqfjLLox+eP0fuL96C8mNhHHYCZ9nrxxqy2NQWYUnq
R4bwXsYxcsUxofTtvKi7dLEaWfFrM3JP8vE7J4qM0j9VK933y7/v2OeYv6zphmAkKKFmRxlH4RcY
YHVW4yDvQznbwHxuv/8kvjYGrA24JfiwHL13nmnbS8eAHR7xvHXRjTZNyOjCVl4EEb9P/2bcdBqp
D3ufmxAb0K8b1VdBJYu7wELCZZ6zEWnkM4FpTBYoY6PDp3gWlQVoRppTsaPTwoa0dhKZD398V3hN
8zDlJ7UqCAYtAtlpFggP6oBvwY2N8SKrChJx1/RBlNAs1tzweRFhoQZfLw2NNTv4TxfpEeq88Le6
HsIc7MhlOU2n1MeSgAh1iALpnvnnIroZT8OOuqYdgilQ+V8v+zhSxJqnIE2XgkprpcTG6OC11YS1
6vOjWUE+EwMazhCGF1+O9a1Rop6EgEA0+4G3SINtT3If+MNohIkuB5kw+PAYw7UiWhq/5x6kyKXa
ct7Sz6bjj/qFa/NzuebxxpLpf2ztKbEcHHTauYQm3IGAkieMrBNgsbsv/3NagLJtb3uHEh/BAInc
gJbgQDio7NMqencVeNZnuhTJYh7ouhEc82TsgqIjCoCV/kl4mRcnhNAzQHbszlkHuy9tHIn5ddN+
yhIj9KcktOUsIlMtA+ZEKsUj6TGIjFQ3bY42uTtNZ4PWlujpQhbVhde0gpHon3sn1ZHBY0Ec0NlS
vIgbCBv1cD4aPS76oKyLFbuGHM2zF3RdHDa3n1h83qZNSdADrDAeOevfb7RwUOPRlflfd3MSQgUF
ElD8ue2apNF6sGaxVtHVKqdBXkTIzTFuizknYgvqst89L89IHsvjW+v+d8vwZzFaSe5vG3qsQD4U
hvSDQRfOuyw80hI0h3pFoe6H9MFThxnWI2x3YUZNBSYQmPOYklDZGqvTWe3wico6vaLsjnXzyZwJ
4zAdiAHDpz/VVFiGORikKC6HmonOG2AG6ozgun2IpJtTn/vgmwYynM3T78iuXlVK5qTv2Id6SGpC
Q8650HiPdNjPZx0X+KN8xCapTiCzC+vxwk1k72YcoLi9CQkXRka6iFWguYE1go8+TMj6qjtHrZbo
yx+6cKEiU2Zr55+aEfk/WVOl39HiZzWo2Qx31C2jFTtwz7J0AZPJgnVkWmlTe0WKJMSEY4BPxF9z
HBspg3B8YWv7/VLy6SnacXTah9ahAx0W6PVrpmu2ZaLNgjh+GNPZVpOA8HyQBTRkl9FsyZt6CoJ4
lCFEgThyS4MbgUa6f11cgfR8K10ZbI70aNoj3jZqYKYmOi6nISu/Azp01Xqoa+xtQQ40I6wJ178h
iJIX0ROM4UkJ0Rgt3O3oJzoefOk0y1Tz3TekUNSXMlh69CVncq7ZMPx8a4Z0OBs8dJqq77BqtXvh
nfPne2dAZR7c/uEpI4kO6R8ZBnvQvhUP8WUZsM9CHPQIYgo5Icexxklhiml4jZHL6OEbqM87X9nx
cIdfdcVT6k4F4LCGUhrOj8DMaPD7OROFojqd2f/LVDL07BkKleKsa5XJH+SDsaar5vjk5BmfJvMj
eiWlKoeb6UiSe6owHewiQflqKIRJ/dOfaBK5MAPWCq2yRm1qZeUxa3KJmKQ25ujDiKk65G2mrDuE
yG8nK/13ynbv3f0g8dOvvfAMDfJ/Nc+8OKFrLbMHIzjvvZL/bFp3tqotMR6jO4+/QglLqK7GW7jg
8DboqPzbHJb57DUl7ESd2Dk6AF+575VZ/9K+7OCnm2g0cDrh0CkzKfYv3vJGGe1lTWCdbvd/Sp0O
6MGk6+9YhVKj21/O6ykSQkkagcHwZpkJT/l7RWovCiZLiuKNpMAMhSxTLziVtIx8sv1bTVXQShtK
OYuoC0N8HdNE4j9b67QvlhO1ALWxtwuEp7VBJiI6kNTqCTqW3m4GDeI34HsxOWG5eMNQIDAUC4AA
VQhktWGMxkRfTd6qYQlaLYesVJHmrOL2ZaGEx4jJ1FG+YphDh7ApYobVcax9tICN2ibikbUIoF0V
OIRZKppXdGTwUSP8E434YWq83RUGmwh5G/nXDZK3MIJ3Bz4Mj1lRgnhc4RDiCKHpmpcLbOkPVeia
lfRbMGhM7clTxuiCj3s2rcGgwmupHiQ65i0pSOjwlFoXBgZ8E2kQBYYixC5oWqixDNDi1EEmI43c
oL8koY6aDf4w0AY0grzFNS+hEH7mWsEV7cwEyTWrjUhkjtbZRZD1ZT5rvEONJP3MR6cs1FdYyiZV
wDZhHXhMVI1a03yM6jXyGdUEQy1TngdPCqU2+kNT8S3jiba4cWfNhmDtSuSwDM2+MnWrlfzvfc/C
smXdOYQARhzfwwW9BfxHL+cRJDKa+dj1pstcHq0uDULk6WCDQ1dCKGwTnHTaZ9+M6Aoeypqq+8PA
ZR1WNbZRY9hivaYygfY1z1v2Q6XqMxOMT0FchNMFSvIrEXLkTLAU+5MXV40/Xa3gWIvi+jpTM85E
bo05+tOEGS+CQCi8Fo9z47ce7rADyTFZ3sastfsHkCIM3sj54ldxo6s0bTeh2rn7Qg0mBpbUe/tW
EOLlRtirQ5CTis6na8Jhhwa3KKbr2EiA6S1Qey+qFeHC6MRyjOMD6eN4H91ovaa9myIKESlCrd3s
Y9cCnGwuyOFKjwSYyyNDbPg0Ibe42rr4FOHiHKvOXOe0+zVKcsChk5Be7bE+leWQiyr/f5S/KTA0
Lkc7CA2ZDZf83B8CP5uQm77RYFJlQvpybSwNHwYkxpO1bKioswRCnGEe/G9luS97/jPy4SMdsaeo
0lYru02p35OcE3X2ehNxEwtvJgU9NFdxRGEEXOXjk7qZLOMSulAJVt9pTZnwHppZPifnqVP7JSPC
vum3K2e+E/gDUDwoovjusjKReyO5raNPDE4Qt7LSLbpIQNkWKvSfC7Qj8EmEKdhH5eKnCY1B8nf7
UiQM1zwuvrX0YYHYtmWfGGUldLD6cxIEFIWdV41o9QPJK/XCtOSyw8CTv+K8uG1gcBPsrCDkHdPN
ScsHscVzWG5wBuIkqaKh3N74PHnGUX4x7b2megEL7FDExuEKScO8Bi/o16/coKEhCp5FEOWxm+zm
JecDdsOLGa57ZONzQSYDR3SP5LsRw/DxXm+nxdUsnbUzkLfkpG6gcsDaoUZixBGlgSYY+QW4dxfS
e+9fjfwLQ37tWhJ/IyrSg1c5dfIx1r3lP1SlLfKngSbN8RulFBe0jZBPhMK22kX89WVTkJG2VgUn
Eun1p6FLKDmUqY+XV6lUkYmbE6PG5RGZOIbNyh6nyOOiXm4OAB43rlM37DYN78XcqhJO/BmoE9kC
QL2DQI2FphhGdY0/xy4+GZ2Vtsy66QsEWCzlkxw3crYngfKVs40dOZuU6UugsOyppoxDyLxzJjqy
RCWuD9FZM5C/eitgPwzbYFSwSKcn0zFL3gvbsFSImaPY5ZLX9NOvy+B+OMO6HI+uxwNApGXq0CGi
j1051QawJwtfGg2ThHBvvlLH7TB4hBLknepW5JjM5JFpJFicP9ex5PQC9Jm0xdpVtB2dLxQHV6Js
n7VF6gkDSb+oxlwRauKLi+WjJX8lmcDHnuFpHcxMz+rcVWd718om3k6gtbrzBLL2gAUPBOGvfdSo
oK14RkaZddMslZFVDCN8FN8GlJzgwY18TE4lQZ59k+qu9LuM44woPmfvuyYKBMU94DHyo1vs/79j
nvZFGh2ccFWwPTIfGTnOo6NIMzxH50/0jAFAHQhnqERc1XM95BEWXIiJ2Bt6NPs+9JWaQ8oB4ANy
42e7vwMrzIh0QkHrTutvFpmgVtzlxae+ghCkWUNXrd5yRTz1UDsfA7yMg0LJvlN5Q56AWhCjTAwY
4e8Gp4OAzDP10+43Et5RkyE203x2cSmMAaxEJw2sW6kh4ziMLf3MHQHxel+syI6Zgex/Q2xEQeZA
a90q8g8kzUFaL3Q9zIiGGKbzlodxQZpZEh0rr7bckHnxNh6c5mk8aG2nl7h9HqslwuAGMzKSg+r5
+8XGLJ0H/W3SnLdoEMtz4j0wc6y7FGTKB/x5toJQGw0dcz9RO1zItxTIAHdBOq9RMqTf2lR28Djc
ahyR3Wdg+TYqZW++pXqG8EUJE5cDoFUaiigQvuhC6le3R2zMBJWmkzwwW42Iqv3BTX5vEpF/LCkr
K/4ejbKCkcUyEtoNEYGnBqWdGNZZaJNApz8ysOTvX3H9sYW9HxfM/mdYExha+vFM8fPZIBBtPlQC
AKqPW/uEYT7HxnelkOnAaf0ukFnAsP1d7fHJGJTMc7lspgC1Vmfoa+v7NMSS7eQ1dCMQFh3AivDE
LA1mXiBYVmpJYha77+xB00Tjrmp3wDLZn065+edXJkI3+fpk7tYukHZlylPC3W/m4700M53Q6JZS
2mYzNl4vLc/QMhseXlDeCGBYEzNUzrVtdquLHjnkIi1fKLk5eo9OmxdFl2S6gJxb/L8UAmuwJwzs
NuUkXuQWuZ8JIg5F5whdb8p6aE7dapX+yFECcRbU6RLlRbBh4OVFMFu9VLZDseFp6uWGl0XXScMY
f4VIMZs0T3+SDeuxGGljy45ooW40ld2RVCzMeP3da5Eobd9mU3dyCFCvCIhY1oJu6K7Rym1wfNVO
W+9qnpyubFbyftOfdYKPivCtVNpE/SWXL8nv1K57bHNpNpvkaEhEf3sTW3bfFyNMrBlW7GnJQDgs
YHcJzjf2yNJxgU81fv7iSlstloZO01pyLteWqg5WerHcXoji0g8Jf/RyjBEiTu5VtFNQARn91W2W
I9gAzbJDD9CDBQ10BbL9r+kzKdvMR5Jf78MANcoYuCBmTZmmZnsMNEstORbDQgrbBTBhird6jTUk
2hkoNfrNvq7EZN31Jnt5aQREPH4+YaHUyUr2PLU3Rx9jFn3XZsfQdL03Kxv7S/Onzbrf1MPGO9Ue
zAVGeUaZhW4UzP7MPVd+2x43OUz/vMVB6yggTdB6M99nT/SERqWtuC44cirP7qrnY1C4NT1zhCUb
vDmZdwxCK9p1JqhXNrwroie/D5SFjI7jaCKmj6zob9eTcWq7d/azJo5BKjgeKavcnKcoVJ195VHt
4BQ5g2wPO2s12nwN1WVmORxcydoHdG8W+c73EZ/AcD/1Eqy5HY1B4Cfa/gaZg1j1a01xfz3sabAn
Z5Ox36KYhcVtEeoYYfHBood/wuVKMMpcZ4TJkeDAW3/AaSt90hUbIzA2hmtD7l20YCPoh9BnPZQ/
Fzgaan3VMTG9ZUdQsWAoT/9GMPlv5XGAtQq6trhYEOHLANa8w2BJaWQZ+Z3Hr6/kGWwTiSB95OnH
Zx8BNHJgPkYMKDtfVIitj+5LIYeUDFGDAmcy2RlKDHabdD9Wr46TS3BGk85YiK1rEDlB+H0p5zRP
q/sRjhJPuj8jDv/Bp5xmsSL6GGwGJ3vfDz12LWLleRi7o2DMypogEUsFwBjVyugOealozMX9xdUh
I+oSRAn2PLdZA9YRihEBEiVQOmJDzF5PTHCppOWXqhyeQCPW1L9jXSM1laxzni8gfadytKFw/s/l
MUsIVSOrI6tiPdoYfFwvj2LR+KnEEC2HLAn9OOTRCnKmvrOPUfZZIrpkXVHt9AqCfBy6to6zTqi3
D1ER2VS0i4vvnOTwhR89WVrrsTSc7tkFiRM2ygMg15cUNJeC2t6nyFDMoUFb09bJDng1/7zH4ZPM
6ZPXh1aKAnxaOPhSacFq2a/Hh4a3hyXjcbcAxNX3VNbhmCkbSRyyb6/oKOznQHfRe2IbnLkM9QxT
W/WUpM7kAUg1+9XdfgR/4XzzUCOXISEuDAs35qCgyT3BkWkUaF0wdPGS8OLjT4ujoCQmte04elmR
SA5Z8Pqvk6BKYFPtiXLFIJdMVtI/n2VAhdJWnUUWKb1nK4ZNRUOoZcljDk01BRyC4vorNwqtXrRC
LSkbeHiX4OxrMxHYqDm2bZ2JSHpXtOLJTgf23ADk9zG6tn9cO0BOGNGbQyCDaMPZuz2nQKfBN/gp
ooWf1J9xHQkqZ33KNLmTsoAG8/+j0n+227eSBFuM2PnyTqqSALJk/ZPuxAXt/d28jdjszlkha+NN
lVytjmzcjON642n+6AaNZhjwhforIp2W9PkHdTPFMt7uV9H5DoblT4zJXbbszoqK9L0YzzzE16Ec
ynTxOpOQ8Bo5Fn7VyOB/bBzTNIflvPd/Eo0GPEW+u3Fkr14NrIgwKJaWgruT/u918sOnjZtGeJQl
bNiOhs6+b/6v7Uc5XfIoW+U0qpRDXL1/nO2n5QqmcGZeShDO2Xu0kYVNe1ShEF41O82sfB5oKXK3
/28LtjsiLyKAIFCvWCZTCynwuWjs8jpLXzEKmBPYfUEvX2O5hYw9oe6y2juJk7QBVSzvi+4snw2N
KMKMdrgBNV5cgFpPWxK0j3JkU059qAsTtSe3slVofeoAW7pbdPGCMjfZO5bVjgsit8Pac9Ebpa8A
+qp0zd8UPg5tyTtkEh38e2PX3VRsxNk3gkLZ6B1y5+O0WihNVsuC6yStlfsU3p+CbxY0dpPL1aNt
J6L6DrnzY3w9kUvYDpaK36UihwlzBrCUNfPhWD4n8cms0TcoqC46OXG6POhLG56YtTUCmtcnnbK+
K/piF9ICZN56PwXKCNVGzVdLDFPCvkTNZ1TJd/gSxYDY6SgOC4Eg03Iw18tgU7Jo7J68ftYujhZh
Rlmp0NDn+hkd2Akiretial75E1Gbp9Y5DdQqbpiDWjUZSgZse5GCup9yMBilRGH01KxAp1ENnrRo
1HoXh0xBt3cmnABwrtBJ2i0wMPJalQn1JSQE048qDNPl37MHYv+kEORjkUVrhYbsH3AuTht4RorG
LRRE/bAsgaNOZj9OdpEBSV2rue1VjSnIa4sqaR4rRqqAxjWLNCJ8KXSq4t+4l00SJ9lpnnLUg+nK
xtJU9mSOScG8lYJ5aZwF3vFclWFRrBSyJNxbtmiTIL6R6Sjo4xcx4rV8hb+JYtPMPCFFeEacsCZX
h0Tbumjsb9fXXHrsf7QDDu5KxLn1mnILHvgmHCvBruRRTnvegPOuioL4/zngEDwQpwFFIzrX3tik
ZwPfaMSo9xqp1QY0jI8HNhNIMKXN1TJTkAZabqec03LtTj/W5omWJrE+AaL3qewyp6accffmUZ5W
cKpdmG7dQCYYbdwRox2g9OHr/NVJUUel5YaAvR3Xpb5/zPzeapfG/iG7YF5qzb6/EWSL5eYCygIN
8FjuUNZJjvcSU4VTgAf1G6cLY2uiXw3V6lRf7RttbFNrZtAqk4O0ZnppwsoEmv/wbjK2ZRlptmzT
0sbtV1DKIjuqZPcGtNkwLK7YTpSyBlVbIsoDufCt/mlTkL2nyfcCBM8apokvOWfEI9QSS3jPCTkp
cdzpJEQ9j2LT9BlitS9JsK5XsjeY9dHkC71F0gk00oeiSuJ8Wzq9PJQeP424hAV3O8St/m6+zZip
Vmu2QO7tX3CSKX3L7fG1xU48rbdN6BCAmsFQZ3wFkEHwwTMjRlOxtIjxzNq4b1XTzKjBnzRhivhq
soGkxnSVn+7tiGq3sBKjujFyvXVIm7BUJMW1tRKNx0wOHr+LiJDjVR33lw81LQRQAKty1XR9Gya1
j6p8KtDIFfn3XESnKn/zNWwNlDhmcrRHpzYNffQFtSzZWRwMlC31IsL3zYZRfigaLwzA7GRUmbFS
TEPLfqqBxG26GFK8DAtp4y2D08vUQasaflwI4AVxeWxeyFdL/zGpnO3P1OX5jmJbZLJ7J8poi+Ek
GPETLH9b7ohGf6nKEww5sxBysUsCe9o/KRFJSBw5kPgfa6Ui3lLlGQ8z7YMQHPEYm9/sjDdowT83
0sfNhWOqidmU4aqoEL85CsiHx2DGOMX5EUrMnzY94vy+Vb624+f67nYC1S1fVHjrCT6bCOa144t8
TrWI7wrXIVI5t6UkLYI2yMJPetG1I/rNO27HmgGiFkFPrcL+B7lXDxUpWvyq5qMTxbngqNuCqPk6
Ka6AwQPcX6byyM7XCOoq2DHd5mWMyPfZqsIDy+yCITws1pZ+nIeByXoiJfSKfa1qmmcf+CuQrlXl
rh/zeQAu2K0oIeNWui0BQx2YshXTFA2YBNm0qS+joa4qgJq16srmMnaLdC+DabAbPZBfKw+emgvE
69M6MnJVlMamSCdi0nfCH/nF0IEyfcIrHy2BqecSGGlrhBwp3b1YvhCv7J/WoiJVM6+qgR4ieOAr
9cbc3giejSlU6h6SxxgVGkyUninpYDUW/i/F36xIb1sF3q/ahElNJWEArTwYgbzfN2IrQbCxcFKF
A6PYZAUolgTlNfp66fImCjNqv/US2Mo/wHHjtvssPnl+HaBwj6zmgoDKWPr34YuwBRvl78K+c2cl
awBL+lBBwTPAyZTpMWt7/0+ZhuuTI5Sxd6S1zagVmpvp2yVfMFJHvaeFC9CyYtp7UKgZ+3gIyfhP
cyyPvqdwcG/XeUOFEKInmNFfTAwrodNixL2PLibBlacUN3JYNYrIZkDt1eablZgBH7C5BoWBSqQ4
jipVGCOHeAgAYEfxa8XNfOgLq0C+0LfZjnoXIQNlMAyCorJKHb244c4ZYKwHmEntxPmriFt3MGxb
EDrO5Fc3IHTLR+lb4z3pHiHUQ4cxgPfA7uU8rzwNjCPBDxouBYCD9E5KjDK+hutT30r5Cgw0lNJl
exizaiuMsVifY3XGI8Z50aIdUx6PRoVQixqQiKBmw+0NtdIS28sWYOz3O+hfCXhyONEwanWgZYUs
qLL29n9zMM/9euS+VevQl3ojqIYrz+JDDVI5/5eKlOjC9SHE6hh0eOV83W1WxxCT3vucBueq3BNH
nK+S4tfU0NRUnFOFppAv65i+j68q9O6/Md8daKh5omHwD/NlizyeGirq3l0PhUpv5Clax3J2DnM4
sCyl99Xvdfh5telj2Bnh1tJfwpg8A+rrgKc3PvVXJAmGsJ7yjjklPT3nCa3lWoMMk1paTuu0JT6U
yTDfhKTmzsfDy9RR7lX0ehVRbF6sl+AGXniD+X2o6rnKQ9/Kn7aX14AzSUv4It9/1G6j63p35jlH
sEcGA98XWGH7PMQuSbFiC0BqK4daoqf1mpwF3PdwlvAciIRDlSQ8bvhlcBRG6z7XEKWcqgj5BIG4
KJ32/rmhFnPEoCq5dJD3iI7MzT0Qp9HkuFtBBXYKEKdNM7JBaJEHRWLD9kB5iRnmULvSmBZDjPlK
6SjL4m9WbzVZdqpScoKDhDKsuggmBOQsxSTtuC/OAlnxrrK1LD6oUZFU1ltA36CP0nim/dNVdHcK
Bud9cLghYwWqfIf6C3/cqhTR6MR0qOys9dgK6Bvvpoh3p/AlZIXZ50unUMKrSlO7zZvw5jfFOz54
q12n4RBXKp/Xpi8DIlyAegjpdO5TvFx2i3E/aL+GQeOAlkhliaG8C5Xhq56GTFmiX0KaUmOFZPSF
+PskyEO0r8wPOe58s4mh0M8NuFuwdhTFn7VxVBxpAmkXwDXWRKaCjsEoQiRD3khfNuH7XqgRV/UV
UxrdRAbQCj4XROfbSbY1kQHg9q3H5qOIqIqhVMWE3ixwWyFiR+A7vaL01ov1cwNA/I5UpHKGwIAb
EBtPolFT55qbolBV1uFWYxYcZwsHnwtY2yHuDAQRPyJ4GFJ4dImmOTXVgUOYQSrkxp82zBLHlG4F
QQctqJIkKOMxkUjzS8/ZQ6k5Gn8+L7Bnuz2rNN52cl4tIV3h2jHZiAMA9jmuGdFHvaeYVghtK5YA
2D77IltalUqeZpxWKpX3hTJAB0a7jwkw2E0zLC8o0MFf2qLJTVkvSq0RVwb2+nQhrAdnj0JKNY+s
GX2KZGlOiy4qKv7CH4hLeTV9ybmzgW8G996TX5Qp5s5Vqj/crXqebinJ+QazK//qg94tU+loyn44
kdBWl6W3ZbaLVkHZlzzoP1BcizNY+/A8+MUPeOG9mBQ8vCjWf15hJY7SlD3ATvRHvixY5vbWHVDP
G/Q6kl95OTvgpfdT1EGk/mXPnhV72hhgtQnP2iIvIjH8jJLPBjDK/3SEsywsYgN+wAvmpROu5tfS
aoUBE4J2qP7EVEA5kNKR5qqKIh3+zzuFkPfw8MTdZycKMnBMQBgPqhDuoGn4ukv6mKbWtOQqkzh7
dEUh122oKSVcS51BVoQgu9qgI8anG0/c4mniF+036G14dl7pRRqv45ae+oF6kAviRUseJLPNb2Zq
+I7RdC2ZZR/xzvcfI9cJWooHxOEtCc8tHOHbicY3pzpyEtJ1FbXufLQtw7ljbAIPjTYbOYczVXuU
NN0QbyZKkpXrtvtF0pdf7Z1mvegVtdwEFjYP0z2j6DnkoSWHhturs91KwU78gmXfZrJYTi0hoCv9
T2yPH3mi3K83dzT/eWNsJu5xDL3U+WTbRMg+iGiqGymzrgdYsfi13RXsgJogz/rt+vpV1SleuRkz
gzwEAUHXNsMgC1tRsMuySsjcnPW8i7q7CTWwZ93uTdHVxnDFG2UOIcFsb0Zd1nG17+JfSOHCqjAR
fEhpL1nnodfBE53dyNrplIMqEzJTeGXf6dpSU+2QKf6Kym5MqCBJIHSyLh8HOLZ2Vl0quwfPHV6t
7CI19ZCunohmdN+3WA/UhQwY6jXDLa3caS/whm3jQ5S+JM4V4buBBcpG7o3maRC51k3FaikaTI7B
haMlbvq0LD/x3Ft8xIG7H+N+51dhCyw+UpXYPFCH73cNaQx3YQz4FcAElSlGnQq/0SgnlSaIZkLb
9lXTrMRz3ht98pnApTBUYj2hz4Va1pVzEZi8ZEd7dGMWBvV85OtM5zTL5jLKCfFBq+faNhO6PB8N
Bmzpc5N+dMw10fD40oy5NfNrtQ+817YdcVZ7MgY15K6wMYah67kH4kpiTg7wfYEKh97NGtHUlCsp
69bMBCg9sgOX1KvweGLmPACaPvrtAuBP581RlI+giJoAzIDCH0kshklggR2Kf1iYZ6tYkU9VazfN
tg53oW5fKHpnGF1iQ2z8oCugs+fL0KKpW1Ha9WMbuounzIc+owDMUF9gXy2EP9Wl1tW5paMqvjcN
q2bLE/ZAQ7kpzkTeXfbgcY0fz6+zGyVdYPvgWT3WlWoys0lMQOyI2wzDbiX97A469GBUp7UllEdh
0WLQHzise0VCuP8xngcA5ESo3azOZW8ZpIXQiKhHjopvsng6L0M0Wy4Mpy5Voybf45KKzd+8MHC/
a9vtW2AA2FCoRY+xvQPzpLMMjzdNNab6yHgFaRccBv55oqAehIqGnFkAbexTS0HnzFh8RmDX7Sm1
v04lbHWK2n7iCwHz5sTY9k1f8oV4GU6PDmq7qY1TSi7Fbj4TEc1gXENhLaN41iSLmlD9DW2DmzuG
AoKulboaCy4NDgCqFLXRqVFPhRbQ9SWpAVZ4LWGDxCwNIFGZOZJoeJ/bk5GJ/neEBIcr6yF80tow
43JzVGFf9HIrUPO7WZiVVZyOEQScd+eswpNrAj3vIxEZoNDY2Hh/fdvi3ijOqr63ErVVGVTgs1dr
y/Y9bFFy8hmPlnFyCNqlZk0ixzTrkH5QuOm7BtvPVsOj2/uUivkMJPdMNkXrDc5xRZkq1gQppQLH
ntlwWe24YtNkm+dK3IzsFAWOX80weVR36rmetKZgEmnXCwkqmc0FZbqNlehlN/eDnB5cEey2BB9K
bMFFCFMOitplp3koT4P2Ey0p8xtmqBuXcweG5eXpfF6lQAGmpN1t+mZRX9aiKhdp7lwXr1vaP1Wb
PSAVxcCStT3Se07CqD3A3Wvd6CbomdCLJLYfiP5wQPClvZat7rJUt/FBZbPULD8A2SlYglgQLsAc
CmgjUFV78E+7ZXZf56+kYM2VZtuy+tI+AyEHklpNPEATXSQQEE9CBb53cqak+xrFOkl9sWfp4BIv
WM1jjfAwGkXW25XQWlANnrAoFrNa58HBjS3ZlY4CR6azBXA5Vg+vmyyZ9G6L4TZ9rqH5JaS5hVVP
z7UfvRxmbglGCVaJZ9kHDWvHBxSm9T+hhYDePjmh+39HUK34nhxqrOJaoR8rTZdH0NOCGfWkL0M9
sy1CzUDo0XZ4QhMoq/hFEKbQOlMrONSYylpf21OtxXv4WyFG5uMW6ygz3/D6z1pzgE9+LlHJzpt9
X7bc3r2yQL1efwOwGs72a5CaVpAEZ/ysfNuGFkwfVdX4epr95LF2KNR0f4Hv3IJJ0klejflKckrJ
tZT/f19NCFJc4SUkR99cKMfEttnDDJ3cmlmTgAHyegn1vMzFOc/Y0ewAG+K1bJxDiwLH8TYW4qbr
qkLFDKFUnXSXMUcRlxolujgXbSX6Iwg9E8c5kqIOQG0eU0fH/5ADseWNWe/6MgJxN6AnhtUP05WV
jcFzp2xKeTA3sVNOEvpO/bHZ02c/1YjWlMaW8HLvyV5c6L+HpQcGY3pG1QckpP2xqiGJeoJrImk8
x2ese6PR59ebp6MmDsBtHwp37mN3FqzkV2zD5O88oj2UOIln+FBDgUQEwYl3OU4Ig0HAEqoWx7zw
iJYce2w7YtZULgb+qDMVnRBEWlaHUXA2scWEkGtwxSY24edjk43U53xSYED8bhKTB1FuMNYS6XOK
XdSsj3TEf8QZ5kVuMGJGG5Bg8f8DL65+Zx97EbD6geRqIdnvJzxF7lg7YsEdd0W/uEN40otnRhIr
GGtsePX03J3aMqTCYvFM9giRsayPRyDBeKrONBkTiBoP3C7IdChBWVHv/z89DkzkOMohX1whsQiZ
GNM/FFGxVD7ooov0gYClu9c7Tc5Kh59CUJ7nWuCA1whs6Po3s6yw+PhYfdEdGRcMBKbKhVLoGLgD
xO6mWqfJ9htG/LtV70d39gFezUNouAfzg/Zh/orrJHicixP1vdj18IZPbUHKlZC10yp+i+kPaVsc
OiZdU0Jf5fOhwmiFII/v/Wi3SOpkGnTjIgcieqkFViKYg4KYunbDqdZNa2GG82OPdIO+Nxo4Cjos
BMDZXtO/+uzg9EO9BxUF4QdT8j6N0DteApYdfIOzNtnT56GtRaNPErVFiOyMwpyn98OV9yZJKRsJ
AGYQQN1rkTXSoK1hJtkUdxUjlKy4xWw0GVKd2wyR8sjR4Axv2uX/RStb0kAVcSxZ0OkQXin4V7is
76rTj9QPOnJLevVg2lUk04NQ4N0grD7JKiUk5uGiwi6kBliZbrGWGK/0dDgvxIk3iUA8ftFw8Qll
lsHkkGyj7lYCBSXblXplu4ct7toVd3sEUo24jahGw6kKTt+RfNtDpc3SOHkO9EH4F3Xbqqc1Yv7h
3PnoQGUavaz386PPHWBSfsvKEJXnWTc0Ifiok3Q2P01jSKHKmFsykwebpJJ+Qqb47QlIBa83hMqK
SbwuKFc9Ua5SnM4M1jsiYrLEI9ZSbmKhPX7zXKAh93wM1wWIm51Xx0X06zrFbheW3AEIEj+9rtXa
/7EamIRSPK3w/I7fuGsEtQ/CwjZC9pHtahVQrGSYENhaw2EaGuX3ryHbk3wWmJcINnKcHXK7i3lo
5C7TtHPUL5gQjsK+bsj+gMP3LGIPsqq4rP0HlCJZILHCxTr5P5VRkDR7rLuXkJLrnuUiMCz2mviK
aeapxkPwSwGJzy6UoJp4e1DSxVwR9epplzzDt61n4htA4K5B94xd9n+GKIImYG1F+GknDnJsESI8
tfuL7lZDto4dJXsS195Q9ZNmYFpMWtvvzPL+JGdcsXWcmkydLAgNCyc+8+lro7pGBlPoTE/thg/f
Bfk1w5sr7RiHZg5Mkkg8Pu0zYUekJXkbBy+ZiCMJKjg4+kzHV66q1dNjMfZ6URBr68lG0eGyhhQd
UsD4GevwfnIk2V1n+HHVhSJuyIrODnK4uCqR7kSO+C1cn8YmSA0t5nk3vya70ydCYFKae67hJnV2
ahGbcnCRMP23gIEMqRQSbiA9VtxKBcU4nEh1XyfwL61iEktBqM7nVUuxk9FBhHhzVh3ND+cyCJh2
M5NaYhUGQU27qQztJIFPeHjjf5ty0D3FRcNcdPhWWH7ZqaYg4AON91RORx98EVeDzxwKyGdl0SiU
xaadeEc7Tr0/OHjm3SyyW8FFkTgtgfT8AL+TcU79z/EQr6/+0/fGsqVRNY+9QjbD4y0SmyjJ6TMI
ESTNueTXudMQqbTB4NjY/73eAcT7I98N6pg+MZlKfOUWwJKBYqScqUsPscmwfZxUXkySXwMpi7kB
BpbvwkRzE9BtC1CkeG93qHKNC+X4d2Dpe/5HOgPrCw+JwQ/r6yoHDTsdGEYYRFCTN6wd6T3S161f
ZQOnmBe7QQdwxnXiOSYfhHTFwDbUj2z9M+5kUTYeGA5863pfaZ/FuzEMUiQybIM/jGjs+9ZG11Bw
tatGMNCOCtMlYmMimG04trv9fe5PPuleSdLBY1MoR/fzTLPf954Zz2DV2+Pq+/FfQzrTTHneegC8
dW/8DmUEBaVLqXxBS6XEKPky+YSm5YB8utTprxxZVsa8HQgJz4Wwloh38ochJAJDPS5KbYDG9Ct3
EAY/rN4Rx5+JgARbn5QXaBFuKaJd6ehGqT7mvsgedQpLY8yiT9urcKLxYlAHZ+JGVE6aT+dzphqw
nRuYFHlHM1f5PL6D2d7/G+BRIcdhUawGrLoUILcYvQlSUHqbCHm8GyP96R19gracUDdOo8Uww15e
lQoTi0cDdPgRRdkJoEF+1V8R2IXI12yEHBdw5hqLmCNYrjnpt18HgOfeqFwDNmwDVCmFsMpLLddM
YytpwslQqMQUf99TBmGnzrUcsf6cBrkFtRICdwofVNKrJaZ9aAUuwSqIvYQpKIcl5Rwvoxy04cqB
NW8h3v1Bg8b7s7vVTOjHNZSBxaQ9rky8W7nrZlHKrva4ItpQ4mQcGugvjXKrMi3noEFiv9NSIYX/
4BLXgktgJfcPdK3+CODAyDq2S9oYd2yENiYosXI7+ppOn23OU4oT/eTIcFTLIKVLqn9uyEv1HRo4
1U7hDJtHngeh+ieO71YdmNr5sTsUIA29si5pKAbb/bNtTfi65bYfU+e9WV/6GG0gJhFpTDbTKjoL
RFeSa7tZ673utCFat7Ui1wfBDix++G++cVafvN65iRTqkurivmVclbN6V/Y4d5XdOxFiZt8ouGLF
0YtyX796imFuV/IHeu0wRd2SDtvJ8LROSoYjpntcX3iLWoGop21DklNaBmG4bOd0k94/lm+hnqhV
kFJBtTegA3Fw1Qwh3EumEfQc4kcaxXKp6HqH8hlg4V4AhTVZk1FmLuHyopsUkZSIsfdnRNB4Dhyj
q4iZhE4uTGEDtLlD4WdcZaZ0aPsehKrQQCa/+gSpMzgEIuype4qCfcOfjh51A26pHxaLvzhuABDW
dgPXKnbgbysUirqoRZxu1BqeWjoQqBsC8laYJRkCUpPm/1s52dfceXTZ209zpKJtdHvraHNNLkg3
Ys7k2eVqJBqYVplG06H9hFd6shkNZLvHxvD8XXZ+0Q327qucsF91sPsv7KTCrU0zryshVrjQi7AK
SBZOtTlYPDYzE3gtbP1f5gDlATn4p4DbsEIAgFD5Ux+haj79wL+O3wbQRBd7NGV2fjcP5pdeZnMJ
9jKHZSrxoYgLpcIFMzwJSzzMNJvlHohLWb5Z8svhjfElZeLu1zvM+bp9+f7zKlKjoXSMczc4HzRA
1a3Hd7Hf7lBs+ZzbjW64Fd+N4EUocBwaMbUqm4brxx546k/0Rg6BvlHMHlUedo2JOq4KFcZbKr/D
4TOG94NFkl2i2EE6lyfJimyQoG+9XkdvX2+PqViHSwPSXzfDdHWotosHC9YN7bJrMUqg3lmycXN6
nwh6/pT+D1u4EUX8M+lejiI3oFeSGFs2rtSba198Fha9oiHVuJC8jBboPYg2XgW3q8/UKkNoMdaz
TfFm1JQuBqFmAA0RFkKvvL5tSoLv8jJ/3ZezSl9f2ktcceqEiInOMcTCK1qv1QCfVfN+AEmvO0sq
0sb5Mw/ohmvtyslYqfWPrsNtYB+i3LyYNiYGdl2UpBdF0hPi7pcjor9Y8bBR/59O5R06lwOtDCnw
K61VJRM5lF2QpnxWWB5HLPaKDn0ZxHZRTAXT4lqFAVkxqL5wtaFxyZ6PbwWVCEQmDMTEXVe0mU4m
yTSBonUO5dc83BaWTXOhg+yBkFU32DXq6iDY5jETjmKfkSy/ZkOQImyYAlBFH7jqdYOWbcrASSGk
nwJbOh/Ri1v99EixdgN17qld3tSiDNL2pMs/RF6D3vOEFwo8td7lAAhWhtgl2AY3xALqBmDSNTjE
dNE1CtdjrXU9fujUbUTIubzNyflXfHx7gMe99fGhzdI4uNjXMT1FNnqVjpbsa5DwKRnqH5iSNJZd
/PgqAll3HGNBh/K4o0hudLtmGMyVRWnalGDvInTYh8f4GW2Khb5zFb6xJOM/9EdfQSSEbjJ6Haj8
mm/tyRvt2n/0Q9/hjLAoXK824XkJMrvwq1jvETREz1GLkJviHaZNVZ0PftnZEQRe52PQIwWdBXs0
3FUgNhPLJ87DhtUfBhE+C5HRh1b8gxbN1HZXAjj7whKMwotCmlGHtWE885H97tBGq0zOT6vmiHXk
BkXsk2MdMWufM+jZAyGq7Ytznjg5g5+H2gpK8kpqeqOWpSCvyGwOtlo2aUHOUMMrPDFZ6JX/sL+2
U24xkA0Ds645Ib4MRH0oUaWa998IyIrngks0ZcykxuuaAcmQJaamxSbLs8M2dW1KVD3umB6YC/3+
07LaDjCRmzplppT4Rw0/hs/NkFRgJwlt/KxoCPktZcZP+OixR9+jo9XYStf4hcy0qDRWtSyWxYDO
Bh8EjvwPcJy5OwMvcVIw9SuACKd6Lnn58S+zIOjH2BIQ5R1if53+867BZYBcoIgylfWOcI+xO+JE
4BmWiG58SeuHskDk91/f6iCvenie9+GNMlAVL6N9vWoYe1NdXnPDFEgGpT1CbyklLdC4N4dkAlHt
mRykBIjFKUpES3uNxW2RXlYhD54mmieWs8F3WHSFZ4lUkDbR3IAcMbkJzu5ZE9qPGEm9zjyUDb6T
2UycQJGYyKF0umOVqTB6RVWHs5d/c4e/UMCpI7f50QfcGZlCFioAMI1GUu2OwSxIE4gAflAcgk3b
+gthrcRI7CXW4MnKsVB3JStQ0v1R6LiMf3BKuRcGns1QJTKvuew5YgDQxvxjkldbJnuMfUcV44Ds
Fm/ZjjeJ3lc623ok+ec2Hmc5pfqDeVEOn8zIJd7tjD+/N6zgAfPagXSWwvRL+Mmr/F5R7vrtYg2k
Ce7MDtUowXEbEQ5HT6Ak+xtgl9Nt7VeUVA1Cnu4Uxa1u+ao+ivmVpOvENaqtZeWeJBC6MuO211M1
AQlD8dgoEZ9J8iFd2Kcoo1fqiVNlW3s1w5Q6Weq8xFFH61uFsNJ8BAmo9JhPIhmd8micZXntIA4K
hiagmceCVW21iiJD6FBUH8caGg9o2r3cCzwmN5CJAywxW0ozSQh60rQ2F2683C737Adc5pdkIooz
uoAhuhRBQI14tLHB0atG0vk3WsP7t4UtRk+HUU8OxDDq6/vlxKCQ1n9ImW7TPGfyzu5Xa40MCzbs
9I2FdaxXv8h5dNRQfzWof5xpmTjUWrzly8vtjNh+BEMMTVRqm62iUqu7rPpR/rCSk/9xtp1ai4Qv
eZ/0Z1BU5z7OoAxo5lh4CfsT7574ejzjqBB6OucmN5b0B7q2dK7rjp/+su6CxTuHlkcHLvGUNtX0
nsJoEm3XH0zrkX6J9dZyG7C2l0efjaVYSBapJ9KdGPzpo2ID+NYizVDSTzbBFcEs0Uu5VdRymyya
fl5B2gmLnuDLz1wo0/T/fpGLjtd5GTL3yym5TYL5JnuJm7O5BfLwawfPAahyV8ctq5w3+LzT0x4R
HJZGMvafmVovntWtOhISzr4OEwk+wd+xR5uveT4Mw1ErrYUPoQITD7hvVV72BM6zH0g/ZN8MDBn8
guYLWGCVO7sWUqCsCMkWYHPX3K32nd7L5Xv4Qnu47FV3EvYeq+NCj+D2kI8eQOUSZddrPPF1qS3j
s8u7Opc3Buhr16Cz/z2QVA1c0FWCzDqw/NUsCMoDbPr9jez+pF3qdjH9ApJ2vfmSRmCJ02KElybq
9citvRw9mC8Jjz2oqs0jTP9sxZaCKU+CqjsH3YNjUvMgMRX99dkss9UFgVX+VUbYoQoRowSFYxzg
savxD5aDJ8Nh01NODqatNj+DxZKTGBmpHakjbxtXaWxwaJnYgdgAGaPih3k/M92VH78jYUXJ9Gka
4zZ1M1PG2UR7WZVTKpnNZvgTCAXVjJz5ZoCcvDrmObpk/BUlMmgCSW4lOCtmTjK/aUgHqR+XOICf
oH0ogcr77cg6cQ8pilW4T0HitiIFlI8hNGhsEM6FZMU/zMVYcJWXCTi9k0wQvxUrAx5KH7xYZERj
3q0ch+Ng0DV4Lw+i9ax6YV+DwjDYNdOJtoSYmoXWNVPiPyDPPlBDEQQIsLCcaw9l+XoaQ6ELYoRW
mLsrjPT6dOXa4bAk+hFhOAUw65ImFmn2rDLyz2OW8KikvaIyURyWAXf7Xd3+WewvR4m5BXvFzWCS
7Vep98SMlIOk/rrTWGCu0Likmx/EvWdoKjzPB644SfrX7kdKnF3y4B22JTZUoTK4jVGcdZuLR1Ax
TAzhx1wnPxIElpsuDcCHL0G/Od7sET4WTTAvXuiTPqd/6gDzkIwKXKrCWpekfiKt2K+PNAMj9B1b
c4IAZhll/LxdPFvni8NAp6zO1m0BPU6o5lDpvQQTZAgnaBuM5bfVXTDENMU5Qmt+AHPWzqYg067d
rL809byyCLoXZDcMtE5ddvt0Dcja2iSt6BRBSv/IiINc1xwlk7T4nctRhOOkmJXk0YMvncUH1yoW
Nwa8FG3hLjKCAHqPkbdz9B29nEvBfNMh79ma627tpe0EF6IwXj2Aw85WmuBjXKNhi098URVnJCXv
fjIeL6x+ZDb6dgPdysbrlp40+CX6SkYQKs9Sjdrl934l4r7pMrqaJooKKaMISbeyKXJVr6P6T8yp
S/L3ZiK9JSeXfZ78AQOjcusJsObCsA/Tw9cj+k555I6X8GZESFkVxHCQNy7EHUY8M9iV8UHziqB9
EX8D3jEselTzSSxUn59dZSmFfi2cJnr6zfP/9stIXFo+Wf/HHg7VhlkTLvjU8FkAkACDd25jGKWI
GXoPMv2tVa6P2UMqYOK/A6aDldxjWMxXeSMK+HJucsrPF7gYBspw9rY8xEX6awrOjsMFlGPESFr/
Iw/UHqVoJbm0GYLZZz8KlL95kGWzwlDeywZE2pO2580A+vUT42k31/YqV/4Sa+slhAdIn5Fo4MKe
o0onobfjRhE8HwCwlZkSbic2Mn01dbrrF6jYSZsfMiQAj/GXzRRxGR8Y/lbJM296JqWbtiidsFvw
JpL+uxfwuS2i0+hGzZLpZu2ukMm+GVumHfl3tJO5VQOOTraMmt0FAGACp9u7dBJs8FA23GtMY77P
i6/RrESQbjBMsEWmvoL/0O6OWwYlXI/6BJqKtsnwRzfpKo9MXVXbxR2azv3eKea6CXH4cn8mFeB+
9XkaHbAY8vRVbQDHDOf02UbX9bOjGJ+eO13+RS3moSuB1RtFVCQFvszE5ixwOkKapC3SFrTwEyaP
f1DYoo+1QnZ4jFac1x54Kx1EL/B0bfBpmXNFe1hHezBaaWRLnrQ8RfKiuQVMgoe8Si3N4jhKHHLE
xwAsxt0si9wHoJjLMXIEK0TmEXC4C6IkcptlYqYxDS2wm+C71uZuUU/lbnjeHJVXjj2TeNPIkx1D
UzWXYhwN0kzSEyRjpF/pQSWWUDPaBQjEQYguEVF9L7RPssgg20jPuU4gPKB+V0LjLslZYllgR4sA
R1cmgKdPcaIrALcfOuOZE+0O7frB1R7x4mqd5r8gxapTgFSefixvCVQ29D//U/IuR6lJd5Ze+V0x
HCrcikn2AG/7MMmBHv9b0fgpV8R3SwavfhpPX0Lh5vAj3+IuNfzDCk1bkh0Moek5yQC5AZaDM7bZ
USJ2cJ0WkpcXtOLqRNQz3tAHfgX/6j8dylRKqRSBmVDe2L1kpZ2/+JWvFn6NnvvZVOTtFmQiIUHF
+UCGmyt06BHsYilOUGdOhOlyDYhxYvF3ml25hgLSJJjEDo8uEEEzn04KhfkHvcc4eFS/Bmne4cM+
HaFeTQDjIGXTaGQIxOTib6btM8cKLaP/AV8RRWQsNXJtcH0ZSLYb721lwIEPLN7q5PjD8x6ivjON
0SwyPEoCH3aN2yfSaT1xI/wXw11prWqIzgX2cRBIWRZ8kwTKdqgWvKuWNDRkLMl26HCx72jwP8hx
FyYEDSDiSSVTQpHgV8l8LnzIC6RndZMRTN6HTChVZHY0YqkuKewirQL55m/Fr+LMpZLJOfcWCATK
3Lwwx9t+x1WeCOlhdT4o8GszdtFGbvHAjQsXxWCjDDQuDgoZOWjh2of28PBWYL4lY1xud2yKa985
+R+psL/qb3+jZyinq5VAALPDXaXbap6RyiKY37pdSX4irmx7HYfeoLLqZaAJ2RgCR+/JGvjD0Nl9
LXZBWxVKYmM8c0aOFZaYAJ0xZhcRdXtVKfiLwdhD8IEpt5kb3taaOjqkGmsJ9nx6vExioH9Z2f3B
+FfF0ngGUNS/ggXTutk4TjHqndMqmWojO9bO72+nscpeuoDgY4aGWvJgzjm90z6aU60MZLZVc6ya
VrlLz7UHja7bOTyXlJjFSpvZh49GKz8dp2WUPMalSYjZnvpHTOe87S+s3batvJ1JJFKvUH2QSrt7
bkmwh4FhXv6LXq4AD6ikvc4r76vSIRsVvEv5Lt+wE95Py8C9YAsuCAxSgAYWJYPwhDjn5Q9mJIOs
/ZG7T7gOKFG3xxkGCoqjZvcfdBZ63UnsiI3ghaw8rAlIoPQ86jt/KmaIPpydozoe5gxK7MQLBoVi
GtT38egn/Y6dsNsBfK+/Ay5P4P8aUkyLf6IAN0Gh6Qle3HF8U8Q2TOhi7jKgD9sNlAotucOk0dqx
GSJDVemJevtpW+XqpRmohSkFesqbHGZcC0DQHgYmvy9yTqryohBO8Q9DM/rAzcAjK4U2NUQ4qXTp
XVkKo5oWTE/II+a66q9M4y4CUcJ0rirZByV/iONtDVg0lLefQ0LemfwDqCc7rJ/BH3cPzMnY2ZGP
V0yA26XTbM+3ZNZfpJx/yWbXlJrgD9ybHqwtWcpSvmJJ9t2rKK1Q0epM1l4VR+z1un/2wEG345z3
nADCbdrs6b44MssuLSrm0auWwsN09WrZO7lpnH5senCLlkWMH+5YfVbNVtwe4ih7+g/2fu6BHv46
IEzy+kKGBCQECYj+/Wa2Zf39xp8KCe+auuOJ1wXNJhoJryV4OGDZr41Yt+WG2ghX+Ov6wB/5ttvW
MvNg1xyS27v86Yqr9BhxP3uiPP95Q9asDOvvsaT00JyKIsbtWor3yBRV9ya2zqT8LF6Zulao7w9J
97HYtc7aYISjP5cP6P2RJbVB2crPXiaiXv70JQW7FY9XlmcU4NnNF7xgyA0okB7xkrrijshPo0Xm
bO9HpwwfRoGVN9exFFP+Yk5CcVSgKjl7ZSiYW07wEyyQ3oEN9QkjN1hmeh4Sd1LzmwG1i4ty7C+v
7hXo38ZQ/oAWTDyVe6uxWuAyo5ajfK1jL2HaAanj9dwjGWQnFu8YzndNXpLUgJ5fjvM8fwVluPcC
JJKMoB6Zdxp5n0sjGYrOoak7pIx/u0GwbI51hwFjOQMmzHJEK3urY7Db2M2NsL4p/+9xNS9bGEi2
EfJdEdS3p/1FK9XLTDuWldG9JFrMEuHxpUYaCQqpkBy5zcf2ZI7btuXnaIXm25utYo3XviV4VThx
TgbEI2h4mfj1kH4hd5Atqnmhxi3hFv6BsKQaUCNIicS68tb4gz6YSC956saIdx6IDyUF6NfqHmQc
8y/dfonJ7O+nZPN8c5EIs7uk7uj5rUYhecwreguFEvhM0qAWJpMg+d6AUIH5gSmGFx2w/AnZCFnY
HOpc/KHNaazWNPPgH641fLcUcDAqoxWglCxN0dBJ6kC31nwtDQAa2Fn6i5za8iHbMnqB7uhZ20ft
Nkmvj2ycQ7/0xu9iyZ1w01KgDfvpQf9SGpQ9xVP1IuX2JXoCWYh4J/XJtb1KS7Sty8yOXrlnNx66
A5rsBHgaVHKBeo3LguAeAo54AHG8qcDXh4X8HAIadGXnYeDXA/WriNzL9PHBqD7ednFhrWCVQjYD
PBacSuGyICxLzstvz7R1HHn5iBsQezAa6tI0Pvp9e1az7+juIPM1CEWjZMzaXP+CZxy0at0F35kF
+Y346MtfKKiCZ/e+Prr58l/QFHiDniUhprF9daSLioTgv1KKRuICcZHr7sgh0trzxnSFun7sMvof
xUKNk06JVft7loMFC5gEU0xqco2qrHt/1JWVcybC8HH8YQBTL9+vnVYPQ9HhHFlKdCiOmOY16hdQ
xkkytB3p8E4tSwWkxe0hR6FG2UtStSOul7rVObZol/rIyKNNZDD8fr4A10VT1ScXx8bFD1nvrcsd
cBrPCI65B0OWaRbimd8nGYOcSxhxHw7DKBQJOUVCXRglLGWzV2DHHjPpGJqcbet2Cl1vgTsJAbSX
yfQTYoqT3evk2wOHPp52ni3w6wQhSMzXPDOvxCwBtWdjUVQZrQxXz/cIZaovsyJWao7JFDK/uEGV
+2rxoSVg3u6NBNY9U4YAtRs99P6YCDbLVMFzTgliUJLbVciWZcDCfXTfHdMYgIPg9tkacDOoRaN4
6g2gHFdo4/VU27d/jOOc0TkxxGePGnR2d6NQ/EA7293Npmcy9UTXx0MMdOgMhTHkp00m8czDj8bi
pmg/XdzcCRrHV0QokMC7qjE3XErFIp8mupp+ZqSlnA8GtQJkltd+fanJDfyMuVb4FOg4yiv9F6HG
5d2dataoE3d9i8AZOPRjeyPvXD0R8WkiGkSemELoUEemXmU4f2cxq+BVkSdGjirnHSFlJDUeraz5
i3zWxbWJLlSxfS98ii58uvZc08I/U1dvyFLi0jtSttG6nOMkHW1xKUQNywQrRdEiPugiIBiS5iX9
JTsTNN4/7VDnbRPS4Dht/MsmLPqhTNS4j1sR1uiI/+PkwPiueQ7maCnR49WGnByyMcyHv7AvD3A1
+NLgjD1M2bGUTTm6xa1JDa8BqHzneLaoxcIjQ8ezd7aJtFgNh0cnsx3vKILHq0lPCca0CPvF90/M
CU/eVoj8A3acSuz7NQjt+rcd5jDnB4yGjyijreq8iOiMo5Oc1V/51GsRHJLX3OYECFB0pyHBmYa/
Pk+WufBqdnRZbe0Ss4UiJew3EX3XF1QEv/rloeA0f3v3r0ECZUgfMb4hzt1vr+THMEJ3z3k9Qv1a
Mtq9ta1IT5O2OQN69sQSUUoRg3hxy77c7pnigB3JqqxQ/AvbHPzWIauZaRu/5CL2Cn4H++77YsGZ
4L54n86fTtL3WpwHWdoFmEcoWTlnWMCZCK14+b4Tva9eFlv67XEexC7us2uez+35LlJF2WH8o2Jr
aShFvCTb8+0/2auqiuG3qyPGcWCIyUGb+hZ1mIxlVQH/fqMDiIdBmpn1kgqN1N8TgL5rd12h9Vgu
CfteIZVvNXSmn3jyvEGfXICcCnjiUfDBRh1Qxx2EaWxkLNv130WFDfeJ8gp77s5VknyTplLIL/kL
f58n8v4JPC/1BIZr6UMi8UopEgYWiWN/vDscaZqAEzvfvpKqJ5uXQ8XQ0CNcUiVd1eNK3JkEBjx+
vUvUpNz/HobdRZKx299eNJKkC4KLQ14+fJvl03qAw47nKt4qff0aMQJQI0ZmWMHazglCjM+wuACl
4zM2U0kNjpTbZhHs7aes3KLYIkpwB+nRGddrD8qAe365MpwMgJ4EYCCPHefnyATqtwSFAgH06+6T
+jEL7t8rasEXwQ7UNZm9dfHZlipnhlFAC/+b8IWWXzxC04scWXGMub6bCdvx40tCSc2TtMyx7+tc
HERXr5aLLP7RnAg6zrD7qD7t1ez6RgRiKfiAlhaau5nw+Tp4sMhho7232smK3JHQ+PkG49kM5SGW
cbV5RupeLhvMvlubG4PCAluo4X82J+nf+Q/XEsUSKNVKYddakiu6341Gr74QLj3rh7HzlPccDLyN
g+gZ/Gvm+i3o4h14s7VGCyyW3/6R1yAbjWt1/a3Zb6Z+cWFwG/+Wz4X+B2Avhp0+y/0N4NYql8IJ
ax4M9Cg6fJhRV35YHd4a4FgAQEqePLOV3On168O1TYXPHY3Ad+9if/MwMLqf5MKr6KyM0Xpc9irN
FMiewH5WyoGTxy45apq7ZroZkRb1whosr9pqJzycP6w+dMZYHE1aUKSUlEtf6j2JJ9XdrKTnMtT2
qfBnKfjgRvqF6D3hosDIeEIpzF+9AUR0TCoIM/1dSX0b3o9Ot5u5qcdZmfYMjb7Qt1ObZtIv9Am/
Z1lFy6cyH1QQjMHfDWWNrXacTZlJvMVw5a5AHd3SFAY8e85ZJ+KmRm9b5Ly5Zu+A2HwlXf/csQAH
Xg6wOAOXMA1Qy3nGEDDzdENppu3wFooV5G/5P4yFthpwQXnv94FNhpWq4XaNCYk6m6LC7FzrWOol
UgTfrqIkIIEPadcR5xRaLRPE3ME3HJFChRAL6X+xJxaWuu4X9BELy45SWtJzVTuFbAQRbqAn4wr7
3ZF8N9UFEcMNDLvsgStPvWBSx+XrqAw0wHlDL+Zy1RSMjQA+6ak+UbtFQd08LZyJ8S5FoPG+cVS3
0r4fdeLaDhZNFvtaoeJnTXsymFLyprsOt72w2qDBPiioYyr/3vhn/JF1F/NC8RwFmeGKcDWfHwlZ
y3xRMdHe1YZAEx4RPRfdUvvml8nbXGPbxINpj1gOgj6fcvyQ6876f1NyVsfn7RVWt5BDDew4OcYl
IPMR8z8wC2qX+8bXshW3BPR7su/THtNhu8u/8BuUzsN7cd+p2/kALwUadUDHg5s3kYlre9GLP7ag
7GPWtbWg59Y+uLl+EXjj3K8UNs7io5dYWdrkV/Zp5/str8Y3HASSIBt5MI9on46XACt/4kjqIyAU
PXAxWtHDXzAwQBr4V7+sKFzeNq8UpMFEW54yfjQCKcUB4XlUvkGt/OnKRsgS4Pp2FXrJBSqTJZw9
P/UEe7OlQ5i1VcGPJeGjcyTiuUK2T3HRJG4KK0wJqbTPi0PDXOprcG2PAeUseuhtPzHjBhTLPYUL
q/MAyPNPzl11h3GLn4Ap2bNFuvXl0Q4PA2jgOGeWm71hpiIEja4noWqTG4aakgBwRSOc2JkoyV+R
YqaQ1EpJ5dpe0ukIIVhqaaOm3St22LLnNWf7NJO9jXHFsCoY1+vliIzpr0/CAV7pGr6z9ieGSlAn
SKVHScE08LUm78Uq+j/g8/ckAKGYdzdfL0PlIXsEUXwLBNNlFZD/rFBiL6ANQWP8RKrZuNALF62s
3we47jxp4sJQ+LMAKgbJwX21mBdtpyljx40yBUVqdH2s589EniLYOyG+Zi8pFZ/M+H0jxZ8O6U7l
+w4Du1aolsjcppMG117ovnp/kKCrY7TSEkkUMx7Fl2UPuOtxsQDBYYyPp79hVMqrasxugEtd6i5g
ArCEZJCo4lT2U1y4CTtR/I8ngDIsQR2De4+wV284Wq9E2zWNTLiRouM9aR4DRgGyGT6Xi3EtqkIb
EBZ+lt40x7DzOW1o+ukRYmXT7TQfPU8h/39/LdjeVzwduE1jjAf3h5fLvCZviZV0ub+2LESDVTe4
WAwDZXTA0YdEKLrFE6TZa8IVUXi3Z7/Pu4t78FrKpM6zmyIZKWTRPTXED3R8zaPR5elCU8iWNlU1
BoPBdeIqhvvdNYecnFdzyRVnRSrtlj9epwcZgotNWfOgnPkEXM412QeCORGwtSJwQyFBjuLGGV2j
CT5gxevlI51XgFYczu/JP1Y1Sq105MiXWiYdkrHYVPfWz6pu0yANSJ44GhJ+c/e7ALxehhOd7ajO
B9Isz8zumRB9KP8iwnk8iWMhTECOKUO/Ms+8DI0Jd91bS4ssejmHo3leb15GUdZVvCLYMiSlyYZ/
WMunx2ubPn8GG7+FEn81SemAiU27k+pEhsRqRp4eQ6YJH+TzKOalik+l2+Rc6uYA3VJ8sLB7ztrt
0x8GTb8oJcb77Fi3vrc1eukjtDBiVpsJLv3Y0/SIwfHJMbf+jMUTGUeeVGSRsD0qjYeIyBJQz3iA
J8UuelscV3dHPWRH/9B/A6MZUp49kjxuq5Nb9Svrl0o42XCPwqKMUiZGLno37yWT1iHe5Yn25p4i
U24OJn8nOwfSvbvjLxRIkJxo8QNg2IYbYYSPhT7xVLuC9PsQ9G8MsBkyuxAGM89A6rvtCYbSiRwA
Vt+7CHgozPcF9Sm7vFkxp5POYCwA9V7dYPRGl5ax9lun4j/bdVTVC6NQ0QnoIkcxyz5WUy08MzKu
XkPWhr1rfNAx7BI+JjG4zCFNISN3AFDEdirtxanPYPwqlLXHOxTUkmF1YftKDyOr3EvoSDxTb5vw
Lyqvxj8bmxc4Bfpvn3nv7r4XBuiQPMp83XEMpEH/2mNSjbvDaP78Sx5nX2Vho3TW3fkKotyBe/IX
I8I7p0AIo2DHjM2s5cav+3E7nqU6fgIYvIvrHJCdD+8NHX+v8KObLXGDL7bcWZzuN03Ncg7LpPa4
eGNwhyIdk/RlcY6Nqp2+zBYNWie93MT2F3JkiAZP9TQQhjTiG3Uklmzzi3HuXBc5DWViViBFjCLI
eZy3v6CixXTdi/Djl4v4HLPkKUP6yAj203UxhUXjBr987KeCe1ttGa7/sJHIRozx7ygcm/CYT5QL
tPEHEvO1jrWm/iOBcwNXYYu/bBw0EM3IuB8H9QCQGaNfMUbtVB8yJ8YPZ5g5L6XlNoXcijU8X4T0
yH+5bk/r3qJPusZ0/ad4YP7L88PGOwe2nPJTEWi/GCNFyz9VgZ9trvII2NPSSV9hMCtOPyjwQ2DG
T1MvHwSO/TWF2CzANFgVahd2T4ZXzyCSsWhR4SVXsDbVgv8spVmfO9BGedkHj1f6wFQWxlZyanzG
qaHcpcngo5ZrPc5+cgthS3X5T9dAetLAUyXmANohJiIvHs+dRO/7bzKRcIBamLl39z4J0GdeHntW
iIaj1+jLHlOqfJwAtWcotgefb70i4u7hABsGn2lLSRY+cq9HAmjR7xxcOyWOAOkDvZ4B52f1t0JX
DJ4bmsKYKLsf/iLAUsSONXhSGLyHxBeIJ+ZwcfisRuYYn/CGMKpbd4JJ/0fJZQmYJFjcd9KMCCgO
pSHOY/PXXgx5J1SB0QyDnfdWYifXOJxsjcmVRcC8fr4nYvZQpDTIPlKFszJn9ECrApif5DGtiZkE
s0fUsSnPcJAS11JV2tSwvd5X6iDpLGZ9EyAUfncrEmcyFxUjVWyEo3fTUczYA4Yl8468K7hEq7XW
ZJlxRlA9zc5VNb/bBlk/bVskPPXKBxbDjRvsxsNMT+QELGK5BhAPVjOhv650wYlw+/5OyakzQjHo
XMWViqQddne1jyv4y2U4Xvl4dA6VdERefmM21aLT1khn6lvXIq+aMOMyljzu79lkN2LgEuZJQEB8
iqrSCAkL+HNb0uIfYpmeYf0NxjiDXV3fjJMRRHBxtpeuY3CcVxaHnaS14KbUZkisVLGcCpALbW1r
YnV4JjoLsSTG2vgUvkoiDIKj8v9Oj2wqrvWnfCS6P2KCMyi1tPOKM3LQFdIBlEfN/sHSi0ZvjbJ1
Ph8VZXUghe+3JnOBGFO8W7eyxe9AROtXUtKkilkjWBaCJI8KmJytzHncscGGKnc98jgQz5fvskBI
bhXnoeKKUIU4w6RQZ4/eYoUWy4n7aFm1DTJ4BtnFzwAqXa9+xgEJPA+r/CSS/hWyUC1GsC2uJEy8
TLVaCyy8pRj6LRPLxkFYaVS1tuLZIw+Q6vkeKn2zROBRASHqiGNzscrAtBzNcSIYKh4sOImJ7cKI
Ud1xIuzHXOADih4LJyfQz/AFA47oHZ9FWMgMFEWe6OGw0Zmz6CVpVq59q9UFnmLzxdNMEGHcRTy+
vRM5WyRDrHuarp43MokQZ3d7EU0pMPwVKark6Z14YBCg39qO1a7pSCFz/5+TRJPULLaPp+Irn3ZW
L1eywD143LSsnAjhHAyuOF4ncgAYfq2gb2miuH03wm9j3DROlcsLnlmuklZzcm6cRJNlC3+/bJrV
zxzqUCQ3+7L5g6gIeqVgUjklygvvSY62pNg5qbCwAOI7ajzCl3lAGowMYncAd8AYwInT2fqAxqMf
SA+OKu8EoE/gxLuj6iWT3KpCCcFOLVx69urzGk4RTU1Bf8g2P2qiGGhC+us3VmU94HGkuKcisWwi
KmBKRhsIKsormBHxQcp9vdke9bHvKlq41/AN0qZ2wEDn7GQ0Z38GP64906QeZKqwvQf4marABq/o
GIV77TKVQ7AJiHN1CSc9ykfgRUoOZ3GFzJ8eRFmci750Te5x0jVkRJbjT/Zi5ZHXEaWYUxaq0olt
850m517ZI0G26rNrvWUgbqLFbB6HHh2aheom9eggVO1RG53Spbrny/o+Dp/GPo85vVyu5rLHOVwR
G65NnY9tdhF+j/rAu+nzsI/o5wSbCOGzv3185FhF4bc0QDJcMBGN6KbYXx60qMt2bDt4bQRI+oKX
FQhdFCnuDiLd0z4uIvQqOr1m1pBvoJ+3yKtKs9t3tpnkpJRsNniVTPp+qXVAz/MSKlVKM375TZL4
W4X+wcjqcALbLjpR32nbSqbqw6ch+uTbSp8c3lcsvGVx17aGGcPyJejFph/8ZvX22U2AMbjVxPqW
zicbnsLGIffCulwu9LHoxy0LYhG8mHXIFuLPnRMkkTDF+dtWXRZLhWygkP11Ia0N6ZPLUISzGIfP
viqQGEt20X/P0UHo6WFSegc+95OUucv3pAagXJQ1nens1YAD20U6YiJQdNAsFACWvtfDHQCDETZO
M2Z6wrt04wM7p4yiwC1i7u8qQnybDxfsy4bG8OTfIl/qA7bq2fU6aE9AFgMgVGWVicc2En4KD8xe
seQ/Acrr5IMGJ6QLdsSfptOE13Xm9Vo/i6mD1MQ5YbdpVjldaJJbK21emEZo3GTtUR0s/7XD5/oO
w60fd5ivZ97Hgr1/l29bWoQt1uhNm7oM0Uzqp5d3EcKls8BQrCl0Uw6vuLI8UJeYpzib5TH3c5l7
UoEdCG5S/RT8V8QtS3jLEZP9Hd2tTXJvAKxfw74+QJwTbD+Tup+VnI/QX01R7hCm6CkQ9tSxSkCZ
en7FtySu1ZHdlDXnqlFPeGEjIDiM/Cv02GkYCljiBrB0f/sFyift9WD2pPsK7vKwGLadJxp1FsAy
lVuQJTiOjXuU2x+hSzkHMgvixEGMmALQkX4ztx3zZLC6Tlt5l+nvO8v8lE4UZxYyIuSgGMYB0Iqj
WGQhS0Ht99jA6kzwWVZILSGnwjux4+Llhm/koY/mDl7RmseEJ8sSI37SW5B1zQL6sCPV82RcWAMW
q/2epoKZO8Xs/3Y8ZivGO/+fJMh/qoruHqM1Vdz+e/EWONrvK1G2A0aztU4i+atLhvLuEsAwUoVx
Otv+uqEGvpiD7l+ZEuCpszkMWRy87GEnvyuWfCGHHuIapxqa6zLPELKQaiReo7l3+wccVum0LzKb
aMlhkvJ3cXkip6tAMsxpWvMjY5RoolYRXOWKuWn6g9UPaRWvOrrAslqQeN9m+ACfc2JAIlmG/9Nw
gkVsHOY03GO9FYNYX/YqoZCxNH2Msiv6ZcFPZ3Ap25AjU7PMmR8v51cmcQbt7i3dw7Ndhr5YjHEG
lXeFb1A2MFbNfkLGnZnPdzC6+smuFBPGnWHVOJ8hbflTtfWqm8qGwYavQ84XDPfqroz/SfrFr8b3
hk1uKjdX10/q6Fw+BVmQcYFPNtzVUfqUgmy9umBjeOs9CulDqiIBO5lCJ3dr6x0fG4Vdzqrg8uom
kEZAno1p333w3YkGfdBGc3bQWlnNtd+6A0A04UgRuQEQmRbASORn9XUH9Sl7qlIwdoImLiwGFoBE
34mIC2IGm/1bhoRUr0i4Vk+mk/txb6LOab2Kj1P+/AVcEK2WRo+78VT0m1+cg0gJHpG3tD3DlaeU
4IgfNe2n6ND4WjvtZihXClThnt+Y5YfPL+aN6ic39QBwhh/GzrQWnuSVBYn+89Rmsgon5njndo9A
9hCyyysdhb2+AToG6ugraQTdmRdu8ENDW158TRUb7/FjGefTgDy1ROgwOPTdy5ckbr4B3j7+3KPO
7MrpXm1jGrA0nGIn6k7oTu1E4h7bXsooO6d4zmT7gKeZuEQIhnD0xfDNVki1qXLz4T5XfKN+KFdO
Oc6AclbJ1iMc3ozCgkXq2oDaS0b2r9rkBmqT/2/4TBMtX3f/7ffuODhlry3+ummVhOwROUxkSxnD
WlSDIIWKHIf178ESN6X6pW58vgbNA5ZRdOpZqtA1n2IkaTPN8phmy/lZ9OaJ+DGQ+Iz1cJHGgQsb
Q4wsr0Rwus2wgcJW/oOl5A//iUQYoSCYtn9/ykzfhEDTSsue8DVv/cm61ldrP8fxtggML/MEPlFo
vl8sIUrBY9tznn5nFhpYleU+JG2rU/UAbnrQOfNBHIb6rfzATlZPmTFLTfuSB76ngjfEFIsuCP59
Ub/8+mxduzv70Om70aZN8PJ9PSVOCoJRcqZn6r8sqJYzK3qv9dSdSz7xABMCSUXB35P2EE125uhh
aM1GWL1ygZEofCBVqBFb08yMJ55GmX5htaMghHx12jB/d0zV5xsTcLCPCySv3ln+lSXRZ5xt0QAy
ZwvgdlB4RNS/GVLX6RExSZxmbKupPPBW2vooeoJVnLrp4J8e2KrCLZxKiXraQ+arvhs8d87ZSh5b
gqL7Bwh5czRnw4K74jE5Vvzzbl2/Wxmz/smqy5oiqOxaE1uj69OZuhIWUPzaDSFQS15GXueLulrx
R2BT/h1a9ZtbFLINgq6k6LA1Cp5jyzoxFwjgDFOIukTmW7k1nQxYh4VXORjfWkb5jNfzzzwy+16p
GyllcPIvtLu/AqUy2dId7GuWRxxxjTkSJ8hI+MOm2+O+xAM6kMEUeavEhj4Mdbv/trwPzcWiCI0v
wtOrDpU2errQlRCuxLuduquIoagyeOPQl5TfRRUPrdLf/A0GcxV1sQJfy462ZjadKgU0W9MTM0rl
62aQFNMyl23vQUn89bROL1B4CeDeCsLcLq1Sm+Jm0y1T1UPN4CwE6IbWtT0lEXZYvgacNAYi5ZkL
QjamE8S9l/q346DF7adovgkFu5+qHsPke2tUlwzUFTGcfm4Z6IJAh09XlKDda2VQg4oGoGq7vr9n
dLBE+z1fnORSFpbOvy79lUdiDfxcddRVMJk54if0auaQ2Rk8ib0yJA0q1EpdfBRBw0ro0QznDJxr
PUcljv2gKr/1MMsueZEbf7Ep5IjkyAzt1bOh2P5bV1HUS7+3uHg+mhZEDkNLvwFVL1bXXMysaQVE
8KrHovukoIf1MynrH3mJsU29oqRdW25M6Y0GmqDUbBj2bfgU/TS0a0AKEGF3jHkwZjRsGKa8rRdG
LvJYBBpbG5p43w3KYkcYltkoERe2Vip9yHcer/ZpYmt3NTgjadJLNUiWoNYFt/Pzy5RoHRIipUCS
+u18aPDDHidCmSm3MkYM+CVJoHO2iBiUwea28/mj+WrjAzjCzRY5ogl13CJTzkmn9g+idhZHjqYj
Y9KOB9w70dJ4RRKK/HXz2z5HkixASmbydRHay1nVZYDVpSNvcsrC6f+vCV5bKB2OzQFOQ5sRsa/L
7ae/YJEdpXhm30IWO5b2XUJH2clrDFwg05ssHeRuxWxw5pC9N4kG0oddQ5h+4UmnT6xwQ4eTTPpQ
pMbjKljHgT8QeR0RYyoLTJH5yVn4J8TJnsGLx7kA24vxMm1AORnPvMsMRHPyBeAkKi+LctGQYOl1
/NKjkMAreNspeveR118NDzAJkXKsGxq25UvJgRrziMofnDbL0X0iiC0ODWayt7uuWl9uZdC0aFLw
YE26MoKLpWwEIhIrsiiEZCVewv6igtDS5IZxPmLxiW1xMY93s+xkGlGU69pAIVxq+Zza+b5JSAR/
N1OldmV3dFrJrdZJ8h4Ga4/Njd9//MtypKxpDn3xH21lAF8NKQeAfNApMXaVxv0GeesCjB3zQhxt
u/Cj+EMVNWU5CdvP4K4AKIEJlSt40WMDzCaS8xqoMVofBgvpXl/P2781VRyRzhOkQDzVs4P3E07Z
/gMdWLWm60J2RZbKIPjD7xDAKywBhyQIWLKF0oPaMfgx4EAIuvLdKd4nsxxwjyQEw5ksy9Rnkqwa
8r3tDjp20fRmgNlXVaDrzjlEzJiHTHPhZ8ln2eFZGFUIGnRtELL4fhRbt5tmPCDXQqkK+zMFdAma
V64J5XuWp4wDdE9g635v/V0vY/nmc+jAWl7FtezQON7Uz+P4ZVeXuPA1vRII343YBqKNlMrof2uJ
CGHtqSYv3NURiruKzLYduYdMf5H7SfXtft+UVlAzIz/KlJECFbiMFqY00IJhCprT8szS6+S4vulz
kau/ur33pJaf1tazLsVHUIxlOIxFtHjrcgbx/Ksu3pPYIT9VSMjPOOKmnfgEv9tMdWwRH5+PpxaK
/jxaMS7FFhq3pPKTkvrOGAIaK1tlUNMmYvFD/ypEsxPv32ReTuIQ/f2aSlFQf0S+TrVwoovbZ3l+
HTEoei41xM8sv+ROCTQe/+845UAU3jJkSfKouqpf4UY7JHbSkR9wirhSVZZ88Q2UqZqNVRZ3XMSA
xyvKCtrinv5B+96XULkLzCkn3vzki3sQvamrVnYeh7shcQt8ziHPqjAe/4iBtlYNYB2Db02/5FoC
0xl1WEDMJLNuPigqovuui8aqV6mTfHxYL6Oro2qL4drXgQqS1jJCDjsgMCwz64OI8/IbIKvXdnKh
EBrmMfxMD+KmDrFeZZXah+/ItYpRFEGNIVjRl6BbWchI9jyODsbr8iF/DLMrkIZUhM/mYwwt8Svh
CYGV8WC97NXVIA+SHdS7Arn4COL3XwzgHNXz0G3ln3/X3P4/PneRc4jw5Kn5hNpoB7TObL6TefFY
VTGEB9p+7oJroBDEGUaeBGslejhtUqBuOwaOmzPACN6Wqk/SEVVHzQ19BRAHW59uK4cZhaaviCHH
Yhb4tU2MYYwqnZECz7JPiZoy6OY5vBMsFY41uOrPR0dyIzBd/nR1gKE1vSxs30yHkfHnySkQYORU
T1MMmJ8Nzil/hykW+C9OhqESxBP6EOc8x9yfgEhQqfg8fPVp6ArToRkazyZ0Iyt/+rUW6DevMgDv
kNPDm86NgsISHevBK/fV5lcmpM/NPHUY6pHy3cMjxTiBMqooB4W7mA/TzEJpg9RnyHbRBLPCXApP
G1XVirCCRPyiDSW+35vIcQEWXydusP2rE8bMHElLpZvztZu5sIIjNYR+U0HWx3YB9b62VUdVwrBC
/og/bNdECe+l24Z8lJTPFrlBF/hvi6UQuC6MeW8rx6jPz5n1SMSfuMkEEr7AX0X9bg+E9enQtpOw
a97ejqfx0B307isciVYaAXgNOQEeVVVIDWIU7Q2RiSZe+ccMF0bZct5I03IuSRxFvxDJnl8cu8je
nm/bDeA93zOWr+UzIT99DceFHQr8eyK8c4OaTcdtspFSwHIDDIynpB2SLGb1Oztg63Ugl4r9aEEM
JM9vUrkgza52JxxxRCQ/+kyRr4UbjEhWy3RZSE/LN7muKXAA0qacLBxK/KIyR401mDZPmf7DOyjm
tQnyjWSLESoN/Yl2vKEWbKNI6PhqyHZGxIDxS8VTKG9EjZOYxVLtuzIfUH+mJinmXsrq+VKtTqLA
eQozLb/z2wlh1xA3eehVApmRlf0d1pBbO8vLojvw6oqAb/SxmNNN6Z4zrRUDWbU5jnVNdmH9VkVM
+T8G6Vy8tVQ8SCxEtHevEJa0cfX9qKPyLBQBnUB4ie/RTtlf/9mc2MKJAZnoJ+QmPUmmy/tGs8JN
9ThDrFwTbLVA7yAtmDmXdSWN3dOeZFj2PMr/UfJ87PHvDiMLpP23qTrphInC6wzD5vUaHjLQMid/
q6hePpHbXhpdaTjxnJJCNe12k1YO4vuDZkJehUKSQzgtCwkrjMDXsqro1+otReD0ODqKQWd4HBSs
/ytglSIxdDLfWjhBQeyuy5wLN+k2ZfVuvMP8m8bvfpqxOl+JtQmXjeXXyDaK3RP/vvPwBrP73eYy
mXXuWQ90GBfw4OdP5xOD4FDvEReilGmBW0g0FjlQlJrRJlSEj3R3nclNE2H3rJLesYUmsQiFOvUT
QTZ5bjUU344s9jmlpqTdxZCtpZxFxkpe2MwolU3otlLPRKp6mq7hGTtuH4vnaSFgEClhCaMpcyEj
vtedB+4r7pZ5t0tdlF3iFa1MVy/E4xfAQebx/vRrTeuv4OjRmMMbi/M74nqSnL9JefkifbDdM+0y
/vg6I6eTJw6sdittubVDHh66DlX9EYH5YMhGre8V4kV1RPwh4oYmerIpdjh5S/Xz6p5Mytw6Ow00
H5q9cGvHZAMO7YZQB7De8zuxg2xcJg2oPsgySx9qzJz7HT36dFb1YrelI0O0MjyE7Z5RhZWrKkq4
Si20EMSJpUda4LzBklLF/4gA7CJt6ZyYYZOHTIyPgT+7y/b0kdpVZJM0UiRRqDzzNy6oLp+JOu4p
REVKTE7DQsgdpulrk3ndx7k5vt6S+ii0XrVZkAPiV1h3skJA30jHJCBMw5EhVlUNQnlh6lqJKZ3M
JmMN6hBCHAOMqX3cWfm9uzLLNNu+JaFGrvAoDMUlAV96sfFi71J1+texU3E5ldXhWpskNYyI7PRw
2yiJ8znGKKG4ddSOxNE2Vbs/hpPvVe3F0h2C+CpmvsbJCP5dBwxaVUnQrBtv5mxHz8TgiD+PUj2C
s6jpATaTAPQpaibG32zJX6tJILB37fAVJjzwc6aGyPE0J3FKMwBxdK4tcZ/xM2O0M+7B98Vy9tPm
tjwkfUM2PLqMe+1Hygcd+gqE8td/hQc/bf4BkkN/AgVq5BdI83fE3TEL+osr2Aid295vq6Kck5rg
oT5mGgFA69jx6QRa63vL1+OeskfqJPysRwDrsPRguV1JzbkO3AHAHrzlJadbgpB9rwu3jZ3S3rhL
cky4T37/ckIDW91nD9sFn2dkXLsBUHuG/Tyq/j25cv1il1BCOs93Jhz3HDAdvhhKQ7keAxxoQ/aj
1qy7q1pTfAg+q2BW3V6pWB3hu6Cfetej9jHjEmrwD3xfsZv9AWRHLtuE90uFCb7lDj4sH6wRhLcQ
+HcFgBPgoRgRD2L67F7Kbe+NU0Aj9Ykayiy9tdBCxIjGzLVz1FqdvLrUampbDelW976/iV+pBgo/
cLIukXFg517Lqj2B1cBhgWEq2FEVVVWMSDaO+gYNSTmC6hIwoLii8zmsXdHjDL+aqQjxljUhsz8k
jnL8qG10HKilCBfF3I0ipYWjJdwPNFfDmz9YBc5FCNTHf5ep9aaPimRyaqr0GOquOQ2ZU3FhBAku
nUyGSZnqSLEY3NRN8pd1F8BqUV/6kE/LOneR9I689PjAaInWysgFcioEJjmeCsHev+HsOWr7Cvcl
SVxR1nnf625oIciYgi+Ak5TGXyuvxQ0pfeja42QEavRyG9TP78Y+6+VlFbRbIqNdzgNa8pxyOLf/
Fe7j0Q4EmkHnpWsetOmn/IaPmssr+HawkU9DTjyiIl0dfLzi7iOF+m0ONpALQAIJOzDj5PymIzrN
18ci4VsH6tOTWSUKb1lxukUf7EhWpWqpqTy/73qe9Qen+UMsmdKEJ8wnHGu3krSYaUvfa/YE8R58
ie/61PAzcvLfXvPjYrGNYO+5yiRvdjruyBjzVATxJB6qvuFiC74YG4mBOGuFjPij72M0OOTKGdTj
vJpoGy5boqpiK5l6cfKOrfi3iPOzhCQ37r3C27z/pzZAb285P6wD/LOxGy+Jde0NRy3b1SxSiSpR
9iD5JdptpTCLd9ere9UAE/k3flJsaT+hYnqYMynrDfyVObkR+CHsjxiiZpNaYeeS1jjjMVmViSg4
hG36Ejwt4q8UPmRfz3OG9eVD6Vl+Zn33hZyxQuAPxRwh3Qo2v3W5OfswpUs7Syx22TI5LV2B9BKJ
61LXEtyUuWbRox2xULoaW6qpnoTLvlSwGXx1XIJJjxRq1dBSZvNRB/hh6r9k885hoRZwILdinqDf
EmOiKB6hIMpWKE2o3+eAV6LQ0nCtw5aToletHCgZ6PrNtvrwD7dIjkmGqX/v7g+dQ3o4tFHPKEkU
m+UumKW7yJNsbxQ6QNl1dEyphaF8fgGIOeD39Jn/0Lt8qzvFbSTMx6bH1Zd5jQdSrDeETArMesrw
c75QPnQJ3trbIBWjlApnslWXcx89wH8Qmit2tC6W3UKzKv75b8A3r1PYjNVkuZr5F5NwB0v04vEQ
0XIT5WlGzTZkWQD5IQP9sF43kRsse/7Q8Ls6iPfWX9HZ7KCEFBa5yio9Tr5k6BKOJoyOXvLL8AxM
S/qMy1j+iobCfmmKdc98qEu7SGuPRl47TG8pv9/E8d6kTa7Ph+c2GtDxyvevPJo9sHu0MqHBDmq/
mM91KXRdrgpUQ1iYJZ2qjwcbHT53Qob4cekL52jQbQgRlffyKJ9jPCeoBmoRhguBJQIMEYWDB/kd
o/ZdYtd0Zaa5PLaq+9i7yqWR173FuwBCEc57AvohaaTdK7AfMjXsnyJHI+h0OKSQO3AhvKksVFuk
sioGqCG85GCM+qDhzbyuBkDlsNQ+SMEXPUldnqtUQX/Q/0NDDJhcw10OeMO2AbYwtOOY1gB+UD1r
KleOayz5Bb7R0chI8sXWqKW4o6gtD0Hy+SIqJ7IO3CqtPeAGG/bhZA0EHQ7J75b5CtL8mRk/Ac15
2WwTI16biKxKdtVKnHINvWrNcirq0K7m/DUa5fg88hGfA2jBQleOWW5BIm/4Cx5+Z/6pQy7i91Tw
Cox6XJT84v6bAdvBAXvuUXruTtVvrEXdOvAAUApMOjx7aYM51W15YmMY4OfNKWCG2p6JNNR2qgc2
/601NY4tL4hkU9VvZY2GJKyox4SdvKXEIZnKVR6EljjPMd8n9yVq6h5w4Nafe0gN6FO/Uk7K2Czb
GCkc95xGQe+tcWgmp2ikc56SUQq8Bmu1GEQ8EGG/+8wkKHGpHeQ5jzcOIldND+dS7BZQSMtDfgWP
gwvmyC0nWGTVMsyILFKpQh0HWskJWXAB9q3wqMLBvRCrkeuJ9RIMBh0YgEwu0L9Ada9wXue56/E+
1CYZAXhsaoYUCyTaQWcaHgtss6fjd/yvUFrumEIUXWn1U1i8ikjutczmmQRXZqL8D1hSqCk/vCZZ
JZGF8bmK7UwyXmQKgLL9Mr1XnLuUxXle/OPJEiQhCdLbGhBD1zT1yIHgDXQH2rcXTDyhwyspozpr
tRch+t+QMO571erVHvA3A6pD/g5X154R4wBXCLn2Q9H1P0TyczG3h+abUAQz5AiwQQ2T1IMzT5Mn
iwHMnTly+XphLTYt1dWCmFVcO2X2A+fwB8XbV0G093nskSxfGbcXli/etiGAcug2bfSg8vJXvksC
jBedq4VId3KOhvQSCQY/xYMrEUgi3ZgAuE3N/b++BobfD746YgQpmtl9swtDUIzLz08JB53deZOq
8svKzjEQOELP3YaqG2JS9nuoU3kpVwJkreBkoiNed+ildn2pkIBXYgJ7TMkFfbPfdtHc1jWjBvcf
eQbQh7009VpwIUD+CAzteAxSSD2wyrU7LtSdGbffmwCNd5f1dnJpNs2903+925Eu9QJXuhSFoygi
nr0YFuvfqUevHd58eKMEWZOf7iGnYFZA1nFEOb3z6dA3PI4+FZVnQWb5ERh72sKz0/zCK/nZh6vm
KOCe+FsRGZDw8w3iK5eXp3u4gBcT80Ld8mhwP2NntForz7QEZbWdR9Sa7+JsNH5P10SqEWHAxcP/
r67msZmRDpjO4yZaiYqdWOcDvjy8qLa3LONPWEDDH9naphv+8Uc2Tk5o/NIyJa/4A8noUwX3g61t
FV4F59wczWNvYr4ngO1Eeo1U3lrlYkpUVPLP62EklDXm3K4MokHKxN8/KEK/lvADD+ctlRpKuGEP
5IRWUkhiwKUflfXyg9cZAUs5kk3bVj2IP7c42EpylJPiptZsxkjuegN0438I8S9pcjdKeIe2QFkw
1mUY2O7vJK+mvhLLWY/TH1thnB749WmO+YK2/f84nX8Dy3GfqGS+AsJKccaETpeZSTJuflJmb7NQ
J4sASEemYs2xlnXWwi5JIYGcQNS/Q6nTn4iyDCjYHLbYJnirBlFek7EYIuyV2dF3ZDoemo53P+ON
5urmLkcBURuvDq2KB39RT1bjHngits0cEnsSUVSTFYkRBnHrZyfdlyNyyLvfbnsdJTuNxytMMDCZ
lQHlNzFF8bZXSAhfftfU6JiyxjR/evHPRlvFpIHmU3G2yOmcV+9z96S62sfS8tpAzKY2xxaNLfKn
relPXtA39eLuSRBhsDsBYGrGgaZO6U/vdNXOCKgLntPmDCovh84XG/r3IY3gtYLW8k3ci7syAQxW
9XCa8mq1MYXTyDsl9XJbAEf6QPZbsH+tWxFcNgknHp14RJzRwFBigMaXbmz9BhT59X7Amrsfe/jB
IHyyd2WFZolE6+EUFxgsleC85J94BuRQXX5KfsZAQFySzJiBh3e5wYKu8BPSo1709CBJ8ZXmNJWX
Qf2QVAeyAJxcH88O4OXNPB0eh4lbUs4cF5inMosv5rIAX1BEhgCtV80v7ycEXVkumwJjD5uSQqRZ
oA3RYp8D8yhgvBKwEwuqEQtIqquMMOaf4FkzX+0FBaBxCLAcWDLpn2wJShsdJ24wO42F/2oXl6cZ
qz650jp92oOVa2eSQ4nhe3OX0uexmRhxAgzGC1+5gy2dTHZamXF/JwdACTewQY4mmgazdnVNuyNm
5pNL5RylWaDwdLE5I/khEecA4SOIz5YuSIBmTqp99IBZW6vQ8y2Nl83P94eHIhYFe3P6umtewA7I
SBqI2xIALlKX+Ia9ok7G/Kp5AJj0BJMZ5ffvxysES+n+gq2ByacLYU+pUc3OzESKpi78ufeL7Jwf
0dvnXBPOUE1GMyGbqhsG3bIRc3JlqvSHxW0c0OH/errgd7PHp9ZuQc//1EFFpRkuCEpxCMkPKj9P
9KwKabmVXZQUygFmS94AKLdp/fqUEZjXG1miJ6GKeQ9JHyJJYjYd/S324VSUprrbWYqlFn8S8CG9
ln/MSGnnK/bhDvhHu7KTnuSyZCXy6txqG32lIWxOsUq5q0kA0j9UYGbZ6r7/2v8smAaDzz3jddaP
AjQ798Ns03z95PNeLrjRj/4MXmUUfZhX57b6IvJJl2Swnj/AxoTfKarog4RJwb5tZeUPXl3Bc5Tz
Vnuc7oXoHI5XqvzwH0Y6m2o6OVW7/9slAw36E7JCklkShZdnQUxZHsaz9MrghmEUYQvm9y3D7Bgh
f6ZtHK6N1BBNcL3bE+kGwB3HFpD8rzHhypa7Uo6tPbI9aZeD5qSJm99GCIrMYTlpMSu+EE49GPgp
JjUhRpTIvYr8y5m+dvz2hRW+ssEgeEb36RO4obDIE0hYHfCvG6wUSRtX9f6439/6qtYclLjJRE6m
dIMJ4vgkZ4PV9fuXsql0BNTEFXHBKXLki9R50IHDfHxJPyaVS43kUxNjAmkcLOwbTiXUfgFy53xf
xT8hWqgwGM5b55X0PCcxkWt3RhVR8fevqA88K9+6h7jP5jVbImNxHmQLSyiYohsFKtgck7xkOL5I
UIuqBaEJNmjGr2+4YIj0d/t8FoBWz86H0BXtzbFQt8/mz5v2wm/zJf91AAcPOlHPnUYTJT6Cfi4G
9iwjnw4X3ipIRNJNCZt0wBL3LBcejwk4zPqt1VBb/xL4nJZHWeOOwJhIO7QEfpf41TPIdGJGhCMX
JxusWGnN8AdwoDyxuxGoCi2vuyH/qALJqNlbQ+MH9ABCiuoGtQgvC1dwMVWHXefaqdBXG/Z0wQpg
qwoGJTKKk/7N9gVYfJrfinTFLEs9DotnJ5n8PtgSiROdfUsjfjNpdjOFq46da3JJu8jJLXmhthil
NcPBFMo26CzWj/+H9jLKUsRJ0YIqJ6nQkX0pYkeprgUTqpCKi++jrb/d8U+knBc/Os2eqEItCecl
uj5IGgnV8dH/mY3bg4/iqyQkiqKEmojrO/yWUCdwRGeVe6KKH140quVRkzPoXFWQqjO6ds4fMeVa
9Snxev3L0IIi0IAQ2sMOHnGwgLjsmOIntK0c8H4koj9L6wsSR/1pf/bmuxQy3HRJQqXIetRl7AgG
FKsD0y/s5G26p4aHMGSrJwEcWqHChsKb6EoEYKQ7WOLquVnIPAZHza4HSIaTEcpgdl8lq366tSl2
oGOTS79qlSDfnzormZwlWz1/GfCBaKFYkXnHaFS97cgxbaGfziH1MNcXNE6dnHWb+JH7PEws1pUw
rNJrymjip+fP/ChwfIrZ5L7ZXNiZgXgoMvRH4cdD52Vz2I7HuOz++jGZrwufBxpa14g5ho2bOYC8
wUXT0o3rt65RmyvdWglcmnozKoFTiq3PUMVuXZv6CtfbXb6JdyyMU5nX3DpUmThOB0G15o/XnBuI
m0Oy5RMf9vSR1NYIp1sre/C771KvR+Ck0pEL7toxG5mWOz/TGDhBORzUFE9KFOh1KpEGMGdQ5DBx
nrTIXFXFGlm4aysUCyeMbwToI/yuiREI6Ivy7k61G/QBh0di3G/vKRGv+VIlW3EBs65O8tCqaEA3
VIfooHPjgpx2tVJtRovRgg1BLt0o63zvEne3+MD49SctBJUGuO9xaVHWL7hGE4hKN/ekf3/7z7qV
AMTmbSPPpbu+R6MNMJEPtIaMM/oXIHcTj553FJMzUBuiuA8UTyEkMB/5aFGL3suP2SPiJdqIBZhR
b9CxsvxfIcQF6xW1l4WmhPpSfELUSl8h4hYwn2KFpIbEsC3rXJ/qWJcFR2BCdaE2rzIc+uJJ5Hb9
1aEs0ALodboyLFPNkeLCpyPvFazLICOJLqhl2RszYuKLF/kNKwoiF3NdwAx1iySxpibgox4XydyM
IFJ55CNVhmxGYnD4u/Uor+AfWF9H4narU3swgvnvtWRQNrjDNUxdHiXlKEptIx5QBWehElI8JJdC
gYp+TkCxyXNxXeNNY7CzhgSQesA1YHE3CI73lINqus0Esh5mmfuH9Y0FRj6eF3fSpsZhZPogNBNt
afUwBWq3V4BF/3843Uhw/CzNEzSkqDk9ZQhA2gySScvuLsPWAl0ip83A+GDOFuf2DUmzMQMLTUqC
/dq8O+s7HQltTXrJ9Q8PFoO8/6rGcqdbBu1SOZWAUo9QOyUwN3wcd1Z7TJE5XTa67UuwB2kyw14p
XHgRDwlcQNgS0hQm7rw6vKLvsFNDK6O+JGx8LtYL0VM2osk/91vnkqNgD8daewKjP12i7FvLGTQQ
lhk1Nz7641kER0auG64Y+uy3PXr5nCsI7gTgbPA9S3eSw/p/TdKdcqB8XlXPMwOoOAUWeG/DEEhZ
IKybRfhoUTS2Ga5EhMa5BbOSotbBVTA4G7Bl8YL5d8xd+jgnFdaEzUSsGJhn/SEPWwdNMlFL/6Iz
bC+qD7Ii556UC7ICWxc0UUiHJF9ZV378wYCuRWD3FMproCuNDuuBVXgdSg9qB0NrYOfftuaQlW4h
gdfnjsyXIuaZVr77LY19+vyzTeip1NlX2MeIvNHoxyCsekjK09QxU4o6h7j2G3TuTBqbxCmYqgfu
dJcY2gjvYN9/PQZcG65w91XqHcKj+S+RUbXQFxNs3aHCiG6haWDDPLFKJJD4gU1f3B8PelfIBvbt
3k5cbhuRebe2eHkS+cCbJLP+bC3kpc59YDnz6VfdR9phdm0YqqtunIyBHeiArZYW+46dEUt3BwIS
ia+CU7rbHV1NlJPdjok8YU1yEyG+U083R0hMbSviKPjAonbekWW5rxloBsjxPecYyE2ncpGALHKz
ZP4XeAmeDrNXmg0FtF/U0Gtj86nwhWJn0OYJkUps4KWkRsFcHmB7SrvHNX9ctN296rIt7xWmwlzJ
z5HVNVWOsPjsaBL6k+Pu9Yz25ZKR8vpVEjcU61g7LtnvqOH8TmAcE/MLXCQskoOAGNnLHj0ptAkR
z7BWt3/q5uiTsZaftODEwarDGtXV+baPNDTQl1EU4B//rkTvf9IPURaVExHeQOvvbQz7KkZ3KpiD
LUhnFaxXN8c6++KHndiDSF5imUdTss84wMv6oXVCH8K0AFkUGqFCm5pue62jSYhDzBdye4n6eyG+
/sL2L2srGrvoWAgMqOnmLl32P4futSbS/Vc53gvF1M+RiQuCdY+9HMAOobd/E0WDCeVfPs2qm77P
eBHdRKBmQj/fZ+cZFTFgO2AJNvf34lt0CaBdZ9H0uYfqL9RXUSPOjTKloVArfrI0mi8PWy0wOOaD
VTFLvOPfLcMsXEX1qW8fExfP93R/U/2Q9bQ2txlw196NoMhyyt7uC0Ay/I3RflMnW0HyYNJvpWDi
UCgEi6Ko7/WemgwT6+prGwdKBFAKQw2rZnVCucl2NoM1VH9LcVP3zjdWtD+JNWnzWEbcTGtND+Gq
3uBUtf59MwAsFkfHrcfIzI/2sLeCucyzL+Zu7l2YKOHVyZlcgRTw4hLvqvwF4xcFayxnEL4P+ehQ
rWHTyk1+dBJMHDUEMn4kNbgrcrsKMiYW4wgTTEJYphNqr2NRQho9pJyPaXyMKQUUCKBEueUkUX+o
lg/dFHiO3nBmt7BfUhSevW8JXdPScOWJUtEWaABsOr4YOnhqUf0jPhHqCpU7hYZPDTTaBNQP5tEk
ZleuJ4pe8URK0ubEKl03nMsZYeKNy21BZgUuXrsG2l5K5yQdgcTLF1QelDQIQ3FpXeu7+S+Seui1
QfhvwcOkeJa1QYX+oCcMPMhTVVPcjOxUV64BnoB85L2NgY65fhenSeLKMqhKJgHP4cwc31IqZ6rq
FJxpKqOVukfMoGvo5Et41yCrbp4kS4MYt+4kgOoMa/0O9Cn4RCAgjHIq3k6M0iHpAVXx7iuWcOb9
TMPoneWMiMFOzvOl/0zvrSKBT57dIDCFTaN+O+IzzCIb0fxAdB0wfE8N5vdpQHp/f073zi7P5oGT
TKpF0RUoIC8h8LZ+w++Mt1Vqp45myMxo1cjs6HT9AUBJAQG8Yle+oJWmcSuePX+Z2Gq7LyMo71/M
AWSFVJkRiewJ2jRe89YVMXAXZBzWDzZXPqe4cl5xO674qYmy7UzwXIlksXOIY3Egs3Ec9b5bj2dm
TSuSZmWniBq6+iOZALXbIKox7qnqbli4IEX9x7aCTHHg7+7iuquz1zi8y9MCxy/Wyk35MHSZgtIi
mI/vejeYfh8kL6qmiY1biItFndAtwd0Rh+AGay5VTXukcSdJ9bH3w9bpXT4peA2K33KOtJqqY+i9
FwE2LuNOW8DNQnv/vrHO+h7L/flKMmawflp1RmY1DgtbTbOt6Z05FzbmYRBkQtZdRINVDvKZ+ubY
M8yGj+6LcSRVZCLqwvxuBtQZGCsUyUXvWbPnmTthBhaa2gSDTZeFBMjjKI3d86J7arh4KLcL3fMF
3FCICs30S5Fdy3rR7yB1QDT4OoBhFgW9npdX/Ks3Nah7xoFdxPivunUOrpLzXRlXzhOlOmD2qvlI
uUMAAF+LBcdb0Q0jgbeZ3R8CIEkTaxfi/Pwm0Yv8+/LGZT+dNc/SDKz59LWRriGyJI23iqt9R6L8
kSgvQRJdR1NcwNdHBsAXfmbKMIyzbQOtsIiwN/nvqGfdO5kPLnMq848qdbS89Xj176+QEYLEEzKV
HbthvM2nUFm9vVO44ilHE95sT0xZEu5NDfZz512RKeozjGAiXhmhdiLEka/+hxVB7MXMtObM1Uny
4o5JRaCFvWvnbofl0MsA3utCq0ZVPIYLLxrY5Zboi8S1POqWKwSRenXOsYBe74kePP0AK9hegVV9
YKAqg1Ha6ZEFQqZs99OoC48YAffms5M6IYjozs0goMb0FPXsupSYfYCqmdAn9GBYwZJvIeoBxe1a
kEKW57LjcNkDjw7ZePCfeXOeATVCRbGMjwtYKwqTxrNcenVN42beujgUdUm6IH4HyY1QcPG1xzQh
kFmeENl1/QATpWJHOyK6fPVCwUXupO7HQUWpBqiGkZg9oRK2Mko/5AMJGLWrGkEWgymALySFMOA3
qWVbfboOn+yi6NDzqPQusGjSUxPnZvrjG67A3md8WnB0zN6pYb9eSTrhKC9uB5jBwjEoIhdEHPzT
M8lqGoOfQ/H7OaE6cz/U+nV4ARpghSK9TdZ9iTS/bSlDUBjh0TK0deEIkw/BrvKwQmzWGael6iWA
HOyRuxJuJat9+7ewHHUFX1iT1RXiLSNrJJDuyRjAmvo+BtW646PqPvcU7xGe3/7alH27Mw0jwNfT
M6QnvWZ4KoX75RrFYo1EPuyyLSod9pjec0rQ8z2Qx4cwxNYic/5NIh4+ver9bqU7OQFpecwKhkT5
3Sh3JCHXdu6+HhaCED/UKiQDxzSP6fr9S8TYu+a7j1Uy2rkB05dHczMfBXM85DmNdaGQEYhvb7vI
/MrtSSKCH2jsr7AzY4zASgBMjmoYAr7Lp5MaZsPXoo1Zbho2Sc3dkAzLIaaNnBohRvMBgI0SpDhJ
JUYH2pF03qdtiMAzJL3OnKqgHchDD/giHE4mZ6PEhNEGGqOhESzQhcI5J9WKJYPQJsKZ0NKIUDjY
OcS+Lfigbr97zLptdKX7OP/D1GtQasOmZnUb87EoeNlvLh7c5PSPX2+1K7c+F4MTgdA1JJbbH2gW
wzjxxVP6llI7LwjzoETOWlMBhVhUQaKfzgApQJQ7gKWEkCtPJbXpD2wNFf9r07hhSte3peenV02B
3K9IwH3grHKX0w0N28jhXBgcJPeFDRwXDsHYWjwex4YQQJOnX021J8Co0E2ddm4DvjGthOREIl1z
/5GNedxRZrs1uTO0LPOQle3vj0mQ9thhKmA6YdPWXBkapD32mQDxUD4pqWgtlwmBGDik3Q432DO/
8cNdxAbrSuE5SOzb4uV/yrKqAJZMnx1CWP46Q5jh+D0t55Bll8rwvTGOWxBMuUuXBXjEqzREtyH1
+U+p+Ur0bRgm3/noOBV+VFlYAmURAvoWIQVRJ/u94xFakXNMnkK7r6JPNz79MCnNcpK9E6H3qg6C
es0hU63sUbzRcgemati3Oh5/U8ruuRtmU+ec2v7tsP7MH0vKmdE3zeMEt2uW7us7Za7y0EMfzkBi
fYHYtcKFjoDHN2S4r75E5em8gswKbdAnLW50CwgfEHXh0GwTBHdSW2IYxaTMyvX3RPihAaVJ4Lb7
pg5MNW12wAvw0v/uAQNEArzaub2/TZktxhVULHw2CgQ2dfJccLbpM42yx7uiTQveLmCaeFXoaZ1O
c4JgBZ45LPy6Wc+gwmweYntQdkVqrLSddvdiWExf5v6Y8UdFUSEc1NGzDz1dg1SeiplpnY6sXfwk
F7o3A0uChId+b3yhW5F2PplArJkJy4S7CuGYo0xTSoR9jA5bDSZOgHoaukDOlsey+6kI3a0zV3ge
JnzVLVPlvjr8X63OB16f89YenHu9eH1Lk5MATOjZbBt9WrwVHdWfdCxA0WasJQUuINtyZvqpEof4
ofO/7S0XZwXmFW33yMZya6sWgNSEjvxBZA/9kaIrrzzSSzZcy+1QTuJSjP1mk+wsDO54YmFmWUVk
eifQO0Ehwqkns/4U91LrJsXVYAuZNivngYO5xdja4C+bAYjzpDxsJU89RtqS5LHLDUOeQWpsjweI
N4Td+Ym5vUn/VqnzMsgUusiasXYmJVpdQDCHlEVjIuWTukeWpvAXVKbSbjK8KErJe3Zbk8lk7evL
khYJNa4C97bpT1yVmWyKNS/a83xolGL8/XetEuO4m5Clxp3seb6VlLr9PsyDzAwbzLH+ladErIdS
P9y28pbCQcNcVIxzTZ2dKePxyKuy6OEDFg2L1e8o+EXC97uoY9vy2r8LlSeCd4wNQWDxXVWVH/bn
AnlwKBo5fLgl5I3FgVLnFORCx+SxWNXTGIPZJEDxm8tH00cvtm1s398LbcwBd5MoyeqM/ex8OgHA
MADDF2y9oN39eCDOGuyZJSQSkijsR0g56S19z92CcuUQHpjDrrcfi6gdSLuY4bVmQFD9at3Np5pF
0d1TuupUMsbReQVvmp44lVVGWAepPP5NxvDdfd2IWzvT7WS+3sn5CvM60LM16VI7arumFlXvqM5j
i+K4sLk67Oi7YK2aGN+gyq81lck8nhnsRNRkFGX4ckSn4j6ahtVELacqsJ1nYXuM7eEHgtIQ1t4B
gzgDobhJQ6/jquKGxPQ27JsEUcquUh0mRXpdoFZQuGOeVgVFI4Hc0T4/jo0M712Qwe5IxQW7Ni4r
n6qW/r+7dy7kY8RjQqau9v+SjjlY2VHRH7MJgc8KnHFLI8vXdgHmDu7PWKSXiHc1XZhecrluH+YN
S1crVlHa4FVSPzksUZHKLETcL4/MuZuZG4f7acIAGZL6g6DiUXrp0neSAKwZh02tK3dvpZL6gvRn
GYEFEPTwMRxY2j8yyLeRqcGzvJR5OfLhZevE3YPH3NPA5LI6uev/9dKlPL9Hv7Q8gwbOGuB8hKwZ
dL/+4t7+/hVKw6fcb66whLplU9bOFFe4E/7felGcJiTXb4fKxb7eE3r1A/AI1ShNvqrnKyA4F0yA
B97tRT8zn9diAhFiaw9Swt9imecF8Sydgaw96cA6FLhcyRAfa9gTfLm35P0tXpnVNZnrDHcB2r5J
Q2dMEARnLHsCM3Ww6e/06IEq2pmr9wlbYuhEh+JwcRKde+1Q1G9MwO7KVU93ajaoUBFIH6YslVw9
7zp4cHZyprzByVsABt2yx5ytlAqkooBou5OlZkG73hCB6h0Yf5MUck6Yj5Hze2LD/wfsZPDU3oNF
rQOyXHKEWnDY4SrvIdTeekaHtXXDv13RFBnb/JhxrBbROxTqsOPdDn9+hkiwoOAmi1KONsWIQf82
M9J9l6ewSGGdy1BC9TaL3tX/k78MxGmaZZIpYf/87Vl01skv/tIxRxN8aGjSW9DdN5rN6g4BmX+K
ixGpcUWv5YTZAXEzozdbTPnoAVUTQ55oAO8C1B+WvWJHHB4ghhxRxNDvVK+HGrw1XAhjQlnzeffk
3EwEGP7IzE2ToAhlj+YCLqYV0Lgjv3j2JlGWOHS9fFgpXSC3bLmEVHxqgCx41OiW+gs85ObPDBy6
lK2jaJY/LczUVAD6KFWP41TmkOqB4essuwxRc0JgePKtKqj6ksP534uLE7c4olxlFBqbM4zCg53l
xjC5Qeg+QTTQKr4OuaBwmBVKHohyVMs+OBDiGeZ/FxzM3wBfWrryqn1UHehEkFgxcls8i34BXBQV
T930WN2R28hRc1GhUOmCyWCvP/QFTEiWG5sT7tNaiz6Df71+vSdgyqkJFl1autDtcusyN7hS5gkN
+m26HqsyF93izNO/Yu8Z5IE46p8Ds2x6EORbd7pgOMfs7yugW7HhR1NbpiOreZDzr517aIx8jbci
8qCdJ0gNXYqlCJNtZWQC7bywK/eE1kTQ4HE8XN7pGW0vSG/7XGNTzcCaOO10eUKvEYCd9whSJqK0
mknZ7PbzVKyZjhyYpeExNdZR0Qyba++SGtdoneKiaC9xZ5075SUuMg3kvsCN65Bv0ZNiIi0TjcEA
JoHQVy++qKwodvzB4ogF0CFGvwpkqdtmTuEue+Skkt3UB+xyHpF0d1/05BLUe6PxOgE4aOOwA4H/
+rtjFlZmOfZzImVim6Z+OIzQVTp58aICC/5OEAu/o+jhbiGLizmBJbVJp7OXIg6M1q1JXle3G8SU
J64V0zBuhLFa/KwP9mUXryQTMWZew1iSWtqDd097+ip1CfrhtAWhvanRvu+oEuqvjcUQpdOh5KNO
sQAwFLlp6Wcms6WUfAwETU6Gn556ncmWKdWDzV3Zq9DaCuVt1MXwJ01psb1AdipJO3USHAr9BU8Q
IkTg7iAVZirtkWCwT4UJ3M+i+ZOCl24TMIwCZHbR7v1wJ1DUiMdfpBr6EHu/3a66+G+t5Rg65lFx
yYsVeVkC4ScxXonZpFVHnHL2T/DV2915EpvwUjdPsJhCf8D8PwYVewfAvK/wP25/zvW6NKolPQk4
Yj18hQk9sZqjKveHXDuz5Kt8dgqNT4gWCk7D35JlJTmBMGR3mgV9teXV/LiBNrnEix5alh1I/Omw
dEvvdMG+sRV31PcR3XUWTaVSmuGK1lr/fHeowE+WG50abowhRYBdau7lI5O4tkhel3GfyZuUnqJA
8eLfcKxh27FayZhJjdBo1L2ltNybX/xZ/z2zRQHFBTD2HI102XuPYfnnWnPqshUYJZPbv7dYcxbH
PjMVIFJogtPLBP9wslLau/5TmGXkcxqbPLjYbh1kHv1DbNMZjqe+Ue6+BLsoiA8LnEKcVZSIqW4A
0n/YKgx9ZD1F+uNPVr+E9Xb+kBh5xrBzFt3MCyzu2tsQ1dmhYMK/58ZTScJei3JIckTbFngsmNJf
F/WlyAEMSwKfXvN6tqJWxUZXec7Wg5R1etP8sCUSytJxs3uqxM7wHUSkVRNRghKRR8HEK+8cyD32
0aMRYSgrdDFtPemKNVQo0DxnjtaaxstnMLjnYDb0Lf3YOEL4o3RdDYPMBALxlol0Cz+wfyJLGh0S
IoC1TDk2op6Lj+NhXD2fOvdbgcsg0TmMfWFR8adBZx2f/cddyv7W1zMZfDukSksFOVoUELW9Mh1c
PeO1cUHUv3xaPI/lqJ9FPiuzZbFqPzVMhXVdCeC+xMOYi3nv4zTAHEELn01Xd/MaGSDRPv/8Hd+f
N5Vs05fLTqf76Wywfl8NbwS0lT6y+Vk9pOgvtlxU0NpuYwgyZBEaVUr4bEZ5WmFQdwD97uyT6QIP
5ewxHQBabU6+HhWro8ZRSZ1MqKHtBcm49VFhEx8c+0XFHHoZryote7G+vuN2mVy3hZKKwx5zfRq9
rjBSSOFRKpZoOa8C7+mlSA/UE7JFccFzaKNAS4WPAUMDtol7H1ArCQhJnCKuuhma0Pr3YDhXvm4T
g72Rm2rNA1B7pVs637FLjGac325JnR9PSDJOuMIdvR7Knip/RZOjzRd0kKVXSXao41djOYl4lJ13
ZduBO2PIh1+za8aYWTEdLfqzyVxa5PVIplj4eQ/q7x+LjS6r/yF9mFMpDXf/2OBK1ARi6ntyen4O
JPHSwle8rSIyYo1jF1FH3a5kDEbSvrbPrlpKV30QienT5Zy+DaHamXmtTZrVVMdIs7Wv5QiP90Ea
pMvM7pW5RJqCjvBqbUbLyOljVz7800bfdEgqCL/WYED56BHT5pMFmUHJg1LVks9MnxQNTKWR0FBT
8XyFhkKQKuScIwpxh+Dz5eTGgw+hcrl4j6PQJ2Pk/a0pR3IY5p3V3KmE5s72fuXJrLccaTaA4eAZ
jrVdEwUY+FB3bL241NubWDT/qhUYs4DjQcF2ccBzH1U8HjyOAC3wKJVAharxknjbhW83XvIJqfEL
CNw/NpsFJl3c15XTjb843qhWd473ffmBRjXsEIniSPZZAlFHHM9UbHpMjYmyf2T/3whdXx150Hih
j44sI1fvdKxksx0E+mVXqBpmMN+XiZdjCpVL8aPNpTbIWqeTnXB2InJkZRfcrN7Y/AnVnzGem96p
wlqNuM3rIZSYAqZd+xYDUgzwFXCv0yWninjJzlxiEHs5wCrlwqskGkFuxo5CIRTO4Y982UsXwkkB
xe4b86qZabmVDCT47b3EVuA7+JAhm+L7tx6NVLsFY+E3SAWQ+8TBIvNR0FryyS8qTKqZeJ26XIe0
GTyGUjYgLWO7br/qsxMNWAejYsPz0v7mKiJp4A+WXBv6rdNNgGGdSP5KwT+RHL+uGevRO6aOZ6Ex
6FLiI5bPswfBjIZ3TkfZHM2uvCHghdig1R/EjWwVqkw1Op/sGJCx3wr5bqtG4yuo4F0GJe7hNWmv
YoPYcxZDiVm3PqXC8Z9LlEFl8qtdCzktYbyxYu6XDUpljmyQlPGjrgehMYAF04+nKAovjZYWZfFR
KSzeGUoikKI4s+haIn1rRVmqEXUjVGHACoyR1XUdMOi2gXDDmzlpyRb0JQB9Tk3k5K99toFYcP+I
D3sF/G2uSXcheE+rPPUWlvDeygGZ7W1DNaH4GbotzvagLjg3KfHgvaPLl13I2Xjy+Jkn5NufcacC
dBqsD6Apb5bdwjuJzeB3OmsVf0/98Y43rZRBgJLyow5bPD+Z/+z+qdbVAZPQCXX71jqG9jcbOX2j
sDQwiIG1svsDAGiTc8AM5k/1BqToh6V6pJvbXTSLIupZL7gYUPaosb9EcFRvNeuwpc9kvmZxVBfj
Vn5m8sUQCeObRskyRV+n5jQvij0V3Bcaq9Y+1iyV/M5bqR6d4RDFVRimbluMsb7iyI6CGmrENh/T
iryaC8ASwMSq/ySvnFFORV4ibwbo/NHiERvLUuPaS6HgUEANy/GIqlYwSOCuWVqTh3DxUBVuq6t/
0u8ms2E9KiiYas9J5e8AOLXCZ4EpOobMw4d9TMHtekCVPtNDZD5gQ+VGRGL94Ynb4/CaRYQXwQT7
wj2/jvqPGpUdAKVSb3g7dqFfylWYzVhkahFX6zn4TXP+dBr/8RqNDIPqZt+kbI2P8CKcRuHWS3sd
j/KNuP8OUjTxI/f2ZiCHlwIU3V+7dfHKYvLOYFlLgx1OIf0GmCmDLUJM2OPYvVEbjaPdCcuCNVGg
9Y31HXcyQGXFi+OEzunTuVBVZbfXPx3UyZ4higGHxoOVsLypTqMQZXmPkuS7AERTquJS9HvZex/c
GKI9Xdt68tctCc/wGokHmmB8kepr5VidzQgknZn+Si0KL3WrJMa3IT0eDkvG/J4ZxNygR211fb1/
f1CfLA9tJfmmEnNgx2YGjD7AwVXyAyRjhv9Osj+Bs1iGS5llCD977jomgTkM6ur4C46pk5MYpKkM
H59r7jgsEdbvo4WKHA7fE+n5ezMJt4Azsc48EgU5QHKhhZ/v4s71yBQX1+wyINxUhn/gdyP+DQiu
wTR929gCLpfg6hyVDMa8CAJ5JFxfSExvZWg8DnLx8rlHnUru5y68G+m2D60KJxbHkgXb+7fY8MAz
+kF8EHqQaZUV/BoXrtX6YOX9MPjQi2Pb0p7H4AIS4+q7lwG8nsP5TnkCxp7IbfdFKrP0BUlveNFL
kp3bfnJdEHZNCa5FRJvYF9KR+ApvU9+FiQ+4IsQ6UrXFLLc6HNdseADaDkRV5aklPlklzxaP5gHQ
bOF4MtVFZHvtwVli01Pbb6UsKE0pU599Sy51QD/me2XCgppWP7uATRrTWowkyyNR/F78ODyHtg6w
oWGffzuL7TQfdfCJt0FvlmRZLnyO4dg4j5qhHDjj99C4w0YmJrTlqmc0d4vKyQqez7TuVg9j539C
fIqntP1fD/O8Umow+UpvjYO3+a/Kl3Y4AnGDO0F6dNnSvOoJq9FCHzB1N8bxvsCKDCn8Zd2PrPcJ
RaoDa6Rden1br0P8HW3u1lyaqBmoPJ0HnHydZQeizm7t0cNH60jFMRjqeprDQAKvnSSyIy5GM0jK
Cep4/oUmyUZd0MpBlrp7vO0s1+z+rj+j6eCt8RED5qOSSncR4+EIDpcRQYNjDiz2JcqjzmBzDMb9
cQNcHGaB+0uxUgWX24yfGqyb2AYMNhDoyNb9tXPpm4Zp4OaSGBB4ebzvPrJlOPUMXM5QnGOK+hkX
BKKPL1hZsRuXETXyXFtuYpP6SD4ntgZ6n7IV2kesbxTbpvqz6OwVOFopd7lFfVhZ6SDDIEAGjeRj
ye8QhsJJ1Y3sncEvdG1geTA6Poz6dDhlKYKkmipN0lZSNqfLXJ8m2hSjaFdEmqY5hwcrADkMaBvR
OwRIjZLpGRpdhx2CFNRS3n4XAMEMLhlDPi+qn4mssS6P4R/UbpsvJ+7NGst9219f/gAXIO382OIo
rUVSs9VwjOBZ3DKBPuM62d8+2zMz0tnb0yO1GGa8ztS04H68iO/RBaXl3M5NB1gKqiH0dIpNNPJE
aApI6rB2kHZ7Jwe25tJKh1iuR8pc/yITLyNjytV2gLCZHX3tgbeRRivFPZQPt15QUGADSzTDQLRE
cpdgSEBXkjy+BXd7cF2/utnRfUB79ghLCNV07O57jiU1XFq1RjA89Td7Q7y/fJngnYoOnScV8qEC
gcaD6DVT67yAmrjdY8E2N8BQ2gMnQSuV0beUqC8Q+j+ajJpJJbZ0F4xsOLTS17e1jCTm3qwDGMA7
r8g+SAZdOU0ZsjNX9i6VZF9QwKTRyJCslpZkiSxstIv7qiHiJ8qpvaQhl1cSjO7vRxxlhE3hp55L
3mFmEWQ7gN9oNgYVcZSHGEcZqoqycIfgRyTz0Ebt80XcI8fnCzsFSswE315+Y/w2vCPn/0ER+lNx
IZHBcYhsxeAySzd4AOZfxhCA+5UWLQtvJlpWyFTaiBUvGqLeUQK2ixYTkm29VXlwxKmToL6DM3GM
nEKLDwHm7/nMnUuqP1iuWkoAF2kR02BTRrRl6ST7i4DI2ebnck+W2INP+GMqeIEvmslzJ5J+aDQo
AjC6drOqis+0P+r5WUTyQSjvalwaOaoAnf1TtCU+t+n50iK886FGnszVRzSGPl1VELpI8YxY0qfW
NESTKmqrumaSvsIi9dq6ZrVA3EsLvNg8U8207qUvLAtuNDtlNmxwLHf2xxmP5EdsF/4iT5XOuy+5
i8e56uoJ37jCyaz4gfKOoaTb+WXHlkvbD9jCE4kos+GJPFg20CCSbfzwMFjuogRFeI9swIw20qwI
avoF3ZUrm6aCITd30X1zZ3tsj6iARvTY4QwPkhvFtsTdroQZEg5X4EWj4uVBwqqgyqfIydvCqTaR
k+mFuHTjgGzXRSPKGGwbVm3ueuNt8LmcXdeeDcFRwWcayZ6jLRyPhrXW1ceqeDWRzt9hyXRF1cn5
9k4jT6blxgcorL3vZ7rexIb3qCxFbhZds4z2wM50KUa3aKIc34bIxsrujI6KjzRfOiz0XX8pZS8U
Nmv4BaV/TGVWt7NUo0Ucl/NVO4BUaOotr5b9q+uRgNWWQfDCeIdf6UPsfYkYUzmZxCMXTkLL9HAu
yVlI/fe976wNMhArc+TyffFcbIz+JBCCRg8dMACp2w9tJ4lydDw+LFf56gp6PtHXuqnn83v3kwE1
jQLztrO5Bh62fQqm67M3SOO3OxUqLcRfhSaFc92ypWUY+PDjEH42de2UyTYnHmhW7BApqi/JZGu8
a2o+xbSnvN8CIhIKMhYouFpDjBA8J4rhJW0wLETOSTr9hUM5dVXQ7IeHPVzDFt1VVAj4AEE4Rrx8
lOEIJpmO1b5k47t36iMoCaZks4UWMhX2uEWEpIwlBH3AAV51AelxT+or5jYZhyJs+TudFREBuHFN
91GDdsjdwlkYqI+AUqhC99Xgi4m3FLg4wKZbTLBKiNHsTkzmfwKsJX0jfbBlbJWwGweXQEiPp/0G
soGsHvoWvNHJ3ynw9JtBQnKbBY4kKH48e6bD5JlJJPx+oZokikxJJ4VgRUzW0BR84MvOp/DOJdzS
UqO9KsOxHhfcoxaybwC+kjissKFnMvmSLiGKB7UhfP8aXH2zyZqCi/7RbGfyAasddbX+azefaY8Z
FoJ4NHX/Bk7Kq95vjKKOWOCTHkOsPko+YZSRMatIgg+Rg3LvfVUL8yFypXCJnqyPVGR54Kx1nW61
Tm/ZaermKImBvCY68uFuzQNqlanDGMgc2ZWvRf4dk+QRj08Kn/JO4Jq2vG4/jbB6V7wG8zPHHJ7J
xKsn+JvYV6sBX19K75ZfiC4X6/NdiYBiPZzUFJbNLhh4MOx47C7WGnSrbrDTybtJkNn+NvLdzWNN
rq9usL6EfqKyCzjb5GJ0QOMkKrUGV3a4QmCFq9wOmyVWdUDk7Q2TGky85HCbxKaGSh8hgV4yFAMN
iPKqzEXK+M2ImSjqL2VsLUSh+k02TG8KR4PznuCbz/mNI0Sq3kJGxnuGN1RsW8PomTcL4gXhq+MH
u2aG3zUbitY5yJ283O4fcb8msmXbsOJUcHoz9kJu3lB21/gXvnNTb+EGE+QLTaKaJGl3x4hyK7H2
CJ5wbGHkfuKiwMj47kczYwucjRLFRTCaXuFoycUjNxp5F/k1SiImHdvCdCr+5xdGzDuHMCJ+dVJz
AZXDHyk06BQU3y8Aq31khN43UWctdLRdsUnyYhRqwp/kqr+J60ZwTuWz1nep6Au6zzgskTgsdDDL
2a1BuRUIGNUhlZK6CFimj5aiddqYntzq6A7fZDaBIQzEfjCPAB6yBMn5V99GKbnn0fyhFZHcw+0U
LM7pzvRZ0f/uCxir3xbTdAbUKGwrkAaJqd5uqZ9Q7r3WmtPZSY5EqnAQzfT7xsrcuuvmjOFFCIug
KVgV1QKQnxJwtgmYaB7KPRcq67XlN7CiIg4R4/EJfnvy9nAppTvpD0rUMnZvLPEE2kIA+7MmfG6/
tzzHsCffUtepwSHtDqnB9DWZJY78Ju9FOUkPVGLor18AnFtmqsM04fikPHgsf/IGlzsRFg+4/EUn
R3Yk6SOQ6aWNxyIVg/MpjBwJuH50BIwbSHXjEHgFSR04SuxSE2YLXKXO6GVxikrcEHT1HPg56zq7
sB1XhWgkgSR27S+2WqRdX7b7GjyCi/yMv2GrZyKiSlwYr579xX7aBiZbjg3yucvAEl0UCaqdJxo5
Px117ErHlLX8a8hQ9NtBINmI8fKGYSxySum2UfJlhkN+bASNoophwNwupZFVh9iWmoCjDN93oDXv
nSQzxC2KShdhl2AyoLZXzunA/yWd7eIoVRlkzBhXLAm6Gf+oDzOMx9QTeyLtJY2+BkDF0lDpGJuz
YzgemEpVnGcCFpghVFXF0EywK+geynAsnLacCW+eCK6Y0/EXqYA5/lV3LcaxKhI5e5lE2A9NGAjY
qG1Z2m3GaexcW52BM4VmwkJwTR1kS5u4RjwpdAOW/qsgFVCvd2zo3eCH2+hukDZ+uKySby8f8xWZ
MkZIrUJstFetVXAWpfxDnWezKgAS/U7buHKCGRPAvcl0q6qXy99VtVvkBG09HNBXsBgSV1gd4DDb
KoLf+h8r5EhUjmCWb+LzBfF+KrZjs7MamtKFgamMVqcolyUlU0Emse16M93Um+Wj7lf8maKqElxs
YY2a1hdcDrYDxLMhqEhnbD6+p3k8LC5xQt+0l9s6NUHm2mkwXBHjWgzH8qNMnrctqGF+cTJCtOPv
9LNYVuw73RUqrjeV/9n0NGWBfO367bOqvL14UEiFNcnVKG2zp0hDO21zMJmgCaTxSbTsNRlXbgpD
yeOzI+rTMCQ3EZT6gunVnOU7Dmk5fnZgFwqV/jsPUVmoWfyfmFXqQnWpm8xrAHXGH5C7afnVLjOI
cu6vDeoInRZpoZyfsg0oZq7EJpzR6KsKSlmrHkNFiDMZeFRErPPwoMradd/Se8S54bNSI/QZ7st0
Wd2NWrdc2f4lwD5uhCXrP/kknG/s91PSq/lY+tr3HC0ZS8JujXqJ4WJNy5ABoXlIu5J/hdOnzqpR
NETheoYwmB6gkYJ0PeaPfjYZWiHS4FiEZRAw3/NIv3DWcmdMp98+lnlD56ZC5CwGSIppJ7gqJgXC
slLkj/ad1T4cH9t7HLMU9QB3F7GsjyDXe/gzOoxbECHFnf2mw3e0mke30pURUYM3Zxpkbc9Q41uY
J7/5Hf9YyRU9VQAkWbMIZfeG1Oe/ALb5W33+olKOgE2lbbcLDHmHRORqVmfoBfT5inXKShLW1TbO
UKZHqa+Exp1LlCBs3M9dhTfaX1eg/tAB8LfegPeNqjApcviEP0X7vFOn5AI3ptL7cSZx4qtvl4Zo
dL4aBP+J3ssfipxka9TpZqdXG/pzHwTNIlUVXyYE2sTl10Z/G7/eDBQYyhlii0dRnbu6R4fTi+YE
UK4iIDjMFxCk3o2OLWb2f6D7cZGWiCuvwqZ+/Lxw2gl24La/sqOPjoKZ6TMAsYYunTCiNAf1uODH
mM4FWgX19e9OGhoTixK/flZWNRqcBrfTcw/RVK1sDYmwpf4BPfPPVw7y6Fy1ZA5/WxKEnTefG2Y3
sVgQJHRIjHuGcHRxyre6McMgK6Be15TACgvwv0Q4AME4fR7S9JTTqxrOz7MzQSCO2Abvq2JPYt4l
qrkVSKnHNDok4lAULtjy+uhL11mIm8RMBuS5VGOcDi3Kxvyx4E4wfGcKG+SrscnVWivjug9AxVW/
Ca3wxcp/oOYqVHSSB+7S+Jz84bdGZM0JfszYxUPaT4VSoDb/nOSchNAxjwk43+VePJcswn6hPj3w
D+wRSQMpoGommF8YyZcbfGtK9KgpO15j+S6CpPWUdUSGdRtQT49Ab3MritcancQ3PO61vmNpxcXR
ltEDfebjJM0PZQaKDOtuNvPasNo1CW5aEQIsuexrmqTqRvPW4oMOkt1voUhVPP4kNmadhHVqViH2
DtRcCRwZJLnzXE8tY/3HhgtmzOUOqkO+vdiyDQqADMKuL1wTyIjaKoDkq+kFhel1bdbqCfJT1PLb
W55YoQZx3xDSnpmI5VCqelDITmb4+Fp2CbDOa/J2pfzNrLTsdeQUmJfxsSzDcIFpl+Om3hhpDrBH
yctTkIoGlMEyhupsHErxGcbQZSqBH/EWXp+zT/SKl6C9CQqP8ZMDLje2LR9C3ZnLFonTKM94wodQ
PKSiR8qiNw4C9HzvplPW7hZXrnRO5OZmeM9XwHUtqvVRWBAycc8p2GM2GJ8hzR0RDWm/LKjalAH/
1HvhVnJZqaOalVC8E8Upfw4kwSugIz3yKinzCqN3wBNxAC+xYbvmGT0CPogVtmCL9dUVwoF3ppXT
9YZM/qTGyBSxi3KbR53P57T2+bkAB1p5URmWHedPlg+JmgnyRaG1vD2IdG7+7fPSXg8HgYygtQKG
itVjFpi8cILfVcE4Tptdf27DMAtRi93DCCTGhyXDGMQTmQbTWMbk0czmJNBAPs088tVvOTLtJJvK
c5nRDoidfMaqQtVCSRf70PMHGSH5U4DQFdH12KK3dGeWCQtjF4pwb018MEgY/29dlkV7HsxP/iOi
Z6Xow2rSAT5g8wCL9sX7mIXyQhoggLCQMEYlTCLiZtTzmbKhsNAe8HNaqekybvROjOBy6gVG7Jdt
9C5cSJ1HNOcCK3vEm0dZ71ZYFF+rCp+wVk70liAn47w7Jl51u/jT/g6nu6EWnGHeBA7lwgGW/PPu
FXvVhTHYTKTL3+5C5vBLM419D7/C/L02/KKEgaycsempITKGFzMoTscQ6uqQ9vOP1ReV94aG2Cl4
gjydEBzxt5lcJ0HDbltIyyvF5kA8ukoN54UV0mASNGFoGyq4d0h4TXYywV/DZqGu5IneXXB6ranm
S9k3DjE9qGegHrdN964CHnYBdzhtaW7k83L9vBRvIXll7cK/IC/v4xWwPVFjJXCboyG7Jt0m7Ylj
/O8EgVZY8Bd3Ad8hMqIlzxVwe/0mH8Dws4sMsKVJuxwb4I7nR/pOQqliAG9v1xD/6J6DvS54wEsX
4LVS7+Y3aM6AYiigcELnhPIBsmQNYSMU2BIP4cr5QyL5syhQKpoj6GgOnKBCrG+9gxVNawzCX2Ul
q36OnsQatIpgzcGfVhX73j8WvV8NTYQDF83nGE9O4HGN+z3ZsmV2eZwakMi3wuKDslNWrqmkgS6l
VrPTzG00d/9347hfr5yC+9y4UIIxq2YXc0GWaEdmphyNfCBlc4s1f4p5DKo/4taXp55MQ2/iAEdk
mDV2HcwZpZKkioqfsXbKuqe+WESAuvYLItk6XOtIccvwYmmENk3Ld0QFZrz9uta1fnI7YcdHxIlv
9j6/t3LbUUcgknTJbi5rA6zenwPBDgixwUftzMZrN1Kkn/O1Nf0B35kqUYTx9PR+W0y63y53+Jg5
MJ7LRfdi0bZlmrSKonhT+dppOpBQsCUSIykuDyHEX4UvChiye80QbMKz1hPTl+GI3vQvfRM3zh1G
3vE5zwytoEsUgCc1wHNLjcMJ8rrOewVrlmQaZ3Xye9O2/6WWXlSiHCmMypSc5nVi4wzgQsXReA5q
Fz0zbzAhTd8MU/oIQx1gHhHpBovaq7oMBCo2q4St7IZHNFYc4Lf3kIZKAMNw1DdryslAl+oGdT1z
d3GINuRnld82oxvg2GQGdOACHXAebaZFab6sL3uKqlTiYPMjspE8poqgi4l4/9tHL4t4/+3ifHM4
xvvaKSOHgRv/1RSOGaUny97DbTLlWA+2CRfJQpKC4vPtL4INbplH0ZpGTVewFNCJxKA7SBkCaqpL
7SDhdsdg85QLA4P9DnfhkDaUZR/MKIU3GifRXrh4M9bnjQnUO7+9nJwTEEcxfWaJbcAQxWIAy/R+
/eiF2S33XpcjGuzz9731Jx6Oetc/wAUY8LM2Z1nArCCwY4G/GxSh9xPakWmWJRK/8zWhXAy0GcA+
2l8vYUHmkGl4mK9jUX6e+hG7vHK5zz8lcXQf3yv+A4Z1fZu9gp8AwXHQ+KXTcIoM4TAf2ze7xf/v
Et/VAcj/kwtExt3XnydalbjcZeiTFVYqzCj7VqHSV8EGPl6hBnuTSueFhQkYj6IhFdRgWDsiCbN5
w+TCPCruE9vGe2IXn/lV3ql4H5g5D5hJFebf3Gdrt0K0Ew42LU9bJM5KS/v+UUr0yuugkfOGtrcL
oN5+zM3F3+M19FK4HKVx87Ck8PaMEOdKnV6FjcWzDVdarJQcyYx/ONclum8obQg/0y0I0T+SdHVd
2Rpz2Md0bnEPZ1hysU8o41uPw/Am7UhmcE12T35HtekJGzkgUelyPFb1bCfZYpu4eK1RjsO5ggip
QRMVsoOpKW/Jzlin3vgPCOI3Yx6K2LxvwqSeYH1MvoMhJ5PolaSAPaN0VvDuaL9SpvLb5zcUzV2J
YgqaiD0HQfjZUGgc581rgldtZiT7hsMh7lfwtbUd/w+YzsTBFcj6La78IFqTxNieSNRu2Xy416zv
ktrjPL+XN+6hQYP2mSsllV7tBGjUlnHAnK3BY0UPV/nDapnkAuYPaC0YiPi+ohkmHc/PzT258xHX
sB5PAyr0Ma+JrKOo5TAETkj+WcA6bTFOzkNkDualAwYQC5trdVGLvebEGFHLyy8zxsrTsH5wuXkX
FLVho+qh8m9J+Rb+Q7p5iXqgfRmqqvAm1+7tyLFX5Jhb64Enm3uNP+dpokin0WJN8cs7J/ZwJMpj
iGx14dY6u0KntW/XdOo+eQo4toYyPZ4LPYJuBCOugdXBVLCO024LlsyiTv/1IpjgzOEF/oqsLIVq
VXL2vgRNxsCMcyS+C2b90RxtrPia2IAMFjcZmNuh0sGUjPGChRZYzMV/WXeZkSV1HQVv/520K3xI
EAmEY8mP8SNsSYpoAdaaAIpnat2ymfMcMWLTX+0mCndTHNTg0dHOowOhpTSUYGv0xI6tusMaTxj6
ygPMuOYsNtq03AnWz9EtfCErkXs3SsGyQAUdGIRugORY4tjkn08ApLrt0bh5/0vy8otv8Txs2H9p
HO7MNhvxw3ipq+AKmkc0/XeqiezXNIJBRwZfdt85q28uOBk60dUHdNIQyYxyLw5wk8Lh9eyYs4wi
wPxUnObn4KIWgbmkUF7P5X7ne3z7/qfW5qrgDxeCM3HrEqLl2+zPvTMZbC4flTHr+p/3c+/BJbwy
03M51WOObd6TSy3JK5t7pHTCKHPbjpVIDvI8Wd8A5BOG6FMl3dyXmWjrpiTHfnKrLV5mF5NvXA8P
6dgdG1Ma95XD3tb4AmtnKsVsQZ3ASQuwNN7KwoJp/0o6Ed5Mi1OrR/qElkWQknRagxP/7eSR/YTE
uKc/eeHlMIofzonUVMTEOG6Hx0BJKgHgQlkVdCbYsKlVhgCZTIn0INVWGEYrFrNAZhgrjYH5282R
sgLrFi57NP5j3pNLO5SBF2drE4tTZ25uweLtSXfNyDeKfzyKH5NCZmRuQh18ePwPe1h1elvYCW31
2Wpkx3kVV72HA3Wkffb6Gf7z197HEdyeyZkqkm53mQuBVdkdjDF+yJ+AjV9rHhx2X9q7oSif/9vU
7f1eoOMEKGSYFBf9BZovTdWjgnEnk+sURWviqwbi9x6S4eJeFiUiLuTx0XcefBV5QH46HJPrbmOF
Yn2tiRpkCEYFaTl64ZXNHieGZVL19vkeHgYg8iTr1EgxeJ40ngos5wpZ/tOt7WToPEpveiwrDb8g
koBzbjiqEkg0B6f2xUZD0sqPWPu91h2IWtdnl5Pjgg26wxTteU5pa+gyVBun2O7/Ra3afomD15/j
Fa42GsUsJ7s6yTlWEtUlr+a5Sf40tT8mUcYi93+v/DfgmVCuGDVze3xwIEvLmerKOhJWkfWsGOs+
W6zC+h9zpWNWFqqGJrw9mjGdteoHwabo9ipfna2Lbix/TNKaBwHmB355k0NWWpu8GH8/Dcecf0uv
vY829T/sJNg77r+rm0a157O5p1y3vA+6a8lkKJAcugehABfzDbZfIn6xNEuJKGp6qcdnL8nsjzIb
RDAZqskSPEEM/LX/igtNGskg0UF3D55QSfuGiXmDIuUm0bqw4iAH478rDdSJjrqDfUnsKOdV82dH
6pSZFyYt6YVtTUPau/CAXBWEQbYRV2a9pXyDpZmwUCaX8fNNTTrR5Q0qcw1iSEs23HtpwGow/1aT
T85tLdK5CaAhKkl3AiFRn0kEucz4ADA83B4nURCFn9vCVnpcTQn3DF2fXOQSZNNLYjpp1Z80VNCx
TNdRMztb9A7mZwdu4bbTy3CGsmc16/fM8wWmyzatB9FwnQvBTkWk8VPZnKobM5wUD2sfJ3+UjZhH
WSj4vxNjEuHOKlR7Bx+mS4Gf2OYTTQM3xDU4N+U30XwpGXp2FtWADrvzLmNb7YtIaqUrklMth+4c
h0dsF+OrgbNXRgUD0DEQB48ebYjN12vs6WdcvdSdo7CE+XdchR8jksdmOV4ESvC4XdZGtIfJCiiS
h9AJ5nf4A6S4ffU2ZE1DnsvbJlFpvO93eRUqlr9OE5o2EoG0yZ8WvU9LHM+jYHS5RamEHe/Bc9Lb
w3zPULnKBDN5H4c2c/MyackqtFyfwm1WHTBskZb/Ft3Nwprdy4NuQ/q3aeHOYov2qx4iojcPYCha
qarZEBZmsE057TiNXffZlMuttt7lCla4+UGrN5cdVl1GZXnUgXeH8NLjpXDH1ef0ClSut63qXQOA
ofp4rwVwcA6EMkch+FENQggfHMrnPoR2KRzHjBclQ39MzX3soPZbcEuDDXxjyJNi65XQfi3o0W+B
oTW5J9SBAYuVxzlvmlJr9r97iHGrGE1SdYzsmxqDErprKEST5OcP49qJ5ZfqRJy3C9kBABfVSjSb
5yqHf+wTwQudU+8O8/p+OMjZe7F8bw+fAXBhpcMkuarykK9ZMR8Qc48zb17envruHhv7MdeecqEo
V3VxzTnkKUlhkqf/XN9RMW4GTRY7et3oGuvyejLqecVq3U4YCPbfKQS6UuVNxCgfhvp6IWcKuI6D
eQ4dAJYTTPwq94zO2G2qes3fulF7wstcV0LYkQO1cslvueP33FozgC4hXIasVkwQ7F5T81ZfPPSo
Bvegr9Yf4Pjq5XqyCQ4cZxUxhlEY3hANLfO5B1DHqbMpC4NVcYTCBvNwPbwA4IWPSDRY+oacIpF2
3qFZ6PHt8KOyDNjN6CTEtv26RTRG3VJyjdrr1d/C1vvxqEkpm34qSPJX/n+HVlNJokkw4V2ZpWgZ
kDOURuHW9brC2ukpJSBAtUY5fOoItiwWywQSFlOQKz7KeO3UUkXveneeK3242Nh+Ck4af7k9OE/a
Len9kyorVRqfCKQMOmTqMODD5f8icfKz65IMsKP9go/nr03Mq8IJO1OEtzl309cQlkA0RDVKIN6U
FcnyFhS0u3q318Cdq0w9o6AO/BH0VXq+W9vaGOORsl1KsoW9WMuIhWJ572qSfoX1GokkMO/ffaX7
G93/FcdL0cUNBNEnBkVli7k5pZ03kVComMg5PZuSk7H6OxLUKJiPkpWprP88y5T+GLXeyBC4nNhI
dBIprYQ9FvhbmzodvtrcUJXdYFoxDyEKUkJXXPRqVrWfZD/XCzopaAeXxrO+3TAhhWXiV0267jeC
xiRGsMr7ZSEtLen1Je5nyb0gfq+gkuck69siUrHSiUMG/UGKw1za4vJTtvHlzKN8iHDo70IHutvv
XFJTbh5scn00hdAMM9lZ6JApVu1pz7Q8GusoFGssS8bicNYZJUxtFjqy3bDJxOw0ZFOm02hipA3k
Z6BlWCY1JvBNy3+WWfKLULpzeh4aIfmcDNfqwJMcYJOBcMZE/7/71Q8b5IcpwhCPV6BVxoceHwaJ
WSfAJjVe9IBuXuM/aMzpmMh0OrJ7KFJUgej91tl9sS3V42Tp5fiLvOkyYhuew7pXrWPi3qe/amVS
0fSrtGvlPOfnIhHIFi8AlJAVD/0hjSgdxvV9CxwPfbF5daFq82tqOCI1K4CKMDr//6m66TKXEBP1
IxlhzG3ND+4mnfnCN6Fl6A3EEAoUmWipwW2FdbKieBWqYniIR8Cav+TAq4hdOzmwqRdNgyEZgVZV
GfqLPFd5+kyWaaR7GNS+MkyqMPBGee7Z15swPzbjk9mYq1Rk6Qn4Ae3TcZGEa9uG1but8Z3h9/1T
cItAqLak/xOtb/KWL+c5A/2AY+8G9WSLbv6ogpPvMj+hgVV3galFrVx8p17mhQ4q+FKWZq1ItrGa
TkAiEwWPGzHiU7aQnj020aQDiNs3PEhJmZCGs0Qt2dqOREFPj2fCSqd17mpz9bQ5yS4xt9ISAyyD
7B9rqF0bgPFlat9X9t2PyD5e+4wnZLUUhYRMLofsQagZmIO2qoebOZFNuYBn/sVG9FdEwHXg/b+1
x+3ioWqhPX4UyIuGlZHvLwUYARe+HzbCmCgjsKraffJMX7It+AAU022lEwatwyqRq/GNlQFo6Wt8
8GBwyjiXFYryl6uWwfCbzHBg/98R2+sF4SX99t3zlJANxTEObc8NQdRAquPefVxebljQyyYMfN2G
y0294gCqCcy3NbXFFaPDUTez7XC2jU80HTRLtTVwyh2ihS8jFr18fe/6s68iiyq9EbniLRPoZeez
ixZyvKoKBYp3Lc3fqZUVO99FDLRnzctQCiweKWPp2mZU1YgsGdbSlgOPfVToin9tTO4M4D1abIkI
pI8FquzwjeIdXlgq/dmar46/8nX06TcOFYT8G36MkIxJocG0l/YoN2A5GMPkXgvPm4SyCvYvN7Gv
lnbSki+b6sWa5zSrVUgEvBBHKTU6mgesIv8Kve7zb9TgJd1DJ+U6S7XGYnOd5erisO6CssRG0KPB
RW6rTQcvUCOn/7J0c96WsnGlsK9TryCx84vxSVeBSKXVv/QifAUjpnB1yKDSlen9C0h0MExgpEEX
6cx/7PK0HKjayn+TgEWc0reqyHP86sGNyH/VWoOKk+QeP+hC4t/4blOf9fLoSGbl03r1B7nXR17K
N3D80hoJj/C+3rGWdOAjuS/sY7XRn7rxaCY51VFpP3GHb/IA8eLkIsmF2WTh+QghpbfCMN6rHIc9
vOEv5hMwUcM1hH1KeqA4BcCXuURgLI+gPIAQLMGUPW85s3ddBSTt/yoG62yuuCWqlatEkUqZG74l
YZET7JR1XTQECysAf9L/68KXm/euE8rV82Nj8984nLLln3afKl+Tb8SD6Hrchlr8RpuNP0zbBK+c
qS4lb8ajnqC6RDCzIagJs6/k3Zq7usS9NKP5tPs2Kxw72kHFfLoPCz8Esk0d4Ue3W3Icx7+ctey0
3uqg7AT8ETUuSdoZwIcnir1E7br0QIXv0M3lUdF6nScrt+QRC3WotVD4FZvErPXZ3kZSv7yaF7dI
lqZ/gWwtcUwaImIwDFX/kLSH7AqZUMIh8O6VxGUeQgGUj+VE3aAeRQXLBtN3gNoJkSshtAA7etM6
gJEELwMT5I99DjWI8kMSHkyxrNJKGEo5/dv6JawAyPOaVrhZLL/FZLAtZLcUceBVNIlLGfVbQ/m/
L3ehdlErDIBdTuOSO3tOigAMOPQzPHlxznJp2iq/ozn64tnMKM226FD800ycOqNrft5IHZ1HEqsY
xejXPfPqCV6y8O8dJAsLm6iWekg7zLL3wW78rkD2CxLjXIhefInCFKv7SjIxDqAVzkxgK1u8w3Ow
TkGSki3pT7j5U9/pVNW3+IoCW3nUG4AhT8bnV6B0ykFl1Y63fyQFiZt0vo0Sqyqks+5N6wiPrlWw
izT6uwTpf5rdDbGJJo+RBn7JqFcEsavX0FeRzvbEKcW/dmtQO/j2DtHq07AUJplPvxtT4D3k4Z/5
axEm/XsDw8eJRLbt446XQxSbqR1w95HZ2RKh5XrJqgKDrgtwLluh/LKryXoEBwTdWidK/1ajpsK6
5R0aLXBoT1KSpLF3F1whOD+gnZfnpj47TJcTPoHPtH32u4fvWl9hWkF/fNe3S0dEcUs5YeeOLhPW
YfdbHfYyqQeu6esuTo9YHDdinL8hHcuaUCeXrSh2498dUmnXQx2h7AQ1SwTPvLRMc9yhM2WumZPr
HnWi4UGUaOAMFiMqQWbUAqW2w8GKaJ6jiv66R2Ievg812Hh5tOe2M+skogoJYt4H9OReh4iiDJ9k
vwIpbF6YzqGJ3UwEw9lu2WgIcXw4+GzwPXRrrB/R8XKla1PRL34gl7O5F42BQyaJRPUbEuyqLLOZ
Eej7vQ8dt72coyjMbUaSYcSSOY3A46PWtK2pIO2V/XdEmmwGYcRQ7BXTET4BDJyfaCki8SdSGRSM
hJfJwdMT11ypxMb4pnHb/UqepwNpN+Emq4YHldQYHxYNoy1sw7oUJnBqrJH9/gw8K7w8cL6UbWeO
e2+rnUvuU4NkFSvjSr1E3KnvAkkInpZESqWWDzs/614WiHW88eX7vpUDu0+xpjb3BYeOdoEcbGjP
lIchdY2VO1A+r9KD0j+78Ew/AVFGJHQr38N2qsYs7UpfpHl/5ZCuRRbzyzM8gsIsqRoyRyUd7ONP
AQOS6xJvyZHV1HWSQ5RlJ4sWSFwXkss35SFdwfi72XLBedIxBx+0B+M14LJskdPtZe+5pJiQfk3d
a8DrbPsSdrTdzuc/Qq/omRxoBY5OYT9nbb1RK/OTL1ti5gkLJqg5ok2wvHjTchxUWedH5NzWszF+
JYYTMNRp9UhuOuEppn2EXrGZMLoiwWFkGajp/Z9xDTODJgdMJpOPOJ5tCqNk2uFUdn9mmMWVj2gv
8TlVXZwZnH5+aeQaT1Q/7AL25S3azuntonXZe/XWWQKlJMYFGLktElhFspsNl6HH4prPWZbZ3Mrb
CYHPmy/F1IXvlQF7hTW53Xgxd8/f3UR5YdEJp3h1dVdVfZo+gdlY+TJazaDP/jX4tnq2p1hoT/Ud
t0/O+9ZjHvFQIE5USiRu1safcVxZb486ueHdTzQxwm0vhbhdFuaT2mbffn1ZK5EPRbVHAzd1xvBu
2gILg+Dj7UX4P64K4006vLYLa6FfRo09S7uwnLHZMwn9Jz1hd0egPNrLMAgO8wNm5/vL5KZQsrEL
KpE6atI5v0ZwTdbspP+ZJ3DVwpCS6+rAD4hW3fHY3fp6p3oUYc8LbZ9BH/2rzL9DSJLiSxrbQMuw
zvm808tTqOXTAi/kFMk3Hv5dxGKoIw655BFSjmO/y9lgB94sXcXuvTBnVT7LoxVSKO1pAL5ZB4/R
LcUu+h5XiHMsdeyNpxSfOyTu2ClwCpUi3bserA7XKYEzoXfzxrFCRIABnxgXTgxzrDk+L571jn2j
9HToMg+dXG8En7HBtx6MJjuF8j2E+YeUV18poPeG2AXgCq9iV2104Ud4SjmGN6/iw6VITA2cabJm
qup4IB/AwOUd8MVXRJ8YlZBoohjTdItkT5kv4hzAz9A1Y1gWOOXz55NH1Ab1QnBDkytcUQrWNkmS
GjtHEbuy0KifZQCkfewbDtVqsjcLVkF5YKJ4yd+Eio2Y4Be6J0fMf5KuVyvOMQ+JrHQPtLR3x7IM
889SjIeuXt+4PPYl4GtRFHF1RNCLGMieu/Jm+c5af6md1JOiHkBunzCay1M6mIS+oBuRVlIYFQx0
3RX6EINZD3GMTeT1ML0DzvlUVI+7ywp3fOBA5T5MMxzJ64r/TlR8bv47ab9jscVNecX8vKLY0grM
wN6cp5gu1YXdMW1cP7EyRA8fZ34biDiQ6ym7az8x9NbYJz01xC6KTlDyzT8L75MYxd2zlDV/mCPr
1ALH2yCWH6lN8jL7D1xCTpj9jo8QCrFCpoHyRgXr8CvFPGq5Ul7xEOpIzW0SVPdJ9QrblhIxJMVz
BL5SJ54lKvp/Ft2+7aMUkPW4FpCwfNweXIGsIR4G7g5hIuWsrYysLrKjyAa+DbIBUuQdGEt+/0+I
8BRybBB71An2uZNEK7V0g/9NaAYWquiH84NJ1LmPMZsAOmYr15rxBMBOZB52yCufvxzpTw7UDX2+
kYS57AwzE5p9gw9oov/aXLU6jMylFdNNHwqHhg/XJnVg2p0DZzJbTni8QZg/7xNBbqqtndlLUSJ4
/oKSNN7z3sLqID0lUsnQsBsmZ5n6E1RwfjUxaU1nbFZ8jF16VSSeOWWlRpoZXnCdh8FKoKlhzWLL
UvAkgr+RQ9s9OKjkZ0q6I9jpNl99dRgD6sGLap/UZIwp8RU9xvs1zz1Ok0S9gqtkgGAQTeBWpQ1k
EALc+bEnyU/3FVhSj1/T6olCv5VBHjj5Uob0pKn7XrgPdCaNp59s1nPEzW8DNHrE3YpkzzZcuavR
VoPbp5fVTBGtOX1/smsA+RKvmI3w+SZr0OjZeOH1R/JjE4pw9tMBxj7f/9zRCORkRGxxMfauv/il
+c4wyeRO+KPNSc4iDqmgZ9PkaWARjrPnryct0lWCYAhpoYo81WYSDvlLx9GQjY92GLc948hGQND1
9bQ2H1iKlzU/3KwLQcwnm8yf/vrX0Hp8xb8XGu19MrxaXXzaSWwPeEtDUFNxvfdK39byMNKyediR
iWCppXmS6PIZTt+u5GdnfUYvW9Sw/Hb04YdObBiZTsqOKPpaNwdH8HpJRn1VgA10b0GAggfXIusr
g3tISl9fYPLLpObID1mLUtPsR946wq5QWnw1gWsR0ukMetXwG4BzrQt1rGNfp8UOF+1s7IihI97O
R5S7N00Ou29qPWoVd1Htk47Lgm/1os1UlgQXUlwXD5WJUMX+ldqQEs8wL+9ShNL8TA7GWQY+3C3g
+ikvW4F6PeJ/Xfw11sKGQsboyukWf18UgfXeZFyuc11Ais4l7J4wOWCRR9AuZOzaKEwa/dxBxXsT
x76H8LtvUg5lRfW83b/m8/N2R3b3Xc75HJ7y0jXdzAv8JEkBGe+kWG2J8DMkgWrsKHDSiHrRxuGK
BAOJ/gtGHQd/yC/gO2BdLN3uyZBPaC53Udqn3s53RoZGl9FGrZr9+5QCMSbbVkEB7CkyaCr7JrEg
faDhd40E1QJNJOvd6njBST7qf6ySyLzJHKCsgKzf450bbxhHjL3DHCZ4SZjbIpsZ7pnLrJ6PlDdu
1OgOgzqTGS41fGhGqamSjWveMyDQkmL+HcH2GsdWRveiONySzBnZ6GMQd1SippmUscr7TXPM2JSg
arplLUGhGOqFMMVkUoJn4UnME3M/n/TscNQE6o3CC+fIyMHXd0lPC7DNQ7fKANcQF43Qo+Za8Ldu
hX15OuMrNj/m5uHehmur0Pt95sdC37CVdTiEMm7QENDxar06i6JIWFpC8cSzuweiFtCoDPZimxS1
eGHUToy61nKGG3jCgtfagbGxVA0oLAjvlm2lmwpr56FKwXfBt1QaNvLGa/TtU3x/xdwFDTrlCZeK
+0zXgxlTK3jXhw0N58ggahWAE6CpMj5X4V5IFx6y7cSqLWFGBA1yrr6+4D0mWfvCCOgGDDPTpc4z
CGzN7c7Em3TKfsRREsGcTxJxYAx82r+41Sbt327PXg8HE4/eseDYDqlN3+DnuyNeQDOlkLJiURB0
JoxQBtEc8Y20AvUltZo3J3xpynQGPduLh8AXQjBlNtJPKRHXMY2vWItSQ43DqWcfq8EldAqn091z
KX3P7SRTHyLEnhE/sPWVZQFE6oqhUFl1wfMDKEM4h0swm5GECE9nFqjVi3iS2jUyut7nD59HUxr7
ZeYusWWishtv3tfyRNHpf4Md7BoV2RexguvDqe0jwJCnuVEdxeNyZrL4uX1YsqZztUADGOeeSsao
Q2JhTSs7H8UEZZBAhXirnseRMwvBv5eWcrRXalGVZ2Yb683dB7HFz6YilgeiybcjvuhPzRcE4Kjz
YqAcmFIuInGmDh+q/fiOt6J+IxZ1r5Y3PFzatGOjxQRS4xg2VazBjpCFA5JGpgKbIEWY0PqmmAL/
e2wRWoSCb3+TihRxMNcgwigQKrE/D7MKm9Yjw06dsvN2Bnnr3X7Ch0w9+55eTzTRK3j++DxDYqOP
Dk2qQ21cN5bC8By2RUtpdJlYoSzAY6kPnte/11nqRlqsYV4X8Dt+q60z012ZxSibM53YM0Pri8B2
dz3ZvClQC+hcbm2Xd8ctZD9N0NL/Re/yEUwpNfdRKGnoDcRNQXsZQg65HRbOCwp5bvfGmwf5W3ir
tTivJsJqoJ5fBLDIC9YREz5spWDsWXWc1eFcq9tQ9NEq8lvY1JsuJ1pU1WKkt9hRJH2gtfUS8633
OGUN7mIp1iOMU6osTkh1Sn9Pc9xr0+MAL8xCJE+l/ayksRZCcqGGvJ8uKgTUqucm1Db/Dxb0ZMOQ
oeCVCxzlNDut51G1eWlroA4rlcF86kYltiHeMZ/1DuLK02y48tziKiQv6OKkFaQNWZJb8bX86yY4
ZaPk0zfWb764EYo7+IYwAXcoz2WIN8yPtkHxq9r1BrylhmypmuBQrLV4q8CuWKW/SCxV4btLjOPy
QKWKnpy3yFjdeSadfQX6Zd9R8tgcbmU52o2xP3nZ/yCCLyY1zKUiikpIY1j4sYYxslwa4lr07bUq
btibz3B7F0g+HYMrfdw2J3hjkDltWqT1bbUxK3zcsUPp3LpIwjyA3wZ2MTi8SZhvr12O69ztIjyc
fjoS/Q4nAZvtiEYiVEFybl6BEh2JGRMAPdXyYh+fdYjiilzBC4+dI52Yjwb8hFA+XgvbJWjMRLc2
ZARpiRbHwJf7+7mBmvf6Tm/eBkakNytbG77qnVIUCeNGn3p2y0f3bYQ53LuB4q+C0V+xBnC4ejbZ
S0qdMcr1rx8APdzKHuIFHf/24BQSuLhF1kOzs18Qo7Qssc/eNI+9ksUUMldtTPuDfZUoAbDTT2n8
UwGjQq84pGFWh9YQpTPehQJkrb+kpXa/8FW8yxJh6zheWySjYPqIzTdSyoYMVkO/kzn82WJQW34s
2zpVIO7Vk1EhNSwgiZmrkyQ4XnbipXHBZ4ADkPU6Kvn2+SIl3zGrgrooDVf4IeatNoNBqZFmF8PD
SSr2gQQmLX1DSdRf+JtosrSsxvXpJVe+XpcMBiDbgPNnc1xP3TfpOQ04Cn2zIfBg5VhZ+/XKOQmo
OWRuNvsqXdWrepv0536SJ6mLulGdUWwon4bdy3lFjRUtumlqvuCD6sTN315Pntf8c6jHZkzpx5HQ
f+25YubJCF5hH0h+KFHbfWCWLS5/hDFhKD/dpGWcxYaTE/heD2SPCY95AweGOZGccm9obNP1lSJo
AKN7mu3scMLW9z2C9DOTBm70xseimI/9vFy2bgd2VzkozsHSeEGDPYn/xxs0ognRVU4ux5wWs0a/
HNRxtz8kEoFJwNrXHHqYJCm87hAvVJIrgFntz4eEUoCqTfUwxivsVIcwRXeN7HMHcjzCwHmOofhM
OqBOVCBzruSnjdNRhoL6EfCShdq5b3dSQprmyxajCT4FkUN6/LZRDbUq5zebxEiZWoAvHLtBH9ag
16ZcvId1eogPIERoUGPedLkONp149wcTm54LfRyyf/D6220ObHVnTZBJkOSEj/vFKyyJYLmk4JX2
3O10BdpfiLZaxqS49aRhAhZ5UYDvWRLm9qGg1n72tYBJyDIv6po4ug2/NzvabMG5U8xP2wRYQvc9
4k3d2Fd8E/bzNNMFwlozfWujDVorgJMq4YfpSF1UrfTruJE7rb/6G/+qOUXdAXOtd5oJxhsYJwUH
gPunOyJFtuDxXaklDQ9h469wz9nvkWhTj82Y7YiidNcCGWWqRTRGlv3uPBqNvzdMRI1OzpeBKR1f
B/7VRN6GQyPuZZ7W9bRWlQncGg7VOlNcnlcF7V1uh+j7Tnxy6Am8AFc9+1F5s9eSawroRmu7lM7S
W44Rliey4A41b7gYlCHuvfa5zawC4JGkMOfXkvBf/wG5+nSPA4Z5O8M1CaMMA/IBjZFi+yacqn5X
yrA5AqrR+nFqYzgKpfbwKrGZInWdBzzoulQUs8YX3ih9T9nrnM70xCA+MmK5tG/mqcFMAMWbz7SN
tmZu+efMLweJe4SUH+EEXsWYHsuBtHMTx4HkxpSVP57IOIAjex5FnqcUX+voFav4jKpZ50XO2y2R
F5oVysfZTkDUAX+C+cTCXBv6hWH4EqhODG0AIxTXcRBzEAvLs7TUtgVfX6Y+nnDTCZTWIHeQ7Tc3
+iSybwlGrAJwfv91wxx2psa4E3+bUWTmCMw3JSZm/4toNYPsgvTtchgw93r6Zk2R3hKCWdwN9H95
ZpCxHFNJqMiZ8rDtbwx0Km0NwnWsCywSeauUGxEGE5i22FKPN7jzmJPOpmV6e0yMFJu7Uooj4UW6
JSPEB/7C/Ax0E9YMXQwcX4PI3kfjsAfQUwN8PUpcDJ8X/3S47WFcfqbXIxI3evs+iJXZzAkFKmg3
UaNvj8G9nND4qb/r1iZxi3UcdwcnOoi0wB3sqG1VMOPsM93YWjzGlNDNuyKTNG8cyj5TJe2ueyVU
qb51OwQ2AJ1JyElbyxUzQsqjymWIughiQ2XFBvj9dVMZAhsO6igh75vGoCVXIcWDtJYkmCXE3P4L
HlVuiGO9VQAsr2OL39KhDxXq4BAL60BMp5qEP+ykzbaJH8Did1rnH2wf677M3GRc82dXBdumdguH
YH9qy+i2G26xVCBDvJIwk/jDsXSYFBj3lfiYvYJBTOOjPPzqW6rnhOlphi6pN+9j05HBNpgebtra
+7RAj8kjpQK642x7jObVYztkJdia7+Cj4CIaD0/G/b1p6GMw/NpOgEj78xjHUZHoNSHkhScFgH4m
3ZPJAAkLT0XSM2ppU/80/R4NjY7UqY8DPI3wIg1o+9JIvtZtag5qh5NZXJ2aobtWhHABzmBHJdcf
kwSOa/rrCXZWqa2OzqzDf0esc+uB/SxkULfVKKhYj94InQezOiIRUMHnp3gBNvu4fKFrs00v+5t0
dqGvysvavSNHUC5M+uAxVmQt0OukI+hwXSzTFsaZi8FZ7JVIvh984EfEH/HrSedFDSGV6KpxxVB8
bSglZyiWKhWgoApTEX7PCMyPIfEhxs0zvJlP4T3vCFnt5E2j78mSplbK2EYlUcSX2HktvuNFCHon
CckK69zoBfqpAOjaKWkvrNQ3FsofmCP4t7pG4nNyUAvhu0ow2XqsuwhqCvXIPUfpdj8cEogatrYG
lo6lzeEiCHudbR45Yu2a6vrpeNXi+steb5FzHKwnPOAQRE1JkZenA5k/qWO2WGrlJfGF6/AEPQs6
u+lIwDu7IP/OmMG2lU9bIexWRyYa4s4k5eAikiaIJKlGslwmV33KQA+HB0KU/bjM7odMeCIbYWeQ
RK31eoC2HDCrgBL6vLsI6kkg8/LjlAIv5pb6XODMlzVYgRAk/SxgOgEUe3+ia3H6YbGEYtFq4VZH
JmS7eZ24lia61LaCa0ogxlv6y6RuVahdmVIibpfVnCXyMoLTwuMUuBOOXwbdr2t1axUZfHHU7YXx
zuVw4Cxbbb/V2PT7DKjtNvLKgW9ePExakpexLLWBv7NY6owh2COKHVEj2mdYmUPAgrxigedxw5U2
xpGmtum0LDg6VZjw/eawx7fSOvQEFtx/huONP3u4cnihUAsVyuC1+nq32AEb30JrY9Yy/RddONJR
d6HVKXeGTzOkJ9M+/C3B4DbmoaTqxuFp1jSUWBpiD4mhg9pdsQv3wX9h3p8jWnonxnJN3wCLSAH4
u3l4UIqjeUXFp/QxpWlTNsVc5mx7GD61ZBR9+wzzogoN0Va/EQq8TLEaAcYKrl7K+2ICmMCodW2M
2fSnet/IT1FJFPq/cXc4SPZXUmaWU0MeSxIRq8NtTQMoO+8yshvECmoDELt+aSjq6ziaYWK0knyP
YCPiRJZiXMyDJz2z2iNYGz7UGM0cxf6jQ71rXlLtC+s0QAnpfacDKuocJAarBetouCjKjtPqPuBU
DrOTXMLB7ks4b9yMVev7DesDmEB+6ECpvwznhTmiuSTdk8aoWuDL4oDOjOote6uFeXdrMGN9yNO6
d+5GIRj3LDusJWV+cSIIkWn4qzvHlBMpGxDUabSKW7aiyS7coXhqnPPFfFgV3FaTQGjaFKvpDEcE
JthSQFBQkqVF3AO+KW5HysbGObFRehVw4voRuauTFKCEptb58vqX1i2GcOqtHvVainTmE3nNnIWD
jlbAVJAW5YpRcg+ECJEhGt5OIpZ+1fs2RNbDw2AUpJBsBKWb7aY0ra3w4uXdHo8Jmoyrm7x7ALM/
Q6HiOpbn3AZAQtS+P9/kDROgJm7Ny3QT9u0py9oPS0RHQQmFSieqC/BHPFVf/qu/tnv9iIs9DYnZ
xYhIvNsEGZ1kHXjrvyIu8TI9Gl9q6mewQGlz6PrpfbSV7+9wMk+A20OEKa5sKRnsSO8lqiEW/6xr
9rHrw2RmTj8UuOqqgIqGQ2FCirl4II3TZg+vRgpPozzPoboQjYTxkhejxqCJwdgrXYN4YMyb/Pen
11sksFjE0nHoq1USLvQ/nVgXkpt31HfoqAEMPWvW05kTfvvX8xyRCiOUaOOaDi2R1vhpvy3c+9Jt
eKa/q1eHDzmYEHjcOFQlQnhh8tV88KSSCwkrGAiz3cO27adZ+lsawbh/HL9H9Kjk8MxjSwinr/i4
NvufNh5YC/XQfUWuw1GfKFHPm/GmMLk8XBGy1NYsjnaB7gh7/I+r9yM4CakeZccW1JF4ocLKffCJ
JfM95CrszTKRm43fq/v2gUAfNmD/d401vIWzBi3BTEgrhiodrOsFDDK91zCep8ek3ilNZMc2mc7w
Ko8/oTHba4iwHTePpPBGwUz964YA4OleoGpvoAc1BtznPhj3mIDzh9GFI4cq86uE1rOVRKKsVBJx
SbkA6bw0lSTPCwkfXGm4dc4FhpbCgHvpiVDN/vTvZ37nAp9EntMoChwkrpB5OBx0KqvT6fF2YQCl
7VX1TDPSf/VoES/2oeLXCCD5JmAQhOfxm39x8W97/le3PA7N7DMQBjcfXtyiYR0WGiR1OtmlJL8Y
0pkn11Mv+nJB2KcWG5o2A7vh3ZOXLxt6fxQfvghfVID3MotTjxmNw4PfvGfXvb6nQrv2Qv+qjpwM
C0N2AK4+nSGcx2+5GuReYS8vY/hdwegIfxC3xpi0wCZXEUxl4ix/fw6938b8bwEgZ1EMDNRa8SKH
ycaq/aYq2EMSw2eBCi4+A+G1GUEGd50p/tii0FiN04dzHbJY3DyybKc2cUl/JXjrrX09HOdK6MyM
8RLOI3ehRF35JZcgSLU955NVYiKJUTVNRtPqXMjJurm8mBJBgfcYgFNf0SECx27HN3qP5Biqy3u6
dD2f1BEJIItRj3YGh4Q/FO083zhoQnpOzP7lsz/6MI2KzIWW4XhF9cSnMB7s+KM6ph8Ku3MwQ3jI
DxuhZ+8Dr/KIRfXigTUEp5Wl1HNKQ1MZNfcNyLJQE0qaA0DuTShMn8LYhH7FJv1898+Yz+xX52rl
p9dvi5ePZSpR+fwJMhWok1uiPi4M7VbIbXnU6uPjEjGW4jCO8fjPgcDlvc9PUtc+pjx0SHXSGgIU
yC74xLO2viDtIVxyn1Q4TxE21un4gIpUSqDNsSHPxerxjihQJKRSRdkJvs0jbzCV0X1kpBy94NML
quqN1ND2dz83orzWjgqQmAq2U8v4viTzqcVUWTsgvMnr9JQQbTssfpSxp3vAoLNB37qkbCMHGOcq
si/olGZRztGnQ72VJiZNQR50MUFZUkJc+zEkTqjueDpZx2vCOwYVCeK4y5zQDCIke/A88H6+dpmG
8hy2AlcE3nGKItaQ/ig7ApTVRP12hikGXf0xknhVYS6t/lLnR6Lvp/L3eAdJN7m3IJru0O9M9Nn/
IGySEBkhdnTuoRdk9vdrrMVCZ4CADRquwId4Ba8lxk8qtkylun9tP0Q2GTvjqFmXZvOo6xgPDRcH
zo8djjqD/cQ671C6/cU0SH2gficnNsvp055yO0OERo7QTNn6n4nzHq+16PMWPgOaQgBIrjbNmir4
vgu/6UcGNB0KWKhHgtqSDEgqk96uYGQqZAxrkVA09hioi9MHDHvDDJtvCbjp+6bq+zGakoLdp/ZP
4w6SZgxqCZSlc785/sXybB8OF6qY/961qoi+JfvOQlb4/RKWKpxNkDEMq/3lVVZQCs7cDjxzsEbS
3pJY/fTi6VV8pj34RtLwuis5NG7yOhT+tqbSCecMbM7D/Wdf0j/G2lY1uvtzWD0wM9FJJf1ZCxoY
j/ZsBxMb0XyQY8hmI16B8LC91r9UM94jIoysb7olDYc1Br2vU14wwOFEGQfsfn17rX7hlOPmi1Cs
/4lKW8IX5xu0SmFADipjJNSNlRwHVrB3xZPwv2zMJAocxtm894ZV0v8nt2ig+QHsqjmMM9LOoTrj
sDb+IpQKHTEsSD84WgGBNk5vLoGlE2/BFxanPtzIuaOlZMODki1oFTESThINoTC8Oax9F1wpO0VB
OlpZhd3UqOq/0V/QnYftJewhoN2LbPANel6qDi5RYTPvw3dDGi2oAJigAridPL2FIJOHprfQAlO6
svzSOx0qDXvToi/G+sZvD1auJQfLDXNlQ5rIuU/XUBjmg52nreCkBH2nNDeJlrvI9E8SRrTmLLia
FWOyuF7QSLP1N7uI4zUIRRlwEQwipyuvwx5ApN/GkFEepnhQV8CWfnR5FxGXgmGzf40dgUFtbWBJ
MTXkwCGAeBq0hMTSDVNBpq9F0BUGeVjRfj2PmoQn7TbHdFsBmm3iaAbqbLJlyNeaohz5bnAOefRM
j33dup7TJ7EnWwanWimXZxOzYyJzrpmeCo1bjUa8qFNP0E7c2JYVNki1TDKCTKRptXxYq6e2Bx22
NRp3OqJxTA13aVjRz0Cqm0eaWYPOa0pE7ayCZN12dh/A/szQ5LcpT5Mfyu7n5cPMyq0zxWB4N4Wh
A4vpzADEg3VEYCI8jm1SbVpYtjBSW57Ui3jL2uJjGTDg7TGrJiXRQhxLIm1yl1USptp9p3OIgbzc
pU/yhUkJ9Aj91GCGANz8EG3LI2EN8jHhreORET+74tQ+NdABjxXr8MdLpKXG/Fl1kjmMj/MQ+Z/N
667YtCRVYMnOFDroLsxIM8uEpMdvlczaP6Bjk91UOrS4npGnnmOo7U39dLaRyNWokf+PuMys3Ivy
P7FvFcuPLx4MRDRrr0aI/3F6hySs0XXgCGv6QgC4f8tMr6OQFCT8zbA/fj6GCwYGxr8mCz++0i5f
X4dROVQPflX0IItxaclkfP8vpMopWeibE4pm5NSIf5bUvc/SbNLplgAe8div7gb3EuyfaS2yArok
8twMQTckMzuju/VdXAlj1CgV6c60tFLLuQRZfGRCW+45ZNmyisIyk4sGGgpQMywmX+AZUDFxwDR2
polu+uCOjryiA2LyIKorm2q6aMJEJA8drQotG/CeY00Ypo90C1zT3LCEl7rnwye5lB+6FWzXWN39
+n8H665jxSjjqLuobhiySi9iz9Uk2jDNjK7/8keYxGuDCzc48RevlDqV85RswzaHTgEwLaAS+Fet
Ma7WBjIGtZnsto6HUWiLsn6RyRwip7gCklcHWVdxerrEXAJ34Z+472Wow8r7//ES5Q/9VcEk+3ie
KqMlEyL791BTsJiaM9PQYSMuDu2IrpbHQY1ifNP0YY8+blssH6pXGMtHy7gcKIMwJmaepiKJRxZW
Fi3jd0sZcCfefh9aF3KaJJuWK5QHO3LLgm+PexocVr4DFByeRGO7+6dqYgftcRiM/VArm1uGfMGn
SmzYz1UZbX81nP7aI7lcFdMt+UO8kU4IOsy2lFOszxmkT9eQ8eJB79CkvlUksMogjZaaGwgaM1Eb
isq05gyXEllN5QCVQxL8AnD7l8haTG+h77p+kUP8pjnZovTMRFTqEoxFpF3/T8AjbRHH2sU2xHqf
R/c96AIl8Uoph6xwAQ/EBDqhCGrN3pugPWjdxX/+QzT0FC5X/kG1U59lGroVkQXWZi867uiKit9t
7RGi130QZlNOwH5WqPvH7oRLYS4DK+Cw/CQoT3FTZBsHr2VoHF5JBvujT9zAEf5RDlx96c+znRM8
HzPk6y8/OmBblQUArZr8nFTZbIim9jvURdRzRIsQ7ImVKJkk+u/+SK7jSR1ZM2bHjBOSgvpIaIQ+
SlXsi+O3DdCwNRwATPKHnabtyuejQuW1tVCqg/LoKTOkKYq6tSIw53zNjlHZoRGQ7shUZg77d6ye
TJ8QohwfGRYg6BwPPxTpaDUQ2qMXBqYg0tRWgj2CeA2EijOXk7ePGayLyQlWdfN4r9Wg2dEcMnQ6
IGQCIUekdfS7q438/L3i2Ie18e5P9tblZJIjlJRD135TWkjBVy0srC9GnVlTOogcWF03MCBEt1qW
DGwhV0bQzkea9UZLGazPLFOWxaVqU+5fWApRq0HOFNWq4+CZRDzimzsDj2gdDLE53tfukqIfOuIk
blVb07yK7O5sf+eYzXD4v7Tlv5Amt58s9bBS6/RTlAqo9rM4OJTYa+bI9h3VCAz45KDzJxHYTB8q
p8qJUFwcQk3uc+pPcazP9dUrFnnb04sCaMu0Q6DSQ3Q1UVInpJI5bfZXtN0PHz6VmGjoZ5NabYOT
SGDUVfrECA5Q1IOo8205bl6JMV2au+El+xQ9KvbIQheyol/JNlApRrHzRtvhveaCy7v2L429epfZ
WjdyGmdnqYxoNs0LPUs0+6VLYCR3CECcQvBA+iNSGDbXkacxXkey/wG2SaDl/PbUXD2esOZ45Xij
DtkoaN/pHvgkgyAuxxthZ1vcW9TlNE2kdES8qpSe2Tp0GGN6eGoMweEPDKv0yu++nF0KGf2Mu/2f
Lrh38N9/dvGa7N2UCtLCxuVj/m2I+7D+WgcIuHUTekD2ti1FfT4pBJrZortA5b1jYDBgHaRHjfWQ
+/uqFdJM4/v9NGMyKO1VRaccAmXEK7yDhYcEKyLrktLhg1JDHFC9NEm/r6LewfvbIXRTuJ/2X6Qa
bpq2pFkweoEjdNb9boVz9wyxcaa2VtQpTr2H4X4rjIR3MxL/yWH1m3whYzDVsqYmtYAGc9H4uqZ3
XDkG2Ga0jD5ezfOLT7ons7ii4vQvYEEZVHnKv+wIjw1jLcLiQPb/fKM63njpquorS3LxrfoyGSAx
0720vFflCV8dPgyEzo9hh7fie2YY9tW/cQ+L4fqCoMEWCh+zWw6SNOXJ3Wiw5JB7caeHRyZNvEn2
6cRyHxx+DroWhr5E4Ev2xQ2xiG2cASUmHf7zA7SY0ljVxcFN9MIKubZv1yuW8qVNa45HHAHedTA4
w0jyHKo60IcPbzCk9qgteB9BsAaShn3j5mAlaQqMOei7m6NJHh+ZvCYT3YEX8oNmFp5DXOaLsdy8
zWn13mqUekCpSRZeT3pK9coHSTP6DWJC9RxTp2ycz7bAEW/4sxH+dcp3JW0iEhH3Yc6VxQWTL4b5
2MrRbMFPE/6Fa0ioLvuhqiKoKwO51hvKF843MtD/zLdJ4sQcjJOZCk68eSY6jwCGREinZouu6Lkz
OL2SRmrG9NjG2eAQjH8aWHF7melcbrN50jCHIgGH9YXSmzNEjTiYtlKpmPEBjgxHU+s23hiBm9Kw
8jPqTDEKf4Jr6DZjgBQXhe5N8FWXSuZkM9mrMj+EnSb12pvYEmmPnpa0r8YSNFZtPAYs7kIpVRnU
/JNL2WGlc3qtI881Cotux67JSYmzrcsfxa1McUTG/PAcBlOe+MuvXQFUsFLC7I5rhqYOAQY6NyL5
Bm1Y9HwGi+IAoDMMTwWpwY4iInQVkOYh20QveScObKclACbUxCgFnoO0SpH6y7bmMo1fZ+0tyYid
P2wsg+yf84Q/Fcf31hwhINYeGsdz8S3gPWTnKD+/vYeL+C1VVijrP1AMm8+DTYCQQvaaZ+EwCZHc
Pc/h+Fdu2/2+7nqHwayqwxspG0sqbhwIgfI1MclD5nqTYUq8WM6oJNldtYpa7q07HONLA8Knwjld
4NeSNXuLPbOq8udzWeEjc7SBkGwExI331n4PaUmPXu6Ids2Q/meBmNf0/1sE0nTiCqPpGKP++N1l
IvSF5A0BMbS6Z7nzGrqfJXMSmydAH9IVztfuDfl786DUvjYbwNWhSeGETYRf0c/RHmbBoRqwwwPU
0RnXUXArMvzv2IC0YigKBe4EEpwwKpYgl9h3K8ocYOdG3DZQoAAiZqxOW/9sRyxN2HFkDFsbTV1F
ENLyOiI3C060ic9ZfLcHtK2mds9wJgzF7VxD5+YLRV41PFaGQ50Ytwk9Dge3tEnKfq3bXIrEeWER
dlky76zMIrJWJ3HCe6W9T9aTmVrjJCnwrZ2Ne4yMWh77/+0CcJVbUjup8nEhaNLtGs+r25rxOr49
H6dG+Rjfbm653ah6PZfNE7pAzhofSAFKlu0EYUEDr7HKt1oZM6eooSprtSFQ1DomeWv+daSDgsMI
dayxb0dHXAsmwd55+8A6syafhZaJCewg1OCepnOTXNmtp/o+E+LD8Oe58/9wffmdfiRwXwyQTwKW
kIJQPA74ajPxElG98sl/1Xoi1TMmZoqfRbNg/QrukO1CYkaMxkX7VaxFQZlmWWmMcPjCXJbG2L+8
gkXKaQqpvpFfxHvZZcMTUzTWozTlHXUs3p8585Zzzckd/ZqGXKiZoeFAfDhyhk4jafygeZAWrvlD
RhUQkEhDWxIxW/N/j7Bk30Od9bx4C/nd8odjJO3XHkXyjYo4GJJWoKEUMlHuTAxJ0ebq0o/QyuaZ
5p4ZR2l652+Zd3URQycepq7JQSGpiDhsiogBcMNZTp1+ae1KouirmnVCUVBfdaTaKaAkvck3+TLn
zTEZkhXWyA17fNVxS/VqV0r3o6H2ImAvGZu3uD19BVcTQHpk4LBoTY586UV9WSg5xDNhytzdWnH4
lYVREDKOReTI2FJQjrHDHFBzkHwQICLmiVlCzQQwrLjwfl+W/1duBYJE937+4HqH4q9Cri3S8Zjc
VFBNgAJEI+FPzacopCLpCSoAc9WOxJj1NqCQyXINzWjBfYZXoodFqdNzmHpMGgy0/vJvoXRZtCUO
9hQA/JU/pPG8Y319YFKwM4Xlt3/J211Ap4M4Z1Cqu+GL+usVjV9QZv8YIkq5Lnh8Wmxku373FI/i
r80uYsS0SW1DuuKWX6vJJMxYWcP05PTLrsHIJmS65ro9+GRMNqJ8wD/LD6b6obcB3tJrBipSoTZX
HSMvVQVOq2kvFS0FmPXwhCX3w8Qagw0C8q4i7zSuaEdWaXMarCjPfD7BxR/dGw/7WGbFYdbJNcu7
cHwXZcKRS1JT2iOmVtyAIxAxRkVMXQg8hAr4EB8mRKq8dytahSphP0QMO4718h4/IcVXvOdWrSNq
ab6NcQV+z9Y0aGQa6JgyqxK8vR7xWU/P1/3cyAS+oOPKX+x8zvh0ut5KTxewIn+WIcfrcatDdmub
HBf+4RtvviVuN/u+aR22NgeTYToNJr8OQgocW0qzZlAwQ6UQ378va0nFTeEydtLRyrTZeGFyaQS8
MXq6bVVpUK01d2pAcO+mQsDGWFjIrRarlslGROnwDRlq+s1pObN+irlB+OlPvDr9GylDjyR08NBR
zcKYWR+68x+gH0G393X+zv9YSDVtKPSBs5/3/hNveiuh9iCbp6PvXX/qQMxWhic64Dgfkn7HWNmB
456PERdikpQjxrgDcrdWwGf52sZlC+JyUI7lq8/DWTSTQJ17Ceg/1JeKDMwj0kvOWDVTUPKuVXKv
3J+WQaKC/HRkqK857iex6+xgKkFxGV951bvws77VpNRfqMtcI63CRyHAAHK8jjnAnSrGRsJT60LM
Rb4GYf9frASc/yQXMTmtMrd4p/BO1WCyzQNtGpOcxnQuAgaYfVuVw82prIqXCyiCsay92DGqtutU
HjRfU65bNCr9SoMq4h34wfn+H6H1FFO3gy/d/NZhnEvqHLPa73VcHdir9Tbfp8cW95aayUKEIiCc
uGZTLf78ZQFe2D22u96Cxj3E26HA/abdQr7iJ16mM1qLc6dHno94sF86yh6ISuJtWPBbfoeCXkcU
W71ahHqHdR+DwV3gYvlgQ4jBCFfHwRhlKGoy4EVJ9xzqyPoZvvj93YU6ZvZE9S1EKLu55EyhqrPj
buKFmxcxHivLT9fTcuhG7BsvG35PN1zFjBDRAFndgLlgF5IGlH6XAd4spdHzNojwJEMz+xWtOTIC
yukSX+lHrQN/r3KlsjjfV8R6a3ltH46IxTRKYIRhJdQgB+53+i/lLbYR52qyEv/VcKmAcYf4Fhpe
5bQsgXmTfrBQX6kbkAg4s0Rs/mWThtBW+0C0c+P7vZP08bC/7jhQ2v0ZHcu2Cqzm3mJ3fClLGXAB
O571yiTFc3RnX5Zz3TyNq2uWy7SIVmU4BmbnYcrCyxj+I3VAlZ3wKG6vRYh8d/ehlW7ppse/pudc
A6u6drYIh7oBPGg+hRt7SNazfFLxeoWATwuGY88XlbsFxZIc/Op8pn4toQy9enev6dLNr881E+Zk
5eRE2I0ahlLRbmtBX+s8fuo645Q3I9V3rWsVqXVGhjOO40bKzObnxhIc7qvRmNHNPeRpj/GtH+Ss
/8FjA92jXXkZoWZxwiWvlYCHuaxPb13CfZfkGzWAsWLnbbtTjapN1MmxURIFgNeTWKRnDmoOJSPR
vOsqRINDYgZEOAR9+CD6UxIPtNsqxJZ1XN5FBmaKZjsnL1YlbZIzcStO5Z60xYCQrk62cgzKc+CK
HUthch1TscjgaPonTQ6flYnUCuDCLB4xKthIt1COnuyTRWvoJ3OFZaXB8pWQDbNte/W4mHI0tYM5
7YwVYZA6jyB1Tm4pC3sbxxoP715FqDHD+RjEc7M78Yd/UDN+UBrxtIoZpBOVI+49EgqzfKgdntfZ
ZiP1B5yBLQqG49/UwcxBExFkdGSKfwoD3Q9MkJ88Ki830OX3gJAkBqZRGtjn+l5RDDaUPf+QHuHp
6IzEUg/c7BtLaPKvLMFShDcg+OWTNCbuYhPRWzHDsi6thMa9qZ41PjxruXbFIGrGDYrGdHn9hGr9
W2zzeKwCGxGIUDO8tAL2TUJyEo8dOoLkwQoIG5ATetCekOPWCK2cUb3zC+yTO+gzpkSppu/Eis78
6g6aD3fScBxoj451u4vRInCsVdF4u0+PkVus35SbcTKBSVt3zXpEcCbjxC45Egn7KWrr14B3zlA2
zgh+a8kT6qXVI9NcJqMpEMEBuc/cP8GRjoeiJdI6NzDuGSEHD/eSnHA6qWkVi8LHkdsVnpk5VLgr
SauFEJxOdolqIt2mS6I727xsH3qL3XoCnGwT6pNWR/wNkWVmbQWDl0Z3h0HDW2s3Yzko7cPaht/1
WQmKcABSDrcTyZi1HfZ7hDk6iDoXmx9x+0aYZhcgI04stngqR5N4Tn0/cbKzf0l197bBALn5VBFI
/87JZO/CVqd9HzHZvnLSa+J1XXvBR8Mlfd4TaE08MaFkHH59CZnP4na3LLd4K8vhtQ2h4FWV1zDQ
EWlxdPBJ1fM+Hut0vAuROAybllWrkLUVSAPCPKQH+D2pIIe646jtU8xyZ2ar/Sdh/BNLmwbIJEI7
9qvaPdnb3oFln64xZs6puYIlwbJDi58QF4wWrQPcbD+G3dq3U/crj5p+0IP+4oJVt/pUm7HJ+E7u
2wcB+S+xjKoDUjcLkwldX5J9FejcNbmFW/bSEhRZLadO0WEngVKy7M6uTGyNob64slBUqUwHKp2R
CQYfzBPWbe7hjrDbamrqHKWYcB862rRVnr6inFNwuWiQz4BVh9remW0tHrD8dJ0u3JM0Ngurk6/9
pO5VdhU1jTaIuXq1ErN3B4nL/B6F0ExOZfMuEHqgX2zCntRB60T1FUlQlh1D51Ilwai1CP/Y9OBM
h0I1Dryhr3KoaMKy9WK1yMsZQGcvl6E/zNF//0LDtRnI6s1oeU0PE+yN/QbUu579zKAy/PFEPVBl
FaBq1oOPhzucQHbTIyG4ZZDea4ZiXdPmnOrsO8SaOEf2hBu7Iv4SgiWk0CWUB2eAVtdhLOuOM5Rt
1qTaC5S/DabCwY0B7JQXunAYD4TpkJ3ZsxxfybFf6jNnm3aS1zf4PlkD+FVCMfrp2fdURMq292SZ
TPaAtrXO/LsC4rE03iLdczZWI3vBx0JM3POKpO04ZHR/kt2ZFKZza2NsTsHbq37lXdJAiD9hvdGh
oG+gUg3of1xZy7kaMjgoT3rMbMiQ4iNKXW0koJpM9gvGfg6ty1wLdb/cBBTmyjU8Vsud3eJvRdbF
IMFe0lfbYT5HhDmtB0slzNo66qu9e0lwdWzmNbg8raGl9FYrE4rVGQfbVvWY/5HkVz9/lCXoqvmD
Silv0wxeKgyRgaiIc9iZ9g8IMW+r8kbxISR+oIllUPNgc3ekTiLvsRFejSnES3c53QSslKcDY1Wt
shaeaKdwZC+VyZ4M6hqArfJ+gCqJq2U566h0iq/UR18lD44G9gzjAwFKuqfoXYFRFDparY3Mz5E8
pza0Ldfl+rNuWPsUDsDWR8Zo7dAVvDsPBjZgEsJ6bLLCd3fUoHuj0IUP7z91tseUK15mbiCGh4BI
OGJxZUNa0cSzkR/94AXs5MRWJcleoWNC68CZkEYD1wCoLL5b27Ckmt0Ju65O3BgvHUocvHo8rc00
N+NK8Wqep85WW4NjTb/AmuZoGTnq9H80ad2XB+6pGM3q0m3bgSoYOcz1OhVtCxu8bB9/bMK/S02w
5ZkrBfQ7TvhZORXof12Au6Mo//pk+SqNaHvfP8j9MQDNA3Fie6gh+Bog2YTw0oa5MLF0MSZHtjPA
QQQppT3RhBI03/griVliHLGVdXz22QPS8G1o0XGUVPO+r6oYA8lcW0DqBTTQ64gSxOOUyfUGy4D8
ZtS5SarJ3YDvFW0YJyvClmB/zfKsXFqmRJX4vB7r3huE/mJ9UPhU1bzfFDqgWG72q0KIgoV5QR8P
5LSutOG/DBbDGuwqMAaCJuDG1O/2udgUU+VfpsvGelSCRz51WCl9korcQg2USkQe9Tn/SU7AtmN0
E742rVFouqCZ9F3wxBs3YfI2dyJ/lnB5uBfLzGANQGTI3TLWrWi4zwIanZdztrsVfrKMTN0AHHQr
Lfi9sqlis9BKgO0QpmOhegtlG59VdSjGhQEdNrUrmH0FXQwOtM5qN1O2m3bt2uYI7iifuqte4RcS
uK9kXACPgudq+OKFhMvBCqXnBTI46U9VbPYdF59osoKqV00nZL5kqGgJUj2wXCvq9EWDPdfO+8K0
aFMZcxOFyC3E8T2xJzW42cM4eQDgMSTNUvj0yO+97yMAXewA2AUnAhg7tP2Gj4drPMoV3dXO8/LY
VZ0vxQ2L0FU5vUCTybiFLx+wzFohQwMybHaQgpb2bGX2ba/DZyRAIfYqXcvHsXrzS0kYpKMKdChV
2UKK+TsONdfAQzj7jE3O4rT4K+zdEb1nKbPnI2mwJhpvwxdRSkkEE00pJIQyhpPEksFt0w2VJ+L3
pp8tkk7B3I+D/Yl/0Mei1hG32v6GMl1HOR9rcgtt6jcItr0Esb8U3qyOj2U0ryp3+Ui3ZURx47QL
kmY84KOp/6PWrnihZzXT7ZFyyLa3e3+jEtB5g7bz/qqk+FJsfLFKIMjKiCUVDG4LilDq42FZxfCO
K+HWYK1gOL3i89Misw27DJHz4r1BvxI24V/cRUFjUKRl61Op6RcHGx7a70L4CExbqLACWtjQxiGp
9DH/FKysDRD2rUxRME8mFDTD5PQaVBTXpWBZjbTxwWQxy5vfsLHF+i7LxbR6VMnihV8WFduTK/SG
MzC9OBUWK98+TXBya4GfqBAImpgtmw4K0tYDC2wiLJg4cguff5eF48PvwxJjia0UucmgnuW8KaKg
DOLsbgk7pBiK57R4j0xCVmkO177m95J21K5IdWan0YRXjatz+9E4b5tDsXi0cO2hPBtiCw/uNFJN
2uuySApjzpvySeh1rcwuJy87p+UPedqPZ6h9r/BQ6M20J+y2vT+WLQMoWEGlUBOuQ2rVBzGZ6cdN
mKJpUZV3Gq63A4eSW1TH0LQKIy0CyMLf96KVp/RXlFc0gB8qI9Rxga3+t/4M58ye+Cqz6efvnjdx
0rJfpXZejimegV7FlY7KQ9CoiwYnXZMOukSFCag1JVP1Szk5gvcAZyEexxCR/mIpxRUUYOVXsHcL
9Q/KWOcFPJUViecO6IaEvBGMR9jBm37WY/4w2f/2AgCZnFCje4n5Q6JA+0Y94Fm4a8SKfKLx67g8
9294JWs16TR6k32cIL5+rcTWCnY63rFq98FShshC+Tb3t8ZFC/r55dYMlKTxufqh7dPv0M7ABqoR
lgFO1f2fBPHUKMr0uQ1Rgmx34JfzgKfIjOocunL7F7eVyQLs3OR/Lx5D7UfoK9LM7RkZ0T3r6q1n
KJClRTokpT4J3QKO6mrDv1x77TM/80ybWTd2b2CkkW6TETR+dO09iKaKnVoUfq8zBltp2E84MBGm
6IedqsUWcobjTZZOMcfpDJIC9NMbM0F0DGcPhKO+sUWIeHtOHb6pTSgcP7INUGbx9bmvr0KzUx//
4IaTjm/dkRbsul+z1IbuY4C1lUB/wPVLkhK8dQXxcHK8Qbek70NGsBaRE1opacHyeMbfDutaatWL
zBH27c4+AL/ubkHhTwg87K5dcuabHtgQ0Yqr3fOwP3TRvm7myafeEzAjml+kznfDTolci9I3hj+C
PY4KRqJqY7STEyq83lSrlORogp1D63z0vyOqci8EudX+0S3NLJIhZdJB/epAfHZkvHhyGAyc0pcy
X+BrCLKXmwhNEcx7t1fgqRiQQjSAAl7q2JYL9cVtdTPIVnJCHrvSCYoknkrOOLapcZjJsOZgFooO
kqSGXr+zsHpSA6V9EdME0s5l2dRlZEc2sYyUp8dEfGWvkaOKCPJ02z9ff8fazyMzicO2hlkGikK0
dNYsKiqzWnm27WLi+S3r4I9rWiXRxqpSg/LNUQavDm+PjFJuWqXwSEzBnajQlz2mg9nAEnTTbiET
p3pugRqe4+hei3P4r5CnwDUKBn0KwacNYmRQmwF2le/BrL2UuHTfE4a4xa78tdYmDqZJbdJ5VHso
koH7gMHzap45JSPQWSR3NS/izRS0awPmX6OLHzP0JShoFnLpIINFvStR/crt2wDkTSoEKsjD61Wu
zCPsDNWDozBsuSyq2RUYQSJ1Byljqnwb3zPGWvyH8rBUdKMXAQ3WLqI612OmThrBi0Fkki5pNVTb
lpKIK3WjTWcMJnu+U23J2oPxypqjCZENlaG2293KIu/ApV7g3wgI3J51tUlBO7jbnOlD6lSQZUTM
wYn+qy7EiUpwvcJH0XtDYY7Kr3vBLT2vIga7b9QxxOuVHOXbL0/qjm26esCzFBrRoeZNoDkY9rSG
VGh5sY/eqzoiguwBE4cOmwPOr5iuonDWvuFjxNA6dWVtVoH3eWXc3lR2G/JlN/rfex5qwOpcQl1x
p2uH/HNk5LHqtac22KxF4t+qmw90Gd88iq2PBjTziiXTUpqaXaSvmdT4VSl7r1O5JQvkmoXW+gd5
EanyzY0eAffNbnRlMPCx3vGi/HSGef/yiOZxGe7rVDPCXLzmMcPZkeRneJ446a1E3xI78f1ZCtfp
Bs25BzfeQ3k4lONnO1GxRswqD/QafnoKbo4rAFcIdhD5B10vGl7KzqHsxN9zIODw6YGWyDcLr8V/
2ATi+jh/a3X+bkJatyVwZUcKsCZ1ZvWNLruo99acfFIJzKIsbWKkrIF3hoT7jceq49jOiOEQixpk
5VPykycbi/UAlBlRlPh56Z4qX2pcp8s092GmjeRcDNTdWqzp4YRLQ6/D1v0iDIkLg3c4JYJKt0vf
73cDcZUXwi+mce5vMxJNGA8YwMGfnOKspH0wZzxG4URaUD4cjYY1IKUs8jSJXd0YfKfY/SPX7LpN
/XFbqRTpnJt9KxQJGj/P6oOGFpyEad4y3rbiHz+sdr8QAWr6f90YBnNVd1fUwMaJ5lDQzpLOYAiu
IP4mRfYErMC8+n42z2aY9QhlcAX6FWTKNH5C98UFN5nRkA57I3fxTzjAX98a8DUpa2ece3VKc8Xb
JIr01QsLnn3US8WCuJ3iX0ixjfSRXKn8FHxMUkozMRsPcSVw8xv5+DoP/C3uJJ2ACK9szTJ5TveL
+VpMjYcW9g6SJFuLHfPfAMIwp12BhaM+yM+uk6GLfbsOfyqhB/KADgrtorCD1zLNDJcNlCg37Mh1
9ohmvHhRx+xd01oNqxmhVngNjbcOwZA96RUAErHZOu6QySQW4sDCVPaYUUe3mTyaj2sGurmeexLD
u7AZ0L3k4kVbBwrtX/ZjecizZAommbF/MlmwCkJpi6KgcwdRUXiczruj20JwqjJppkKLzCXyKZxM
rsuxW0a/rqtOAYFayL8TrNH2BMlRLUupsyY9LaBqWClDFDY+EPCfEYt8RC1HtUUId+PMme9ihJRc
a6G+sc5SZycYW3OXwyviSrkRJ2j+S2QG6+x3chS6CVqYcdrGrE7fvWCbhE9dsCu4LatpWqH4SrTD
+xKzf6azmkMVDFEyiauWWxuVFEhzUL1ZLgeBIVYFnvjg4tvZG1L/MLyXmhwTyuyfX+hp/GtxOlMO
abrwhDt+Rb78Ecxr4nj3CN7UMpKbc8zQiyj8eveONcpwDvtnNYAje1kS3GaKh5gv0sMmGfBGO6Vh
M+OjgbnaTAmVC29iYCMfhlU4tK14uuAlgMMeDsMkVtp7+puQBLUEx0TbRIbDF3AHHvHaK91VuZ9L
78SsFsHewabCdQ+7igmG3wAGa95hfkf061R4IpA+AiVf9hoBGotpe2Aa+GxlRMaJDOR/317AG2tg
ZVkRXXxnX0gYiFpQ0ao3I6jrRKaHmzFq5tI5m0w5gq3awo2dfV008ivJU/keGWLWA+Tx86XeYtUh
AzqBbOUWIIwPZBkc9PuGUtvCEOeid+OVC9FUR1GFNf/DirbLB4AKb9ZXno6PwUMKz1UsIJeQpYYJ
KTICHbPfyluZgPC6CAoYrpyhRGOp0qdNRK1thbZLu9q02KxTYlfH05/xeam2WxymtRhCPC8rLYF+
lTuWVK35Ybmh3Vfv2ff4uq3kASfquU5xJeJ8+GO7qTwm90FgxtgXrjYiHtnrKQVecR7oNanPrh9U
ijAb5amzrlUJDT1Yy6dsqwJZVoGXl3OEQCmPyD4d0JMGNOsVFawetVt+XbWWVEPZfU0KqN9zd3rg
9zIIUMaRmZ6978bPiVIgdFkMvCE+7FijlFxTdipxBJWySMvFxNKJdxjBHcrJZybP1WbmnVLhzti+
5GalaC7B4Q1Ces6YDmGbu9ZTXLQ/MM97OBt84DwfuvRv58MlPdqWjh03bnP38Usl96ouDxyUnlth
5nr2gQ3kwojp5pKjHd3vPD25Hi/PRMDgsqgglPGbLCaVAVoBENma10z/HeXqKNYH3xzMM/VUYi0C
AEKJoKJzs6//MkaAY5DkQoZtnJyInYjFE0VclvC1OaldUeHMIPJhTYAGKF/Fsk2xOgRePQ++b4tt
IhVeJdPg9bcwYopI/zRWoVw8XRjW0YAsiIX7d5zCTXYPh3wxO41yWOTHECrEltxsPMSl7eRh2IzN
ioQhqQQxUs7noBKk87GmWWPjfM6RBIvabYosNIg9Y40znA79sHge1i0xboMKqrBHzMB5TGEfOt+a
PbQTGtbxPB9sLQcEohSIhSBv7HiQpzYNkuHXJXjeqUOajWrupcbBD9gsUpE/7f6dQTBJtFMLmy+s
PZIhIHQ/B12r84tpaj9FOizmL3oLtBW8bYL0H56uLCSiYs61hhfjOGcTWSC7tOFqdUHvbh7hMB8O
8nwQJhg5zoY2Vyr8+DeNNQ4PjUQOSqdoTTI/2i9cHoKvU6Q/G7ez6OwllBux0XRz7ZlecGogs18m
vBt5fYXP5OMDTpLMMM/NvCGw1UVh5ZO9b1kmTWmcuRCr7aGfYVQzyowtrZYrUwa5Ej4TlIg2Bazy
YYqdL4oX4drWjS1RDGq/bXZcVq4ihVgHKxxePX53d3GYcRLiEUX3sg1BAbNDGCdlgkuiPtybfGQt
tXoS+9kRGmVRSgHeR2gBPTdemmSwPo0q43TEfXSAD5gAwxnOsPBIkeXu4fG2ncRZCO+StPCPpYKQ
LDs/xlnccOxYQFW0d7nlTBvqCEtYxGKvEgRBgLDRhTyUxt9vuZywOgKbiPAhJ+3tc0YgFiZ8FHNU
9TYgqOnUFds8ZjA8W24E/q6V/XnhEBaHVSlNgQcSNmeQaqaGzTzwOjnzVzk+QioDJ7OfZIcze6Qi
qjDkIl1x8WRNRavxb7U2srjf93rc3YIVOV6s9qalIgywaq7fV1crY+xifuYSaSeS5NqGaH0aWos4
Ic/qo7Ik8Bdxzw9x6DXIyjBs7GnCW9vArldKSDzcQHXzpiJt390+R255s70an/v7jt8uWf0G3Uwg
V8To1EYbKcen4n3cFq+Hvjpmkh/jdfo6iI1B9S9S9CE/n1/KiBRgbv11pSMoTeX5fQbhS5VfCn9a
iGWys3W3l22Yfi0zGPQsUj58NaN964g2yXpsVn5jkoikI1kCCGBQ3CvJWz77cP83zO/Isfp7L88S
tYzE1lvN1/q+2Iq+EhyDGBZyLn/ubdO0WkThnxsAmmb+B+tSTNromClDcP+O0Q3e3gDBmQRlx59z
s1b1PovidDflmMOqs7hqnJ4VZgd/aOQhon9bdbn5PJAdBU0LPv8KAe6T6HlpTJxVgVBVdzP+OxPw
VbsLr13TGAwMsiH7vf14mzZIqTPzkADxfrdhSSDmIbTXbBIKGiAGKumJ3rqDRqUSRmnOPwNbpoTk
tJnnkXNxVo2R7i4i1WASQ98iZT0gFFlhU6t12BGUC2vhLKV02feYjoS8nrgVuDC5WdoBlw0i2NGo
p9nQrL7CHMMGKuF2bNUqxzEh11f3DYcJoKr987DC+mTQmQ00Ul/jwXsVlG2vFI9xU6Qu0CYyseFc
mEAcJ2QO4fYccPMKMJO4h60IdhLGsAagN9JAcvKBzLwMgAedJvln9DNpqJKXJ+WPyv3XTiD6MX8k
TeBk6SaWKNl+lu7RMmpjx5NIUf1XRTMDXlg0NBbv2lxLNNttBTdN4qxyFXr5lPuAs4qCfIR0gnsi
awyzt8UQ6YOqS7HaEMe5+Luw8r1hVu73L8nn9RCY8SU2RtRpPbItwsN86CAci/r4cTU7++6Z/C9n
/9j6nS1Sjx7v59+hJjMq58AFuAL5p9bf1O64v6/l+11oNWElbbRmUT9Juvq726xyZytmxE7XY0Ii
tmnYU6juy7rbcfVKoOV/7xwS/KP6DnrpBNWQFctwE1zXIAARHnsLL9E6DrulMR02TVnPEGsw/Qt6
orGovCMJh/p0qETOADiZ1KhhKE2XRXL006xayL67SuAbnahkLsfs3deOl0aEIf+vHn1gFBiXsa8e
MpZ7HAdzM2eYxIfOm8K7e6LU+la4z/d+lHHrvauah9xVC08ZlzhSJudVTWsjExtVO+9G3hFDKX0t
wwQ2ZnN7j9AQz4pJeW9mIfRWSsU8rfeB228IjmEH5iCOjrJxJdYCeD9JtF6oXFI4O3s5PqwMDKVQ
vffUI4yFlE//xcv4b0rS6R+0oM3MwiU2ryZAmiqd+kw4wjj1dEVQzp5qfLJoS8Dulkafif5Mp4d0
Za15mKnKXVhjNW9AQMeofndPPikAaN2M6ajd+TdKRtvSHwzXg/s9qWirhAV2lhEIGcYPdxlMOFKd
hBYp26mRJtSWPgqe+XG/fuSXolM1whKJFfV+lddGvJfbZCTzOjtfKKrqxPKmClW/PEOcj4ZnnqgV
aMjY1BBRrmopCfjkaNy33cj3p0WGBumVjC0o/Ft0e+l3OZqCC9iSfLBTZnEcPW84Kb/B+jP/Wg9R
6XLjdt0zNeTa2R81Qj2TYO+Pzwd6+z2xofrNFtfF9GmYYlLXg3HSnApDNDHZnOMFp74xZTdj+dzt
/58Pe8GFIXQYXoLblkLYK8EZ0Z7j6u3ZJxFCGoYaXt/zhUn8qzql8F/OGDCXf/pfaD+Z0lrvHuwh
0hZjUjcga/+U6Qsehkrw+olsdCXx35zVYsr/zubPKu6lYCEE3XnRfK8b7/vVCqpbRkVuT/hZWkuU
kLH66Dja5RZtrxCCY5t2DLNPnmVXfNGX7izdBRbO8xuu+srHoSkgVAAi3+JZXVau6bvF3Xvnr+0m
sLUfLs/BwpM6rjliskhaOPjmICXnSi83/kRLrIOnEHwh8z1Y9ZWqs6g/4jGnuIOD/cBheOg+TVqK
0y98XbAKeuRHHBaXDEFy5L6D2RZvmy7GuF7fkSwODabn31nburlWtrRsNG7qi8ADEo1GKNA3HRiQ
wbBPcVH3B05DzLtQnv6ZrAcd69M5wgg8C6cfGu1o1UFCkTq9qdVhSrvDL87ru1RuxFegZnpoT6mF
5p7aZ7B7kBczSfnbXYfflS9UAfcubtd0JXPT6Aa5Pkf8WvJtSI5Qc6Iz7yidFr9BvbXkCWUzKwj9
xZ7DBnJ9+pdi46wXbZayVA/HCRjMN4pkbiyT7BUvQac5oHII5BX+oIOAhkx/bCLELKe77w2+6eRB
Ji4pVzgxTbt5U1CMxV+W2LF60wnvR5CqExTZ2JHd//s+obVOxlBj9a3U7nMahctMD+wZsAo4fR1H
c2d1GLixn4aHCmLJrHFDgvnFVC6fB9MBONCNbp53dbOGLkyXY1SANzDr7Ntc3VPwfQcP3yfwx4+g
zZ7QDCcjKn/zvsJWJCLPsXCSl/BW1JOsPloAsSzTeMwU4vqZy676wWlTw67LPUCcVcPie47A31wy
GXtMuqliLnsKcgjF2Rj0nLU2FI8y0PXf9mKx7GZicK7GgdJ4RFAbJdJ9YY3Oh6C4xU+nHL3Mu7gl
ADgg97ov62DrWiBfnIKIJ5NkWJ2XOU4Ok5VRPqfLUvpMVoqsUS8KkYpnK5MGOwdUa0iaJ4VfVqrl
gWhCYqqCSuZZ/puEllOr244jzxEtRW82Uo7YbYqYnJ2Y61KkUmrq5TcWaFbdtws/G3aeNnWrSlDi
gb5TdJagullb748+SfIJ/8CS0PD5ZIugAiyOUJDCFLtKtUYeuAdmOBZKuffvl/ooC1Wr9kDSasCO
GDRzXDu9Dbkf4WEXgd0WSILyf1uoEQDXUYmy6Xu0I9OYBTsbJL60qWlBzQVTel1B6LuaozyRYKvC
9BtqyHSUhm4nNW36Q4BEvnwXjJpHJMqWAScX93Q4v866kP9wUHtmXC4AsbwtET1w4YGjuhaU0WMX
0Vmy3OBnq91WiQ05//R14B5iyocR+PED6trH/qkG88dn10OaqSzHbrWAQ9/TgBkKGrsoi6fyeOWs
3yrV3m2XLyNal5kvGzr3SMm0wnnmlaXIaoMYcOoqUaLiBqk/UA/JaEO1YhP6N/a3gl+ppbrKPr9+
My2/q9euL4y+i5ByVw6VYVzfPI+hOq8QTZeupNLYRPhK3IqVXiRx1kkFVfxMnEbt6AUAECHjgw5e
b6Ycgsx7dcyvuB9iESd3qOQEdti74ZqsUwPF5QwFnNEmqZmUG61osWN8aDmNLVF+GdxCJh1SLnom
tltTPdzyWh8qQ36Jj7LhC52/4Qh+0ATWKSEo2gbra998Hjwh0ev7ToN45h+opVCyw94vOO2XM5SM
l4M1tnLXj39LGMQq48kFSN53rkk7Xg4ziChZTAxzQsrbtEUih+OxU/pW/05jQcway/5l9aEVFQIk
XE2uhWYREMcMlwsIEzdYh/YcJKeAoX1bhGnENJ9GkgFammU9Ox0tNm4UMC13g2pALGwpdhxhG/FY
o88LnTDWmsHyHySIK7txPkLEB5E9nCXq3MbEucCzP/yyiQg5QZ6u2NGM2vDl7IvWXNKWtghwH5C3
FmA8qe0/2YNKAU5QkufyFtTiixb/N3FBMI2rxqwGwte4DjlBiUC4dCF4AYQKDNJsd7P64gquiIhZ
daUc7sSVkzdPYRrvIqeDwwWQXZSDyns5Ly2YC0Pmn14i3S1VEZyKhPODPO3A6PGh6FtgN19XsnLX
68Fx3V1yPINe9ID8Df9tgMYRGwZkBxkBUtsgATbwCWzqUYea96rdxKToXn+M8KSDoFYRT5Mnha0c
2CgAJmrOg+v6dqaDrSBE64sJFiW1Zs0gakEG78IJEgRCa45u0wf/uAGFbP84x29xCUxiI0U2/hRo
1sGK8HKU9RjV5FTty0PnM9/SLyh14sV4aoIYYLwTixdBZeWzM+9zsXyK8pwtn3qOK2vZBHAxroTS
9kaZPoMF4WGoX6CLzUf469i5o2v0qwnnh5ciJmW/bjGTAxxu6TiAU0mOqQBwGIe05ifpKjewgrMO
r7Gj+foFoR2rWzvZ4ogZ1VT2qq0Ppw8bXHosoGjmS4/c/RTMlWNJ2kUGn0dWTkHMjRGrOEhlT0sF
S2GReMn5bHdbdVRHD+FWd9tCqWiTa4bGntmyMuTAbM4OqPuF8SgWwMgsYkiQp0Zd/k4GbkllDi93
pQfSkPNszY2d1XCsiq2aDN4m9X3of46wxL2NX5P1xQdJkSXOBTvqrRIfebjpvvZLSFV7tcmjkgPr
7suyjTKkwzgnY4jFfwUQ4b190raoVGKrY5qZLgOhNlgfaxJ9GLFLplHvLoFzIqLV38mkNIbQ+M9s
9GTpzZwQ9GMzx+OA+pOpQqIDzQiUw37OMdnzmp63le0cg0Hss1gWZmWr9GUnev2tqjvjW+iKHrB3
QMq+Jt9wtyHQ8QuJJmTea7UDmz+vD1x45B9DkMK9J7mvl1gziBlQ6QpR1stScTfoYlAnhRkB/ORY
Nga+T3+3XPvaVdxzRfpANqe5batLdOEsW7KIg4rqqsEbHof7YXDhnA84h4ieId6t05BoP0Y97T/U
l7+skwoP5BFk4+u25tCld5Zf+YEtiFT+3/ZYpw/3eZIKxAW+NMdZuU6BzsfZ4FAWWtqHr3uMgivE
AbPFMxPp8HPkCwyjK2vVaBAuAaVxy0h/64K9rZnnKrP/9NU196pqh3M/uzUZTUhK96P1qjMwpx+w
rngeFmO+k+LvDrlb8nIGlav63IFdWXF17F04YNiPwilHFCxlHh5p2TixnO9nr6fQSRUGagWyvjH2
SJjgBSu/Z5TMqFVePX6hcmgCcwSKj2kCpBCZXYwrLoyLXaO2R+f+Nnq+MD4oVLrovUuAzOH8WCX1
OLzlTnbadOSiHG2d9490XpYZJ//ZjW7eGhdhDRJ//ufBgrNAf5/jAXoKLd61G5dRl/BPdHwmI8V9
hvCB5DwJsENDIOU6SgXFh08d0/J1MDgTmGiqjiSH4DQuzL7zYgllmlkwWXnkjo3yAJygLUPBEe97
m3SfSsxs/Mj6xdNZXWXDWFfmDjdS/Cxv85tsTCahYs+Dd7utlGyZvuG76JiZGr1SJy8iRqdDraj/
BmQAjor1eo8NioubQvLNyD4ZlJvcLsX4KYT88B2y7dle7kCR3TTm6obxECdWAMhVMnil9FW+gVfa
1+5fgKDWJcHyXibkO05dNaYVUni3V12K3M77rtBU24VLnnWqPYofanQ8w4sgRivZLW1ULBETiSiZ
c/T5ijo4kEOm6Lis1XeHRpV8TJxI9Vd+E8fiWyGfBZF2k4hIA0oU8ftC+jg0fSkGXeGvoUkn7sVc
kPi090vP/WyUbYVB8LsDj7QpyYcSrelZClGITIwpYVwI70hF9a1AxiqxTlvmt8MaKdwYABY5TPFS
JckO4TDaJYCSO78+fFK5PcyD/msjRuTpCFpYEQh190/B5VuzbgEDzr/RWIsumCznHmrG0pV7jg4o
tB8OpIONwCSQYgcDI2uGxtrR18Tsw6v5ThKq/xThAhrblSZ8UBCycNDIa7LkQwVRrHSWSgSwaNZ2
O3D76DsgQl6qzO+lc3rbq8vBdyVx6uALlOdri0r9eTRaJTyozZX6G4sXGlFhJRsKS6ggR3cDnBmz
MtANEiFz2QPjlS3KHJHM2YrI2vMmSMAOWUGhr40dK6KEQhWWAZBq71ahNA8Df7hxtELlcapVUVVZ
vG54qtewXpP9oAabhh5LYOTSlOdk4a4tl9GQfrHEUoTJM8hcVyEWNW0yXF3+9X26k89IFUew0pxq
2gDA/llQOfbqSORo9QZpt1NSXW3R70NVvQcQQpbiDvwkWx3SxgFrQMn/hwFTwykfOdVE/JyjU2+d
byyUfokc3jPh1NWEfIvfnhKhX/+xAB8T8OhT5wCIUz+2dujihmNEiiKdpJDW3sohBS3z9zdIw4Dj
RiKDRSiA7VV7bSmGV3MwVD9Bm5EGzSJQy27vzTD3s41feKtbqq7YyiRfVdObX2Oj8DidABZvYGti
yJ/HBQRjUSmS483Mimy+z0kyxhKiBTZWXn3lRdp0PYPtmcY3wi/gCDnh8LzcD+E1dbzSUY0W5x83
HX54nDjj+LqNrPypLRdEtL6982VQ2d+MPiV7YUI/QkJULo56DY0dOs7koy9SRcBHqlUhG3aOEgVd
fjTf3eKLUkPvNC7cM+dpvb+RJ+vE1ZbTfIlLupWJTTP0CHTGGQibuyNffOIHptmeyLyjUpcDYDjP
rFWKJgAhfvVxz8kMal33rVt9epRzEY2JrPrGmXnL3NnhhiQTMMItJoeu+P5+YGDH2GR33/u6pEmz
iyPpDkNl6Ux67r85cxoNQoilsinPcF+xM2K8IPd3GNGHdUNfKPb1HBozqPpTuLNqkbd7qNIeZF0z
Blk5KrwEfi4MiXd5kOjBIPBXOBOkLPOx/XekyDPW7SmpQoiySE5cTIJEt5GzJ7OPdb6oBb8yfZ17
0dCYN6VkvjJjezmz8NOgmfblRq48FzIGIpisUY2fit6m3cnDz6+RN+gfMxhpJ+iWQgffygq4SIXl
+bNKcocvotR27x2b/zn7o3x0lAvV7fdifMtWz50KLWE21vc0BhXLncKuetpmHNqSXRiOa2/kZKAm
G0XsvaVOZuuf7+pKB8GNWOSZAFtj8NcoMxttgaG7g0Yyinwr/DOD/L2JttO7Kjt6YVi2q2wQJ2k6
4icAOTpGPFKwDqzpCrLh7WoEFsbJlOqRBKHjDdZihu+RGsqyT3HqWo65aDvyIELXwsDdujGRjtzH
IQrIpJCJWh26AaRZdOXihlfGk3Vqhn7dh40cgps4tjFWFCmzT+AeipBWuDl3J/nXmMW/KUTniiW6
yhoys9CtVl7wmRY9wRn0RIIxUACy1d67Jiy/3Bu8lz0lBBJKJeTRQGQpqThMaGOKtXaUs/8uWwaR
tB6aiVUbIGHX7cF78rYTMJxkOmxdp9isMpY0y+V9wSDXDoef2ZfHlBDI+if3IUQ1EQH7t7yQDo2Z
H8w+qJawGDDKE13IPxSQUVKzbAaobzQgAmIbXgqCWAdkqs5oqnWbhB1wmRhXHUFQ78DRDrSizL7s
GD3YupPiqoSbU0vagZmTAhpQwrW74C+esTVf4xo0DWw0ZpXbFMn+gYlLscC7bfhnMo/Dtzp9Ze1i
yGevA8D0jrfYjpMbiCJsJtJqzqoHi4IeKWTnWhSOfrG9Mg9exIaGz7k4rXZcqnULjUh2I28lcmAK
95GumkB+I6O59S1ELOzL4mcSIuYM6ej9akCcxEfSef48RAdY3WmGP3yULTtP3YnY3tqlAnc+R6y/
4R0OhUx0DABNbVu0goW/xMqVf5L4qL9Gl7/AANnzoaUxvroy2wm7pnO9DdoCEF0X27wX14wsu+jM
EpV3BeOZZmuGV0iqGK0ALicFiWUOeiYoo8KOGXvHhV92786hpyOH6z1nwXOMlnebvTZwWJ5bBQap
8J69HgeE5QB2gSApzD/JxnM4R+Iq6KY9MpqNkkPIwSFMqKKjO6N1rSg/w3xyYDouz9O3rg+ssYTw
+R46rMArwj9ikOLmRVOQXzEyWXd6YCgdfIKzI7pn+2TVedUeTRnGrpsn+nvQi3WH47dNihmEdGC3
uOcMdSHwjkiNpYvTjMZqsltiZc7nSveKPbqwjqSPEVVtyzglvSdYdd868aCcTzf/ebUJ/N1/clOe
ePUYlpk6B48jsKiilgdF3D4O0iOG8aPkGoT0ulYEWjUf3Kl6pEMcSeAq7Kr1+Q22EJ/CNbbAjNj9
p/tjBqZlrEv7liGeGoQHq5eeoRX6t1OzYMzl6XMfnWshIU2SxpL+06uG9l5dugohKE0AxNZXRn2R
4nnVEFSvvLHWJ8equhWN2lodw5+xWPqY/QQbqpDusC9K3tx4/ec1JQt36LQBcedwslOoONSp1ImH
F7F4lOV2EPDLROQFrmsG79ESsciMPbxc8veFqwpRtyjymdhcdxf9f8NYJjpEvo5sVjJ70SJck6Nc
Z211R10YdebtMqqHGX1cMKEkzSUEzQsHdiYWpb07idN+APsbaEWq9xU6D9SO5I+ovfd/ynQJXpzB
R1KG9e9CizhhMrANiD2E1mqqVX+H/caJOlS2CJzKhgvF3YMyQdVFrAMR3sdw2mDZVme5BO633htA
2ky0UDhgmibClmO4Sxgn7uxLT0TlQvKY3avJRNXofOV5Gntx4EWSm+Bd/MG29bqwyaz7EN6BV6ZS
ww3M8iE6CurgaTppVs3v7Cj0mFmJEynztQfpJ0v3pZlLUZLeCTOiL1JsduaPPSTh7voGKCQ/QeCV
hSuUTdvbIjEaWzNMGL7tdVKIKFFPTj96p4v49c+HtGckhcASyu20sacISQPEcxxQKWSJLxY9X2Ky
mzS0F9ITDrj08gPFGv8SsIBZyZkGbLYWaW8v34/MaXxF17EqRQiSR8r3W0T0vQMbNa9Nj0RsmW4C
dYcNQrX6Om6KQzfh6uFWdABpF+q3adKt8UtyNKeK2giSPajSaUrWbDj7rl3FgMdJla1kEFjMPS19
Y4ygzMJaE+JNQlp2U6g4yuCfaCgd9Wuh7aoh4GqFkD21q+WYj/iBNk4YwCDnusLLQQmxlmhV2D3P
9NUUURRexEOONx4MXySDJm9SJqBIsCLwyurbpHcx/J+ADVzBrdfVMJmof3vNc/dAHoKWetPpcgZF
m7nhU32tsyC4OLc71tSQc7N/dGjnm0dLUyxoP90oKUcV0RA0eB6ksIFlgu0Bxzt8323YJF1W4Hw9
JDA2YAZhuWxyUF34PHOlA5Ll3YwC9AJG4YtCqa3zARZAuoHXWzOvn7FoMUGu6Gp61VH/WOltJNNH
sTMC0I+ZhNQQ29W5AqoPcGhvSH0q/m9iOCwxhSL8hmz27tmNFgZ7bzVeAdGQ/SPH/r9bJY7QuXWU
3T8FfCn7UZ3JvQ3NNafQcG6SpIqaWUD/+ZdqHgyfmk6vCqLAYVNBc6RMiDpu4llgC1boolY8kSs9
7dXoJDS8KAQ7X7I2SR4pHfoAqaoxJNgsGtPztEAwFPRL+8PAkwTmpEQM4c/UM505c1dCEKKqRHiX
PWyT36Ly/wWlfJfNmC7xF+ze653jhBEpckNxKb11dnmZpkgcTaWT2CmCRjveYVCgQgfxT/hPJz/b
+5Mp+jVMr10c0SvS/poUJayuNZac0fEp5HfsxG6RKY/Uu0aBRwcz1bPw0vKKWBU6gyurW0VQ183b
rLhvoYBwgOmHGpWoMJZDoMCsVv+t9aWvzWQpne/jxjOFq2hOqbHXYUHc3EPd2a9+p7aVIiBwElk0
dzcEDMFUW9Pz9jxO6Ig25jYBPAxpPgcqqbW8bTC8TvZQl3WcN4TrafAMHSbMk28hTDCR2l1vLWbt
whqUtJGi3ynA/98tskGhvCFFB1KuRh9jAICIL0+R/afy32OExdH46B7r98nN/2iJk0DF7M9Rd1v8
4Qj5hirQJNjR4fegPweLX3WEkISSXcRUMVl2yELRjbd6iopTo6+0zAMBBYRZnqAWK5YLXphO2ttA
lVCECM7Z/zhFzfb7rsCGYUNxP/CMWcMQLaABc7Buo4ZCj8EiQkartsIk2UneuOag0OVE91O4rQro
fWD/q5Nq9KPBuLuP/03jZ3FKJuG4rVNQjuILQL4Dx5EtpFC+7EW+kJ1RDqgntxYfC1KhNFF2mkVv
WeE0YbNX4FjbEnWDGzTR5bmll1+iadOQULYX2JCPMqxfjlnjoqhK7BwtaT4wBk+1dxyANbi/bEM2
AMajpInFif9WmCYp0HBTHCAOlalryGTmtt0ZTktXOFSD8NW+HBq9ceTItSM7o8/ESw25XEHYO33v
OcSBKhgplaikrvhlpvdAht1+c55JaXrpzcXg3KnBEEoQsTwFSoKfcmxhId12qcZD3FeaKXJuqncm
iFIVkSYdMzDM4l8Qfypfc8IpdsXDxobL6EZ2DpuPSuPNle1kzmKnlbUWeKWn2AKjbBykNRlD/eLc
jL73PYV5eR6rLBxqurj/wLm9ROvN5um/qrFl4tvQNfpcwPlVRE3oq8oKz7LGfxTC7YRaLM4/RzVe
5Qv1aeSYPqL17j1rWiaOm2LJYjbdeAAsPURclMHlyjSPUi1r582g02TVuXTh3wxgRtyYVOLx6rlW
POrqxLL1s0tQBuQYOt6mDjxqSFeGorXVgqvl08PLXX2kCE1KpLqTjGL4klBu3c9N7djq26TkwJw7
mf6TqHqx2gbsFHBchUv1IYvocpbD4j331bl55ccMZ8ZwLm4Cfo366IDjHLi8TJknJk3T2YEHlJ1A
i0XFRceLlW/KU2H9I/kmTz4QYLeEJU3aguuTDxKI24pevX5dFjbt2EY6+iYZ5Mg4vRcUiDuBERZT
jgom1gIFrXUh8yU9iEQaQrkPYgzQZ427HSsQ67+H+EdpE7LiX3pjh/9JuRqv6FZOFpA8LJJ6Wqmy
H+uIGiMnJl4ixsCw2Y2nZom6QqlvlgHUuqwDfSlB3VoLRpeWhrBaunzwgB+aMbbrdCVYesUL5f12
xMKlEu4vRIipT15toEsnhEE1PhlKhj0DJR0MIR+4cfHrxpav37YzZ22pisfdJIxomqxC8ZaWosBR
5hwG0ausLYXm7GIlAjyxCOEmkPjvncs40T9XUtQuzvXxPLGWR9ickekLELmxSVREMaT7k3gnZM2B
eRPMss0HAq5qKV/Jdx/rMeSk6OTbW7pCMpMJ1WUohOjuYIK4Kq3/f4Zj5IBqmhMzbYdgBdNRUsEP
5Spg9Ok9tI58ti0QvQ/6CxoFcPJ05xIWdGm03rQHB8zAfoysHOWSZdbxgbmRWPBlZuT02uGrn2a4
JNTvg5a8UWgbgyjSZC+9ZrFdJmaQZk+AjxQMVJFdr5VxNgSw2TKCR3gGttIFXiEK+yHouciiFZuv
VS+KPAEd7dWfoRYQTZWkcUHSP+UTDXm4cqV+ssqtHQsay6IYEqh+Z2FV8BUCA75MTPsKoTgmNT8y
NzCwn4UH1t3yyfotcXyxSbJ0EoHqE/MIZ2qnbd9Ybh+7KmvFHqChgg7kYv8Ga+mygi6wAbknerxe
6EL2qUiyR+ylwTiGmVQ8d7J2xCuH8iijPvni6tDAIuA3U8b7ecrjxTvJiI4a9eQ0tQWH+yylHfJD
PdzHycL/0hxMYD0YwM1fEKnOQEc1TbPU/+i3BHXRhgPo3kEQXdNrilzmZqoa9LylYpJnHU4rPZTM
bMsqaczr9eyFpIu9NaJSpcg5gh9QpPAQTT+WjRcX6Lb8EAskTCXrlZ69K6S1nneQRVw2Rg/eVghk
N1w8iNeS5grLsT/RRdTwVZGp2KLGSZI7GCE6sNBHo2W8j2tS6kKA+y6r3jKFEwJ8jhhsDvtjBf0e
SIZGDBO1FTDNqkjKPlc5nB3GoN5VUangM59afpHSMm9/xOurmmliSGDW1Xj/UPHJ00xDtO33ZhZo
23MqScQh87TUS75xIhR/Z6gyBlfXubm2PcQAWpzOdgkRwUBpBxNgWkkWl+vFGovdjoOxllLkQJUy
3bY4UjDXSwIzG54u8Jp7MswJ5hfwKby0hYDameKi6kzHE/6ikp+CB4u9QXGeAhrbzr4o+RIgT0My
HbVjcsJXhTHcg7yvPbzMhOO/a50Abu9LVqZM82tM3b2PMFSjEzekxTPPovDOHn7yzv9dZEloOesB
+mJ2TcVfZebJdvWOV0RHj4mYiaXVAgq7zrqgndiCjbh4SPID2IwYpRSDz44lkIzZ0i/H3T1pKaSh
GUw+Md/vC3mHrJoDwc+v2GS5E/A0J2kQNm/ZdiHKuyaaCIw6N4BNrHLwGTue5NXxA5suIRUq4aPe
6UNl6jM9cipwHwkBy+TeQGXNiXCXsE+g8iUudHDfVTrrWHRZL0Aqk0r8AQD53bgm9o97AoiiblEk
dOPcQBhMCl9WFkSCkcHSZBcmZDBvwJDND3WhDrN0Zj2JVuKmmgZdkRFPnifREORmUonExcGkz+bH
0kbyKVqncszK+3WO+qXPZLFDvJIvhWVrkPC/12WCLa0D8AXBbQ+gRMSr7bxmex7B2UW2YyXU0YTs
b3BZch8W8GHAEF8OwpxLdavH1RGQG6WNFWNa8nTm1mlOCIxy06Mne7KPHeVLl90YKAwc5UXiIYpb
v+Dduo2ezkIVW2o0EuUes7ka6SrCTxkAhbZPv9KgHAR7+g+vX32MRDuYaBwVxeg4fIrE+PGsp0Eu
Usv0rJ5+M/yuTV69PY2c2R12EFCyzpwTHvQmEQxiQ3J1OJ6IeQpwdGXP6qayR8ckmholoG8SVajC
se0Mb6XfJ3CTJOoWCoZQOTeiJxinF+740SYvOiZzOjEx2kPt6AK87u84eGkeeOkF/AiHUM/8zSL6
6DMQ1fBIFkGoKDUJYMJXN/iADqL7bfabXqhWlSmlbM7HuSJThtxh3+9XMgqRb2tSzXct+VtxvMcV
ZRsuKpmfZiuDe/ZagLZISn7AvOHlLgm1BnsIbWUBTIDGzsCs1admeqMEN5d0J5QXg5sk7Xk0wPDz
c9IQCCPQrxanNHZYjhL8VrsTGoGIF7cwRvsP3N0VXg02kb7PpgJB3Q4yiOy8qXTU+B1Kt5AK6TI6
nKaR+0P86SRuTAjWbQf/3sKZ/DalDtqfEGI4Ag96oJ60l22Qv5DeuC1C6wx6IgMtiR2eP2xoEWBs
N1nL0wVFhTZfctSZmEhk7GG0XW8aoHEifafIQNm89LycMTKaVExdDCZVsI6ojKj/dYKydl7ppgJK
mqItxSFwn64K6T0UC2WUMt/qYlXpzg4cQGhtGJA7eA0to+sG/Ww30CPsyz1iCV4/1EC5InEGJcDy
nMyL45+AXf6n5mC556kuTUABUkBevMDjMycVs6Nyko371XSsP6rdtLKsycFPRBe8ghVsP4av+Ulv
GSqZABSeUGjdYLfWu6baLkTtz8/lGUzm6LwrfjyAc5/3ABBmx2bdN2R9y5BOXmtnATBpDwlVwkqG
VmW0VAmloNTWZdRgHCBVvbfSM/fysKg3cus+PMJfWN142pe1PcPnkLN8KS+m3v0eEpvMrh/p/9XN
4gfwZVQ+DD0+GRrQ08kd0vOP1ecXvtJ1lq2qM8tjMHDyd++Jbrk5KcanWQvghp2fbCDbejlyDd0N
ixQiL+40F3+BSqgf2FzA/mq8aNX4Kqui9j9WVP7s+TYZVnWFDEGlBCjCijagd+zv9GGysWpAor3H
umNJm0obo+vT/ad362/HBXZXWCyaFiyXfjleygtLxC34bkHQkBBuFcLy9Q7PU2GNagdmwM0inloa
aQRTdHCwgYfg5tvpCAdD18NTpVq5ydcV01wqcItx3XqKZ4/lN9pw2wMjd4FQGZ916ElG9qOnQjD6
wlKRmxVuPos1UwCEcYZV4q14mlXvZZrOEiksxOJsO3MXxAnPfgKyPacAGMPMEvg/nPmXD6eb92Zj
PrWUjTVz0vvD4MibqYxfuxMvt2tDpVaC5tLoK+8XTKbrozonT46+GZXeahceHxQEDU+QuGMxVPFp
wcXf1cmuw2laWFVbd2YsMHJe04/aLr1oHwOYPZZCWJVUpkt6vrVzcUfHwgQuZTZOpgWwNt2YXlxG
xXniXhkORSU1BB6zTImXxeNrLBkC8KAjod7XjOpT/bF943Z5g4y3qQrmMCltGc/4l1ZnB51naHpA
gUBFNFTLH4UUHbzDC9xZbhAjwT1lqQ3cRwjOHsqdPBpDHZ78BDndkcO2wQP5EPecNiAW5U/ni5Oc
KbQd7rdCOQ8ywDQdy1s2pB14lhGNkL84U4JCAigCGekegKDfT72GI2V5XJWrb7BNICET/opPm3UI
li6Bt8tvAzr1r+H0/uUlC3x2yB6jgDbxLZdnaYY0bQwfGe/oQdMYgSuTxFJNAeAPik3mqebvDPw/
44m32aaNhJplHtgJhbIsoCYZV5MOlz76E5cfamT1fj+ygi0eqE44pN4Fsqr/aLAMoaFrPXAZXW0/
SmAZ0nFTceLGqe1GZqDIPjPi4c4iP1dWf2sxuA9PRvsIxOAmWGsEg3qEfzlaHzRHXebuJ+q6882Z
P0VeaexP40WFs9PgDZTnt9knzAbW86GMs6vY4GeibHfqezpyotTOGieppl6f2OXFb7npW3p4cSIN
jglm0kbGrDgqwAQo65hH8MN/b1FNqdpxBLKCw3JsplVN6JcfLppfPYmUZVwyM9J3v0IwHNoFlgCL
TE+OZIGVdmvPljqR4I/H8lAq/8hsMmMJcSeW1eqktsUOGLvAbM2zwZgPcgbLFiPCBOFzcWSgoZ46
CA9VYuHMtR6c1UNIcUpBokkKhjCB89HAPifoN+Avu5jWhY8O8Hot8E6mHtf8IvrbC7uk/qo7ptrS
+CKS4buiR06JF2L4De4mf4qTgS37Ai/NXA55d7+yaRQpRbqxeDB3wiV6DS5csDvL8jbtIJLgL2r4
fAgwbSYBOZjXgrh+GWEWpiDtK/ieqYdNHm+c/CbA1FPgzVztDe7f6lFd/fqb4SFVxGEFRAHMwezy
lpy6BDXlTO1B6+jdr5rzYSNyXKrQF1Z6SQngyn67pcH4ccFir4LAEeh2EcO2Up41Qsc8h0QMrQco
dbuZy5n98L80k36avQbXx5BPdN7gicGdkykPlU95vyPRxT4VxvSfI1exHGXlN0/WdAiIuZhTVwd+
iipZW3OuElZU8y30DZXzs56BpHAyuaw3b8llvJP0SUR9c7RvyMDEn8sErds4NVRbkVrSHbUZTgHd
VeLuHSrvziNcfdEtD5L5F/h8iJrtrkXj9N+R2aFg10+otXw+ZXUIlS0F1tbzut4dH9jXnMv+UdOF
h57y/ZHJWyPUnH8a1mmG9o7bGdrlFmsbUd6U2y0b2FiAxsJimiDeGfExgEaKv8Rp9cOtDFM5YRaE
Ezi53ovWejrOufevB1i/LG/cj7uX+SaaIJdcaoCO+7gEJP11vdLhxzkZ/Wv5KnkNIgk2ShSMgVeX
y9NrIW/QPOur5o6SLH4bjuTiIPWPNxoI/WNMiI0JOXQpKITsjXJG/5d2A1yYp/1xipIrTBbM2i4z
QgWjxoUSJFfzvOb4ShL8asZBsSvXrTyP8oLOdmuhIultrFAVoTc4g9wGm6tNRr3WJeaHqB2tndWZ
kOnHUgCG0U0CwyUcVwy8ds03lvNhGBss9PasY24gsFbTkzWocXpsQ8E/zRxL+MspxO4CzLqsn6Iw
y/+DahLWmU1FVraNlvjTRO1X89cvqid74zY2EAoelWEQ/64GVar5lm6ubU0yJuAv+muo9lBqO2nk
C9waso3ZzVJFe/S+wOixrbdZl4N5jvDjks7Nja7NfetLrdPC7AnhtgI7acOJYMqrsreZNy+AyYb9
CTK2f4tLtHxBtWas6hoFBhzVD35VVlrLg0XQE/ZwwIG1cJ+9J4SpYKZJ6+juglZ8sBclcqa3sxXE
au0HPFYQL/xkGh07w5HkofZtIpklRqK1wq/EP+v1B54z2/atBH3r4hw5roMnUfOMmo2JWontrGZf
UyEC3/6t++2HvJ51PqWoVRBx0RRbpq+OEEs9WjxTDxQrhEWMtegOdSX4Y3IpHdZ424SZhTCGsplK
PIBagIbl08WSW+qxuEMcblLAu+jIA/R1vHbwbWtGADkFqjKwWsI/z3FjQ9DOOqy8hQzz7ZkVbGbg
JjOdKB2us2WEM9zCuiGH0+zeCLM2GSWruuzsRIF0o3sEVwlFX+df2gxIpe+ZeGvXUbKKgafaPS6y
KonhnmGGWCED9Tnyv6cFn8DMDCDBUtcu4dzb8E7Am08kK+etH43+TVFf8GooXQdrT8vDMPY+W6jd
YB9Njb6EdR5rMfTH0PflZkkSlpLLng/ZPJzzpKatuWBlKJ8qotIcndJs26QNKlBck75H5vf8yGyy
IQv02eEcPO4Enh4ZLQxHDer0NkQEj9C5CECAP+/gd0YT8UmJX8m0zbmKRNpSaMU8uNk1jTqa6GHK
qPJTNSpHqZdOQ7ka7TsLfbr9OGCrmhblutlBN5qyy6CATTUD17HZ7QIs0bNv77kbyVfrnulTdOFg
UwL6GdAOcA1OrghVgBY8S7EO3sGqpvBXWPwWrDcxe5arFcHDif2OFE/gZ9LHIEGpyd5sN8/1uzNq
LvXF9c1i0n8UmY3zw8c90/0dHPbNPyNT68m0e3DpOvZRQcZsih6Z89R/a717611/uk1DN0unBXz/
5eJR1bpZZizfMKjNH0A1nngwgalY5jwXnQot1QcbXR5/svHnayjN4XRMmCeq7dBVmisjwHP5RznT
O0ojRy5U5iMIKdbiNI9y2+YtHxNuimmSZzSYYALSCTncMvVggcrWX6u8w+yHM4yMpo8rtpVPI0HM
uo7aph6QTnFxIxDj9bZjlOWg2Ze5KTBhO/vo+CSvw41LMpIRSfKUDaYkKRvZ5kTQERuLBKkVjB9Z
2AeGVczde5jUvMZ58DgNfpb3BpsHxPuUMMcxXxDcLBA6IvL+JFsykIKUYciprAW4CAiPPc6DMa0m
5NfD67s4rf2oBNy4snk1s1jntBEx3+0delRynRS0Vfl21lvrFMGimIsl2PM17hXXAr7NQGEeEz94
8/dmtw7Q/gciQwbIKbhb4S/17RTSzv8dBdTXOI9YL74Sy1X4Oj7tqc+qgZk/eBS1UfXh+8Eu2wsE
hz8hqcfWazpmQTG1VQQ5z8F5Wo0GWrcqtsUSV7hRBmoIBic7U+DCoMGBxIm/fVkOtHi8nsnBqjHK
MTLaUjBqX+IeOASkfBAfgo1qFwbczcC9PzWNeQNvvOKoSj3lVxTat+nWD3GeQvuVNpEupztF4iIZ
z5sDZZd8oZY9r78RNRdX6bPY0kg/wsX4mkSk9BZR9Lc/H9yjCwrIie+tFBg1ihCK8KlGXkROumiD
vzQ0l03WZ7V6bF1Hr0sTDJF4vJFFRk6n3QHBXBvdlENaCSjlX6eBLJycQrp+wNwINtldWIdMJzW+
rHxl2K0V9hsWdD5yCC7kvjDofX6FdcNxuAqGn/RmEgPpMGvq4+OD0DlR6U9F3fHtDasKSMpBdTfm
xSBBosUANfSRVdGiNCirKBX2ElzCwVii0UbuZaLYWGdvygC2t/Y7mY45cgv+HLXHKWuVSA3Ys+4o
v7783bZaLOTQNgvSMubgVSHjD50RjskYCx6lIKMdWQD6B1DyvW8YCUEOKuQxCqTaF5hl3Fv7qhTL
O/UqwSxn1rfVAI1TzHJ8Y/AaTuDOqmPdPI2x8DIXtAImJfIN59L8CFXGB93KU/Fjs0VkwomhMcSF
Q/KBpiSvkXAb5S/9ZAs2Nqne+PZymj8M/sW0DBXyIjU0JcRJIDdK7JJrSKSqvNzlCY3lcgxRNebf
wHuhoK1ZFb6W+0qoz/78iDTyeT/UX2GNBP7UFXv1WuLSJp9uRANaxdLpsMIpuiAPJ4ecImIJ4aZl
8WlyYqYB0ZSE2lrZUWRpbGZWZ0n/IYjeJo31TqP2kii3Ox7pwAU163B/rrWGfK4rbOXEC2myqv3Z
Llf8/D0kW54TJuAsZoJY6uDhhmyB1SYevCkcGWiiXacDKqSjrX95/L9blAv6SP/BGT4pW6W/caiz
we3VwKA6hSwLd4MId8nzJuYfwQmU7DwLchCE2WfdyTekWzTdEK0tZdBTRVlry5LQ6CM0SafJcmzi
5k8xpcJVEWpyYtxhnpO5z7ke8kk/5zNg/cnxr2XfPZ9xRIyht8MmzYWqE4RGTLTYNd24epYeBEUO
mDgdz/KA/EgPaqAKwif+HH/tFjhcto1skyfwPdYsvhjWOc1B0IJDY/XarOY5cYUM4R42WmxL/2Jz
7CzjkF+WVEh0Ntp2vOdBohB61+G0x5ibiAePL06JiBklIIjxdI3UR3gmvFosXml5P1rTv2OMySWA
i9r3ajMD1jIP+WTIJPkp60DnRTXcK6Qmsy3tWe2/Kfmb6uBzAS7uEgvn79CUjLn7x+1L1IYCJN43
APFUpJuMRA0SBg1U7G6xd7eZkRp2CFsGeUZpcaajO2VRuw/f6w1wmAT4r3bdfZ5bcHNiuLpmwVD/
TH/7gBNxWjLkfwZA6ua2Cr9E0RkYcOiMQmUkx4bQekqyJJjwSmYDe1UX+QsDrYOOOsl7TGnPYbrn
+rnO5umQ6MyJOLOSwrrR5fTPkWDK0ygVek/OA0/sJbNUUHa0Ax27QGPP/ny4BC2tMBSfH5BSMWMv
efpR4nr26nMRw89ZeGt6AdEFVTMP2TzyRRwZSHjmeFjbk9wgRIh932AzFBX5qOA/U5ahWKxbckre
zEjXqgp7gEE6jKSiB8md9fmGY+wVaNUTYqDRn0sahwPVD7qXHqAHETsdaHoj9RK/gkc8uFkw+oJg
4SJkzGjg1SSpgC6zHXabahux3KTorcyeUtRaGRgpxPlp7IxXIwYbr9R/sViIs8MLLLSHUakwTe0u
eHJpnG1EaWzqbPvCg7JHq1a8B7fci5G18wq7lDpJrk0znbis2M3EfLGMO51e5WBzi+XCvsOLLGx4
ePAH6baHFn03oitHsjAesyb3XOIwslqV7t8OsifPOH7MzE1gloD6YhI2/wZcG7xtbXc1UaZWA99P
N1eLQ81xgAYbxm866Yf+k/FRUj+xh5bGp9OcFUwvVxmp6Fp8FCx+YyzIovj2YLUL+Nmdk3e2Y5oQ
sew3aCsO3wJCGaSNq2mfLMiRX6U92CFGzADZEzl5/sC6LasVK+ljz3ujCBb4aDM7skYxnTTuwbgs
2RfocmQTngjJHyaDbwcNCmHprJCM1Us980iy1vV1KneRlJe877EPMB3Gdt8nDZDLY17lXLGER+lx
sVFUWGTCG1CR5V9CMAhV4oZ6xHnoP6tjfLeHA/JJAuql2ZHJSu99N4sdBZaew0s1Ai3mPvNMGteP
R3JC87T6Ah1BuDRB7G4f3y6P7MIll2rN3CiSJduD5SNrLBxuHjrKytE3acv5JL5jcs+o0yCQczRK
EtxzC5I2YmwGmtPu1+o444cjDjLJdZEPsGjXpLttEghT6blzgQ5Y5NSbgTF2qvDwFWTUDtHkuZm0
7HHWpqKV3baQSxgy4oBXR6Wa6fJyC2juzCMdnlpzja12iGqgfjPCTuGfNBNS4GAV6bfnl1pV3B9a
RxcJr//Kjh1W+MhWEiean+g9JZis6/zWG7TWf6+cvcbQSjq6qkbDPjij6QXgC5WvTSAg9q5goZf7
nTGc5dpX40rYzwfB3MkZ16+lZs8iy1KOCsUETpiQbYQCcu9qJOcSDGc6XhWiQIXkOm/j6v3nX7SH
JSGu/5C8kbo9sM7xpcfVp4qCUSoxhhrbwpdxFXC8v4biHbFcA9J9Gpmxbez/QBXeokebVpMXqT6+
C4oOur/l20fmdzWkEKPWcoGBVDWo1b8cKhJYTsRSi+WXi8JFOv2D17nVTFydMOE1anSq5jYbyyAv
0voJQ1yJwgN4mRf7mKA7Y6Op0ybeEkdlN0MCzFMxPFx+FoNIpp/8WRAM2zpdzKv3ZTKB+M7WwqwG
fI2x2D5YTYGc8h5pNM/t9UUGWsqaBwepr869AZYkUq6J3ic1lw8LLdC7VkZID50OA3fvPJbv27cM
2oHjj3OiP0BsL8l/3Q6rrByZ7SWgVkfI4L4YjX4QmDKjhN/dWjX9F/eOjUTctn2DdvASmI4PZ5H/
9JxdnNV+9njQmI2igB6OLZwc2lZelIP4C1YhZYOyhvj2bPFq/4YTmDL2+pzbr0AZj7AJ+FwHcrLo
IYtc2/tVJ+zfJx7fzeI2Eh8To27qhpQC93sNR/0UG0SuEc/VZRqnmDNIKhbIsLSoiwGiN+775ooD
MWjtXJDGwYHKoUmzUlnqifbtgP9Y/Mt+6+FLv7DO060Go7Mm/IJJ59N2oPDGnJKnp0hCXTySbT/o
1gQCakt/4iv3Y45dI9SZzB2MAjLawTL4cxxVOm917uOs2yg+aIewFWTV0P6fuE+26UYob0e0Qr4M
SEeJKx1iqH69di/aOujwnmJv9bQ6QhR3dQ0Y3CcmnSAHnmgMTHPZMYubH6oaP9GFIokAMoLNuuJy
+HYHt/RZOUD09L98nqPzhonwmmuhIMzQBXogKnACFc2egio+HR9Sx9eHs9J3TFH2LOjiBL+sdcOf
ldk8j7avjmwTCAqL+r9/BXunDaiKOLeWhww9gqxHLCaeLCfQK3CIqZHOm9ArA36P8l/rKWX8wROR
YPO5s5IunQgYOauBO2YUrAc44soPl1oXrSTte5KEEG0K8B341RF89ffCXVK2K4eEM4sHFTg4JpF/
0tduUWhSOoTP6HOldmiSQ59XVQFFhdE5BA3CSgxUmjqgOwQ4M2Kx87Krl+q3TEOnsyVS912LTabi
DOmMVY0qVY3Oo9vHoeI6U7mU1IaphBrITyLfN4a6MPpn+HTSwpGLPuCdHFQJzIIfnws6ZGqAeCvX
/jHSTZby9YMjLVV4rG+oQyifG44lLXiWImBrQQpEb14ZSspgKfTM7D93x7dHNcUHBFw7DuMSgOHQ
2wgsg1o0teW6GRn5ZQD8a/XJqAog7i2GiB7FiBX0DaBO1+DH4S3/2Rs0IdSr+83t5P9RXR3YNKeA
/5cZye29KDN1UQdwIelgu1RPQdRIwP3prfh4yfZLfBMfxg64fCzZ5QIpVacDmJ/7SQnbdoIrRZzK
QaF74BwwzflLROJJYTqvTyR4mq4SRsDJxgXOcqEGvRWANR/C9uCF/d7cCuAAXlm4al4lod/UKSvI
b01LcQvdI7W2AecgnPfuMqpLhNQ4MpV0qoPEKRDG0JffFIXAqj4CjC/0HAsGmSyvzMtnY6Ak+8Qn
Rz/69f4iBFzirmGTmgCEABvg7WhjNVtptxCJP2RrpuUe+tCLRgjge2He159oCqa6Kf6ymbWfJOF/
RCdQ7K0ij+9yAQ/lI+OVCaUN2LgpmHZH9RGv+o7fGCKML5zkYiGp1ALEHj0HCqRlzyr/Dq7K/+2a
nivZsf1hMXa5yZuZAsBYLFAkWPFmVis1bGVeTM8J9MWg21XitAyRw1CcHDza/N27xPtIB3ymMFlH
aTqV8VDFpBzaW99dJ/+ZKi1N8wThpA5W8j29S3EpINsb4Gi6Kcbc+fJRPrHTrTMg2BWGr2XX0LVK
QL8sH2gjOR2lcSMJTUSCUGMSVMFXudqiuVOWq7wE360+CwSuwR0+i0bUoSP1bvZM8tDcXyGJ7JHr
peNQda0wr4W8wEUS5VhqCNx12b3mB1lECQOqFYDGyJNlDMml9Gm8+4+jT8UvqyhaPVRSMOs4iBGL
yEKAJhpuTvOP6Wi2+mJ2USqTr0KUaissP87MqmKVZyILtS6UEKU1ca3ccINcaBc3nyZ2qXCV7Bbh
zAJ0TKVnaJT3fmkTPEVrY9ouVRFeT6LCW2Fls7cbruB2IV3azblzov5K1IDhvS1B9bADTVhdF2qL
vdVkRhWzC2jRXOn0ywXoUu0iHhJ5rQwrSj6EYDFzelSniWM2T/9TtH3sAGkMknYQwMDhyHUHv9NO
AO2Tg+HLlsOHPWs7XuRAygvTOGYC+mqSWocFzN8DJaklBJHfc1U9MC0YpW/fdXvcddrfzm4qV3x5
EVz9XRH8A0TgCaUDuDUx2vdXH/1/oTze1x6kU9eo8q7GvG5GHz29d/UlCaGHuxSmZMGX+YaB+YA+
3jLNa1f/u7fplexQgls2cwCGEqTLvN+RBheo5In2NlRVfKuPFXrLLc9GGeFPJtHVe9fi6ExpYj46
3xbZshf5JpgbrsagETAfOK6y1qqW86Eax2rGJDRxaGcd4HIY87O/EbYBEPhxU1bnbNh6bnKzBLfE
C4zIt6IdbzsmGqv4yb5As3PYrkhQ17kFERVoUwzQkQpnEVtjXe2h07WJFigRESRnik9edQPaCuSI
q0c44L3A9OcEtsieJlAwcOSgfEPrFsdEOw8Yq8OXyZzHPYL3pGf/PeJRlnLCY+1wphEEPDGRRe0D
ayp9fQjX78Bh11FX/DLSBvVZkN9ULdn+I6UHhtSprjbaAe13+x9yAw7L3nUU8BNeCAWUwA3eHMfS
SmdH+kmemLc+wNuduIe0ijkVSIPJFjk4ZXmIUMLConL0YqrsBSL7rZ6hgc01MnQBM/ofNMAzKQsK
W0NaxlCsHD6fvq9dbWP+ozCAuHVNDfVUi3r6ONISRM8Zk+gA2iEGI3uGGg13HMKoYKDG2b2EGm7J
CWkzuHXL1+li9jRGzWetAF+Xpc8tb+Dk37/IELLZ0of7pXxdZKDgSYKJnsW4sl7S25MUaEaOSFIz
L5a7I/RepUO5m29GrqYEVG3L/zYn+XdNBuj1Q7rKZCrNd3vW0KMMBoLiuRnbOCn5nzUC51fImt3j
L3VKVD/shsUaYuTSMRX9kP/jBDsPAcNyDtMcMjlxenoSJJktSpzsHdm5fpj/Dc9tJBHGpglathse
qW4ErgOnwp578SEDm6FR6YnOFos1weyZEBAr4qQceOe5oYqIf2Daz6la1v0qjziPtb26qnw3mhuF
omLBa7UYTMRuwq7N3xdg7oqiMDTRrknviE3FmDo/XBSwzNxbCng550vPPCjj0/AfLukASwCskJlG
OJayM//qHD8mkHs8OGhUo9UvK1/bcV3qIrADmWJm0BiGRwci3b21nNnY6M9u5/11Xz/KaQoAu5ec
yX5zzknCMRgIhftntPy59rxeISPotqacm/EzDhhleXk3TNfAmMNjswxZwMddgGRpToMaVJLv7+5B
umG3DWIb2qMjzjxipeUoUB1kcawvx9ZG5DgL/nu6BGDS4YqjS/tCJ7ITEqKQBaRE6N/EJHGgCajW
Asu+q11N5fo5Zg39HMaO0mIEM2eDPD2lZBIqRdjkGO6lWB9AlboQrSqtG9grL9sBT2iOzWd2BGbz
AG1vlQI9r7omLgJkMzwCFoWzjKZZaesLLuSYqQGJSfJ9OScFGE4Q1GJeX+KtggPHRZPHdcEYLqQ3
a1fOpREaG1xBk05gfGMyMuqwXlFT0IKPPWqW9OsxRqfTOCo/oXRBtAUZ7OU1LbXsRZTUFXYs0zWs
+7poUrZizHVw1uHTF8RwAYBM3qZI2l+JkBjLKRn7BZNWoaKuC+QQzt032bSw03CFMSDe8BUPpc/I
odKWNnPejZc5sm3H70B+e4TxCZJG0Y9duW+ujK9WULhBAzwgtPZ3CKjt2W/DDWMJuOj2IxPXuxU6
eT2H5+SMsEH+sKwu10Vl0TJb2lJvrX7ReK1G8HJ5J4pfCYGrqRJx2M87vg7KfRwANelth+71VrNU
sxWD8rYgwwvyswBu6g0GtCB0/MeVvps84KNvotSES3cDQfxbj2I0P3DUWxkp49WhrNTHVfKYBpk6
o8HgjmFTfxNr849nkqsBeFeKEFqR1Z79RyJ/WeUq0n8EyQr9c4ioUlOu9zuKdTSQsmkUJ/n0p/uI
F9T14qSVp/Y4S90TMZolN8pmwSPQnHQYZ6vDn3ge4XKmaAC5EE0dubl+zTXRwDAHNCwUxTeWW1Iz
kbuSO8B0Hfeh1t2iN1iGcqhe5nFKzb8BYot2Em9ybAHeNlWkbLejRlIds0Ek8deshYp4THo8aAet
ZEbujFJKP8PbDfKWcovngjP52tiFYCqhykQvWjKUiJ/kgK5dyp/PPw31I2HuZRRFdb7fenWgXS9Y
U+NS9SqIGJ0MmymbVsBHcEuyhbHoWKx5WgsuRRuqwUEPfvjYPLdSTQ7susXSbSpHvMa1IpPsVWRQ
JlLZADkeIFR+4lKwpfG72q2w9OF5SmFy7GtUUFh9UHPPge3KUMddG1NoYE7sxscbMaWp7f6nUohM
jJfl8bZy3kMyFXf3k09OCZt88Nbd/U+G8NfJX5Lvyc0ARHNwcSFweZelI3Glt4EPTPiSN5KBMFzV
210tEW6nxz4+CJjlL4mM5vfLKMqmWyEEHZZy1M+pTfxuxu+jcHvsVPg4YiBoToXD82qjXZ8volp8
ybcHgQgJExFZCf56u57yFjJZjLaNmkHZqzmvpoP/atUf9YdLSbPr9qDflVzj9PwS1ihUqvZidwCM
nsdf/joKb17aNCuX7Ys+Mx0Cf2agEzkDcc1iVCy7KaAzdehcC4qVbX7bBnQyQING40EMf55Bntu3
EZOvi2LyJG9jqXEPs69U7XsC3fXJS8D/hAz7Ow2U8f0NZxCzr+D37XVAU87oo9RzJazSyHQbBPYE
S947/Z25HIVGYAoQWjFzdy/ifUl1MV7b6gb+zhebq1HEek8JyoAU4rCGUVKtri5+5WBZDKJwmvPx
ZOZe8uYUIDm3JoQZmTb9M8uRL/PTh+Cpy893Ugrrn+Oq1lVx7of27Md4PWWZG3bde8uQxyirzUKm
+1SpsM2S8NQEnas0WSb6qyTqtHqDRtfqumJqoFQTSL09yLAeAvDCID7YR+OIIRLfdfzR7G0BA6hd
R3pAqa5vgHjL5mDPhAE/DR6VECDY0UAnmlJa7rGWH2sHJp9EgpaZJ1QyK0z3Rg2l2s7mLVs+yUjh
s+tQOLBJc/zkpT0vk7b6qN5Eee4ERkJVb8RQZhuSbHzapqetGowuRavm4lFuo6Zy+8N0hB9gmTRW
6OXj3AAzk/PhdBxRGdJGLUD/jLsW1Due8pR1KZlBDutmo9uG3/l4MZbTSF95ZDlEAqQJFx+qfYbE
F9OcdFVo+Q1BHu+8ILb83ZgiFCufabYWQw1Kj9QHhXaLtdz4Fv+FIaWTwMXwvDOLx9ZVbfZzomhE
vhPSryYCj+gvJ5wnpcGbKyIUaneSTWdy31oH6E2pH6obMsmmFEweFPyB5aBFdaB7ZgyJR0y/LRme
fDRHkElt85kYHvtg++MnOyi3+9xNJl4urpuRaPfd0hs/Z8kTuhde0tzs6TFd+cShEEE1GOKdxKOL
CDC2Gzal+TyVTAWq/LLRn9NXCwyKgnPYqqLu5U0+RNDblU28MK1DMhp64BNoc8pOXS0M9XQ4CpKF
6jtmspIzm+lAcHruquq01HXenV0hTyJkln32akMH3qJyKd3OUgcjaEedZolnYq8htqOTfu28c8s3
x6Olm1OTzd5SZN4oEDSBRGcw/smnkh0UHTuc0cSlgZtAi2OA16u/OaAGaz6u48PtHQaQvqWyCAFU
hma+Q3n/RAX5vkl9Folb7wy/D8UelOPY1H9HdRNDW9+H2ccofaM9q0FC0rKvltOAYH95G+cpyfHq
JK4RL7HfUG3TwXyGP2X/sAAU6zFIMkGWE4KKFzZoW87yQW+rNOPW4uof7W2IGx/UD1Xsx1Yv99g/
QIxHNIjYUaBEhxwztLJdo7KVzljMfBmBuoSncEPqZmVyYEiM6dK+GK1FCrWVRYKvk0aqfLD/ggcS
8bbopXSsc9Ds1KgJfGiqtJEFFM1wq8AGOgbFsZwOK8lXFDwV1CS5AGRrJ/gwUVa6hgsZJw9mO9U+
sQ6ILAtTymLHjhBvp7gExQBct4TsCQupsNb19GGGYP13ECwReJcpuqr6qsa1LKOBHACwDcCzIDO9
iNV7Klopun2NoVBs0ZoeMAPvlLSkC4cG4B5gIIlC9ZhAh9+MQpqEgHgfRrE/8JmpPPgss72Xxja7
f+J22gsVzw1ei+yQs+iB4Z0Dxg5FBtE+uTpyI42ZR7Ul27xpXaQx6KHgCFv7FPb3iMuAVoGLjfwu
0Z/nrjov+8NAr2+qJw+8+krFWIAdWEPsw6TNwHoltOG7B7w2hZygs3bJiM1UiIYbfWMqkqk0CJUb
naM4EaRUE4WZOgoYPZQtHlEgzIZzs8Q/1xeArMVya+daNojotiDhhB3FIJhJppBM7z1gXcrhKdqv
8y4D1nhp5p6BmVlqkhnvLa0CweO7esu/OvD7L7II6APGileN01ATM/m0e3EWguoUSaLZXwB8DBRh
YdWwS1C0FmXrYNf5+Tw4+/Xnv9L22HvnZekRGzamillDkJYY5ApiI23zHuISj1cbzr7EgSKwH0yS
haA2JHAghl4jyfx9FMbW9Tw+dNJrxmuyc3b0nFTsTi+f3Po/3hp4Ws1QyoLePupBWKPzriEAKTFb
4mpq3QExXBbQC4UiXed3UWSwt0tA8xfiXlD8qojRPCO2aWEpt3jbFdIAMV1ahjMWPfeIkec/rKxr
jbW7GA2eBhnMm8soc0OCAvVi+Z1NbGlNlKPurO0rpFsR5b7sgiJnQTIEMIJUgj1LryKtqWoNb1oa
BdASwQS9o+VtvEr58NvGHQivVASR2h0R4+TlKiV90LOoXtYRu88qrifNhgKyvNQpJfssJvGJ+fYO
1YlohYofkwE7rDLqqm6RSkWyMy34f1CriZh+wxJB4RKgFLyuBNTFOWq/F+d1xp7vAtm+fmTg/6+2
Y/a4lUXjmifPSOQn5UriGtlyG8djtmNgCU+8+Q/QVcAzf1PSOidP9sVS8FXt+yPlT3kXBYJQMW3f
EgNp44KZwCjF2KC/xf1TcQKJZGmdVrmbvAJerB/4zWt02c8gnwFPLXylTMhnD7+/V3rKw/d6Hwf0
ALDjoPhnW4wDxX8ow+lMy1VrXhCNGcbPA4mCfva9I+Ruy8NRiQdG9C6KpCLS0q6UuI6ph8wifhRf
IrHXg2zDUo8Fi6rDA18IhAQtLkRAGKkWzjzfU9yE4VS6z837Y+QPFEigYso9zRmHi9WE+A7i0KbP
zZ1LMX/7yfVK84m1VreO0kk0hr+Z0xFTPumds9QheZ7bDTI1upIj5Q2MlJ6dfTlVrFHnyu4oTGyj
IGOiD53q85xc+VF8RL/2zYpv68QQsaWX0xk8muQbXDxeNzAgChQ8pqQZmnj4LchXafic1kejwBap
cIBIlkvgH9CpOdG1Int/VkCr5ej5JLQKJwOjdjWoo/+8o7ZvENQAe5Iu7LBYj8gZ2DNESrsEBe2r
8pmG6xY3EiNfdZTlotTkyZC8fkBuPbi4fuPFECwFCAkr1XM1xi6Vz12mNf0k2ryq0BoSEPpXMEj6
0iJPYnyVvAAMti77FmOnXApKr+WZDmMK2NYD5DY0X5mBhW07zzyPni0a50DTCYp6f/KqUFjB87k0
JKgNn7Fs4dQaD9cUspDyxWJhPQzGMeRqs9WIR2KYGkrhoGbmT2OQnAVSUkRTiHU19DSnLu9+DbZh
jBc6NPCDQlXkDcLrME9ccxjEUx0Mv3cLZdViuBfbWBUa9z7OJPfN+1nIiXFIJ1C+MCS6wFazI/Py
ejGpauT9vXm3ohrg8CD9DmyeAiS3G3m0ukgtHRCqHWeojPBRFB0d3AWyp8eFoSXURoDxZ98b+xvu
GqPEodc7c0ZY4yuYZNP+8pIRguq3fJrklau4vIp7wwgwJGSEf1paAbYE6gU0hE0JJB8CbSndwTov
Lp1hsMFw4fnTRYZniNsl1TxTJrFRnc3bE60d5z+Zitk8HokDpSRiaOdSgab6+RokHIej/yHBVH2Q
bqSiZonhLUTChdmhzzw1Pr+MRSqm1CeyOMP8xjq2W3Bjdh5dAxoxKG2H2c4wTgAT1NIdjQM10bVO
y3GWzje71Dymx0dTiWlMrghBXoixtzta/5xJ+Enc57WD1NBwxFxc4c9aRFff2c9fxrpbCGdebzgn
yzlQ+aNSlIUzhhhUzZfmHg7rFQFex7sJ0QD9NOMeaTuTbRtfQmwkSdqKexam+FndyvjQGEBG9lNz
VYLOPorxH4VdXExp/sBvRza3t4Q3zQpoOYB6ISAo6Tcx9whdtpA7Hyfm7luVEgZpAEM5hpYBz80f
nKakkKVc/w16VDrxrzqKAC5CyGxX/0CKdoMdq6l3MMsegN3n+4fkcGV/aUPhW9HAKvJWGeqKxVs/
QdeMWO4ttuVFg+1bizq+Rp2Wsoo3ibFPTJIvX4GVLfnTskPtBnyPkwkyoY33ZhuM/KQYxUHrvjhr
pR+RIZmRkRwnfQs85Rj1SfCt4MXem15Iqo0l0ZkbXIsZZE9c99gTplsbZdcnESCdOhFbXL5/KMgu
GJnOrbWuEOsO5d+xAFZp06EAvBN0+XoEK5ruTNRJ7lvoJtCPvbRHriM5BdstJfuDFMw98Hn03OKL
ThVvCkXiQP3pUn4YWhxtZ0sYUDXJ+GH3LtAMqLFwgzN3x1ayx8YaLsX4Zt5KQ/6k5WrLhvKmnm9F
pqF6xUnbq/l/SSH6KlU/7WiIACFveLCOrBFTjsnpN/RoUtHgsw3Gwc8xvnrf31EhHmAVOWC26qBr
CrqRgrrvxFiq1lXQ/sPIdgVmdyv1VqJynCJOkk6aX98Ci2qPrR6yFZIK11mFGjvvPMmmXM6q14lZ
wz+29idaYhcC7tmJti+RTcYxju1p2fz+wmlk16gWCBj1w1vCf2yHBF5HZ9edmSiMXr7LPJDEYaoq
oCT4vIk2FTHu3IyeQfMw4GD6i4lN7W9anBDweUc5tOk38ySU00PrwW3yDBhQf6z3JMf9yewsuIeU
ZXvxoA1ZvDy4rE5w0Vm0AlQbsHAqSRROvLDMPBsOwz8AEeefpf6jqOO62NbGgP0j+W6r98tlUiSP
igs1k8fiWMjgmSsQMVsPmMXSqgdC51zxtjAvZf41xVK2LbIAE9JbjPkXJnKvIIhiyvcROUwoQ6FM
2rg9yNT59nlYcHUG+be5NsFtaPg1lLfQSO6szMqw0sCfUE5VDCTm4WoyJZ4U2aumQmbjrvNDmyzb
xZAEr/8P5cr3gcVPyLSgAE0Mmyy7etNhNKtN1ZxP5JWZb4iHFwi3fBL8oDTW2stV+K0SkFIGVR+X
6ZPKQDWXPYhrKDkObFhzCkSqjnVlamvqvifgQGqyvrzBBOIMRR9IG11wV2XaQmpLUy9eD2273rjE
/t8r908zQXq7abk7wM6uiBrUGue99jWfT2mwiCjLUEIKeNksLmeelYG1WNM6RXSPlkz6YjCX6H5Z
r9BA6mq/LMoKLDPVUqkac0Ur70ftALSKYXAOhvmA+kvGUTwiqW5g/k6MNiECOwnZBwDYTdZFWQUX
044ps10SKlmp0UZlVNcxKi2IZ+DvNRbOvxmk8k5s3OxDWST3QabCcOebdNOTIl2ri1cSbl3aeA9f
H6sH561YhXymfMQ0vKtagREpBZKhLPcSOxAlh3AxSF8YEdOStMWqYaGbbmgMutmRexvwA6bYbH96
l9tGc220LSzPVUELw/h3mUg0rGXn5BP0oTWejmmp3jI+vL7Ez4xrznr+iLlEGNGRGLWSrk/d6Iyu
/CUplq5YlXJyD8H7c6S6aKqlnuQLSbplDpuuC6atYZPWzLy7KpM2rph/8jzLyNYx5ABw7THO6jFR
aK0YZbvetShD9aLdvHOmKlmERM+ma340WEMWZz6Xj/YyvVD16bXKJxT1rZbJCV5xEmAihzNzbvsc
NkBHammiwbOvXQdRsoFF0iujxDZN46S9y5ur5mMPisn2zCTlZudDgFVhuLDJthDLaQobWOpU2V9N
E7vekYGEt7X5Dvjaap8Wtu9SjKjZykRtw+5c7+1TOX2u9HTgi4dPuMflDCyTe74mZQZ6yhhIkH1f
t5T/3YSA20/dQG0jv3nRcYj8YHWaexV4v9HSDnpBi8HTN3TaiSK5OVlxiHsWYc34JiBMPwliG+MK
WWeFqZJYu1AvQQ0wIgsiGU/YDB0Tqw/Mj1Ec79NBna9kRQHcDgzvqJe+AVHHRWjQsfgHt+D42Wba
UMBEv/6Ot++TzkQawyF8jl/0XTxLHxdJSebqYJG9aj8D63SkYeaHL2je0XK4TIWgM1CJTER97B+m
qgkilgc0xGkmjlKpsnSN5rCK2kanviCeU7+tUPsr4zByYatNqkMHiY3PCnAvTKTiOWKLaNXM5j4O
+5KsjLhfJvdAhZqx8em0skMmGBYbfR4e6boJhsdCcTgVViVhfFAlPnkpLq1mMDh4h5JLfbHgEAuX
aaKVNbvvrQhGtRpxODyrTJpyBAl0cBZByiDgxwkU6jCs4zm59bB1bW7vMLkyTn8dnlAsP05L+qM2
rEVfUWgpjNPcbB6sEykZ9f8TUCIUGt3LyHbROswjLZ1fkv9MqsC6R2RyWY1baCzWjHEh7xMg6Tdj
tkgXueixmmocgY0KwyL2YxGwfXbPA4KEc7RIJk5pDm7uLVRkXAH2eO8EQj2hvtmXaE/X7bkn2zHh
vAw8kWetol3ex4mJFEmrowi8SuWZqdumyihBRHbxjAoWHjyukxroDyDw4lZAxbhUUhiStYtJGCXS
Cng0liR8tNeHBP5qGdAGY6Tn1dGsYsX2uIi0e+ky/f1SfU2HExw9DlUFc9ad2TtrwPHxsgzE991r
fujyoBi/b3+sWD38Wd14/9qpJOrW5gTCkk1t3NAdgz9PeqxCaenBAMmN+Wal9b55uV67FNJqcT3V
BaphVFt9giS1vhccZScdh67mYSR6C3/gCyeDPjuNaoBsrN+eSTP6ghj0dqNyaaFsP+XVwgJiuNfk
kcna9tLZ9RTvBRvqlSZYgMIGWYBFMOrEAkvtem1a5ETLdEQ4P+Yjhsdm3sLpf0ZqOewCCmz2ETkW
x2shq3eRl+SJZ6IVik2tEBfoamPvUEq8bX5JqywUxTAlkAw2/Y3Vd4XLjPa4zlkg6vpenos+Z83N
1g0oaEZYchZn+14G9BWCYTjnMFPLXjX6lfR6TSxlwBLQbh3Dngek1cVXKYYWRX3yn3eEgIsBjwKh
nt8tEk63Yx0F73JpqspYM0OuXWyiJtD8B5mDwNodCewSc+BetStybAxz6tD89Aw5JdDUj/LzJgt4
/FYFGuafnklrZgEYWRRV8BaXA39+2FCAIb0kpIl8Srg/9uRP5Eb99WjEvexjHiM2axzZ4pT3e/0G
5T3k1vzC5vtU3rZAJ0v22JajpRwWvo3gDIiqnY+LmkzzKN4xlE5F+vcVFPvZgF7MJTqKPi1Tfnxc
O0SvGe77RmenJB/ZoCkW13mgfobk8Y/PdF61CF/Ow5Qecik+G6bcK6PVR54MEhgVFFk08FaYyQn4
zwJESjDsThPWyVA3gDeAVwmh5yYjqMRkTziqQ6z5xq3HJqUpfWd51w4DSQIkwJP+UjU6d1asii8L
apOBJD/OMOGzupWyZa5MUGeH9Kn83OSpooa+2q0paC/8aUvXkkQzQy8lc7LD6LHwuDYYN+Zms+Bg
4JRq0D80XZPHhqe5DGO7md6Tejhgeq0hrcgmrpQm+vZoitcuWXaGPfrcS0UVECUvOOc7Q1rpcqzC
CdcpYP9O8xEF6VrvGdFOdK/mmmxdg86SAnq/7++qXNSHWCeFlPdYoxYxf56rWOzxfvMlaDGBmeVR
lILd7sebgaIixpR0EbDC886tJ9GBZSrRdKKfcIMTqZSzABSF++27C70o7drYmDcaYSk2ZRemY+KM
jmHB5fRnAtmMvVp8Q/vPg9m3F18zodDqg18LnPtgVGi8WNkEI6ok0yj/lTs9WFDJgpwnm2wqAwy9
mr9WbfwdRVz5woYAOqpg85jmWhGcmkZsfHCi8MnIA800Gjc2ZCrFOJmm+nfrByUakz32XWNIITiG
qVKxNTkjuI/MGP5AxHJlYST8xrYLV2XvmCX59VbQeMPGv1sgNruem5ZM/RCPywzWmcRlzthj7FEM
TlUAtWhnOVoHWKlgF1vNOeU1KQcI/oZRWtvkBHeSCQSbbwK3RAHrm6R395XU9NMNMallU7jSRE5r
ln/B9PNRP/vZKuu0FftZpWTgtyfvLuFbO9brxGdaW2i5CrUur/N6O3iapbCCDszRejh3TPf3/Ina
I0BiwL40j/NiAumc5jHOEa5p7FsALWf1KWv8kb0x9iDxfFvv+xaiGNJRt/75EXph8hgWdEbBX+OT
3yF8cJp2mIMAibOcOSoMl0AvVP1vGNAHzjvjMY8rbsSGG6DUXDSeEdveqYgthA6pMwtZC4uCYB6q
S1WCiChRIS4y06v2zAQbdLCOVjbL2k1Tb6oQIl+5kOxtAw4n2FQHxWnqWRLQUN8CzVYnfVw4OhXk
8WIEtYcq6h0MhCPjB17E8Os2NNEJFpXivpYQo3naIo0QfqKRlMzKM1xIWfRsuQLVQRv5GBr11jMp
Sda7voEUz+gHpO6SR5Fa9qjfC7kWgJNQqpHUpHV9IQdJ26q7On6ABAN4v0FsSzavQawENG8n/FjG
sHJFqhJf0WkWRwlCKnPtWM0gAnUJAxUu7KZoaOOCs+mubiqwDmhS8YkqVMfxBnBNKB3bXUFYzo5E
buxyOSImCU+quoLGm/wnbijQnqoVTohkPoA9ME3EEeyEg//H4yijHzeSa7WkIy+vjWAIyYB+8dJI
hx2SYWAOJgqN6y5/ZW4qheiOvkkxucz6xF6j5Dcf8MbYfoBmRhICsW1OB4PSg3sSE0lC5aNmlODN
SkYsTk0NHu/3+gGE26jaQFNg/Gr4aATgPD8yU9D0FsY2ftwM8x3NuA7ClHIlJJQD/UYJYu3TcPf2
tIKAx1a4dQcwUJHUYd0kcQd4mI/4JJkYXAyjHf/976eJq4Tu0XZleta6bLfkLxCZPR/hd31z6nQD
kNp4hNHCfWTWK3BnXXnS1fHyGZZ/qy/cJQAQQROd3Wp0IsZ46UvJjBghH64aiRDNZBbAOhwAz9K2
n9Bu0ZkqbduVbdZ903nyAmM0mSJGWjCuzqSgXnavP/voIV/RwryilVUm+776ZNSICLJr1I/3tIF1
VhuNxFcfOacV0owqg5zOSROEjwmxEJXdRKIVnmLqQUoDa9SaRNvvDvWJ0x37UkrDHSGCFGrHX01x
MA0rddl/0HDDl+ngTns2t8ZffIsWZU3VXuoDhzd45Gejkqsl/8SGL3r0v2+Uq2FNvf+pdTDLSBV1
t1WUEBweBYoyQLjd16ivTNZQZ7T+UWcorp8re7Lx6AeTmkr3AgwwwWVD3+ymyMOdZZesW9jWpAnt
FJEFOLiWdAtsUwCf6jqRF1tGlutQ8uRn5PHA780b34HMjAr8fxm5PkeW8/ZqM/JTXRYfjIpDx27z
dwc41AsJAqZeynCklivttRWUNACYBLOb9uvOJdYQ4CQ4hKuX3/W3FbgyIeB1u/txjl32PUhttN9x
D9qDYeDa+hcLvR591ad6a4EgyPqFf3XezllQnrF6S98kay/mmtL2b9HB51U/njFrjJM6h3ZPOrrO
D1Q2UPw7KiP/8iOsMjpk0gvWcNys0EQQJJmNcVXYy7v92XhxR0Yqc32YXzZ6UOUV5nN0Yqozcs63
0ut2M/tqtCf/rGgvCuKyAKBXOwGzYUruYmq92xz6oUjYkLlgoQbSIxYTKZacy3g4Za1dNo2T5odf
bgTpGMfYzfGkt8ZWSjqCL7PIVZnHC90Zx7ThWYdzVpj7XS3Nd0IEHOIqV2U3IQVNk1iLVSrmlp1c
Zy5/FARMjgf7rNXhbOFaBJw2khi8l9mQgQzYjeuYILzqP8hsivEKaDuRtk44jSxG3I8mTh3+SN8N
ipujus+4fCzy8VbPEy0RZVY/ItFlYkzf0GqdbWoubuPEsDjFVJeUBbwo9K+GByH+1LpNjCuW+ppl
bbkkLcZI4UIToTRgfEEheUcUDXvrAOxW4TRsnQRJgTVAe1RI89BKnDKL3yLWf16+D69asxm0btPe
Imcq88C4zMXAnYoG9O/zVhaXMW/u6DYHvMESh5dFzXNdUZp03iBnOr46fDk6xsQ/ZCp56t65jYS8
COMWS4iBuJHM8jrdL4jgUaz1w1QsDqNLZCAKgJSBCVRlUrrYBTHFnTCWc0ahaA+Ci2bw0zN44Jrj
q3M8Wlhsc+sF2nYO3RjCZy0fosCG8HtOskyDpiRVnXBQx3V3PBvNMTiITXhbtcArieONmXiP7BfE
s12iPd6cQlDcJNw13wuCBQMdFPyrKwdL4gtupOc1FjNpDc+Vvt5PlMRDdfbWpb/NgghtWc2PmORc
fluGGUgBOn+BoVLDLRn5lp67B5RdyRoJMXgv4w6wop6RDWi9R8IAQo7w0820fJJTpzT0/Oz2APw6
Mtu817hEyvpnz4c9KH4ys4omcLbFpayMHNo+xH38DwcMR81CsISTH/r7AI1/eAkbFekaxw5Kkz7I
1H648PPKwQLhT8haOy8L3LSntAcQHpH7e7YLeYeY21Ky/4ZN2albkMuteVhrG1/iR5GvCfxo2sNe
2oG4yM0nrBhFtzEAkxd1Po0YxNyM++sZL8LYLs+rDox6tQJOPwaoyxZ0C+nJHSuEjpCX1BuymKni
ziP73C2xdMTa4ibtZe3hzq9F5KiZfaeXKyD3139v7sqiQwk1wnT3ZGqtHzq59bNtt01h62retIDf
h280VRslUCtss7DUd/YZgTxk5TMHaJLr6PDOhdaoYZFcGm2EOAv9Bbk7ks3iPUJTHlqJVcEc+Vo+
nSqg/ujCrB7x2EfAXnbry3B4/xmWI3hwkyvJQwyOuJSg49bd1Xr5z+IMq6F89MMxw3GqGi+fmoZn
2iJTekaOISI3r6y5G8Y2xnOuHb9bLQgkPsdJqoVLSfF6Yd+pg+1fpcq/FH+QD+hBp6raIiwes3fY
kmre8eKyrv27yS++3Ij/X2B9vknLlixKCxDOC54Y2wQ5WdUqSiJ6k5VrVGSzPBA3RFSne9Znr4JB
At+9IsXNo2o5oW4CaG0yUfbmRhWuWqeAPbw3Zr3m4OpHQEkFFKjOQsWKGar8WlbHvNsHLxO6uawd
M2G3v5ikv1+QUEMs9kAzTEwadwCzoIXqh+yVvaDmmolteEZYwHkcvqP28O9LcZsxDjYjWiWyO2uE
rNDiwkKxzb5ddU0YjDvNGdouX6h7crx3Hbh5ihr7Lu1D6PTgImdi77hSPo22+4mOispjPBa/ldpB
oItf3tk0LPkdQIOZ1xtL1SjTLlKh0cYDske78TqBKEza318R98cpYJBEjkeZNkAjJmDCKBIG2VSQ
/1n6BYAihqar2paJw/mAxsnI497bBtwqScJW/8J+CLBFlzp/jxnm2TiP51zHMLtiWPJvG28NH2xg
mj8ha5DfYbzFXUDduXVOQjjWqZKzMi0PsFBl+YWvhyB4g9vkw6Ba5wAW4aorSNoKcGELjSm3d4c0
khxjUc9bvHOpRud853vXCIWUyDGyN9pub0hfet/NakKQmrJsNsMI8VSYLSrA94hFuJ6nAZZdETS1
xCm+ozJby2NjG+sFCOupGXo8zdpj4zd4hwpcq2AIGvQAf1z720ZSPHNTSF+NsXBU+gOaq3bL/YJl
kp+7EPrhbgjt0Hr1JkFrzgp0M/oSKD/cEbRDtRbAC9BAOGMZWIOrfzICdK/IO6NBuFhCL12DHVhq
YPS+iNagkBL2F++Y/b5q53VNW1makL0OSRGfzIOUtpePz8Of15yU4ZBgHK/XRcbMMKrt51ieDQvd
WAFF2EWOqslRUuL/eF0MtQu/O1tuIuMqbfxR0hj3NHdSGeA0aT8JXZ3grUr0B8yVx26pM0cxZWBY
pLZsQFDIVQSiTcz7PLuIQvDP2998OUcYh7T8tvbyAtFA9s9qh0TS4I+fOB9M+hlH7mlWJBW1J9TZ
7kGUwsYNYE+GIgOMesmtprK2cFMvVsC3L/tg3HgWpwgQQsB9sutm4xQaxY/QFP8ReTZOLu1PdOMD
klVut6ag/2u8pMDUjJs2sCsycKEFors7VdquW4idb+wyEgvNA/2BUsvFtFUcomZQESI9/D5CMWAx
dwPpTAzh3/h0Era6zXwneGOscmJH7lCIYbEF81r8UIT7A5eDfZsnXLDcw5n46S7t+KiY2dvBNRnI
tHx5HRfK5qDEWJSBqACzIzFd33Lm+3rxX5qobI+GeJDGbwyAou/hCbUdMZgarlAyb6DbuasFX5S7
ACnbr9gSmQQNQy68iNz184wUCjxdkn5163x8Sf6LOX+I3hzaLF83BZDgVcG2qAmDMawiFBAr4Jeh
/jGtzh4p3KC+qvqFATrDcYNB3qhs9Qxw9APqAxy8okMCbx9Bs60F7OElLxtMoMONIwV9LSynt+WZ
N+T1CZgw88ugipzaFkxUSADwhTk48M094BaL/NPFES/9APrggmU+OPcd3KJQvPg3Km5eDVBOlUSU
wsGwZJ+sh78kWXO1ZB0/UUMOjuczr+DAaRALMVGirGDPsU1iIxONC8hNffH3cZHKlqaRr/arQrz0
apwIe2l3PFWqMxF4lmRKSUCTxoAToBH8tmbw+kanFHHITbb1arkEEUXXJgRqNZKeluCelbnh851U
7mzJ+cuVv6bOTemMtTk3bxlp8rX1VBTo1PrVqrrjHEtY3hnfHCiB2qYVh8aiKPSc8twDkIrn7oId
osXE2kfCaeXbT406S9RMGI9LtlNys7IOPIYOrFdkbljgpc8RnpFmm9oQfxXpB2NBIIQpliMYFbGh
EBBqyrX12n1vr88BT9DeEueLNzGq04ZoOqJY5JjKLfsJfhnL0qAOzUCobZG7MPxJs4VKLkbLNXzn
m56La5ePyvD47NRa5dlbfWUV/PL40iO9enzA5WlNNwWtguhkHLYS/bT0EA23gRmLuBVgeqy/PpBG
c8ZSj9eDhrhkq/DigRcmUk00z58x4XlLyRmVNXrdvQNWCdGqWdIz3c2H/XyyqNc+ZEukx2OpJxNo
yzboQ+D7zggEyFh/n9SV234JD+zK8TV7TXz5jcohRJVfn71xLYfJJMbmkxFwcBUa5lusJqMWVPpX
JPxLEZMSjfkWi4yQag4pmSaW/Z6+me83Es/RL8eeUeLEE2fHlDpILB/9jPRUPvPUX+WKsKXqS+o4
DlBwNCluIRF9ylfeaub1XjWnRtZN8X9EoyuLX9EGhW0NcivkEfdb6ofWHRuj8VbFaCI01S+ze4Vp
PyeJS/+aiOqK2QDA/h9o4pYIaDNZ+A/TVMT5kt8rGMn+qpwm4qcEX2yvSZLx8sQqPMYJ2Dy6zP4H
DTFzvWSKnKB2/85NeHNSOXon3zkgXU4ZYrH+AaP973EScYzJ3BlusO2ol245E61KYiX2aXpd4ORv
dQsAOI4jW+0ZeE12/cYRVi9lRgmDruz08KOUS9kXznUo0obqfD2wp4vlGoMQRRbV2o8wug7dk53I
Ny7l86sxL7yhkTgU1ZDBLx/sVpHsfsXm5bo0IeBNkilL77b9cXdXSQWh6KExlwrsnboeQgYH1RFu
rG6GlqeQ/P3pjUbtO4ZkjDwmRnxkTulsHenP0BgyPRs9YjyosuHRFa9XHejEcFa/402PEZHSS7CS
LEHJgTtu/jIU2mr8hiB/tDtIUhvfYr560kW/okfSqX6gtWK+aYqUMLh0Y+s/Fx2eKLbPHysoMHKN
V3HL4T3LFuWabXMq/qgRM1f6T5I9PynVHlY9gf0/3ABNVKeIVLsyz+96EeKv3ExQ60OatsYWo908
x+/757zbiak1lkRBLm8Sy2NEKnY3jUEiButlNzLvQ+eDlmPm9p2oN7XwouUwNruV8Gi43xXsFi1W
NGX9PhXkRFMAqudyyCtV+ad8b9Cvq67CbIXOD3sGHm8KMygvu8TidwgeXMf9vMveh+3yovtcq+Lk
3yHsnkUFlk8SY7G+y8+2ZRYNX81flI04rDP3QrKYoJtVufa2Ey+ijqMJq/iOFXtmjevg1GxTwxRX
VTPQBViaOBw906v9ETe44K0bXW57oZmC0YkcbzA/vl9BAIbtdkTSen6uH+s0FUwSoKZ5hZv/KABJ
zocQLtNZzvsspeTTH1BT5+hkuQcy8LmuNpEFqkDvXVdbCOzeWgkaUGk5gOI6pgSbFxZcN6AUIQe1
twqPAktopWRIv02yW4nKkBh7KKyiWVD6RbXR9JJGypg/lzyzx7mCnDd0RZXpaJp+jLgFBioOY8Mo
rFSfMw59v9e+OKcvzL0xobGuNifoxCJquVwMkYRhPovai186xgtRuTcROdcvpZoUoz9cqiufdD/5
bB8vrd6Szu5Zt1ozCWCjL/32MqDVdYWBuU05fCqsTKloiVOsWxFdM85DTXwSiVQ2Go5ViksIDOnW
5CoaZyYg3rBatarwGqLM1kp0t8s30IMkmyf249KxnaR789F7vlDPrIbXDiVkDgXoal0zKDlTsEJY
4stJEE03UQSuHVhahwM6Ht8oI33CcnRlw6CVS3/pDY/hw24kivm26cfXIOwEA5yq7dLBxjiwqCJf
dzyEpaqJOJJkSUbd+jHinM+K9t9B8Za0UAaf35qjLPczmzq86G1BwOlwgJQkseMxGEKoYq1P7kFB
+3Z9G1q7FmyyP4wGuJKt5MiJ+nMJwBom0yjR8IlReuPsS1mybTMf8d8mek7xkv7cHfiE/kYlNqon
QRWnhXAWL56WgYC1JedY9NaQcWL1Cw2M2tOZVUv+IFoZQKisUhppQmqhUIOECl3rNc7aB/GRsqPL
PYgugwpWWIU1dF8duZk+JMBqkkKClZ6n6HPP0MsL2FS8oOcbe1Y+CFevuSIgJnaMe0eeNYEmDMHH
9WCneeCpmIJedpRn6ZUGAID+cyU54Cd3aPAcDR0srV9nrpXRlgs94HdLeUsAyMs/FHsl+qqE21Ft
Qa2AR8yLBFMTI1DyFQXYIEAsf+QODAdUkhXB23tkhBlLv3HBTFkvmPlRvt35IQCVYiP1cDBiG5Mh
q5TLIsLPFmQlL3UeyYadtk1V3UmnXWLT43AKvPdxtK4YK99fzKn4U2TKHoBAdjqKxIn6m9qc1yMD
vb0AE4NytTaJU+Szk9mXqfux6DscabteRmdj2CxY8p0F9GG8HqXe4fNEvzdTSUPHFg7nprB1oYXN
jukgQS3AlesMe5BCCTIWCBzaNl4DZ5mQjViw/BZSpbruRnpKyzvO6aCcGPYVY6kgmd1kAiuG60fV
l/ytx5ywqhT9Re9kdAnsN5ArUyZfIRpHSy3GcN/DKriJ+KKu6w54P7b6G8b6wvps1W0lGHfkQ2MP
TIVxPQt/0xsenTLqLLK/zVvELf9hDm+Jdo3L5dI/urDUfRTza06XrBZdQ+sD3eY8Dd4rxeUE2lix
f+YvbxuiLJDOTH7RMEvLvp8Lj1JCCevmKBG+9gqhXppsE+ZxsvX8aXmr2PfUIqfHvlkj5ZAoSYtb
d4q28ECD/BmRB7rRQarZMS1Dnj2b3ifSCFP8DKZjBZFHi580r+fhTsAf6GO/LQvw69Qzy3Btq1d1
rmV7Y2guLwhhl/7eLpzLub6TBSIquXUha5WjkBcDbjIT556u1bFwzd2UM4LtjXGwyTIz+xJ7Lo8n
V1YqLGH8lp2Hbe0mZGktt4ff0ikr8nhrZkwe2IuRlU5qHEfQcl9H4bOGWPlJly8s16PvYr3BJVq/
tKsskr3pRlxTkTPAF8AjgdOnKOzJgGYWKckNoctZi6zeeMBKFjtgh15lI+I3oc6Vb2agIFNlt8Bg
GOsTTOMjxMxAjziLUD2G1bV5IqhbVftO+5kxAApvIkpT4F/WoZXuSeBkB3K+P2UXB6jpt/vN0Hii
Qw6NG2TcJ6bEO/0s5IwfUydMVSmX2SynprRYcnb00VhRUkZosxC7xwpHQLTZxvTkl8vBybBckPhV
yUeAoTvqKbU4ngEXFrhUdswhaYBiOnqd9QjTrEc65X6aiI5C6XPyyMtUPr9D7GooFqgS915NVTWm
kYPgaEj6a2YFQ775YZhvd3dZW/0nGI7NkDk+K2XeGOXvvFxRo2s8+XFJv/DafczVoSxbCkK4iVjs
0JXsFv9ftSPus0NwcObadLldTjDZz38jn7KzhLsioROD8dWge6LjVALzL2MKPI6J25R8g2vhoxnT
KuPudHElQzvAkoKiLRBvI24hF17eZt2X1boLrx0rPcSJ/htx1GIkBwSBYdsqc9LoQf/PVCt+Qqtg
DXsAVYLM6fM1Q31cbqkchAykuD5w7bouUV5dniUrKFXuJzPb8dS0/t0TTwqfw5lT1+lyVTZ+KE5R
RalYBxbWPxfv8oWKkqDcG1aSUGVwPtXCmULOiWoP18ui/CFF6LFUUtURwHCaWCsbFYDym5Ih8ALu
9W9AKjJ0jH2NHBZIxYBNZBId0iHL2cAuZzyTNjTl7rEq5G17J8wMACLy581/bL1S/5vf5yLjqsjS
vDyDXmZegvz8i3G7oNS3+NG/c1wbyq8E07+Gd7ahmL1/Fx8tqSFffNRd4c20MGNpw5MFKOfBNrp1
LdG/F2+3kqfG+iJNO/TfkPAn6HG47kAIymsrDW+swBmzmmEDnzZZfRNRUZAZQXzs9mOAyvkKYxJI
fOb2tikoHxL3KbtXk+2XTcM5//rJKtkQW7+Hm4muRNy+9RGQF2qHX5Mbz20E/K3Jpqj+VdLMf6xK
Sx/dEvIYUQkA9c6G2okWPujjqZgNkP5XrAdXeisBUSg8abAqs0rPQAVj5Y1QU0ZezkBQ5K1QG0gC
TUVsOKnzn44LD5toZW7l2ogxKQMUQwMiWcLiy5aWlSN1qH73clk2QKoSrbaaEEPPXdILIpXGyJC/
0nznd7hPFpuMXd7TILeOGap//95KhKUPfp0+PuM3xPlJ+VVDIIAjMZHWwonIsw1OI1xTMX4h9l8I
Yuh5GVfbuck1FHnRddzdBWao4qbFVRKBzc8ZprZAR3qCxvKTREtk+1bFFIDsk9Z0LNlFVGpkaAL+
6WPK7w+oGQuBSUGiIG+hND6wMZLytp/qUXTAjHeV5GZ0pug1edesXUjym0GwP28VJ8T6uaIDpitv
VJ9hSBLijHvLw39CACN+51to27eQHFl2ehaEU36RkwOjEUnl419sl7TBGGQdH3nepMGC3gb82F41
u0NhLHqCURaLmOz94HVhlz7Mm4rxaOk6gLGhzhKGjFIjoeR4USI1knZB2xtREI9UyA4BX/rhxYKs
DZyaODvLFsK6ghyYPCj2TwbxluqXiVNGeL4ZWjDYRkGJru5H/vP7UuP/jsmjm6kwH0XQpSC/ZWI4
Kv0b6VDoF496P1yQNtSVxRfUj77aFd3nG7D+7KwxbomJp/L36BJUX9TMirism1LvqGF08uQ6xDTC
1in9zB2rZ/pxvapiiGi8OijDuHIxauEWodxlxLUcc82qpLmgdbjdvUp3sPlzggy+U8TArB2E72dn
nSrCa8cjE3wR/bASAcZ+tF8bRtbFWQVk9ch7JuLrFKA1YrDQCDFCSJmpboKwpN8hILRvV1Ln8Azo
H5gfpuG+QpwYnW8/izR/UdjSn240iKYp8XVbS0hSx9wHLLhBfxc3tamOhCkF9wh3kCGNA3QHCWaf
S0ZpFViMXjN43v6b3RgPQl19kV0bSeJLCNiZoGfrqcnxZ5E9cML+RpOpEk9J8QIH9MQI72/LgEX0
ZrdNIhK5wmE+XDaOEg6EtNqHoDvaca0nQtj/nEGEuR0UdGdJsEJC9DLMIxMO1lt7WRfmRt2SbXvQ
coKcaDm3lYzLHlOh7bZfegZhGuNBDTcgfvYX/YmTrasLzbXjA0ebGRBmVzDQ5JVM3B5q2xv9WD9j
TTpCgu/pjf66jN8Y/+ZC2Qwgd2bX9h7azHPh5S/7bOhwmLhxARxSvNLL37eiC/+dBMJOlVsnmcvi
vNbT7F4hXfaXWKKU2tds+skwBCTVI300wVCiDbOtIhiFjifdNKlX8DrF0Ra0Tbu25iNmdLp4gq0k
qd49DEHgiYqWubFhWtpifUxMh5CxFejgDXUoKy64mIY/3lG8weRirQMYR16/o0NpqLgr2d2P4Bwl
f3smG9PK2nhuvT5uyC6KD7/XejoaVgzvbuNvGCzFj0YYeqx31FKtSByP60IgBG7JD16PII4BmwS9
OP2vYiTCqqtl2R9YSrvrPnXxJiPcIPkmKPpNt1YFNEPy1MHVEdD0ZFWk40mEV65/xctn5Bci/3ab
ZngNf2fhJiRGxH7f4Wxm/EDT96jvfry2/NrPb7Q+pInR5YKq6C7wlsJFHyJGe+qAAWMGq7NLavWw
Cz28w2aicr+JX8KGhRtG19WSlR/0PqJ1uGFTtJP77FMORoU1dLXsqyGJzSdO/RRR2RT6Ggmaxhn/
1ZL51jGNYirPVGDkRfsKNr0a46nZ8Hvw2gdhSurpxgVXbH3gRxTl86J0BYSoBNOZX/6mNJsr9sm/
b30E34sdLxdWaSd58qj3z9yWllx1LMTz4Y/ZLHp/8KEouRA9gv1ORS/TVArM+VWmHyCgPcV4n1Os
CB1h00IRNcnkByX/tImiQQXdu2H2U4MCDlXcvFPe8f3EDdXKGLq40kDiZF3OHfQYs9VK1z/8Nct0
uoLoBpL/6EDeq3Cr7sDQZsG2vubi0ek5BfhtVNKqfSvKSuYe9yBZhjxG0VbN7iYtqi+TleTikCfC
qLSGngqyV5i3g/wd/Du8QjsBAhYRvM2Jsp4etfTu7ioI9WUsV+W4gw4Wkr0gfHlA5p8mSTHj8THB
gGeuJemdjbOVmWxjx0A/6eRm3rX9QbNp+l1i3DKlptR3S7BhLQyU/w6w8yz45QKZ+llYmV9AOxIN
B6kqvRsgbWaAjaWo8brmLJXZaAdy6UsI5jsOHQ8gFjGaKDIQOdlI5hX3hD5gSar292w4x6nAR0j/
zWNejTA0oPHipbPg0Syqj0ilJlZ5ubwA85PxSG4ganoBQzmTkS3mCtx5AVfjUpDgbKRxp2fLtA8F
+iO6ELauD04GLUH2KZo0+RIcvyEsB0r6BfO93/gay7gO8F9FUiGEXkRMLsO/nTZVl+0lk0lUanU9
Qmp/23niEvZXBvN5WvtbqWX84mXgPEzoKuzmNIEpsSWNnSlFjlv2+hXvWZqumRhR+UMR6Rlorid3
8rYhm7y8FxcXGMSJehY3ESBHHgGcs5LzxOxhdm9E2dmI6TIvETX4K+LR9x8zxiKG8XO9ONXPUUKP
bfKWq/4ino2LkGzAP547Is2N967UIEmhIBsAtHh8x2HtSOdMnAAaZu4aAEBsho6vvcQEo1AtmLN0
Q1J4O4FK/lx+oMrr3X23VX2lptlGKPMiw6WwzeRqGMWW+3Bu17LqQms2olY3my5J6If4GPXuDplw
gLuIdkIaiTHvziSI/A/VjkkcEqfcdTbyiWnOdhe6TWdnbm2mhXcVvuH1fFD6g4XHAWPLBO1ZB3+N
L/qkrKow/XpsX7QHKIpqiRwyTT9Oe634UWGDKcVzp1ikcEYGoG1+uXYsfTqoebVZF1XPNQamgRxA
8yZ04GecpBnuFhBJKH5iGPUFglE/evkjlm2nS4pWkZkbXsom4bi7pm8KKhCUkvLNtv83At4FhA7w
eb7TFFz6YRZIZ7f8Kv0dz3SUJAccv0bLZ//E5ln012MX0ypJJiN6D1kzRJvx/QJksWYONyEI86XZ
2GoEWpuvxevhD8yTp/WYicSmyNNNlCMBV7n+IladPwEuzMKvi5m72xlkq3hDjmogf2o0MfizpYqD
MDDNBsbh2tnlMTKefUZR75yaBw+N8uz0W1BkFWh8VMnQqPa/XccFCHvDO3ipursv2N2PwRC3rsQH
EvNOXCBQFO5MuRuu50l57Zktahe46fGI1WqrKN6WCAInH78NqmJrOsAfzqLBES5yjk4a0wQQDMBG
/sflOubH+yq0SI5gc4ovXOzJ75CX49lIfhBJlP5cLj3DUaxBwJzoLyiM/HKndX/YC+e2OOq+l7cB
BJb8cahOaSHWd4oTch37ggOxm1E8exYumU3XN1O31NE0+aZ45UBY0U9iXeXdptfVqoqRzVoUpJMm
S5768tVWoKHsV67zk7WpsVsKv3wf2VGYLREQO+iYgcXB5w4qBFx+ze9ky7xnRKx93lJZfvqeE4K8
I1RAd960YQQx7z4RMuxvXORrNP6JRQjk8Iqg+4QIz4JrqVHsS7RCqgPYsMNYast8LRtOk+oTsXRs
4jjo7T3X3tnTSbUgM+uz6jgfPSZaQR/ovlKvUByrotM/mw5adZTFxhf8YoL9mZhJYmcF4ZdZRepa
id2owugdJcbgXDgo9PA8p3PjIWoQIv28aZANRr6E4YHHEZWXrs/DbOQlVcVSqVdmP0WtIo64Sr4x
rRS0CMEExkMmGQaIh+7Dwjf376HXWZ4hxI6zKVZyhUYuOI78JAWYFrGB2HSBP6YvC52H6hlEywX+
tQfX3MS056oRpGULT6dcooRkb7FzGPl03M4vnNGvsR6mxvCV4u3HK1ACLDxYIS2FSxnUiUSS3yEY
BUPvWuRLI83mj5hE2NWCmID1Ol5/ISXFKrEttL+88LQ7S1PQQtD2bHLEXr8zwN5bP1EJ4YMcQR/2
rWNlTx+vfrmgPJVmJ/2dYnqyj0EMZx+6WVv9vCrr0QrDK9aBYSl3otwdkGfqfRXkvyvXrMqHIq3X
TawoCY1XwRsaLTcLh6yzvuq90K6TivX+6RiiFZUu/tg2rBldi/I1dwdGx3mibm3unT8VlY8n3DLK
F7BPGl9h3M8Yuqg2oIcE+kAq5xEGMvQHQ8/khanJ8jErpbW+rFMJXfZj9yJqC52dkkusF+isb2GE
DvlIluR/jxHb0/0wAB8uH1UoOokMfCQ5vzMv6gP/5FxiYvGQw5ba6H34yRhgNbreWT1DupO3EKtn
O620deoaSbtsZ4dkNp44WvLGleFg5yGYaQE3B5F8SO8aNVor+ehKTIRECIvUh9p82ETEjxw57H2g
jPw2nP0g9WqwNqXKOxMEx/53e1xjabZe9UOhuo+9NDTxDzMuK4WKVy4EQqLUclSzQZNics8eFzhp
HmsRmijwdofb0+XP0HbDAceaDWW1XqnclbjF2aviKg0GR+VKY8kzVXHGuQMICuBgFCjBnEo26OLi
UKD1xe0MoEu8Wn5mZ0QTxKL1euJXNau0QI+eOF4RGEq27OeITlO9hXW5oGIE/PlJaPuAaUe/i7tk
e1Enzsu9P+kYMa2DKV085l2mD/oTngh14jqMih0tXE+v+V7HonX036rq95HGoiUSZtEgjQZCl3ov
J3CqfPoZAhzmzPXhvtHlLTqdNIcpoyKeGYlkjMxBX8adsck12NkIolmvGO0EWmS3a9YjVTRHxT/w
RsIVmOR4KuiMDAp5OurZJ1JTmMmVWaKK9XIpP2HfHAMN+9i+jAHiELlMRQ6Z6o9Tt0PTjDmYTKCH
fuFz4c5p2i+RKp3UkvTkwlNBtcS2Mcv07nIRPlq3PCvYiADL1w2qfrHagiB1gOv0XyDQf8HBat/0
64N65HyF2t2wlJJbyhZfAOM18wGznm7PCJsPrWyXwbSzg8jUViogYK/4OF54mF0+6cvZ2nzO2Zmn
EjMjlV7J8qgvWjKt2XBLa1OhpkAuEixCyGtxPEwAl0wZsA6rUgc5Lzod44LY7iV+utbIwbw9bNXQ
Z/DqlD9GaJkbgV5zMw9RUoSHmFRoJrp+LF3DSXvWvWSSkg6ysnB858a94l4Cu4BzigVpaRX3+GAy
mgn+W85P+ElU+dKpJ0NUSwEZBmr5yy0e4b2xyz73sVGESkhDKRYWMyhTb+7JNQtsspkRmMOb2bxB
ByD3tE2QHVPwYj5XyCftCTIVC9EFoAh1IRiBSp36Woqe020GvfNR2rlu/l6WXg+8mUBRIAP6mzid
VZ2d0zF+WrWErdW6mu9bGG+PpwyLymjQSLXRP2UFcgBSUs5KHE+b9T1SKUHZbfruO2SzOUlnpalm
d4INDfgYeaxxIFp7UnFYrKOdzjg1ql+J2g1P9SjJo5eBFsUeN4ZAnuCKD3O1z4cVPPZWYqLRNoTD
KHXbG43uZuK49YgofP6/p2PVYTWRaBlOj881Qn7BAaaJCaDzDDhc3pR/8pw0hv6tTHCLBWAvzSPQ
EETYdQTjFvPw8MizBvkkQhOHDAfH5xvhdyhPC6Bno40vRPJ7bjD8qr2tBvvJykeyXzysy2cT9XUw
cMwkK4kcj+RCsTrumN0uDgJ9lkRobXtenpkmcNlFpiuEuP8Gmf0x0ESLkA9TzxYTNZn2/6s16idG
EYyMcPzclmr2EFquy3Xi81wfycIUbbbqR6MzVBqGPoG7EB0XU2RvTRi3ngxWeRhFOMnzXMzsgLnD
khDeLHV8Q/nTRCXygIjkNH7Gl+EKP8Ri1wjUaB8tvem5fnoGnP/6Z25BUYWbnRRIzvxhd97XLeuA
uZfNEJsLK6vqA9yZQFoPzsUnYqh6DDqbrBM0f62Dbh30h0Ca504FhYI8NJBGs3BNUQXde+TXRqnh
q3S2oWspxwzW1WNlP6zzVcaZzmR70N25G1gSQuLFw3acOpAGxDAdglrnLiuxF5PUt/o1VWMdc6tG
t35adZYRs7oFZAGQUtclhH/fa2UHmv/xTZuVvLaCmIDvF4NKda35G+HONOsarYxjcBUYwrcpiOJ/
RnXYrZ9+bKxtVe7+GqeHIOQci2wRKwKYlJP0qUXb4nmhHI83ap8LI2wk3lhVNncUluFIbW2Nb5MP
sfwZS01p+V3+OXPwrtem1Ke17BrTtxsGChQc8iqQR9ecTxc/r21F53VPb87UFQVOUSS15h6MK/sv
xH/M5A+85gxRT4DOfzj1F59nRqeVAsR1f8Woa4pXjeLSy6m1O0rLwen68175Py88wItNGwkR0c9D
Kne8s5+FoKMNAAzY1rWwXa3waQkq/6WawZR1cQmzMgi9iz7jpj3dIjlSzq4RXKAvrQKKuW5CNPpE
gQ3s0GJ3NACuyuH6NzGv28zmq/iMMtG1fYO6YLeT4gdP6bHWqsam4LgU0X+LBqjy+yv2U56FQqVz
hjcDwG0GXYYQZlWURDScuEch//MbgDYk+20X14tUzoN6ya+32lt+KsfwrIvjjgjppwdi2KxaDyAQ
/VfFR3rFx8UH2xfFGcGRSVeSEWg8HG3xfQOsrts/eCljBb+vJCCpDU4fXgQ5c24MEOc+gaLsJu9x
o0ierZQRbmUBaLpbYwYKWotMYN9Bhi17XTV2adNv2YfWSW100F4+n/MaVCim6ujZt9wmlcTaUqzv
L3sSreVqxwF4mKGGkbp0+RsLipn3buGnGn1+gdJStvd4f5+OXWCCy8n0yt5jF0xuU1gJwzBt5hK5
ALLyjtP1vlBCyh8BzvsPnIlbISpo2q3z3QA3EoqllDqoAI150sMQDcrktdcEKdKryyfPlXwQE/o0
ZTe3ahjp5LNRHCalKrvaYQuJzQjDVGIx/qL0bj1irWWSIgq7qzmDHiLIaQlKNLZneR41UbzsKEEw
3uj8APjM1m5bduntrs5S6aJRbWsgs+igvmQ9OEIsmDyPyrGPqTs5aORNz9nM461l1AFkkFW8HBen
gg9N5YgOhf1GLtJKtXGytmaOsWkscN0DrSOdk4EnZXhsbVXPzBhjPEKswQ5364mRNEsTWbdekeyA
bsgb55p6y5U1KJYXKaQtSR/suKSqW8kNn7JNlCZ2ywJxuu9G+OQIcaLXIG10uczkh6pfATRxt0VV
wmJIM5LteYGmg/AUU4HgaljRzipFyyo3IkqF2FNp0Fk+VF3LbuA+t/ITCJrJVTbUNDDZeltWesnO
ZIFxTa/Tzai/+BJj0vJOZxVbVrez1EAGzJJfJKBkWRUYWLu3nZrBafLqMVt2OhRH7HsWDfhw5arO
HTcn8VEtl60lRr0qNb0ipi1JXVLy+dmZYS2MuLrQeNTRmBUei+HC5OV/KcSOw4xJjPXxl679bDpw
j6ZS0gnUF91NmZvYU7xkc0+06p/MK2mmg3/5H7dtgAJBUKNVKG+NZNsSYSRFDlmMI5RRiCrXt9i9
VuNCNlxC6NOjhM+dlSGvuacLQgeLEleo6gEjHkgbGC+klL10vHW82FL6NocJBOpU6FOorKM3uClL
3K+SdXMvuyy3+Sd9umzdC2sO5RrUz1O3Ih+8iS5DH5zOyHbtGCBPwCNbNzEkyNziXJ+unPaQJe15
lEINsU7WHrN11wczv49jEkc9PyRWrKl/VhLVJB8bULcde57XCwuIsgqbQfEZCDXX6bWokfMQ6pq2
1aPSc7zoetnN58PFVB2/5Zjgptvc2ISysC+t+lncnkDizzw8faPxc5L4aGVIErBkF3uHbEpcX1N1
edOwHpwjLVWmGbfxpQ5w2B4Jx7Ml32SkW01Y3zQvIqTRSyQCVpQOcKq8cdikWX3cfdyKSZ8Pt+st
oMoGgn2olB7v+igkzcvBa467+Ur/qV7CyZ36Gek5+N1XiwknqR6M2TKWOMnkrJn1m0vqiuOR7OIr
zQoRyMvMRa5eipDrtNeHtnoBCk8D5Ur2V2zFZq8OvISHJOPaCJneqnwk7tcqz3F6+yY++nAWtE2R
eDLIrpAHYklPZNcM9fmWpXElodf4yP/GIfdslhCzljO8ioHwZxRQR2hWWrtoD9bsev3f+4XtWEyG
NsqO1d5i4xBo3dQR80PlENfr+i3kIDN6vZ7pSx9yFXKL/QKh1wfhN6uJyPCRxTclmjiZu2lZzEUx
YebV5ROLz2wT88dDLaqqrOi2f415pFrIFEiid0cw1QkUj9rhpnYL3fZ+pwdpaBY1fZ+SmaKaaAg3
k6sf36oSHZ2InGzejTGnm8yENfDTpRC6inO2jHJRxvSyw2/DFIxbSP2e46u28w66lcOX5gRkHyOr
qO6UjQPnBl0eOXRckOjfnJ/+ZLRpVkBi83GtRdt9NCKNN4U0jKt4C/ad7d4Rt1u56vA2pWwfgKW8
jzBtdo7oZyXAUj3Hnx6kzcp0ZeEzZOCL4tsPu/tYvKvQ4JCzzN/vg/FMBe3BZ3ATKWOd5amhjRQP
nHp3nsi7NkIrwGTJT6woZkl3qKX0q2SpD9ceEQGHgWaVWacmRw4XMY+PDhDcW71aRy+ZoTLuex3z
OdV/Twzsw3It3+ZmaLA9mMOU+rK1y4BIsPK852fuJeNfSL+8ualNrGDsoNcgFKG23evrUIfu7IGH
WiU3wTMcTcHgdrPA6lx6lBStqk27lDbgdkGL0Yz8PqhXawHjh/v/WXlCqROFRzcLmGAuuKx+zfZ+
MOrXdDjXc4sVRZcyhePlPrjs2+hEzpWUDkzRw8/x6hITD5BZ9NfpmnwD2ANdygzp1lUL8KSQpofN
e3EciHmN3vzRfpcKFbS+pGyDA15VBK9X6ctC05A2Bb4EAm8ovCsPjjUum4Ix+2jiIUQqUuf9lGfT
4P+60FFfeltMOS3x0NegC3l9hTi940SxGCnruZ31RpmgNIVF87beTFDsKZRkjdNKM6dRaK9gWZyZ
lBIkn5uHm6rKvLczw64KwbrSVhPz588FVdWlUyhxpU82dDUQxseUED6AiU36cO0yiuf09Mt02LZ5
X9bM20Bdgv3hRdSOHvgPuF6e07IwbdYPCKp51cJHTV5GmGaSQBOQYBF2XW9Cx7xN5WgxdrnrFE3c
FjWV9Y6N5auWC38p6KmCbr02gps+Ijl7RL/gGz9HVeWq5e1a8xhAxAfuCClWe5go/JxxAszOiqqa
0m9OHql1i0TrZEoCePZWI8nVOXx/PETCXx/WFvGmndp++Hsk4zTUdg03jvQeN8XxnzbM9+1qrysX
HFJt2JIDorMj+U/ujrudbHE6ZqZIWYrKVf1bOg0Zz9/Z/4y3ZVLSRqoX3ot8tW9JzFMsVWs/vEAq
H8+W7mPEHbglf2WFq9h0YRhka6A9qvP8RDjfaBmmYwk3F/dsl3qB7mtmOwuwMxJhONM731xH+XWt
0lFCinISGjixQwSbhK3owJgg5kIB4bZPC6y75FhKlbktC8xhzmZusPKNAo2Rzo0cI/v3112+iOoS
HtVYtEOvLpn/xu66BfE3mULTtydPhPA2f/x6bPHY96+0SWbXQ9Xl9GDMny2Ea5xQq5I8UCMLB9pI
YpSca0QHK5zqUy8Ej+yc1ve7rArU6Rk7MiP9Lvwb+Ljs48pGACO23njIyzqgFSvMtfC/vKVRpyP/
r7qd8N5iJNRvF1R0hi/EHZmw0SbyP5v1PjpdJ9Tgq8wkBuBRCgAw48Xeux5EvP8Pl2tQTQhTwqMf
9gGbFkE/Bfmjf5jdHNIuJokKSGpznCCTOywc5pHX0HP8Iyr169QvvfZroSdDp0bUeb2rhR+FzSa2
nqd+Vb+hK8mAt+hk69QMVsS3XhUSVoxgZ0NfTDkQWW3bfbBLJIVnx9QKJUh/IpsRx20sWSlxyjd4
WU69GMcMg0tqVbpqxVqOkEpKtMTQKTqKWT/fQLA9XFMNm7g7PuyVQJ8iHMTMKYIea8sF2EwiAovN
I0VEsYsO+DOLYb/swQeHjTG3UllPyBdjRq/mbr/z51TTb9ynzkqEQ/XlwT04ggrwgrv3sn1XK9Zd
6rfjQc5b0kBaGY1H75I7pft/Pya5KsZe3jkXghmqDAtD4ZSg8ZKdbdNnm1SImo/dzBpcbT/pgtjo
fTL00HoXgzS7vU66Se2VMMdXNTwCd9OlbXsV3MfgxYFtJm3w8wYzjTvL4a+Xq9h+wBcOchpwK6e1
s0D+arYzWZYfHiQMpVYc6oNBLdjcZ2nxaRwL3xr2J2vA8GoEQq2Hl2YFJTJNkvda/U0Ye2xzpaBX
tFKSiI2cEvEoU6RXmRg0qE3K6ZIGTpTuJmt0uWr1A/4n/3wJYubPnZpS9Nn8FrLhVZiki6torESx
kTC3ueH/0uZ0Qhs1F2fi8e86oh0sQAEdUijGuvZXwQwiOHzWkpTJIgmL+Wj913tu4zBFCsvJeyX0
oF+sbgRDdHIPsHHlj8cw+GbzhRxiD0HTqisa3vOJHLMw4XMVS7tiaGVDnuLnjDen0/IYkklVJTTQ
JxeLvrnXcmdb03XgxOJzmj/ysvZ57Kt3MzCDPuA5D7GfsTQiybuaOS64DR6BVICgBA606gDHsc/R
Oi67fk6oDDkH7eDm9Ki+P9vOnNsGYtu0Q9Kt2dakmB5mX3hEfAH0z5md0inYI1l5buuOFcB9TGXJ
h+E2Ei95B62JV3G05wZX1mI8g0ixLaF6gOB2XWaHcMeD/7g49VHL0ezWoIfmFFnI58mmE6oCXshc
e7Q+5uQO4V0nzrpY/QCOKZO2NPvGmiGMxiIEYLOwPgZomM1frbYi9r0/Cxy4fSOBGIiWm5Jghdjp
hqOWQJ32AN6pqbyP2ta+RqKiroB33NOBGh/OSm8WuSklKSU8BYwq5qZW9u+jWoYzPKAi1Vjac87Y
Nko2Be0kItMIF1r6ReDIvCOTKcGclaPJ+PtOEFeZbnIEcw6XylpKrDBGs0HZdlcoEiqfMQsOpjCJ
s+l3pxj0W4EZ9D17ZKqHDkXkfEz30SWlFEx/XHd7kglI+fso4z2Kj9Q3C959L4QJTue6BiUrPQdM
4MCh4gvySyX7KL2YVVctV3TZKTU1di3KP0QtXt8m9bH4gPqe3MoG5KcTSjtmwMI0tqxoKvJENsnq
ZIzw5zjvdVV6z8diQz5zFQckG/bRkUKhvr+6Pi17y50qmlYt8nr6ulpNHrLp4tZDHjbAHQgsc2Xw
41r0++IkCqJwjG+YYEheOcnXSYlRJkJE32bRatBTIPn1iaMD/u9zB65n/r6sxb99kOcVkhjD95C5
pm2mUAL1L5F8AhsPwK052l2yyDRoHkUE11nIKfUHR+4UcK5UDIXbphaFmeHxzQz38vsXpdR29x7H
7JA7utlF4h1Xiap1STGoZnjJfG/5y1gCPgThxZeyGuGKQPbmqPrzN34v8iKX1SwLErFl33QAqcai
6AtIH4Lg7lxD1YRinvPbGHZdkwW96LjgXjwPK0abkc35PNNfb7AYisKfhIzEVJduT+NG2q4hAtBW
Ks4neLtYpA+9yJ0OnhgwwBKn4Km5X8DZUQQ2p4oUzfuL8I0Tri1Pil+UFjaXzyShHSY5Cy5tjquq
L2sayUZ/ykigabTTE+7wH8IvKiIEqMrcIEx/L+q7VorZsid1MEYjlpWm8moJZSyWIXDZT3VgBy/p
ZbZ3ckqr19eoODaU9s/qLuzKS1kd7Mo1SFQnu2DNvTbpHP9OaOZkgpAjEE9vLGS01hMsd11ie/4m
bbmK5CVjQ+XupKvQvNP23OYvKnCxsqxZRe3mIhWVdXC5MNnHneorbEJumtIn4KK/Zs9x785mL8ZJ
Iu/6K2BhexKvtgVYy5malETjgMYRb5a3RUyYWEzj/21ouRoxaZhqBM2Wve+UkO1k6ajbvHBqs0Sc
Avhq041QSVqNmEYzbfPmeJMw363/qssaWFTpsprwlcuobCZwjWfOhHwA6+xZU65AyDqbb+7Lh3Km
Fq52YmdGlGS6BVOuk2ioVOV7Op1eo3HjiP6iKo1F6K3eVFpJ+hZ2w8Fr9C3XWWVVqZhW/f6z+aHV
oO2uGHV4uEDkfoq4yBpShCg5uiqSVX0G+hP2BzIeZ06YhpSoqUN3U/81dPYkuMEuS5etzqgK6HGL
xvr4jz2jaPUqO8S4fYZrO33Gf3Nm2HAiHY0sxmV2oNgwOj/+7R8erdyBIydo+1xmdRk3mjEWicTt
xbeCth/sF5yFMzv7dQEb5d9RynOZskzFiXRnettkC2GxENDcF5ii+mNkxQIYuYH/9Kq+N7t1mUHM
TRqPRx92UXrmm4V95YgBdMqtDRL4GOLNCQNjZCfqiAScgSbHTpy1HgiaJExQFm4DZvs8Um1X8sDN
XchEhPsicTwkvYrKxWtjYde0J+05a6lfT5kk6JnMYQKw0NE4dvCqrFF/aS6FW9EvxGOLCsUPsVUf
iiMekqlsk+ewnqvaTpxHhArCEk1XsDQAZOTdlBxtjrVdMdveKg0yW6rMFUQtTS7otyI5DFWqEODR
ziYLpldLSKyw9S7PkXA5286c9ClVJ0GRMbjJXnV0jAj+Tv2/5yB739BUHQjyOmZ6pMR9so96AmRk
xSMftjpdH0vNk/zrtXB3SRxz/ECeGaK5IUV67mIbLhJUu8tJs+KgSGR1selSvSapsi+V7I/MZfhV
vPjMHhnIBRJYAXhnU3qFYeQnhLcCtYm11Q3UPxl7dsc1DQ5FBl7tvOHmrBkDDqtfK3gUMoJVH+aW
fjSwNIXsxoLm4lmZjQMlvesO1AImCbEvPQpmQRh6MzgK752n3TQYOldN91fIko94tPR64ktAbDSd
JmZ/QUTchwMGeAvtqdv4eEcPOyDaKRDd4Viy3NzrfdV6/Z6b7nm7oPhiHvFJnSx7Hz27RwGjEPm6
yydIJG7tU5Vs+jfYfviUEVBYhCjHxNpg3eVKBLyAXhnaghC0NjXER6UCZ5Gf43/CkeT68dUgUNnk
BfOID6KUIfnJERzSu6v0QHZy8sYRjVaVFbFiJjCObOEFy5UpYpBZuNDo2M7mmj/YD42ncn7XTXjH
Nqw4axcxeTE/E/kNTZczcKBK44pA0SzDscU6WP6XsuLax72kU5fDrLRBXtWe8dMYeZ1CGajtF4Gr
rtHuC9YvI1KA286RyViyUKjn+Wmw4SSXjnn7/th8peDXAVUobZwql3bTQ9739+DwUrRAWykTaUBN
S+T5Ol3q938R6+Ow7qEwrZsSPtFOS6aD4wEeD9KvG/mwqVhGJd90qNBs2KFBO3iZ8Tj8nWNDugrY
ynIULE4wFFblImUurVjd8czsClrPG5K6Cnf/zJh03rcf1SNK2GE4FVNJz+ZIHo8IwYiGMUG6UV3T
DlXTLpFNyUQ4ezzVv8cI2PaGJ0LfHza1IQji9102nK8/1nxPwUEOGJHsShzz5pgfD/7GYIjCSEuP
FkxaRgZNKYwqt7VNqSu4jgUIEHfztZjeIXWJx/8SYrmko6OmGTqEyIMhnlr7ttyN0GjFCwg3UajS
yTjeaWGAWzXGjPekiZYgV+1hpSLF9gk1Qa/k2oItgV9N2lD5WKFyUOXs40azNuMz0FVZs+LdeblK
El41ScHUA9W3T2sECUv18aZ9JgiEIZIM8ipRw5wR7qYkv7at12PYIOaSYyUxXx1wFM1E+VTNrb+t
3eVrfKcoua8b+CYnDcNRBLsi0qs7ixiPabKGKQATaK+oDZMeTfHa1FHremB5NDYhwEx0rTTA2onD
knt+NCP+6vzjQ6blOmfdFjNiTh0T+3j+7I1pV8mZ3N7QWe7EeNWvKTvMQ4+rP077yITPyLEUaK48
KKTVQhOCpN6sHgGCsyszySPIn9S+WnFVv+S3aY4DoMUjwytZlz5bvU+nfLG8HtWYd7XwKVm5RWxw
/1bKgmgRyTX4u1qNSmlYuo7w5/gLL5szv2/2YjXapMGHVUKXeNw3oB7nBh8MokSP9mqIac00UHsd
lau6k0IXaGjPzs4xrj9n78GnrW2BIvLlcTjvuy3sIdqKVik66nWB8Sha2fVQ5XhY6qG4RI1FXJlo
IexW5G9NJ0v2eLgyniaw5Ovga04/HVIEp3rMDHty8Vs5c+kt4rX2kR6XfucHyfCYf2MRZ1+BwKfK
ZSytS/fqbr9hPXj8ScV6gv2sy+BapcuuQ+8P6Qe763YXBk5x+4fYj/Bv16pNxPrtiM7Netkkkqpq
ioQGkSisaJz3AuD6BK3y04aXZySH1XFsSCqDFrmZrWjLhTwODAI9+5iIsV40ZxTK3mlQvWVpu4K2
EjN0nxsb313sWtygq9Hxf7xP8yzf+/MupGxfFI8htR5MWtiEMdro8G2+rgebZKEDltXvFbqN7UiV
4WVfyr1F6KyhdXHU3+m/D2+1/gmfRwt/mtZp42/Um6G+s3YHBsWpunHMGNm1t8YCmVPkZczG6T4A
/SPiggVnob098iZQ13nHBnmIgRQLIwyXM5Tjtrdtq3Eqdye7opE/EJQQFWuD99N7JLS+qegyJC8Q
2BKFYWBD+9fjbYTdbfVYTBK+kT1LLY87bpdIDyqGtVk9izNLpJEpNAaitPLuSEbKVG29/rtRWzoo
2okE4OefZ9gKwz8Kxb5i+7q+Cy+Lb0nrugRqEJerrYsJ2EvWKB0IRP8FH94TJJucmIRnEg/h3EV7
jCmFYbhkKBEcKkKwbrj5HxjXkJraLI+xbtTt2eMre0ORyMOuVKqdhQ/RQq7y3x03IfXKSOJg0D9u
y2xDdyxN54B7KvUdCKBvphgJnwe9i6E7b3ciliGaAF9+G6OWT3JPzIfJKLf0x8CMUAo9IiFfgnEx
3usMl6rAxkhA/hCk8MziojW1Fi9/CIzu7TOkqOexs4Wg/L3E7E+TjqAN5nKeXdi9O8B6qpcDLbJQ
68SGf67QKuDG74sDOoLXcXiY/UaHjnDxhrC9ceJXt06MKKLsqmFQXeIRTNxp+kFkFSOqnh6dUa1i
ZldfLED6yC25sA/6j6Z5UixdldCYlDTsp+QQSMe+zGFb5CoAXVwRNubNfwbrtwLHL27j+Yj+oaN0
y7MGWaXvZc2fNNhqM7M0RiWr017rYBbJIjgZPugonwO/kPk1dk8T8sMvWTAONESehzTJ2l2iLVCK
7i+1t9QG+h62/kNfu4mqXnYzftY33X+ENE4MH72T8/bfHCiQbKbOEf+dpSEc9zoWRMP9koMFazHw
TcMS0m1Aol08in4w3uhBAWmpmLe69+j+Qt2W5lexjqWnuH8rytUdU93LjPHHZB9W4OZHgMvc9pBs
HAatIlU4VwmMRgE8NBB20FIL0BW4uJQpkudkQG9vUhaBF4ItWXNj8e5dKgxmemhF7gxWOe6Gl1xK
82/VJyAVvyx8+ESQJsw/eA3K72NctW/Ow4s/FSGTsKemuYP0RC1wZInJh+FrxWPxGD1XPtA2BIi4
0dh6k2CcEaYyx7lWkkNGfZ3ad4tUpgZDlkmk55pyQWa0yEbnEShzAuzjDHw7abrzd/W4BpfzFlrd
3D9+gTbkE+iomjgmqXpxDNthRcA2TIV3VZ6qEaFtI9A+D23IaF4hFVXp6KklSaKFovdqPqDz403l
/dtDc3Ua0bnvkW4ilQTUhNaqoyhhEAuCdyMGZNUVcrPa+LCyyIhcd1LShCsPPfLeLL5fQzI4ihz6
l2MRZ9cmiX10g1gqwjBCRMlvoqcT1IyzhyRmBDQRpqv44QxvLDNHLDBG0RAkGZ360H9RA7mo+G/y
QOk4rZr67o3NYopyDOYqY68ScTsQw7+VOhgVMQlR1vAzxNQs/runeUsqsfAG2yf+qZwZd+92F9Wb
u4yiZrBXkbrROFqPxji3FhBrEC9APfNH9i43Ssw6MzyKBi+rpA/Ws77Hm3UjEpQ2yTriBhSrt33o
ajbn9n242aub+F6m7DO+ZRuMu6ReDR1xKs0dorD7ivknn4tHU8a2Y1L9VorkIxfyzOw/B1WtC6vK
y953T7AIWv1cGnnrsL3B9B9euYANJ4csO8zXIZ4zhwp/0NLCoz5YjeXve2Dyg0s8mxg6HGqOt0Kr
5mlsdVIjyntVe7Q7pOIlA+h37FPe2Qj1aXmzPYMm61EHnehvIIkmDJB9tRJ/zkZunWyms8M2CpnL
CsUTEHq0rA2dIbbzolVcq2lu50yeZx6gG1GdcJVKU+J83q8eagOyd5ETCJWZ+VQpxPTPXdsm2xLk
AAzUaZfw5hRwYVnT6LqZ3rfTyG6xd9Pk53GSklBtO+THTT5VoWg3aikkEgNHK49mJZW4ZZnP5MKJ
5PHlYr6Jn/h+S4GHAqSGnmTZtkVnXUimv1HEZqZvmq7wctY9nUiuynl+s0H2zMcPrRmPApYrdPjA
ZtnLIZdzxty0P0pDShT22Eks4NT3jgrELfVlRU6YfL8q42aVI/Q7RyowCqn/A7t/d8HB6fXtCrtz
8vZLKOeEBHq2TkH1RgtWWX0h/Evkn1EQvOH1tBhIlw4vtAxe3TCfGi3MXxyNhR8KrM6tskV70F3l
Z4ynimGU4YmiYZBjlZmPIvBghKVyClPS/mX2giukoXQb3WWJvrvjn72/h2yfLGiAO0AJ8OSfk1NL
QQ2L0vfoXbft2Sh/MkhZakTXa5buDFUe4m37nP+xMP/11i3wfhObZH1kvnZ/pKRi971gFwAmJzXL
0DRHFGNxlIlO2zz6KhAgKcJ3HxmnSFimgRxZ5DHhONN5pqr98eCar8AfG9pT7RjUxRPqbCDXAi6m
MyNAkDQj2+/KE71q3yV16A/zmNkb4fs6aIBIUU54Sg/USAUplhn9kBKlhO1pHaQ/3ACQAqhFb7dp
9X3helgsfMN0GFMetUYI47DflrUgO6il52MVK9Ed7afTzfqJlge68V46xQn5YXt3QCurwsv3YoNk
zgFT+N7MHaSqhvHFL87s16h7zNLwa4wa+ib4Zr6yE9F7udhlgX4boTydFj3a3WxPPThSmWY3KjgB
3UhoNcFyu2uYH56f9eqe0PlyjAvyIJeaB10LzgHFWYib61LpHxw9mQeRgSZ37+pnvmuo8akUpRrl
cQLbs1A12l6a2R3ft6fFYMpiQ6Elyq9/dp9pS3Z2e+pBCjgsXQ7XjdF2mIX6EpgiXKK0koZ6mzvm
crNwa/iNIXYdx4mNgfQF4MS/9cEWs2DmJZ0+Nmq7jsBKfIroBn08iClPl6JIRvm9g27llmPrD5H1
7Uzf4FHp5JE+ElfXQiZBH+LJBW2aZMNfQEYs7sztcVIA7ki4OwaRHw+HbitnqueuuWM2WWnz/X1s
0IvVJt5/mlajnV8KxtTQnmPClZ5KRyJ49sVUqw99KW6scTafCIv2yXrrzAkeWjo0bkNRdCREn/jU
+SVWWWf0G3+8QkV3yBd62X+fG3swL+0Nl9y0qssjDcFkxXU49NdFAR+f4hxhDDmWyEGFBZbxfty+
+CvWHzby526L1Maggr8Pe8eAbA/w+TrXorx4CYhKc7v232qhJSh+T40bpQh+RhatVjM9SB6Xf8R8
vy4PZ/dKo5VVc7oYAzVwyBJkNSloa9wkKhsvWju6HdWRs6yoC5JcSJ6papScNEYdEl3iVObYs5Db
TKtwtBMhFn7nmD78pb348LfEuiXUWgfIGTcasTJC2F0aQPG6ElRMknHKsOuAJ3V02gaZPp4PVdDf
K5tXI75iNbpG3X93d/+CP4TnyfeVoi1z1W9fbTQhYqWkhmkArVLmE1/yuHHZOQqhmAPu7et13oMx
5+l5zz5BMCpIICf+dGe0W4Q58S6cKN+9YgAdWFe0E/IEplhKByoe0lodllppTRnqZ3aba5SxAYHx
mbhfXHaOyIMLOplFpr9tV835oPriaWXv7xAQQg6csw+f/yCHLGDjOoZvJo+CA0NXXQ4Cj0hEYHMy
GNqBGQVtfjAlfVC6JUZbh4XaRJJt6H54sVaHiRNlih3GflS2ZIcfPG/nhkirVyK8DK5Fe9fNcjek
sBNiLE7Q+MCuuijSgafz2hBiEaU7qvs5mH3K2zIQYzbX3VC+8y/ZPPaopiDwAO51cJwlSJcIH7+N
gX+OM0Eb4gOfWnGgsRxMnYO2Km7RkpSfxh6QK+qANHsQqzHZywfPPdlyUNJVm9IP3p395IxjxJKK
Ooyk5yxk8b838qw3WwSOvUfwD0Y7hEFcZ2Ar+FgLgk4DnfBKWmYaKlSBoTKQHUnbwSc2RzQl/jHt
AgIDxJF7e7EeJgRB4J+A6lNRbB7pqAkwR2nYzPl2Nk6E7oIgmSqlOb4ATGzTLrApcJXRPP9c/Bbg
qItNLshvEyTOds8M6OsurKkzNPhmPKiCJwD41c6YIRTAzwiwWCuJHnty4p9pQ56kCXz4PNpE5IYF
zaQ8fOepQCLijgW8rXUkD+NEZ+sZGOvB3VabzEejsJFC3VrwKRB7BtuixWzbHNI+cS0PsOEvduv1
iHBjADoomjGj0ZOmiIDuf+oXNfYK23mRKr9szD0PAIRFe7obkXV8argUd3m0oJ6leA2u/qHz2jyR
LhZVluH8g0SpTX3DDYkdheCdEdtUj5enpIzUQDV1My8lC7s+6ApXQ2RzGpRoNbq4RGPi7KAo0y8T
uRqshnrEjRBk7u1Ylz9oVbq8QCwwE4pW6g2aJ0PCHlASOZkIorxrs9PkqaJVeu2PSom8Llnztqpw
zMHIelmh3QhvplnSXRCZcohA7pCmv9AgOiRWgZoGT/fuLAAU8081x8RKXx8Rwo+fC+AtmVcjF+V8
dH2VND8XxaOYmW5T4FArmmBYAgAGE648oIMfhdaEXFxXzc0qaaXylD6+bOn3zy+bxAzuZQejm1Mj
qkejWdxybqdaGtMWp8R3C2mgCTdq+yZQXV6M1vkgmg+UWsZ5cHpAqxH5weMf6lHBUwBA1hffOGGa
antWCL6gziMfCRTu8owoKlHAU2fUc9Np7Hcd+XPy4NuWB06ZU9VrjfWWKcyMhUxE6tUucQr9EevE
B83FPy5BxTN2GYt9IZIM5mN8XzNgRw+z848SU6/+tYoO3Edf4Wz8ZUPSyu/mBG6f61BT93AB1voX
KuXKBg3b8UG288Z51w3Y6Hg6X1bWV0NedS2R8OC9weHaWDE3UksViYiz38cbRgHeqljqzAKra2jJ
ByEa+9YQ69oc1b83+EnvwTQ6CvCwmiQM/fc08ye5Imcsg7qdP+7d5oe50NaCaFCfP/OdlBmvajow
vkAhHptbHkuBvGxTPQOjJZ0BdRQfNWyev5IS/erxp4V9S1ZacvrKR65mIXSD6Ptptvm83PGVOmrs
2mHfMqYaBoQ+qkNnS0p9UeoslT22Ly9yIJd7zOgWbw6dODAFZ03Qz4qW7mPcGq5qODQXE0c0gDei
CZzhj8iz+y4f8Da5dUCQ3xDL82Larery/JmbjkpbcOjRkjsL9E003+Y9dlas/fwNrTGL2qj65RE2
NtOjzRSGDxgnV3jiqwW15wTtHL4TiZsTDYQ/DHVUCy8viRyqB1x1woJGAunnbqRaT7Vt4TTDrp6W
JEUXZEoJMSQiE+FMOS72w6tkwILAZmIm/aft7RSvRKZLd2EyUMrRUoKWi/znUPRTDFYix9ZE3UTc
apkchDS24yWURy6eOo5mFadgAs+nlSwflR2mpGu53bcLJ2Xkj1sNApscrGi5AcVXxy7e7mAGwY8a
j/qUF8L4jtBLZhwyHHa0emCX7KOxgwATkFW/Pt0eQCl1iZigW/TrOjq5LKtwTkmvazXYK5/Gauh2
aEhtcEmcn/rUxz1otF6grd/Q6a8iXYbOY1OLBxwWs0sXduGdysUjUX9B0sMyynfnK8nrwavuqyr6
rQ2hFiMHujtLISDXUY0OO8NC4toerGNN5JRivaG74APjFQ8ydvwe72F0UdHXlJxzGq8qm2Cm94nr
TXTqaMrJ3hJ349Vsys9W4lzjZNyMN5EQJkfOSEfSH+BA3AAtYca6NjkoKRjUY0bnSu//Uamp001q
e3fMIXYe+Web6Co8hSpf4gvYYIkz7ZMS4yJXffYiAlRRJqlnbtkjTIe3flltnv+5VkGEw3CPyPiD
r1MiEXEd7hpsRVzFY0jYCDpTfjslYm8G3akgKYslTE5v2YLTcECuBFdJixzRuOzl5XpEMbjYjIZv
2qeP3wbDuU8wgos7hasCPRFzlbhxs9wZe0QhfUsPOyFsCGzzQN82+sY7SOiqqH1450slHvKFTAeA
snvy4Vid+Ytz3LvPmgRhK6m5WN98kxzlikwTp2uq/MCm93TSvPhYH5BVabrKeDf6li/TcKygYeuA
UnDAkQ8PmE0OIv9yLv2pgIYYZ3m/3Nxtj6xPkfE4iC9CIxWXVDqPUxkSLWQj+x4yhPNO1wSINZXn
3PVblTg+9MVAL7UY/QpB1gfvczvzKiScIYBiAqno6LnZ1piGHmzEnswHXcECCsmzMF3Mx69pCKrm
f9Uv3qig2Jdz84qQeJ2/CicECybvtUqUWpPY+Ye9hRNt8bV8xOwdX0KNruGuWG2AOR7NHTYRRxDw
3iweDtEFZy3yMCKKRQKGLWB6hGkZ+L6WalWJRlibRuiDiDFLVkysmpN7FrgYJ78wV0/NQPZqXWTJ
XIskq2VMhVYWcYpP4fZRf9fJkVYNV4mn0qqdci12fr6xxAjC77xBw7s5yQBwtf+HYN6hXPCg8Ytl
bps9pFgr7MASPuuGGD0kDFgEUeR6b2BAnhlR4KaQfBhG1Bs5jKm9G6iYk6MBU9nZOiSgy2ni/IwH
gqJRnK4YdzmMrAuJUdfBKiAonhDTbqw93C0o5wMNrQdYTwqRzxaIJl0jtOZJsL8MLod+zkumTb/M
hCJ1k/mLPgkyybFVJz1P6eZ40jQnb9t/CkKbqMDBjxldZwbrY++LFw6rr/RfGlG0pED/vTrRWZPb
limM1Fba02/6qUBc91lHWXREJuBHfeGQ661szL+tDl+U3bmKoZQYoOTAx8zjxMqlyF1wAaQnSvV6
MCch1c7HQHBtRs5pKHMJgzwWTF0oFpfFww8qSP7qxjZdU0RRqd4WlIzF35Fa13/IsumbjPHoD8Tq
s6Ro/koynjashzu9uDcRjKlSMqoeRkrfGsEh5T28QjOWxClJzocNkHgHY6g3FJ8nQxNqeTQoZM7r
94kbIqCd2K+Fm3ltfx6e9IWcngixR0EngiHfwp7LNXNXYaQPYm7RcZgETk1EcXbaExgyyl3yE/MC
TuvxLTpx2NGvc1Nu+w6EsQs/y1WzWr2Z3/7XmtghkX9ZAYzuttEUjyrbgiSqJA608kNzAm/W1Acw
94cC4kGI9uuVgN8L8qBSUSBjvBWW1HlQ+JhjI4qQhsquBJCgwGBewEyuxsd9XikRiEauKBQYrl7G
81bjzFmOPLX3T0iatbYs39tpTAASQsC9R3GMr6354/N/TN9E/FWvNzdIJBJ/dRrrbEDUOeuYA2IY
o4oOsxa62dbkkco0++XAlCkL74/zdg8lVlCyHxVjxGvZ/qi3TIgz/+M4xOfbHfnUKOq92sgLPdQj
8yNUejVei2D3CF889iV9DTwqFDtojRz0yfYYCQk8/qVa9690zo9nH1OAWoANB21eh4yypPvjf/lS
FGfRvLvSns3BSiHMfzi0PIZm/5KH2VMow411grFpdlTq6XU9UMzCD7c7KSFJgqhcIYx8oQycE4Ed
74OCI2RatUUP+gvR4RkJYtqAudedG1qDDL4RwMJgo8FEXHKBJXc3yXj/h46J4omu9ArEaQd1QfFa
Z80+RqFVLfOUjQeqXkaddauzUanZhdtA/s1RNsFngTLddUVKcH+O1byfB4Z0fLI9zf6tX+TN8Hof
U1A89VLrPFyC7+3fSdcqR8dWU4XfvFGkgIcU0h5VWqlrQdAl4dqxPT2IFlJC7uhLbIbuhQY1ObA+
kEjdcczDTSi9LiY4UK1w0CSdddXLSMvZ0vDZWnCFgg3dLvIoCUhHtqFWeq3hCfttp/bNRJhI3J/2
pMJfT+6rHrruH8HGRdx+SjAOR9ANt1Nhw7W6+7hr9PegFXE+9ai2AKaaRqilcjqVzXOdNlVTq6Fs
+b7ArF6CCfV/M39G0/Y4i3+s6LyH/h2vQHS2jahDyC1mVkYTR3taXnDtgENWAZmFsVDvbzpV4bgC
FW0xaLyhyk69ERgnGYmU+2UEhaALvFPu07GNr9TjSCT4gYMV/QCGKjCbECyWKPq345KYYSdkPYAW
ucHHSkUa/xAfRL4O52talDxcMn1I3fM6YLRhSxZt2CC2yr0aLvvNLne1AUoiVtuXwPRCOPkY2ccB
pQ+MMvwJM/2Gd+KumrjTzrT1t3KMLe6H4sDsyXIiHiu5223KsTXN0etb1n0QoNznE/uiY9jpJwro
KwIXX5aGsta1Gc4OsgkkM51DwhnvCSoQWrHrDNL1IG/UojA688DKjNlItf43JKKwyUyDG5noeoLV
fkgnHDT1EuEYyqFBks/+jQF7MDh83jSDWIthf1EyurbMRXxPZSOwHShlOIwQ2aI9Pj9YRRgdYBh6
by/wuKeUUWB9pBe/JDbVh4PS7tugOnCfEypBkD9C9nysAeJMhhXvXN+IDjQ8snkSh1F8GkUyWvIk
fAEBiVCxK5ZUnt+NGfa3SWZS56ERUXPAO3/5L1jW9jBudrkus6DsNxL88PXRQWufrOf5liNFuSZl
H5e4emH0DOeI9n/wPU9anUlVdXfnPAoy1ZWc2n+l0qjn3m9D7nr1ck9bSWsVoKBJAOL4UArMBjYo
0cMvWP6ogiAQnq5tXryw54+7ZSbKiUvJ5k34dVcp7+l6510kcfJfrSnvXCbqWkUEavaU6ac1lw7i
B3vQh9G92zXKNx+9IO2/3aqOPICpbH1Un84BCXWyXi2V/ALi5IN+MhPCWd0h/ec15kWiDAfEaWFs
Lh0tZgwlawa7Id6+nV78/X8t8XdyILH/EfwfhxpEmtdiZFKdqs0s2GsSiaHb3Cef5KPKzZOMNqa6
xI5M3HS42jx8FOd1mvKQCiD5OdrxptTT/usmYob0mfqo2mTWHpNTWczQoYsfuvDLjlcGPn8ixWHh
DXw+VaDDkEuPruFFJQohXSeqyJ+yTA+72+tQbaS97wDJMtxmXkRtFRF5yPErAXcMjaYaQZBfon1r
1nh5nAkS4vddbkFDGpSUs/vj2FOnCI4K/Ys54InxMSZ8gUWtTP5J5pcanR9XLQXRTA4KDpN5X3BJ
9QG1ArSB73hj3XR2Oi+GK1HMyVVvDLNBcnaxAO2wyGEr2VLB/QoBiaznlqZjef3/bIBlSmr1GTQk
Iihd8HqBm1mkg0inwI66ikLxDKpTmY/dqJ9RP5gasqUL2K0e0p6H4BkZyjPs6oLRjYJjNkrX9TSP
TAkFvXmTF0jexnMLb2Jk0/egAJ8B0BSbWNSozKIJKFzDyhmXmaXx35wAQ6qZ3fr7YhBf047cskWV
2HujTaReU1xzlidzP+zx2MqMRhnFfO13HyFVRV0dVi+4UAyu0IkC6QX0NU6cvoQ4GrugbCFq5AER
wZDHpJ5fFJbC+24riHXvHbflaHNvTmMpzxr+VwUtqa37qzxAFS54OWggccpwg38Jrq799ZlTdBlL
pCLNSb/oJnGhWXEIAiTdL90ugfSgMJJryh3Hn7EBh4haXm4QQgdcVvIfZ1rWz9RzvSUA8bM7rYVs
RlerNtANEzhJ5gkJz/+6BO0actmXcad79Ki+QQlzcvAMT1rxPnzRS5GeOY2O0+Lt8/7DDadMs3XF
S9vc2G8vKHVfKyZOKYYJNPX7/XT04RzUqIT95Ry90PEHjdxcXvdCAaLBfpLrjyhzovjAh/b2ot0w
6Beam0GPNWTKLmqf1F9/XSRqGOVYEbvTwpiEmGGPBrCFG2GP/Y5maP2Ytjv7hX+VcOpBpV2BiN3+
70wKyEXVj0KhvdeB/OCVANyxO7MHAoLWU57gH+SsIElSk1d7X82+CmIFZ8WjZDq70Yk1BSyVLju8
ZeL7EQXOHwrHYBVGpPFIMTRQzsiLSQ5AdfnOsxN1tbpMMzPgWNm90elrHDCPOh18w8pGPncXqXR7
ZW+EZEG0Zd8d3CtsJ8k4sbeiUIRww6TrjHKKSvVQziq7dO/dFPfsI5M51Ei4YOKeuOwDWzwmKPUg
ZlZQCFodwvL0+DfdAFz3GyAgVXfhFgusYtt62hRwI3+BZu7y9UNSkU6U3Z6c2czg3otKUUkORWn5
9wccSGmVXmib+SDeNyn6w254HEz0ZAsYTlZ2e/etD8eLjQDfSn4wbO0ZsrPWMeCklcjPAZvVtb1m
jT1qaw0uT2K0Ubh/BCIbtyunPE1QoIrFHA8HYmFHRQ3aiEIUIybN2fcj66ZuySJVKdVDJiTbidNO
CAWP8fwYfLuwlTiFAZWRJ19t8bHPnExKHc1QhVPUQscPKmM30Tx9uPKixGcp7Z2toSjJNfA9snJs
TpuGHYI0vsVmLxYid3ZCcHJIx+Ht3ZAJXNzWMnYxlX3yYZ7hNGHMocwP22flxMRfjfHX28XchaFp
WdTLV5bbaVFkDYiGOLkQCTRMTiz4iMoXg9iBvwkGOWqbni6uYtBJdN2zyNK/gskChTnyr5WkSF3H
J0iN6iGYSQasL5fCkhrCC/XsHzDUKJ+B7yw+/3mMCpkauSSuVp0qB99Db8Qd2OHuL7WaH94+JuF3
4XnO2Ogqjbbg/JsrqL6U9ziYrmL3aCwo82NnvSimAcnqRnRT7kb/aULepmk+aoBdfSANpAm0s+52
iEmKuKZosVF7g+1NoqMaqzvazEkyQNJEYLYjakxs8e0Yz7GCmgLIPtjsMw93QJ+gjLijZAw4+AKV
/By9FOFoxfkSlO4WRliLPKXnaFluHr5Ofg8HwviSK8/4VWnrIM8skGQm79AJNJDVhkGoXgw4qiA2
7rg0sSn6jerIOIYod2RS408UtdjY8LtqTXm15tqAZL4Blhpl4r9XnNBrXBoZUXCxZUfUhOfEC9st
t+VHLWndz8eH/o9xx6+04MFLFmxZ8y7BXHEcJPifEBaM3L4/nopRKc8oTCj+oCLeLhFT3E4P1NKl
d7yqjqEzYuiMFb+P9xr5QOc1nsVrL83QYXoSIdoqMUTa+s9bx0FfR9fN23UdWTycHVjOZxdtQ1Ph
d+vajLsyiVjI/RiOwHnGV4vWOrORtSpw7qzVkJqtG6j3p1Ma6iQbYNzAY/dY1PbaAF+kxxzcU0vv
qIjItBS2OqG9gOlb08c67BwXq5B9YBl70aI4AJFLfZk1J6wI4eEm864Y2xj7wSnBxiOVOSZUed3B
go4vHQXI4wxo+BtIlHaUtYJdTJ2f4Dv9gn0EE+Hu/JYtb/S2BYabslVsZz353k4o/4Yh8QInspVs
XhxoVoGFjfmv2aCAAn5GG3S06tYUPmQGYNd6RJWcl9z4iA+2VI4D04YEp6l5bo1AMd7sxCfNKQ6c
aXH1Kk/DNuqkq1GcPaOSAoaJp8Bx4Uqyp/rFRGb5yThNh29Jfz2LcUOZUMzaOnc0fc60Y6BRYwrE
Q8BfPVyKjjU0qlIz+CX5cC8Ph+vG1rp+kxj6nj+Xb+feJw3jmPjvfiQVUmeqhrTKSmrQq1cNAvmH
teXcKPOZDGKOUv/4oKZ4eUoZPRFwMEk8GauF+hdOQ1LZ3VMTKBPeEIO46om6EdfQXtu1l6ydqqcd
cIZX2knHyjdSeRd7jtT8p8wNRuToNuF0MC8xd9sb1titrfgw0wVmab3rhZWqvxyLmBzYYImx45Ux
putua5jL/ypgQWsGo0OAzN1YQvXfm4r1LnHs33bZfT8E5NhwNydPiInfI8cQfaVaUhkmyFyl133T
f+05QQLwX1i2NA3e8bbb7W5n1Jc21yPrtfVVpqNidnyz5zd7K1/y9mbSrMC5b2R0sPjmvVC3ryVT
0t0LlXr1gRwJ3RrE5RnmQi9itdrT/ZqDKHm2mLmBPrRUzw7CIxSj53qJAcUMu9o2F++CApvlK04J
//J2tUDX28xCY6brUWLxbbgTq22kd8I2+/EcIpFWlSDoTPOtpy7E8mkFX/yXM6vGwpSSN6tBZqUQ
qig4ZlIXCmTno94DN+bXCaWFUHfEHNg8S8bALjdSAWV7zHK7xJQUCqoc2Vs6A0xI5K+SlQB2thuC
J3NBFlcleHCY2jLkFnhpeeG45LnFbJButD2/7Lu2hHTEYVxXZPkNn++pxhow6X1LzmyA0Cy3Q+6R
WRS7Gv3Vbj9b2N7JSDoWHFlbnAQXJvZAEUOn+udkt+i64zCHdxItdaTIHAokQiqMDjny3lbtCwer
0z1k5WiqgVEuywDOiC4mPQ0Q+udQyBnZ/dEQd6onUjWLf+Cx7d5k2xjqUfg2ivMid4ST8rtG1MRo
ewFOxB4WIacNgG+3J8pbbUygO1Rqtsu8EJK7Xc9rFo7kue+fdTL5Ed5HzJSnoNItNZ2VTYAnT2ir
BW+4Bd3Q8xQ3hzgnUcZ8SjnCQbJ8zI8xx0FZ7yoNZHsOHrki9jsoyXUU1SfOg2AIulUdao4sUWlC
g6SDqpsAKAq/ScRvuzt1JGHIp8oCNq+7K6bxhc2KtE47BRWQAKZmcon4xubylZIS7ZopH/omm/ux
BhhKFi+UVi0oP+vGi0xJJhHZjqvgM36Tnyj8j/nIZJMLdIcQS2RYlq+bVhnYbrl3PZC3G6yyxg4g
OeK6KTc5n7HjmuJMpLVFgl3zyo3KNm0ErXwD7KEWtu9qa7wOLtYX2nKwXaqtUjoO4v0fr3cMnf3e
2ZDZAxcyzTfpszDvQ5Xxanbke+J4CeeZFTolK/A1qgthTe4c3xcNROSFJ1JuhYalSNgM5zgwycYC
o2PC1yxmjTRKSNkcwCx/XHkWHQ9D8R+zq4z02OQjkH7tG07ycCLN6eZQOtR3dMPauoiOfLP3bLiz
K2atCiuOiNpjzQ1tKq3tPelaeYRt0xrMqI0eJFTpOpvUg3NP78ESvQJuD1ljdoRKdBym8Mlm8B44
c7IooEkw8GgHeDI5n+gx4issFfjKtqNZmnVc2m21vz5cvuYf+8t7MpYgMcE1Q0g8PggdTf0/Lc8h
avSCcuqaA6aKq5+PKSPdOdYT9+9MwXRwELqROQ45aaA+u3DaXccw0Hjz4rKfu9/wR8ZKDfYXxz2C
UWCCUltS1rKMWs+6QwDWxKi2MV0pCeCnZvyqBsf0T7dw7mY8rg4bsqnqhKtivhs8hSHGRo+0e4bs
c64VB51bEUta44w77hmceIImssrsS4yIzLOtmuFmSEc6liHJj+9LQKQCmSakvnfEhHir9tb7bZhz
WW+BdaK9tVjErfxUCzMKZYTnRCHyFLqDrexOuZFd9i9Yu+tUOsCCV/omBvQyZv8YHkFDyOt6r2cG
Ql+5d64uOD85FXKfMM08N4WTOEvAEzKx9FBJlg5cQS3VlrBHmil7Or1QuCtjvEwCp9nECmPMEd+m
SLXXXQ0hOcwfQTu7tBFBxy2TaWxAXYiQbnFX1sVr6VbCKZv1E+O75TfSG0wB/EyJ+qWv4dM6MYgJ
5fWcc1mYsIZF530qWcXl7UGUKQ8QYYmc9I7CbG9HN140x21r1iBMibm8hZMkU6dn6oVazAuOGArF
PxpRkIS6Xg+fhZuNvoyzWybWNeXfndG8rFWvzqRzbwEvbtbO3Klnof1/I4ZHiz90tlzqIUChoZtX
FnFm9vAz6cgcvsuxT5n7vCilFawm6zstcGK1tJa8JL92pMJLMwUp2IWEczDkg5qkeaM5iQSo5UAC
zvjisbQIdfVhwOHoYWwlDomzynGXqWaF/9J/AvFPODlmHX2hXi43slCe/IsTK648iRDL024v4GKD
og85EaRPjdPC5bQGXb5FHiPGpZiiIZkgYEhByLPljnDbRH2xmZZ8LGmqH3hSc/xNtweCVYuT+3mY
KTzeZjfGx9bi//roU9tKgn7kdzfh4bI8IbfY/D8myNApdI+hmJk6boO6ycKGStLPUY9fNy6lIJlK
w0ICEc4I0b1HIFLHuh4fIgtSjMuSMVgwZb0Y0plA4RVd21M2giiSqXThrtgDFPQ0aRN3wt20laFb
TTamNOqarA/P7ezOtZ3xcpK+GB6KBoR2MAeOvUTurkrwA9QQDK6htxlp+As1oHJQq1VlaBFnkbDi
Bed27qdMGx+KPd5cYc555qxKW8EmHRqOrc/rjP8q77YICcVMSW+vVtj6gK2ZMA6EKF4BYoZChenY
mjSaM51eXKC09/5JgoKU3ktgQ5U9CeBEkXtsjlZdn+Sn0unpMo8KH/pWcCfuY+oQJ+Qib/ofq7NY
VBNArHy2hYDKb2cwrbbLttAEMj5g6OmqKF9hXjPkY8HizeCgdLalWik3UW8ypCh3AnQjF5RX5sEq
ydCKj3UZD2j11kAhOfEzH9+EgNN5RXYGZFSLtr3mIKrTysSrULIfPjh5NU4uDrAonfPofoThn9p9
a/fGhN7rSAeofDD+pOiRljNYngGMTVAJCiwoYO8DOYZLTxikuPOLjyHEQOHaFlp/KoYA6xW93NcQ
VlkPbufE3eSOYMA4nyKmGKRAzSVvCoU2lVid+3YJyjBfVPYp4UM0M4Bfcj+DEPTUG2AbjBrVGOGP
1VkglrGlubhSgEjX9Vf3zk8adL7Aj2aJi9U0WH4UvlM5530k7s3RkbLcObmy51lJYGrY6+u2uwtd
b3wATVPbaBlmPupnbth/PUkg6cTzTllOaLY8ZBEbL+uRxKcXIPaQCsw32KR8Mma9ebwRguOmG0Qc
m8+AIj6PDsWgI49RjAQaR1jwwNX8uZ4VnC4K3pr3S5eHKnDP/Wy80x6EN/gXDWYbkgHgH8KwKqXp
TLVIdE0Z+/uowzs5Ka57wRb9PujNcDQVMvlqc3faZ4q9l3OeY3AwGTdkW+C/v0M5SdibDjG2dNGZ
GiIuZj8SItcUimE4LQ1zSBUmBCalQzKQwv75zmYp4GBfJEi1/rWSe0AUwXjOzCYQE5uP/hOHrib3
1JVNd49ehvdXTsQeJ0KVo0+U6eC8W6r3GYtwORNgU+Wq8BbWnPifP2IXNiY4A95Xl4p2BoJD3Glr
SbKuR6QCkUdAbYO5HNnOL72Sb/Qx1DFAdnWM7Mi+HrLreBD2hSTPI3RFDR/8hV8pLl+qydMdCbFw
ghpUZTJlfTkSPzrdINEf5xPPcr4CeY2tB4v6ZnmTPB8DxmDaN4nS17krBFcYKQAl1toOsm2nn6Ae
8JeTxejtjVylAYCGUKz+sZ2E4yNkaBCHdaJcxD0/O+7S1skh3FpF+3sipukVDuqdGDWhD05zIEvP
VQuWQxRrbbC4fET79bFwUGEdFmkA9SzPH6F4fJ5sS1zPljwCpJU0M/61t5XZdgbWbkDFUM7FB0Lv
lbMXUpBDGwYIAchCjCDg89VG2iDoeFD0T8ZeYM/oU3uqLOqh4X7P+Z1O1iKwVNtShaTXtcWWmTSQ
cZivvy2PoQvkHZaIGBDwJximXi2R6b5OXZ8sEoakSwl+hPuvz4VaVWA9Vce11KHyfYAIBTk7uBMd
IdyeyF13fv5OnsgCviio+X1n4jjbY+Us/q3qRjWV2U7oWm6Hqdcr54k4qFFyCfZpfJryepaqyqQj
jWhQm7lo6F5nXXyC7ionFgjdcyhsSIAUeX5Sf2O8zf7KaejeMwYKIxBMnOlttmEnujLndW1i1YJV
0z+VQYxYbg5grORtfPoA7MbxDOwR21od6zpMUcX5fsNjfAb1mIqpstiiL3CB/ZDfIdG9gTSMoWxU
R1aBq4qiq2l8q+ltnd6CZsEG+io5r4GQusbLvtuCPduvCZwAsTP7Qe9DzK3Md6S5YWTkMG5VJClX
kGUv99NfIzRk/KKlICUtq7R1QKywIpm9urdjL14UC9It5+rjWU93yvp+2dRGXZy8MxhY6Cs98XTm
URHs1Osb3ZdoMGkMlud02QgXH04QPjcRBchZAtDfwQBAYSHY02UOXxbhFX1d2iannv78acNY2/s7
xhhrW9eDPvxcuH1HiLXKAKLqKeTrDlnULE3nI4XWqGn2sf5bnOFLEn91I8yl4ajNgeCgjKuAd1SD
SFr9Mj5ajzI+ZMCgQDfWGOr/yKGKhB2860+FR2B/d3BMfXNGAchKjkWNffrPCsr7NROOh3KZDSh4
UqLmrmjFzS1VLG13RlygmZjzAhp0iCmRD/rcgCPronLwIMicfqzK1ZywA01oKZc/eZeS/bEAIG9I
5p5roygXyLaMcw5FfEt0b9cnoxz2Gkf45ieoH3fudd5+/Hk7d1BzKSLguRh43kdcSu6vvp2Uy9Gd
KLc5dYdF7yClcnsEqU7kmT/Ee6JXLJxc8aNeW6N7AtNaJZpqPFL9GvvrkTuSmco5uEAMy0r+RlVO
Sx44p4tXhhrv8tx4nn6lN2ulVIOXjmMZUacL6yOvnqggPCfkR0pzKBiZewYgc2QMGPGBgqu9cKI/
f1P319IRG6ZStqBCI0tVllKenpqEFp/OzV/01ny5lTkqcFxnrlBV9hylR3+E3embhHvA3aeo3E0q
7jJLn+JltngxyJ8ns67wLuNKCnarGmjsLokWo6iD37qml3ZNqs7pjppjQPx3vf6r6ez4rx0kqg+h
g7sMIGB/BITT/o1wMeDJnyfJU3SPcNliFuaiNXPlAvrNbL/0e6rv2frtQyL8vEReZ9sU7xLqNQk7
UOY6IMfYy61MfGtM3jBWmUndreMXyWasku/AldcrrPPaiaawU+SjxxJIuQrEl8BDyciCOE7IdHSk
tuCkfEFy++SuNroHnWSza9tAB7hs7Y++H/iee7AvMrdZVW0oLhda5Jh+/S2bKCjti9pHP8Dca5kf
H4DtLR1M/+GIR6y2zjHZ9KQKTl7jhpNUBYmc5viFQeHomH8isEYSiTL+IxZmV2tjyM8kMzIm2b8I
8zWn0VQXcQSPAlMFrsMrhxfGxv/5EbiiGvJvNWvFp0MY4WYk7Gv5G+67qpvtpIQRx8GaG0KGkKYc
V4fMoNG+oKbAT13lEHEXhgvTagHiS6LeyQHx8ssrbRuzkACoNVQJ4E+Booh917Knk0owHvorTQ4M
2Xj1worws9ZkinAi4/v4FKM6sNqnmcimgFpzBOrl57R5BX2Z6rHELROLfCqPLbYSsKY8egTqeHTv
uD91K/edw7d70+gMX4S4fPdamvkDVO1e850NCfkyyiZaEtz6aYoevzFcAxq5xZDHhfKI04fpY/bk
w8PaCBYE3e1BNWW0296yS9bQVM84J+x7afM24SisXKLKHHU+dsBqKJnmHg99XpSFC9WJ16NE9e4e
k4bC24REt3p9JR1vlDfJ3UWjBZ3WBJtiyQl0ut9DXigVxGg8/gitVnm9JAWfZESbAKR3Fbj4mIY3
zGcJOYHB26y8DcigtHumlE0H0rtYc37aOz9WqaNvhAYEUyecVc1EvCCY5MpDirCkUXk7wcS0ZoSf
9eUj/0hwbL6k59bGWPa7Wq5DZvjYJ+zWqU1zTRiW6Yx86F80dYJH7mR4K5EZXN/32CCn8XJkth3k
pvqGC6U1n2BQny8ubnO5KMJJQJkLAYpZNuhZq8nq68eda8njZb5DvLttbnJL4zGfZRyC3KZUVMDX
YK85pqRpOv4WfW7bqPB7SNwa3PKVOOECLg2NFbcypxWCiC5nnjDHWF5PUsMGjVX/RB3rPrMRtEe/
K1mPh1j7SXUFytjqo+y+PbxMu1ZCYejproSHqkCvlKL9Grs7jKn3qn/5zCdPiboQBnjuoybhKIsV
RtY7HKO1qON4A4raLKOvyoLwdCkF+E0ILFse31dMxulb2b+b7gi6zKv6GgUe8DQvzuwCVu+C0/AG
/oHFhlP9dXtwww89G/RCKn0Y1wxzqd45Bpapqy4Fjl/mQX7kiEYjuv5IIfmEfdxX3Wonl11b57EL
xzmgBT1mvaCwYvxWdn+8lLvgpf2zUxC9B92vLu1BvcdlUgaG2UdONX61v2XJBW+fXe4zsV/J7mQu
XEdz1gxvMXx+D0XfuNYQlD5lG/iHWXboOMwYeOok42gy0STl+UOff5VVf/O8bzREG8IPpl6v5kPA
hpt4MSWWskf+S5tXX+I2NH+zTVbaC+Nu97c+RM1qiylc9EfKPQks7K/i+kbA5/vKPyPqpQyfhjP5
tpKjqMtXRfFDM4kXIJH6eygTHfgXMOfXi4FvYSoYH//jAzVv3ICJtR325DSS3fd9YqpFLFnLN+We
1HlsVH/j08npxfz5LUG/M6m09oVKyKEOLtR7Hmh4Ab277ysNlqT6C8chG3a3ZQq1mUy/LcNjuUHn
WHglqKbAhpmhslVHph3+ygA7P9/NLXPmrncAfo3XvNf3act9ilTgz5x8nfkAeZ6zHlaiE3Q3KuUw
Z73b6W30YTXql2/2gBog9aYB9sUQ32rAO1DMC5UhPK/RYVmgRv639NKZVPkUxL3/NLbhzsefUPnN
w5gz6pRiLRTXNbl1w7+vxdKl225+PVnvs7WNYrOLRyWawTkqotgW6Aqcy0qVztBPcYde+dwdgrkb
wdvZpjzpl9ZY5y1r8CJhxgQSsBcRPKrYa+faPrHuTPovt7e85LUU5iEpQY3dfSVpC4tnurrSd5gP
5n1ksvTlRm32FoNyT0wtsSx0BGz/gqrxnW1KXiNUe+Hb/Xo3IALS5agecENzjahLYyLSfEOKvxJf
1/eWm+MQVxXU7Z2sLrDL4ibGcA5v3n5WrkqFiagwGwTwE90I5RLNRP9ZdgYsiVPNcMTiLTy5olyY
SZxcr7xHfCHYU6SzkvT05+BmLIY/E+0JA+aFrlyQMIpcsyyiXO25fDsYyOh98vDzcpSPE2twydb0
+m0AzNSIFgwJ7AQcmIjf1Io/eEYa8C7AC3MDAgq1//2mJF8Grp+alBULxkuB/pYfNknU5UhBwgKm
x190+Ys2KWxK/n0OMeaJ8MiLZIkZfKBJ9BhyOK+pNzNZHFtnCVvYeBqey3tqsZR9OI2P5hi7eEqG
vlWG/h1gPDy7494AH0ReCLELxwsUmaJRgAUJWV6SZIEGZfxX/DXno3yrIs51ljmCfdvm7C3jahjn
4b7Z1VCSgolDQe9+SvGjxFEkUXkbB9tweTGo9LVpQHLdCD+LmEfhUWwII6v1Yg7CAgEl4EHzIAjv
m42AHY4rdNCS1JyXLj7ss+qbkpnNfhlNBiSazcFhXrHTWbJ5UCe7+XU9VYcd9CApCiZ9do8EDRQL
HWO7PloUCOrMOcbbG5fWe1a9+3F9NbCKlk/B0W9evH5L+/OniQ8Ir3TWM6EVtblKvusvLEDpiJES
2U0y8Iaaa8yj9CUPHJoPTTyb6B0GfdzJ9Zg7LJAE1xLJtF/e5PgqPK/smhXG8m5mo50Mdco1otkU
jDZROl7ARlRsNb1hppCOieCjp3G4M9BIyIEee3G7kOESJWZ6m33qDqNG2jNnGDnZ9HmygiaJBFA4
RuJrTaDD1bPL+71Z4B/FztYDEJDtTyeHM15OZTnO4kUVTGNR3DJYA+hTz3rwfVWAJMfo5/1AMjQD
nFFu1phtm5BlqdXbIa+ld1SV+9+QA9HSNADRq3RzZLpWQEf0R9k+jLA7a6o/Q5IYBtW0shYApXT7
CUdwWbqPUx7pyVhKd7ddbmFu/JRV4C+/EzAZSWskfw+Y6FoOZrnreU/DZj/GUjrEOCVQwLUPk9al
F7IMEZg0VWnafnF3/kVJpVQaVhvkfFgyOdemLSnA40+wDTpMAG74KpFx2ur2zvClQ0f037Jt8nEW
T7bxDNFZIO3thogRryP0xM/4JGSNg2LTql+7L9oiOoMElveSS0OxQLDD7rZj/x1AC2n8tEsOkHpB
F8vbz4ELhW3KMlC/j9/iDuI9ir6agsA3vkMBD3qCFefga8+S8kC5La+34QKtvFYvnBR/V6Mjfv65
iEvSgj1JoX/QFiaY4sLa9oLWXcIwxWZbKhJzEo5OgipRRmLZoMuDmMn1fPKms3u3IMtvxx1yKVBB
Ueh3muNJgwABk8WHjph4eXEsR7BwbVs+JVUWxylWXAyIb+6XoW2BfOEW8/2VleZ5zdcZ9LztSC19
t+mDHyTyJEIQdbtlfSanutGiJCMiSTfoDuo8VN223sfTLTv14yUOFXUiALTrCVsMpXbyzzvcI0kV
CGALf66CrqP33QVcOAshcTRSb5UlKRMHrAbak8L4A8Ga10YQlOn4Rw4cPBt9khfYHD8r/mncBKK9
Ck3FABiLMvECTpxgLZKWOChD4NrkcIoF1tiIvrIEPF6iJh5NlHkxl+skrdoQalxdIuTHJpniCWsJ
K3dIS1skktIohAGRDXIwU/PD/QMbQDJ66fIYMFMnmPwTAKq6nMnO8vb8u55qaj+ui7eQ7Qied3ku
jZ9u4A77VShnz9cZFPJF2UcFgEjKVnlqMfbqpxegmhUAeXMVYFmZC3rKxHcBGSmqlEPvkvcBOQxZ
g5RVm64kh/rfxnLPJKdXLpjqqZZbW6fE7RTaUtTwDKsBukLFE22ASujLOuegwFfRYbZvqkwk3gEx
v4ufGE/GcskPDQOvmeh5uFjm1bsgI68rGMz3lUNe8yAkFIiNpg+/k8KtNBLvloOQSSrCmyAG5PxP
EaUFrKUXnBOYVZCDvNQzzWL+L2TbIAY9+6NOi5f92Bjwb2HqCeQZIVl6Igggjbw93xiIxRNzpIGJ
OjnyR+W5KPd16MQL0CQTe3bcAeA6An2kBdbpFp4l/iOmzgPrgeiLwB7kOzgKPQI71J/kJcYmH8qK
g5LR5L42wMXsp0rloyKgezqaBp1i37FSe/Hxdstvv7RejGYyN6ouLLExCNAIl/E2tGlnEMuOh9Ye
KPnEV9RwyJhNo5TNOla1dtjlQygBokeBtL1vC4HAKxqTDxUek7CIj38uR2UcZA37asl4oJ8yJnNe
2Ebh0/BLCHsfRof+KE5YSRkVajoTBXGG0Jo/LE3xTGwQAATakYIzIE2kOllJtt/YnGR6hYe9q05B
ir6gcNs5dw3dSG5ttJxE9buO4jmFkSwYXi1vvxKeq8QULOSzOCs8PP2VRAHGGDJJb2Zw5+oNzJ2u
nrzqjsnDQgNZgbxPkh3tfMUbKSdeyEXNomOnxmo09UMtgMzCPokVPOvnDnSKXGEhsPBsfdmvZeeK
Zn2+VL3Vz1F5KJTrsQ5EYpCvjL6XxvnWR5Lqtdchn3qN8ObUxS9V8YSSO9sW5epusng5JdyyF8AW
wDJdhKQi5rpIvOGM18V6O3/7AJVlSM9s3zqRljVFjMBn8qDIA4v2Zfo5QUNhCDUMBNRQQ/fsIBiP
aetHVrEpoaN7bVaDUfQynL0u5e7rmGRbxtNV8AX50+BHnlR3fiz74s9grSG4e2pIJloEI/pvNx3j
lhEfaVMe0euZUlgNRtEaRxfvZm4/BarXLISBCRcf63Am69PkAPSQclBcJ5LTHHSQCwzhI2glne7v
PyRGmpLyIVhvCeo7V8KttqTBD39n5F04KN1SYRKmjeRHn5y/TjaIDDKbWJ+JVJqLW9qMr0dKiga7
We/CeokAWE8JIQCoBEYHgwvP0jwJ6jYPb36KhTczQdZGC+mI+vkJdlcKi0N0VlelVONid4AIk/B4
ZLJBvK3ZAr2J9AvlEkp5MUuXJbjOyQmGY9QnsLjfm2KwKu+q3Q/+7emGI+18pxWSBaope04md2TX
OyB4cBwjEnzwv8waxbw9+uEuOKsKmLMhNaNQODPFZkR54u2lQ1XQ7vXOdz9q7Sbgo+NHu04fv7Oy
kmxC3TgRSlWR7pvAqqN138NIOIyqXbI19aOCPnwC/461O03RwsewGM16zgjQMedxGNymoMN31h3C
bnZUDLNbazpRwgyoEYtlhxqVNs5eNKyUwXNdcM3ejcztNWcyidqU6gJygbNJ0z0PJkLHnyzOGbBT
N/h+WOCYL8PZXfTFmobXZKYwWdSdCZ2nX+W7yVcYifPylFnuVbX/vp1sX55r88gi5gTHLeNmkQx1
j8u3sH8/N42PpJEvW2ZqOIurbqc+vxOqIav1MICT843fxDjJdaRZ0P+T6+2N75zwNIkPr3bzjcMt
S5JT/yCGANn+o3qdZD4Od93uLmCgBjox3QIlBERCWGVs9Unj1Cbn/5ZXletc+MBKaoARr2+LD0XE
/mBl67ANvt70nQGNs8GS3smnWZDGTHhZkRGJS62PaAzQna+V0IJNWMdJX96YSWQpuYv/IpsiGfVV
FikdL1SNn0In8TQXcIe+gt8sbSLEfM01H+v7t8NbRW3Ri2U3DTkJXrIZ2SrT8sPKD4nBJjFgZ50v
TfFMQN0abZgC37g4vsCpeynSqbpV+BAIPHCS0V/My0600NbYRhuLT8uaPlvILW4LJxJsaiWkpxFk
SWG46vi0qJOUY30/M7psnjq2fdtDDakRRnXjot2eC2c7tKYxIH5kS0RIoonytM1LiKzqu2JeI444
zCzknyWC2nHAdmfuHP0fDBVlWtAZr65d5mv8zksuW7pHV7V8nBMk2/xbGvgEQ1VdpU8S9OxnQ7EG
g7K+/EFYttmtv1ARWVIQcNCK5AyP/OCdddRMk4KakNFW41YHymucBrhp0+MmW9cllk0O9EjL81dt
h7jnuMhMhlCbnEGdfuGwNmx3EBE7+dccQ63+4T5FW9chLbVm8QNqRuQ0kKIn5ggaH1zBbmc7LwvS
ClPZyjy6wovr2M2v57VUSfOy2nnxwck1ff3jqtcgHY+bJpRKPk3UIOedYr4cUVRftWb6rs6dP7Nx
JHSaTRciYoOgtuyb/6PqVcAuvRGumv0fIDlHt15nKiZUxAa4nWAXm6TB4JvmQBejNuIXOQ6YsjgJ
qXbV/83IITAYUFOnBp//zS+2JQU33HLtaKofBwIAwt1zjKN4SsalT87tYvmfWLgfx6nn9eaAIPUb
t1Hpcp5pEM2m8NDvWHfXaXKjou0p/ZYsajELLmxlU64UojVsVStHAvOqrxu1SUDjvXo2WzKBk9jk
kr5Su74BB2hTMBpv+N3tnCzIXBQ9GrfJITXzHpYWDXxKUvxFyBBIGlbmV/Xzs289bLC8/nvGuQP6
g2tb0AK4dI0IQUs911bFqCwg5aSE2YfeArHvmwe7v/y7C/HVou26y61m9ssglpUeCiVyw/CLum/C
dBweoYprhUZdunIyR9BdCOWZYW0kHwQqPGo89RcHWRk+qkR6r9zt5J1djcLum3+UGl/tlA7cFMbs
TB1Rv1BrtkjgP+1WuzNNY6UlVRJiNLAbA5izBUVFAmMexvmCx53O1QCLoYgz2yXw4txfcRpvX++7
m3pFjG40gXqNeG5x2IClmP7njEcZ9EH8O26+ySqpGYD/Y+4vbVbug+4b13wVIzwOTKdnVbKoBJ2R
TeVu2T7qXR98PxVNkG6G20JFaYqSRWaXU+HzWKRbz1jr+W4SI3GVrz872BUWLvzY62Po+WnuKLzv
e8oAaFg0wJJluL1Yk8daQJmI+jkerTy74Spj0hwV3Tjw0kbE2SPzRvtbrMXSHi70BtiBu15olTP9
rgaBLx1M33DLCWJRDWSSeefFbAyG/5YhYbPK7qqjASb58z7ZNUbjk2mGG9et7uCYYTaHeB6kcLSl
HV4jeLuA7V0sDY4I8QSwnvfnNm65vqbUb/6PJXWDBCF//v6mdJcO2lodyfyFo0JhMscLNJKCl7z2
G6mEKEjmrxH4h++J8izcEtXp0qHIds75HRcO6OiKc8GxdXdBuNAZS2//mqpOvrblpuT0IK4dO0xk
0C0i7HhEig9pyq10gE8vdTgrJGIWMiRFNOIwiPleJTeI5xwr9koXYz1OnWDddUVneIkQ3sAnobg5
t+JJe3gpBWEfns3JPbbc7EbmgUT/QQeLolFAP9cBZJ+om0AhVAk/QpyQ2GknaEq2czEivAyLU4ii
7SfE6sHposSYNbCLNVPiKr9zAgEgyXOFYNJQEhh1PZqaLRYmOcaP77cM4sxAvcNS30FEztJwuAMj
wyuoUAnt8OpKqhVCjqEWg9lFZocov2EAKUyU/Er2uRX5wSI8Y68uwfWEVEjQ92LuVbNAnK26rJ01
v8mOjWwbVugJgnmLEUHLKkAiB7fy0wAZLLCADbynzGcrkujYErkdESA8siRTARYlSANBjSvNo0At
JMiutIN2HtWIHY+VPibm2NbIA+Mr2bx2xKHPQOqcRBl+Rt+ImWqmwJUOLz1Xv20Bgqfv9hFX4a5h
TPBbkonnAIDoOHoL3spfOFfcGEV35VdBNTAGAxrhoU8/KiAuSrdzCo8DSerJnfxaM1/hXr9JTttS
UidA4KqCTacPbwJHUOoElumBAa61MEjB7uvRwYshPBV9WL9P2KBu6Nah1codCeATmaYf9Syc4eLQ
MMLOZOXHnPztT6srOX0I/LYIcGlB/+cHdWlLsGUvRBpepY4mzuB9/DwI/qFd8NeHNdgown3Zagug
Z2g3WntIA1581beSRhSM1hlJkReujKLhbypoaCprBhsD/4JEv/IyWeSacLQSoGPCGg9ZUDYwNYmI
HNeDMQK90HoDqqRYoV6jtq0agYnGaGINLGWKBwhIdnEAGQx2cJvkawb1LHuX//KcJcIh/1YHQVVT
fJPjZyZnbyFux2sypM2bzB6+rLBVRo4Fw9gitrmjt5o0oPWfP42PARpuPTC25Fw0U/mONgcPz3Et
znuI3rWHCFJHTJr2cK3BBTxkQD7bnRyDMRPJrtWFkIpeDEoRv+8xyiGjVKVl+56VeH0IEFey57Kc
lszBekvwdJyQGVMWI7o1MxjVo+nWmBl4S80S4yplWxtwopuH7aEMCW/UNnxYlxYwxGjEAo0zGqqb
xopA0CRfnFVBL4SzlbopkF/el2qWrf9ACBZOLDK+cBswwyMc6D4UlLJVwLIlkZCD3y+zOrrODZUR
ggpRR7m8mLmTDTx388YMxd+0eRV6XBQJbLo2M6glalXZ/Umznn5yPuG36EhXWQJvFttwbMiPOUKV
tCpM/biJEiZL+JIrcq8uTjux+hh425UUyItXSjKZobbC9aKVSFDcMvEmS0pvdzQ818aU0TufGgKL
nHGK82tUWXH0k1RpJyTUWTHbDlpUk+DCbcpw0qrqPM6O5O3gZDs71q0mqzXMJCKOFnWVPUDBGOLA
w9hPiNi93d/urmXJIAKtjELqw2q7XtL7BI6le+Fitp1FZO2zjmkWAvfnMLnQnryboFe4kIsbJQf9
Jc5jP0A+DBQI2F78NJot8jBnFy3SeGUHBiYan8/qeeK5I1xT9fJ5Qu+Jy/+svcQLgHPAZNk+vZx9
0zmzhHhudCeHCW/Ey6PjWvppuS+gEYDv4nTcbTBwXk+rqsq6omCgD8cKdZfV//+xdrNNmLxJt6Wj
Cb51Olgo/O7UkSVjsqdwdbtFT7r5zfv/35r1eyqMW8ojdEQPBv64TguwyBrhhGa2LXYNU3AX6C+U
4kqhdhcD21YyN5MPqUAKFxUTLYtLFmdqLLCUR9gfE470fTjAh35ST4L++c2ttPzfGjZB/B+9+kKr
PUzqgjSvpt3krKfuZ848FYNv92EuSV7c5odtEWtdi5y7sIozI7ZwVcjSNDWgd6dub5U20PrfsXsG
M1G+55QEGcaPxbh3vjq4R3GZIuCQBwUkK5iN1YmpEwHUIYqAwkdPTYCpRlDbx33MGSWy03QUDPtP
Vr36WUtHWWIIvbfP86MQr+c/G2irPlTBNh/t/DESdUQElIv+jMaU7irU56POsiLPcdjXp4Tfvzrh
EEjNOi7o4p7o7+DixYy+c5wlP7KLELepkWMk0I4Nm5pAfWYYFTuUFL+c/PBMzzlenjoHcxG76qzl
JgGacf3lVjJWDaZtQ1yw33coRgsdxVA+WM7po+Wh5muYlVRqJyoWX356/i+5KSNG+f2zSzDUsG1p
uS1rqZQtva63HY979nNBqEVFj+Op+Bi5T8w8tXCAC30sMiFvVtiD1ewmHR7lWVSlf2FBBsZ19SPK
fR87R+xvXeavYOC9ZPhjm1UMhzo6t23ZzgPam8467SF1r2j4uZmowya4JzBcMiun/fnOwrvfvdbV
mnaalXv3Klq2E0C8KPyAusVESqvBJwCf8OOyzPiLG2P3YcOfYCW3K4On3YpNpLJcDIYZhv8d+b1R
jkh1zEcR1gdPebB08d4ABaOGGKfZeo6I5RkvEls5UJB5AIfzQrE8fmQRkH9DxKEDTOp7ctXuw1UI
1JMSROwTGZUrnfdqt+L6SaVOawdX3gsoyptW1+XLKymEvqe050bL8RMgIckjvC2IqCmiDdXf+Yd3
YuHO1h1ZafoG4kF1BsZTNVCs8+l5dhHFyJo+OO2bYGO7W71ZTRxzYsgPax5E5YUT6shamS05icKi
XhOTLzvMhTzyFV1IzVt0ZVGpiDcPrkEbosqTMqdwOsOteX+c4MGVDnGOgq19ikJ9qk5asNEZHMVc
vr1eemDPYhwvr6MPkYwl/NGKppfeuRmpkzsHL+FeZrhAkuVkOWJ8NgV/Uj4pQ5BkBfKV1H7bUSDA
fRH1iEz7HxTz3irNbWPDoUQ7as7nCGVStVJS5Kic7qDcg92F8pPqrn6SwK52NDS7Wbng8fGB7zSv
i637GM6mUmam581VF24fTwHRFgQv47/dKskBRbKuSWPsQeI7fnjSBRwy3/XfyrQ6C9lNcGshFKy3
f68RXBWVRkkyTG+ZS8ODGli39PIQwF4Zoeff6OucrQ25tOcFm177sbG20zRzE/YqNnT1hO31bafU
Lt3pU4OhdnaKC07Yh1sZYNttP5yNRSOm4bvS2Ce6BkDtRNLkCF4oDM7pCk/rYuDwU5aDS4uNqr6d
U6Jk4wvmrcJD80QLbg0x4vT7ZbwNiiMqcr9eI8A3omTqRf/zF13P1Fy38rrrYgRQEtTL2PHP7D/S
FMtXpCoQGXJkWKbyK503z7QazuX475QvZA0T9kjm9yqjk2xf/Qi/JVGXRcEPhu68QIEbOMB1/8b3
OEDHJe1rI31eF9W8x4vD3Olli4N7kfFBMq/Oa6gN4n/+A6se3agMrpMivTHRMEZElpsW4Q2AXq20
WL4Sv41COVHUktS2iEgOgYcFmMV1aCe1CcNHUvcwBSkEOtdDWBHzeyg6eqOyVaLeYDKBiD+NQMPQ
cxI6JRT16CxwO7Q8Lue0XHsNsBtlI9E9PHKI25SERBAhaS6bfu7QO+MdVdYleAoM9Rp4Tog0BTwa
kvr1ll372tMk5y+jP1rjKt3KeJDcED4M4SmmmAei2slEEYVVtrU8/ivXwvG+p926eRTtOfE4FFnM
Xg44cPCA8ZWvA5Lh7sYg3jeeS0NuiLJvld6Qc0DXNSTP4MuoC8MnebnYZoMsSCgcPR+aowI3yWso
hzOcs9eOTzB1oyvzdboVhcL99bRqGwHATVI8Z2K9hh3QQ0UsO2t54ujTPeYbe2XJTgVDcQY1QO1Z
4vP7d9KDIJ1t3VQWB5oQx8gAjckH5uZv86gQotXHm7ID0B7F4Y8ZgJiRuv/xbFWXXj+LTFeZUQn3
VoAtkcgg0zXJestpS7kea5ctJkc4vWI75/Z8Wzab4jPxWORtHgUnqRtc/jW66b4/Eb6kFD58MR/0
32+h+xKAG+uZyb4cpBVJ6+f51R1Z6GLOQsmU2TPtWSg4FFRF38OdD3GqkoyDmIRBWBX8DnmFZGVz
DH0i7dMLXk6ayZepQcCzjKbHmhgKnNyIT354MjekX87WbcxvgS3aJwZiy6DaQEe/Hp+Uy+vYeQmJ
h7eXlhgkXBtkVmJ3cHxjf8tY5n288+BdkeKNtnBQg4yShuRPoFfa4RJFuvjYbgk2J0FszzeR5VpR
Ecs1OEbIwW92MLOVl9Beaz1hwPrDoOMhzKv+I9LggMTMu69OP0yQp2/RCgjFb2LSFRp3ZCI29xIH
N0p/lMmkR4C02zikvBOjM+X+muf3PRUdG3SXTnRP4m0gi8ziyo0sULT8Fs2LQEb3KPwjwnmvQumi
YpRIIkxxSDp89WoCg/JUCXcAICT57kqXyl0kKo+cOZRgPf4HuWzr7kQ7UQglVzmfTfS9cM6IAm9f
9ZWw3zkPbOuqZe84UJ+1zGGUJWjM84M3ZflKA14tTWyofWvEbSHJEaMryItVmBYSQ9UmipkYizMR
brvu0shGI8fgt9Yc3XdzsgihZaspKUu+dvM5aVycy/mV9Sga0joNLxuEIwaE0c5O/3wC5J2hpAIz
GPuiePIre1wxvE9M7OctwcBr15a1G5CU305KEB97uIVPoZmHBqv9PAok7Rpkay0rWoldt6+ap+m8
8tt8VRuHpySoAMkTIx2M/ITCWb64CgF2ZW9U1PV52c1TnkwfEcAOgpmSAKR4tOPnCsIpC6/Lsot0
PRyp0bCr+aOUSU4jq+nxw4Rf4gydN6JvdGzOAUWLq+cSDfS/LIbIP/fif1XOycmeVnGwdpxEj+ES
7EY/v7BZVEG5VRv0s/AfsAL82OWcdJrQXzJ66czZj+24KFrp0mgzSubI19ipC3G9jogCGCHbpIhv
yyZmk9NUsxqx+/Ixpf7cPtuisit2jDStmf1m6QA9T2ixKVuXCo0+jia/fr7gNbJt8V/asw+Dgse6
mcu2OhTeEkXlBqepDk9X6Kw3TF3L/DhWUFjVdp2nA0Dg68stexcnDKwkNcOGoddu5kTW43zA8HUu
YQOuWQvtAcay7adiSEEK5JQWG00m2DVn6kecOCmtbXHyYEGv/mkrQVAPnkvBcMbXveh46mmlbX05
X+haOJfbfpAREdm6QZsOfG1ps5r+U1HpQS1fDO8K+T4d++kUBuBKLlkjd22mb1amIoa9chV5RwFk
iXyCMt5bacSaEhc6bHryjkdKfa9GyVrFQcKZ7B2f/kgBk4S+7EHqRX8fLFIGDShB93kkbojjNu/M
emC+VB0+N07Rj5EglYFyfBssmTCEHGZA5900BH7f3GPP7qFgoVOGAjxDVXMefvQG0X5SJgaR2ohA
abOhRml9stB3KOizlQHJMMz4+fSz/RGoCfRK0F67sstM03Ow47wFiOPTlcLSUQJzZHzBd7ZfEcgv
O7RB1K6TrkHYuF28IwtJ95AiNNFuQHyIxA3UsPbawkJ+EPuixByIoQq3rAglropE7Mgbu6k+zqxf
5EYlBiPtHXOIqKjS5U/EaXl3eLE8UnzzY1XrsNDdNnCUGx/j/0L1Iz6MJ8uREDY83/pc88q34cNA
oa0lqOziwZ1HhWjQ+1BbR7zkB7Xz5Vv9Ty12AslwQxsM6SIEEnvtBNUrLf9y1lE2/OZ9S7Er+Ro5
4jN+WrCkWXbZJIHwkaeMdgdFpduirHXoHIdGYkPaxnwbzZK4jkS/rkZRGC5Ox/+RnHVisa4LGrlp
BNL/4W1sU/WT7eNZYxHS2HpPLxMFwVr9lEEBzhG5PfoOVfk1Vt6jcHaONcIgv6g43qaBXLv8iyR3
yVklFJ7M0b7mptIQGjB3F8qcDtSp9cWm8qrdQlmHpaKLupn+nObCRwdeGhHrhsc1s7TblTVPiaGV
jJNMvce1CsyePDJIBZaU1xwDn69Z8bCTgUSctkFuFCRB0gmNY1/+iYuSw4qChQTw72k0UrLBwwQb
6HFh2tlJQausmcw/Y4RBlzLp//sq5M8pFR/hGarg3I+REIjGuNeW/R8v2gDLmShLnQTHIGovyMf0
lXywThGSOL6Q3V7lDZSHR0q4YQ9eV4ftxave8L6UKDRwZF5eeSFzE4ctyv1fB4zK8xTr/YXShE2K
kPHTns9Vh8VpXlhFyTtqi0jeONHYV6rpRYhKiBt/i2+IKe8QE19Td49OHGO094lxeivIFxUk5/iC
0qe/Xp5SCKu71cFXo0PslWNJzo7oHj0QbXiI0ya78nrU2L7SpG8gcnWmeEWUHuaaJbkgfFySBqit
JLXtvWW3nQmgiMEZAeXSn7klqzxbL6qrmz+458POmWdsvyAWUrgk4IXruQLLBP8yxVjdeOZ88+1w
8mLLhumc2u8BxhvLSFCrctS9jTOymTn8jUL/NwWAJNrCJNhgFwf4ZZhGUxAuqfPOem3uMWc5r4IV
C+34espHp0xeg0lGC2cEALs8KKOvPXpO3T7IyLvsdVhyCR5o/m9yGJEhuRfxPJlKk80YV2iKBvRV
lsdB/kemHJwlJWTv3liKBDZ/8J/W8UuVkDAI6symBbXynFC0MJMQq5iDC8qU/5gJVc+WlQs2E9Tc
4oWtuoXs4f795iCCs2tjWvr493hOqIsSBi8/2GbC24Iv2l9/ZM4c3hOoaT7HJumOB6LDaycXKL7H
N7wq3fFhiDQgaCbebpiELTKvPAiiVGG0SOWrgQLvanqHaJB87IeQmHvhan1gWBOomSna8kUkgdEr
rwuXnslpfoouf4y8F5V/Z7HZs95gXevHxTktz3bn/vMDlgtmsDnR/r6QgEzNpR1FwmRHRo+9oMML
bBbo3TcNq+FgEjRNaBzfG0A+5NXaE2OymWGXPdyT9rpOmno2BDXTMXAr7fuD+bgTNxAQDbuzjnMm
Wmj/F2zNvisvRSXvpi29/7C6NrWJRWwtmVZ0EQajOjnW4efDUpgUxzrl5jTHfc2XQV8Dnq8k1tDT
fneME+pM0mbqFffeACcJ5AAb2pgz7eUlmd6Uvhwt0LGdIi6zKOHXsqkDD/dLFNahuZOWhWwOYmRW
L1w5w7JFoFG3o4abQe1/jn2jey5ij6Xu7GWVprJWorXDIY94ndcK0ZmnNG+5ivESSV36F9pZPEAx
PZCsTpnjjrNJO35BsI1xrXLeHPEQGzwJ5dI+XvvOOiX862tZvXW2lA32hA3x7HGlmda+k8tad+kq
deD8uNClxfKU8mz8jkHwmZ5rXVXKwLv83uVpQnLs6LU9l+fIwNyD+LwoCLgQQ9830D7P10ASO6QW
9TLnXVoeV5mi8AGegY/Z3xNndPi6QvlQpXuxDWMWuo/Gns1S1HWR9oeLIH1leE9iDGxbAZ+Wt/mo
VEHuD6J+HbcsFcDN68sVTuha2xYnNj+DfsevRwXYjLCALCAn4m/bxhQSfyy8TOHZv0d7LoKLhHMQ
7pkyVQA0LVDJQoQoq0OSAsXLRcZdl9PrYtJ8XZTxhNuKB8n8hjIiPtTNItDadXuUrtXt2N9xCrYZ
xH7AeSD2c2Sbx0xUHVZxdyFeJm25184Kv9+VT+BxZkOZ3S5xMlvbgU2fR9Vodme7nc9VjPrga1An
+O7KNI0acUxwQkpiGa0z3mU+eDxaPNYVH3l/L5HCiTtdTIQlmo5hH0/aAZxGHRCHgs6DbNTFAyQS
VjQEz9F2LY3wC/PyLtPe7/YzuWWFQjC/w5ct/TdYfYUhnw1QEElfw15AxGncv8RsUQc5ZGBzbf8+
Pq7Cf4trrIQYNocBrGM9REdfESiJkc3uhRer2k8U/s1sRIUIBBiQ/iVBBkR5hR5Io+/CoayBwfZr
qPVd+fvEpZ+A2i+KbJ5lB6mP/cH4btXvgWA06nq6PfvXWIJzh2TeyLRUxtjqA0m5pIVvsWqEWc3t
k3xeHrTmQY7TKK/giAqV328YUiKfVzTBPYb68Hdh93peOjsd0ozedyYg13v8wqgQ+HFniiLAGLnT
phpvVYg60+jUl2bLD4oWp37muTnIURBXgAejrydlPgie9jWYI7UDxvd+7sooxhYxpha3UVmv0cwK
Wi1Ab1UwNZkZL2Ny4FUmcGIERjerAMFXXTdaW9kmADV5tv1hfJXEpn/Kb1nI+YKfFu4mOHURmqbn
fLu9RkDBCY9HKlRUfZETM1pmdEROk3megpqDrux1ZuFGLL4nhaPODyBOgIRH0xZ7kTxfFVy0dbAj
scCHfs4rlqanJPnuDBNkPXVvXNmqWAE+V861MqR1Gjq+OaDvzF2viAPFny11vHhHMbI6HMj/M2X+
p4OXbKbTKcGOrE3cNIttoCL6s+tVF19Ixf8YUv0jwln35pFbligahi6vxaqrIZ6Zox1lbNf3zJoE
536Xhg/lP4cw7D/mWZ6K3VwidEzc9raUT0Sv3q3XGoCqsGtYHgfowa057bPAr+ke3lNscSsuIUue
7eU156jQlb7mqfM/4osOxnUSfFrZvqeLiF9ovZPXAWeA+mvWGIcQo0wI1iGefWNoGgWpmMljr9cR
imEE4+9xXG3gafFfv0Pfz5rNtcz0e10aqiwTC1Ei3aeK8Upa/tVrmHsph7r7m5TcqEo6kH1EijhQ
wyHYFgsYkex1ZYvHNK3ajKjY2YxdfgO7fpQrBEsZaRMw9iHFeu3LxPyq1M9FZLT81SVYMJIHL9GP
yk0Ii6JRPkdElUmph+1dXezMLo1iFGSyPsL8n8xLLXuxpFu9omDfDuPHyHFcgKEsv0VNJf+BrWl8
VygXowUpl1f4oJSpeSTkEIys9F3ikMPVSnIuVp4bB0DOlyXdgPwGr5/SkZkGpm84JvY1/TqDf0Ig
ZRwO8lrd3jp979tcQ87a1IJkpHSMxsStk62HgwByhjx9rULFWG1SdltYEx6O+GiO5tM4WlvUuKMS
r50r538bh/64Nne1pnUGYuNB6heQW5BLy6bl8BAotQQfFMR8FzF7nE3k+G68CMkykciIMEHG6DrO
JlG7bpBF3OajhOy1U96j/C34etuJztOFwLoOZn0b7YQDTlVMbrTiLym9MXObk7DGrUUmr+16rlus
orx2covNT26uIjK9L06FJoUltuG7VZwDJE0Uf86n9e/76S8h+Xmtq+Fsw0brKEyfJT2aBKHHuo8j
8xwqJb50BNKMFpzwO2IIRdy2CNQbI/ZgNEzFUshWefWuck0KWkBnaJfV9BWXP/eXO0uIrZyfiLe6
jQloMw6UGGoK4bLQNcrxJaXfcuuVx1OECCnNyANYwufuhYIgw6O5XDQK5pbWO5//ePba4Ngc+gg3
1zxSNXvAbKFaORSZRQVPWb99CNLTtfatT8BLDvobDgqKOSER1EiTmtN+ac3i2gcX0uP5L+tHIenz
WT3oJDE+JpanRrXdJi710+24TOJ36GjT0H/i8znAImloPXv5Fh0yFHKQhJwWUWX4Xz1xI8oV0deX
P57gyzcOaMBAfvrvT5fgpqtL23FQmvNTDQtsNG9vUHY05pCyePsmG5KuKGq/n5TkkFYWwd33iCls
pvaJ9lYfS8QrvNznRPhmTDN4+vfJiTKXs973FKfHCPK4Txe6PhClCWxsHwjqsxliabwz3Xkr4zNh
qtjZGSUERUeN3lMl/hXqVDhb7I/N7oe+mQUPzlJR6YaVMzi26+aMlvS3ro7s3/jCsosropbJcu+J
FrpRWjQvE3JYVy/fzomDIUNW8SJHOMZdZ2IqB7MApYkyeG3lxEFEOXkoCf9mqMAzpb01hepU9deX
p22U7N9WG7Ze6F6idOfa/e73CCQQdybEMuxnpyJxWqhJ5/Kn9SwWb/h6nmDm4gWgs/uc1cJKxZub
MZrnvnelZs1BYz4WFVr9MQjRxKOEVR/EPzmIzt2X+jZEkgF22U7RoR7p/iTt2iy/BlhulELBxpbw
L5vfVkW1xAi5BzTBDzCsUVhiu39rVvwwUOWzKpCJWW9QA2Mi78JisdAvX9t3seMuYCxnFi35RMzS
AyGKtZygKa66P1C2uFGVxYwhLp14RbQ0FhlOHoLEIvc0HurOGivMVDVyF6qo4zUlwS8E+sWUK3J8
peu/P1g6p2KO3DUuapme11KSf1P+r3OfhfFTUi3fdx0mtOP8aHd+LEUkY0z+KUV5mPWrossrNKbm
WlZ+HqkRTDiIPJ0rRNRF7qBoW6GHdXwQOPWVkVgcYQ1vPR1k3orjdnirUJc5UeosjAW9v79mIU7z
lTPQO4nvquJfcyvTCnuTsLdHIpyx9OXqJ3ooS7lWQp/Olj0QpolPFN12zLII3L8+Ud9ng7kfyHtO
fiYLsD4f8BS234FqwM+m+zYTxoM6rfSdsY7nVuU/51+uFENB/OdjJ1NsRGeMcd5fWNZjolOJCv9Y
jsUJnSwDWw2huEVDU3pXeOL/wj74yp8ciJ/QW/uuDlUkHJyXF3zoWUj92plGDf59m9b1TynGNNxf
aIKN7cGnLrT4l7MPCdgjBS9TLDdqRNPCJ+NkHwVd1hNa8wLL2t1e0KepYQd8EpGo9QAs4st2cosG
rtndskcvicHT8sLXmNYtPjH5L6jKT25c83JufFjUj+Bdt33Trqq9qiIWlFuMaX2wF3kjV44mfy5+
PJDpLHYX65HOPd0PO7/GuSaSoMz9AIrlDPuMxJjpRENsD+fPhh7nwI+KpvCe63MBrr5eN6vDn7ew
gJ1CW/B415AlHYcFRqDuKrR6JTYkBV0lINwG6FYvNqt1xltPG2bZn5RVO3A2rfkvTw8mRYEQ7nEm
a9YIWjWRYdQFY0qUOZEyAjgVimFeyFcAyLA0w1E1xG1DSHhzhWVY9bl0dhsye1C/An0GCceyYkiA
dnXhzJ4x7qWA8BWQtxMQf/enNjgLBQJmFEQpTM3X+w9b3UW9+GLGAzwDlRqYWNcFJtM13Az6U3HP
u8Cm0jAlBd8eWTms2J1vbZQbff0JEwO2zc5RkZV7I00OoxkrfbrP5EoacKIikm2ehIxkfvxdXN8m
4W45GIGoUgWhxwCDq3jS7bY7DQOdOjJ3ZxV661QlWWpDXqHfmEuWkGWkNuHxNpaRqa/5T7Kjmiok
A3Ij7UVpWF4TSNVOBtwcH3vm+v07jDZtVL++j39O7anLo2maZfpePBZ0lK7xG+4XREsmYp5u24Uz
ro4A1lFIalIEGTQVtQahuRki6xcreqXIxVgIGmoluIWn8E5Aq5eT4NWCpeyl5sJEI/DvXvhrF2ZM
qAhLKOUoginbX6OxCEFdjEMeN3ft5QP09s6RItvjJwW+NGZWhxc34fCC0P9GZgfuwpuX9VDSD8dg
Rim3g9ok+tCkrsbNU671bP91kGLn1/k9nMfpXxmD5BAs5l/RTQbcxYlmGx2sR82PbWwY4gUeEXvi
NNOuXehzgl7Kq1M17djOCd5x9rsXJFC/+Ao76L2jsA+LCc8g6bLBJ7KJGaAPus6GUTb6Mqgod1Q/
AicoQpxmNVV6iEWdM4x1S/pnkWtGyQgvnwMh4Zn8kCPeOtG5ybrdUD97DZgLUvW8q3byFkGhdqFs
jkPcIauknf0tlNzqjkYhyJyDsCwsghVHo4vXsGHN8t0GorZK95VQZGFL9kQL/xzvXLmFy/WxSq/P
G39pJ7/Jv/5NYqnhBFPTuNkwcBwVAEePIboSy1d5tXFNYOkjiGgIesYebH5lIucwTZpKQ2EPsniX
7hi8LHWsy6N3o82rR4yAJP0ribFuaCQqTa0ks8J4JlOvuse6xDRD3jgDHImxZ3CMJyn/Oivzbl01
SnpIUdyihhc5zdsWM2g/H/o0x4DH8kEp9wn9N/JFNZdq4CahZxcLy6NUQUq9LmDhso+6JcnjI57X
2qn77cs01rbSzrqpghP62h73NVuGjOXxCuhT1NmhaJPs9nLjnDOUzJsyq3ly6k5L38/SXbypu4iN
1zfNyhjRZI2XNvEOeFZI9XCor0HrsdXQ7Eyxd4iXcYcv5c4tgDZWgKMeCwmIRevooDNASGgvUEjP
TK9d62uxEApAD20ba3rt8B1rg8w/Sj6fTcnXWaXskOluEw/0Z6aI+X0nk98CCmzDF/N5V5HOQs89
fusxQ4qz4O3JV+VPmHTg666wDP17ht/mFcmb9+5ypKtSVvzImjr+VhG3bKv9TdJ331i+XWCXEeZx
JVnjC6WLZyOPVJjmmO60XjlcIPzAxG/veUKXavZdRZA1uM6U1GegjcCeN7Ob8i4HH4J5lhnBQ/VP
IdyKVasn+36TDsbZ8S6ZTWkwyBtOTcXQFVs+g+vX08/YroelnoYNh87OQr44+BhR5M8alRln8CRi
kG7vX5OAxGntWENywenpuT/qeu0BhBdXFHHS4TqJ4K+eBH7AC7PFmYkJFbM1tmrrBPC6kYtaDc8s
dBgJoA4zIJmGRR5tqx3nIMqndlj6ynZfXjtIF3vJbq3mlwrbQTFjmM8w+CquTo9GcrjOWl/mRp+Y
GA74vPIkTpKsGKDVZ5M73J/elCqvndrexRrUzwlZttMd3EZdc0Tr/DedmOOU85K7E+d8HXEQ0d64
c9aAiToAlQOvV+icXB3jwBFPsTMGYnHLUzMoSjxbEWTmSdm25H4qBRvfYwcLY4v09sy5A7FssI/m
HrNQtZtBZgpNb2BhGJuuMT4pASOtQ2WBrrI+RiNd5wrY8DlaRh+SCmYvFiMQYYe8paRXdGTD6RWB
10RYjQ/FEyXGvEJolBw2f2UGxwmDZHncXULBHAJI9qTrcKJ4S4MzSKhYE/s6le8jiq5N9L8qw3ck
E3KuOb5SSJ3ZJMYzXab464I5wWx9VnLWgZTHIkmlP45Pgs4HISTC/cZR8TFJFyUFpjDAxnprU4it
sWA3SQ7dR7f3F+/EQZomtFxWAO9Kt9UeZx7415N9Fv0ycfS9igjjK1Reagyd2IZ7T6hem5HW47sG
cws2NOUGvVDfs4mg+CAGb8cJffqee9maP6tkgbDG/cTxBNAUsrElw2VZvwXYW4Opjj8gOzJgGfrZ
2uwr0ZXS3MIFcvK3AR9vG1VRzTF2krAV+1sTHOaELlo771+huIGziQowaQidDQthnl5Jnmjvfegl
fzWxy3lHU9caFQYrHZtyFawfjVTZwDhC5S+c5yHK0y1cBIMgkqJIpoMrcmxtjBMyKdkZ3vjQCohZ
2BHdlF/Smln98Q+S4/DhJcWOs53lsFMvqucdRXLFPb5MpXkVjQcQSBdXvwY0UbFENCxVFb9P4XkP
UkBevcJVT0V/tvxjMK++RSipuKGuvvqnCviKJfeUgwcRs8mOjSpBhuZvi1jl/ovP1x5PP7MmDgVi
0p14ulypDW4LEzgbKysNhYYV0fiMzHwnvKU6KnO96pKCQHWds0qIKwIerIQPF1ln+Bv9Yhj4Ls2H
W1wrsP6UyxXVmr27ZlVhD/9pJIkiV2hvCys08atGxcqyCi4N51FkBYq9tI5d8rHdymK76DmQ6k7L
zwQujo+3WMlLhRVRKtbeWtMTNS4AOTSQHatYkCkjNGs9GP65iQqApq0hpuFWEAB8OzVFWPNg4Bdr
6Bfpb3/LcHBzKGXEJmHlrtJY/gQYPEmdbU1UWxRcV4Zz8ZgrGFySWVyjlZ49KhWBLqgODcUia8Df
kuXjWwzqoAA4c13mjOpKlfS8Nh9lS2MaDl06cfMK14Pix3JQSsKHBrhlp+YzqgF61oPnwrzxnQ7G
jvI5dB/4nlgDdgQJ0OotgGos7VmRyVXQtlC+fMBV6YRTwROsbkrHz8VdAAs7/WQnk7Dzxqb7SePP
d/nVtSsUw8sLFcykTP9T1dnr2V0CKcdPzjgROU9AEZC1rpiOkpSpZ/3lGubgcJl71Wp+i61S8247
1nUYlw6A7dPAGiO9nZ42fw6vNSdybgaReFY4lCLOVJ1hJTDPiH+DUWd86ZOQx95ecVs2QDlZf7hb
5b1WBEDRLwxEb3xkhLPAre4QkH1oenWWL12wxZoGI4lLs5wwhLuNb4lQwh48W099O/6s71kdfiUl
FQJis2fIbV0w1b480/rdmyrH7QnF4fLh0nq+Nh6y6dUlyjScaZoPCyLk06RZQJ9jtEf9BqKpEsd+
ywoPalTSrA/J7j8qJO8kr1Bohx9YX/rGLRGHqCRTvwTwoe/0fFMiIqxs73WMC5NmcKE4TbTM7QrF
G6wo/69UIJNoUyoFAscI2yr3ih96Di5SJ697tAaogSD8ivWw6plCEvc6t4HgvZ8VPTK84zhdLeRY
YeD7MXAT+NP2Jq6aCPhgdFnxwl0nB5awwdkZycYW89ZyNQ242cptKXpgZHL02oEVGwxisfXozlLl
4hvBkUFenjihFbbJnlYJ8rVDLz59Oeuea3INO5VxQhhHPLzQVtHq9/4jV2zUKI/+oL/THxI1BWXg
lx6i+8xZdmPehBwfrpkVGGtzTqfOnI5LEVNxdi86pD5pY9LvJpzXWIf/twgD/uU60ZxXa2fp2M4y
abXLYwgW9laTDFMeIXXQyB571HVd1lhQhFmQ0TGqkUezloXDGKqMASDhJs5+4LiVxFQvx0tNE/1r
2CRzFuhIPuwcmtK/cPzcxSegzVnmuXgb+h7gdfl+BmW31esJPjZHaGqianmJJKm0U+wDlYlQHtxw
eyyY8UPVPQeNe44EFvFLL6sNhbRA2HhDgmZXVZcj42ltQHkNrqZB0r2mo8OnkaV7H9KSOp+xfJfR
J+sB9jZbIbdlq6LwCJUS8847SUqQrX/yQeL0O4TTH3gfLWCvmVkXwpOFWku5ks3D5g21PLOPBDpf
VAbelLFWziOTI49e9axHvnY6qwgM0TsltUC0cLvveL435wOkVbELpDO9T2jTd4+pmhrPmB8yZyEJ
UBWI38QCIxfaQXgH3KO8gEBtuwC4BaGpjFgued329cSzMvnADyTO2T8IcPsghFHuSaNyvdeyAKM/
01EywXLDUTx2n2sxqBlkmQSvVN1cDSFYedaSAg5F+HPx9q1wB+1wdYm+7YfOTSXyu2UvCZiB+7px
rEKoBGmVxo2rp0UiEMG6fk4GBefQDMaDnOrfAyd9aijY6u4n8WzsxYGlZGDiG3M2BmeU3VITvW14
ZUsaJZsjjvqrwAOV0qdzZKWTGrKWHcoFEfaWRWHjqyjZnYvxxm2vKczPE2JyZAtPqkHmCo4XSoMw
u5fUA3OxQrt8DXuFDB3iVGzUQnvJXaAwURg8yGf5oAZcB+zdmIo99T4LY0gwI3k3h11wR7dT+1Ay
3+xVZAdggQ/R8rsEIbaqgFANpf5c+pteVl2OwN/v88pWsbF50XLi1lDRlZN3hvfY19xRCRswyJNQ
tCLlVH5PTb3eGCqdMxJLL7NreyNMOdS6/Fr7LDVC2rLjFV4Sabb5gKLTnUhIW1KxurnTlNo/YhX9
zipjGHHoa9yufjiqDOXtRfBwzp4bQE0iPNd0WTEVze8LFRYBSxlGb5wWAlEHaWNU4IEob2gZurvt
FEy8/KgkwThymoTsmnHAYjd4gguhoURTzLCErg9UmT0CnPsqeZVqRvYICZh92YDeiGXKFxJDR4GV
p3Mvmz9TbLnATXPeAHERiBvY3UCeXHDnH9Z+bpykT02cfIaLgUy3pL57D55+/6Mc1LGsT2Q+oqcf
IP36qdlI9U0mmwGshG7K1Eff6FQD76glUSpIJG9enXigRssyUr7ZkTfKnnNS/L4TwwFf3f2pihgZ
Kkk61kHQ+vTYSl5PMaPRGxXAiReJAkD4K0v+cE4b5PtCa9eKOoTPqWPDCuZMiWe8aTKe3fGqNqyc
Z4hWevN20DnaxSZNzdgSRL5v9sN/NO0v4N0nTLZcrxm+a3a6CUDbGyB2SLdwlNIX44DyM4SOOZLY
TbcNgP3PS3v/OoCPjwoENM5xSwA8AD3uZAgkcBELxN7xU2p04Tn7V6HIlC4Bc+UZwJEAnCdv3BU6
X/02Fo2ALwP/D2pIQrrvcOHxGd4iP9B9GEBnOC6Kpx8oZ+bXdNPl0SPyRYXry0OyKrrMns7024qz
DAFYxVjylHkp5J9iSjOJLlYSIlvfvo6DpjV4+cr4o6UujYLclYjT7h4cuZj367K4+LjkMFTQAzoJ
GhNQnEjN4/KN5h41A9qYniG15uicFAyk/jEL7+BNHO8GvQXziUySFsnO4Ac5mLPSp8iNC7CZVc4V
HzPqKpkE5SWm0890+LGFY9JWN0H+k+UXGTSgOUCeCLnTqyKzaCmDN3mX1tHOdOERGiufOBlPzNwB
ez6RfsF15vSAxwfoaVJf9v8NR0OmbwuVjPWl29Xnmnmzc2fYWsY/6RSrN1BKbTx+HCvkp6Es1u06
A2p5QAQMb1jqGoShwiF45jKolkHW8j4Wy8tLQnIKq6Mil4ezEqEQKlC3RG1jxv6SOcxknahsToq8
yYdJPDLUrWhYYGlwValUMpVxqotqoPFtEONCQNqln3V7V1PI01lcM7f6iCdrEt3+bJ9wsshGSyrP
K2J5mHNemN/VddG+QpoR6FYqBp8AgMp84wts4VyUCZzM4ilFPMgNTr4yTtCNNj0OPA6mGpNGBlfi
d/rEGz6IjqntjmkzjFPOJm6K1Vml2MdH1P3XMeH5HXW0S/lOjULhB/RffNpg406isDQ3pAOuMlXd
xU0x1avlGMs8TtGua1TZh/c7ku1kCju01RmeJFjSVnuVa3nX8/rpjx2rAtnwTTcPVgxjNrNiz7QV
6EM52I4whe4YnBlfoMUnOpU2O4BUcc58NMsa/AgB5uzhHPHUh+7fPia+SK2TW4dhvRKSnfjvMAX3
rBweSpJJ42pKv4DFhT8K92fhjrXMn4eJ13VZMrZeSOFlyhZ7ng2fQPzp2ingBST46K1yQteaN5qR
zWkyCEz8HaHRO7xwD27mg5CIok/4vNowoopvw0ouH7ttSEWfqghJ1vsJqFOSahTM4ewznMYygMxw
1FlEzJ4ARjU1M0VdKLRS2VokmxKzmZFdy2vsY/0WqAB/aAkzUY3Azx7R8OiWibaelkiuxneTU3UW
gP5wMDMjunGCfctyfBSgsolvOMOPRQpmJhTsMFDBkblLO7ph8JUB1f/r8cOIF4qA2+OP/1P8FXhw
FJJ5HruJ2rYdh63kXIa2HMjRDe5qoS1Bl2mJ0SUe3W2iQvREqL/0R1MkdBsdZlxqEouK5K2L6rnu
cYprL2A4nMGWsGGcUs0TRyq/dIlxX6ExqcbblHa/k6Nm2hXwDsf0BHl2lkK1FxrRIdMOJakX9mcz
bYmtsYuH5g34Y3PJkgKDDyVS384jekxbss8yCD5ZNa6c8sD8zvmn4W0rw9bM8lXwWlK4zgJAB2au
rxZ14gQ1huHTYproUsKJ8ZLb3ETnuao5EqL/5e4gWD1iOKhsC9ObiQD1/ii44TOtt3fzbMflUoXG
cDD5g14KeKYnHx/+/P2xu1zSBXYK2tCMPoPiK/BRZb0DWlrGXXGmunJ5kjWKTYW4iYSQnBSLh8ij
r+OHgabDTozLLe5rrCMzLU2aZcH8NAbvyU7yjazH/Ti3A85ExKJ7233yBpbjy4eFTZvhrx/O7pdk
p2SIMCLhTDNEd+eBGfTatRU8OAjkfUJrp1vdbM2wbJayY+pB4hDIPkgXy2V93n+Tziq+Ne5Th67v
L7UayFiHztr8tr3vg/DWgqxjfK8B6lwXtd+37xnWkEvs6+sCjpHlfk9PGvlgeSPkl+C5xqsNNdeb
7Xk8ctqKuZwKoZK2nqPq6bvmthDlZtCWH7YS2WMArrpnIFIp9rEwoPv9MaScRHNrKHyxhlnZTIJh
OfdPDjTwpksrIJJvzQw6HKiBt/QQhAuIoGDMQXka3ThiqTKXGUJv6yHM+uffsecasGzW85qb+aDT
1kvLaOIwly1/1mOKYogRBY2cvF5/wjP2POdiBXApSfjCOx8H2Ib/eOpseHtMLw70wgBIDJV4PFvX
etrCcNenUhsaAxl87teJH9sgor+GJq8CGfuoZkgIjxUqWrjA37HntDYymDbxoWBGWpqtwbO8gbrf
oSLPgOaksF9WAn1vF2q00tdnfzAKjIrBEvQkWw9r7a0UaSCk6Ej9GhU6DgiLae490H35JySsdpIz
X91In/GJz5VJKfptQEhTDTIDUFxXIgKFo0++R0EFok2/0h8ZILToi6+pZvzhQOj0hV8QOG6UXgQI
GWvTldI3YT3Xp20z6mOSxfMciKGmPTXjFq/Oh8U9eZ/i8tmRl7UYQMqIn2oEOu5zQZ4TzFth7FD1
y/4X1vVE4r+762LiMzXeO76QbLgcTAPgsj3s12W+xzneWMYvYn2ivJ9nk6O0iwnPsi7ApC0wNCF9
hkqAOhIHHKUVjRc35aJrEI5Swx+suCPPhgxHRU7G0sKXtH/7MiEygO1qnPrmWfF84XSYv8dGdIr7
Q0PfGjfqorSNOE/yUpLPZX5DhNhIIScNc7F+j0BLv8UHUugLkT1Cz2b9MEftFXN4tqhh+D+jX7P0
hHLiqm+WCedgh/i23szJyULVF81JkI/Y3B5VApeFnpex4cuKNR3cpFIQKSN/YBBWUYfYDmMeecIh
zSW7TUcNlEn04c0MbUBMdAnEHaHy+j4Z1/6rPnCjfZyyEdy8Rzuu60273XQGpZTD1FuO+D7sbEwJ
q0V7P15ux44MnjH6d9s0oDGFp8cVW9sxilbH5GHnnBAxKGMnAtjMsKjie8QaqTuOrkUmnDEuoHiY
BjRQC5Z9KEfqUfOpi0QNm9DUYWpN6vbmPbqdyIrVInnwXHkK6J/oHw/CA49iRLXW7lmSwC3IiTnZ
TpN0eZMbG9qPftTJJ9mqKvrf5KnKMAho3zofTY8/Q2dF47xKsKyx+Oan0dYJriBv8CKF59Flw70+
yTe6SG4Qcd9Adk/KbrXjklKLYVutLZFNCJfdApF2ZR3AB+H/p99+zQFssGphDxQ3T4NWZchbsfwa
RcyUTEV8E9Bdx4FWGTMeiAOmghvh5CzxlGMM4E/uZIeBakDoCujTN4LQBcHPTZyuyt4Mqxyba3Bm
3Gtu65Omk1h0cRjjkgYWBoFE3w/5prc0596ozqu7oLumMY/O1R9mClSE4dgcTNLHa16He5ES6QRw
eYeXfFuh3d7IRWHp+EFd69z8Oyy8aVo3DS+Ay7ezerSDk899tKAiTt3PjidclLN7E5LN/LGYYlTP
Une0ft7vekqUwzmU85J5muU7gAmyy1ePBQzS8J/uEcm0lhT/HxXxOS0Tx6tX6oeWhsB0q5vrCFJt
7ZnHl6rQd1viz/FbFYxW8lGz7r8jh/18JdZ58+P4RH+zzgGF6QB6W9FvUyKi4ysP+O3xRerkSlPa
gbscKRdFgFOXFjXuB5W7b4n5+I/GyWi5be3MtmJjvOHOdAS4VoCg7jHKT1PehEEUuIvmcpAfkEvN
gviqdwLPuuzDGSv5XSGruUml1AK7lHb9pJFsmOWdEm/neepBIycKxgsRw8r9YcDw03F/RFFgUH2o
7XsOVUGQ5vw/xR1b2N95zj0xXlFA+K0E951dChqDJzd+IKDlQ7RLZv8pRm5GgnUEfj2UDBV0PgiQ
sAxPNdhWt5M7ss226xwNjhD04NSKi9KuyT4qAxiy1xxnhvb4ZfHnarSgc1URL8qcUFzp5i17Pocp
y0thKGZumYVrozjT9wjndCMwCL2hNgru/3oyRrh0IpEaVoHWJSSPo30ASWqNPmRd5xAMg3Rc5Jx1
i+uCd8zBCOrOWit3oDjHQPmvUNIZP2JJMmbMh+4mA8iA9Ooaj379zv7rhtzV6dwWEmTHigjQQTwA
70FuMEDNbelWavebj/15VK8Ac7W26yI5h7uXYRtqKvykGnZTO5PQTmCPn/Xt9Y4G18rLeAIzBgjt
cLIuTs83Qa2m1YBhPBg6/y8jjl/uuleQRWTeP/GdQoEuyWwV0FpxOhUzyC2vZr3Z6ApJnxrWFDPR
OIBjd1Bm2GGhqHvYdXdpdf6TZ2NSCThuISx57fs+aY21TPGnUX7e7eqyQ1Z4QLSkJ/xo1O9PC+A7
vlXSV+fzKZ0/ny+ggh5sUTXVoAjxLHSi63LhSH2JUUiz+o5CNd44WjUTrwHN/dg9FzXIuOINc1Wn
Z0Ngae0qdv3H4DfCjO8bsm+Rhgi6831VoYImYvADYgpfi9+N19GxAN+cu6BAwUHltzXxCgZTzoo1
gYKoJl7eIO2qjqOvnM3TmV8iuLM3l7gXm30Vb47AHf7qJXxyYBI42q1Js4SZUTsIbYulf2zQ9uLB
sdAgcVeLjFPHatVCnUNLHGbVI6lMbZjxj8W60UfU9IIy9ikiMNv8jgdiw80O5DdZgbgUvdXl8q0+
92vKUDL99gc5URueCFs5vMXoSOwKgEGmbLytblf9kObXWAe2zf6N65eVX08zY0Qgu4UKL89e/RTF
MQlpRuWVmkArBNmGAQfgJNYdtqJp5ahgoIXS0/YdoKpjEO9/KUvyCpILYBjlbE36rijj+YEN3F2l
Gllr2T2FEAOBa+RDRaI2a2njiixWFY2A+36syWNU6OMFeNFxSo6J94vqQzsORU+vJfAfp+7/00BB
AZTPkWDBY660GrhsrIqx9xuG+dzq++2E9rEesvhQaQOUZcnxFWJlFY8glk8zXjldg0VYfGyTPYvI
k+5e4u/1Syd0MEZva5hLev0eNkAYR9Nsnu0njbtk1jY0XyiNizpoTE9zJMglnbzaID8bjvGhBxGx
MRBGhfpbxeXxk+Sk0dX+DZPZKVIYmQOyZ/vtE65EIN4NWMnWUDSbC6//WSzFIOg9zwKVxb4jsl9M
ulUvoUck+JpB7dtJ82FT/+XEzdS85YznZKJfeesJ7l8iIoWSDkZRV+oEpuC4kqyzHHGlIqtJ0m13
V8PCixZif3roghDiiGJqpNiw6kuJ5U7Fey/CqbDOacPp3T2KjpOFmsjowyY5wcbMHyZSjQzecjFa
hf2v0NjsrXrPLXqhJUHJjKp7HmVmMFUmmJXriDjTqVTnc5JaTLmcmtKoydnpsYiRqJjn+AJJlzuS
wkCU5ok+rw/rwXrUhJ32LBsrgUUKimhQOzKvpnw8on+SyqHIpczRvhZpzC5Gyp2GeRzKVyEpUzUu
lOS7bjLZ/BtHRDqCTLiihRZ7wSGixJh0d6Iojl3FwhBnqFQ6fySmfpsTeqK3sanweVawOqWjFqa3
IJIBomEiqm/b870/lREoYOq/q/GgPrgURmDm3flp7ZaeagVkSh3AXP1f6D7fuLXq79xu8JZT+lDk
tGhzUNbGhbawsGVYZKjqcp6mmbhJQoJTXAncMw38bFIUheiSr3iVsCIGKvCUWHRJpmrlkkjM4gLd
vnfZQtFsewS+cRBnPqJv57xP9Fg6UVY2Ohwy6WgfBDAKpbAyZLvJm+WH019vVq+xj7/aT1CwGqwn
PrFY7k2USP6V0qlT5CbbzAj0E7JsRhMMCxQSFLyNDo520h5pl89ko3G2SZtGkko+l3RKC9zTrgwU
U5vxTLrCMgBosKfL78CB/LZC7VLDJxrrU2zMhEWE3cH+Rl4Ar+KaLakdAbp/2ZZhdpr4GECJHxcW
YhUcWd5RT8CypNvO6Mk3yRIbu8iYuDODfQGrwFQCDhZHJHUKQdmxDxly+ILbUqTp6i3A5DRS1NwG
L6aiLjOEtTgoWIH2hE0hX0/x4GeMQvR1engqD/H4p+fkbsXb4rsDqbUo5OwXTVx5jLCQCWVAoi2F
zuHmWIeyKHTPnyxNYrX9XmC2uSzH4z0AEopT+N15hSepas4cXuz3BdF4u8VnrsV7jdPfb/YbIMTe
28fIjPRUH3HUqJb/3ieniobvDb+YfbkOIIsMB7adRUI2FgEc8BZhGUXVV7hAsz7n+pEKTwbZf3Tr
rOfRFLQROHc1EaEcgm42LTBANQgz/UIuFZ0glyEFdDzVQOx7UIE2nimvy0iQDAR2mGJntOpJqztO
Ea3Bvhn0WmPMTGsgz8Kl+KDGoHsVkcvD989UfD2LRn+Xw2tGlT+bN+N5Kcrk6GeBnC3NTcpkChDL
ohQaoLhJFvMktL18yHR4dXghhbekwu4NSJoVPKaGj3BpqcUE4qWJ8jyPDwxibUkYqxe3hXP+iPYp
IMSTqxMOSLHQSwdlEqTczgHlEuJxxh6ZZB5TM96G1cyoDNd79i09qnV78IIMFeQ40zNGTniC/3lB
NjZhOqdJCgGHJm5mWcnAeeBtRS+R3JiK5sdmjPW1oWktkt0NiDbZ5gXttijQx0455lgesquIKPR1
6GU+NiIfXckVVZJlsRjBV0viujmMbvRW+W5F6ItMv615tOauQFq2AVNnSu4/19bGKWrA/ycIZy6M
y00EiWjNgMC08kivUgebIK7jrHJz5vrqugUqMj2py5g83paM8DsC0ATj9eanfd1JEOyl18RxuH0D
t9hjftCcP51n2inpmV/ZJbMP8S3+mRORdeC3YofCIuS0M8PfrxCCAZfJi54Y1bZq2XNjAeqeP5Nm
lvCMvlSZ+r9Ywid5PGr96ded4+C9vgctQJ/cPnjkhAUAWhSS+tjGzYm/Rh6r+o3S5Aaj8vFYZHbj
J7dezUhjMQ2QCtfhqGFp2beWM5TkR1kMKIUEK7P2dZE+3WXLj8hKvJVeZuYokd+MdmRmNba5xXKO
7w2JQtWxTBVDoeDA41u1YWdgFAEC7d366+v8UCxXvJSY3iglwmZYBQPRQTzpQm8Qjk6O4klBmjKT
+tzIMhWdF2+gcAmNEegb9fRWOoaQaY1+WvkK3Qr+oDfOTTVinDad2ZOafUOKa/xgSpNJrQgcERKj
/0tlG6gaqTmf8MHFmEH7H5Wk/f9NXwOveMlH+9pc0JRKxj02S7SjoO9yocpmhxkVyzTqlrFGKP7h
JXOM7ppjBjlmg7vIikUkvM8GoE81W1Mo/3OmSYhlhJx0XULStIKbvoFJ7RG8XLo9QRba9Umyi4Ek
pZugUvB0AS1DFjJSNUcStbJzITSK2bj56ZAO4bslpcbHDDrDIOOhvU5BAu3Kbtoh859SSdQ23T7z
URNV/iatB/Y2aPXWK7mhmH64IelN9DlNRTjSodw0ssvrUn0ydhgUSloNo4eMsbZgJ/1ZoBH69SDd
PFE5dvIVFKBmdYjMIoWktkqPCvIoxFAu499cH7YuEBrstHdoVDNiFliW4oV8vofR2zo5Ql+zdegF
vnX9kzZfANsd8u/FT/e3hlX601M3nL5BamnC6iqfptemf2YJOoU7k5VFIuKTphYodAv9itNFqnjK
J2c/Q2tITWqEoKpltTnP4WmC1tAo0euchwQc0xFlPcnEcPFvDsRS3dT1zwFN0czhHTcxm6vjtE6o
AKahw7kE94soq09io99SL/GPb6pRT4GkmdOaZX7620yYdnGVMjtH81JJpFbFvrU4ew1iQbHSuGhs
Vodvscld/99k9YMaW1awGEygZ707N+oXbZKRyHgUxE3o9Yi98g10xu4nL20SV2/a54r2WzD7zRH5
W3TqQh/GZFmTfJ3zd4LEDAuNzSyzDRTNhpxLb7zx4pNSej3eogEnqCwTL+mkO4SAlinyyXV+WiDJ
zbYyhLel0e34/6O6PzKM9fuxFy/VBjnSxZ/1mPzMjjNTp3piyJpu2xO+Of/CR8A9c9r4JswDXIXp
SguxY5jaLIc6og1J8qEYsIPBIvA1Hq3GTnCITfrM8Fqw3jsSZCJqQoJVB0uwDLGP19Q5IebvzqKM
YdDTEeGJIbpLB+EFVkgmMJNF1De0YedqwAkfchyBQ+EXWaIoVNYF4b5FBKPantsG5zIB0vaG7Loy
KwhN3MVD6bbGljz/iS3Jm3Y9SxZVN2l55RbWVNbUK/nWCr+mR0grsZwANSpWAP+O4NIRCyKKHWL5
75d76mI02ydOzvyllyAPK8xt16Dk+5MFbuDue/BxK19qUZQpFgUv5ys2bnIDSMjSilyoqCusGjr/
4C22es8d70LVebZiZs7CldHxpKc1Oenh25Qzb4pKFtBRe52m8nV/DRL5j0DMbpowwwb26t6MBKK7
Tk8ZC2zUyr64luRMScqTGvxnxloYLB7BpDPrMAyB8na/s/tlYc9IDSBVgR1eOT/nfFqneQp978a4
RG4TAe9wRLD3MoRk4GETXDI8ACB+NF5Je5RO2GTIGCWr/nfU+7buRMMktHSoqntKde9/eIP9KeRs
gmLDnThVgXuE3xlaniAp2XrnqOQS0hRU6bObHSezZbXAI8PhgadcAvJ7zVll0rNf3Tm50lJXC+EJ
eWWIDATixXCXzUlSacDJE+sBqGT/b2Do5oKkO4PCOKYbNzTJYYqItbWTqjFvk2wr07vOfqudCxWA
gKpvfUnqLIgwZfhmQzyrpOjP1YtiAHTF46Gy64+Y/ikbWY9NTQsIBri1Tv+MuFHz5ZjbaZZvPa9u
C21wv3Yg9s8aMwd73sHfkKeP5Dzi7RDNcEJt9pCooJFth41Q8k9dCFEllY/r7BVc8l3Rl7+Osav5
C661oUA1hIZN5LAq1h0nVbVxL2TH+Gk64nP9fxkasBA37PaZpjU38B50/oMgD+K+jQmxf62VD1wj
/knsNyyeLfX2A3/BPAYlR/BLcCItdrri3Knl1min04k+60besC0GYP3QFCWeghM3nAotSe8O9BRp
wBIUTg7axXdEd/LxaRPw3FpH3bLMYiW3FosFzmW44pvmQyUzg0MnURMbw6IWFitnklnaOBslO12W
kR10PlIdixm/DmO+8u237XmJPEh9QHRerbohL0o6viDOAPfDrFV4/x24Z/YUhoKJszmLhWiLSjJS
GhSy6RC0bKei6ab4u6LjB1zk6zixoewTf1sZokdvBj4vDtnefm5nzZNL/4gVTrtg2c7wIvCwsC/j
v+wZ/FPn9iChJqwjMjoUdUKNFcLn402Uy/NNTkNnBDCWNCrt5mXDrzsm7CEulxRTvBahiExUO0yx
yBj9imh3Terga+o7qcZugcxD2aM31dgwj+djZmoO3xQeyPuqpHrYNcpLJIqz6TjqMd4qM+rZuooc
jtMzVmzRa/qv+7k8UyMOI2xvSjiH8TtxAV+Vc7Q+UL2cpqr15apkH58ttHJOEgw0IHkiuIziZHY2
NiNPZsjf9Oh/V4QlaK+LOcoaKm2Kbk8ocX/a59IKTcPmKLOJIbBDsRajuI6g7zBgWymGmA0dgjKz
ev97zdvRbizunBf3JQWs6fT7FTrOFJpqwr3qcy2Eb1dybkxIQbWwfiUoAGP8tDIdSzDyICs8Vzm6
K3GRZkzV1wglNYIyYW/Pc0CulQfPUW1v+6s42xqi9VNXzJVRWIX1myduYjSWgJtM2POl6QEEo7mf
EsDDzdrcPDucJiV3UTa5CaX+jlIkTs3Y2cyVJEpz8dZfFa+lMQf9v9kr8+otINuqcCnubBSDXIjF
6z/6hWaGUp3N8Y2Plu3NAF5ziAV45QM7ODorw9dt3FOh5vh4mJnwmt0ESm8EdMfOGFRpwW8Sd+97
OSZdOPvdI2eSm33ykstjIL4qvXVg3oldy6D5FHcjYnbE4Qz3CtnfDarwJdS+9YURymM/VItH1+lH
+pV8z6/ErNzAxIJaMh/L0SSfnkR6obhupKIf0r5tzRly3OPCJ0ei6nHv9qnK3lwgzF4ilvhhLfr5
IerAI80CrVUzLi0zlOvW1lqqUq763mMv2RoEUcek91PfXKXzvT9/2bdcEpOyLmgXRIMXeqnvOpzF
kczr4YW3yjvPtyFXZoyxYOiaBocSnHVEekqawbcdPMAgF6RU6uUDrZoN0xYrMnYB0tVJ5xDEXrVw
zq03KrY4yDlwNOW/1Ew11Lh1fZ3DmSzeEjtzYSlsp+ltAewajHzJG71md2iYbNDnV1Q5P1/X1aR4
Bfxx6rjnDthn/pzzta0LPsZ75KUSmGKqZZq/yWowplEckoeYE0dxJQTpJjC32N70f4cwaHVOWZC/
bCMXsQnL9sJ4TAMLoQ9ZfagDYe5QKuhJZQQrJAt0NmOmEQQMiBkJlygd1vM+msKcrC/el14PmLki
vNC0T1C3hC7SFwbzYJO09e4dNnIelLE+VDMFrhiZyuaRBfQR5B2Wo63wRqjSR62VxqgvIMrSxMLL
QQJ5U25iorKBfuSosaJMyzfb393VwFBjm6KDAk7CDNtztl0gPuIeYyO921EE0g8AMWGHiTFquM+7
jpGmZnn6L6ElJKeJ9aY8T4Bzxq0snwn1/upurbCSsJfIgYyMWRo1+s0kjTvntCmKPPEhWBnI3zWn
lyHKWBWWrLLiM63KZ5ioFV4LPQv8/Y+lRAGp1du9OPeR4rhsKtoNly1ff6rz4SHsLYYirZcVEcCl
Z4ObQXsKdjVFmTeGVWe7irEbiXQbUoHHRa4vXJCtMkymqUB0RtPRAUeqnAu0PdVv0nv0umiiyYjj
/yQh01ArA/6O3vJ7Uq1NFo/j9RfPRHuqcR+zrnpSK8of6EZMCmR2cvI88enMKUI/Bd7I9mH9g0k2
rw/CGvf+bUNUrnnjFKn3BwzrqQP7FyfP5zIR5YHRBWAwh6D8+pBajMvo7s0cdZa3va51iK397yCO
gdGpN8xT95YbmzMlytvNu+8dPcUxo4sdSP263oOnaQ/sJGk9cBNdda7aF/YbgkNLSXmcI6xJc8sv
qsKsuMFp+ugAUzONW/zc9KTDYdv4mMCBGE7aCwDfLbqy7Vz9ND8g4bVnB0jBvZ0p8NyVt2rGgaUg
dsaC3Cr/P9dvLO//FHafJa2lzKGfuKVE+FTunZ3RPy+owsoNRQaxVK3CFl61OqQeTeMDalF1GwEq
N15wFXCPf0QE4NS/O3S9TMaWN+FHCXzBh3dlDDff/4VzoFxHRwUrVZmNJkoS19m5AgTkKQ1y4Ad3
VwkbVrvTljWO3NSbS3i40Pux7HoRnY3jIOvk8ReFsLgJy2PZd9V3Hp9TdLGOxdbUk18EdXy0WqLR
GUi00De3FhGRi3abho+hRDIanz2Ss+PVRiG/nVn34qRoXbRSWW9JkSyAzJldLdXSCuEz4kbqFIR+
ijoFHHDRpAV+2OdWBGjpa1lOUYAyoRKdg7AZWeZMFhQoiB9ygbzq93ayOyULNbUF+u+ZoLIwRaRz
tJtNdgvufOS8prNfse1NFn84pbs74QBd8r+7KSFWGnKQQMdx63nN+iEsVniuF/2mm0Pj0cgPDo1V
afFacYc6wUfZFCnnV6+FHbgxbIE1g0dwTBkwydqXL1PCIXU/H6owWzlvjNm/3kHN8fbiPtLziDtR
Qcg3haRBfL1u5rbA/9pNbugT1OmiAFQQvS5jVnEKZP63woBnS42mXXZiPoK4oMnkEH7Z2VopJCrL
paf5wztp5dh8JP7+t3gSrUPkeTzalGh8qIhp2I30Xc6IoBGyYJBJ2fwrdvFpd7gpoE+bhW2TAO3j
VLb3oLUCB0GSUwAnuk1ECNYH0Rxu2hncqxVWARKSg6kOlzRam9WRBQHWUvuJeRfsuNvvz/yqPoZC
ZlbP0/otjBv//AT/FhpJ6DQdgixcKaam4jHktqS7Enh+uWbp64oslUTFx5LnQ3hXGhS9uyTBMxfK
VP1x0BQh8+DC+ZktwUN29qxciuXt1kxt7VX70uB4dorq078iEmM6Zq0hjM3HugtFhtSLMQAvQfW8
5ij4xzGGrxQzjkIzzOyyZpd5UO4EgrrBOhdoeYeIRyUz0Dum1SNKXcTHTBLwjdZAmG79mSYJHRKZ
lWxnSWkMA+INNM32fgcxKS3egH0JQk6pbZa+kEIQt7yOS9lupHk5ngv87+ms0rIHDbLn8src5zTe
min9cUY6ow0HclcIYdYcuaKRQ/FnV+SPa69V4r6bLqEyuybG2lsrhVvBdzUgIzj/YZhqDQYnRrjN
2+5o9fHppL06P3oBaEBK6K4qRxPbzvpiES6Whar/HMODJE2fxZ+9YRw8GX39gHBLGFSePH1txNN9
nY9c/QBt0dYK6cSkzrHY4j/BVKVtckDpNjWPQnZGYJGwAy3MNjv6iSWORtjX3CBK+AbAVJ4tm/w7
BGoyRM4Ubn+2pgAIunAITrW6LX7OtWRDvkDp95mc+1SmPlpryVgvbIAwmhIximGPPLQa7Iq1d2kZ
EBQF4PJxbgx+hBVG4yE2ai1DITLjpArUNWp1B6t1zt3njXlDYeXkPmWKVZ/AWJBY/cVPpoLv6iwO
ZG9q23zfGsSdVbn6grSkv7ls4d4RkswvIZNWP9KfIarN2D2jHP8PJACrI0pVJH05MQ/M/tOGUq1+
q1FL1s+tvXukukuCaUX9UvCQRZWHcxpya5pIsZYFfTcEknEJ4lvpp8ie8tmqhYrdAJDgddiB2GPy
i6YKNrmFlig4plBns7btWeDsp/SE/PRuyPEstRtXZslUDnQDGoKm6zmJ2yu4vwxrXfItjNFjOvpn
5T9bDTSbdd5Jhm9D0L90T4GgjevYGDsExlV+Lh0JAra62E2Qiy0XD88lDr+iiWS9OklKq0Pg0JIk
OEbH/LPxZsiIO8X2kwIckFzuk7jp4WcztFPGWD/V8PIj2XcbGXgPbJ1rzgJtW/VydjS2VRlcu8Ss
d6MU+rb7D4Gf3ciHV242RaV3iFABYQ1UUVgHtBsrasFTdLzxJEygUbIjjXMKyKybyVS+SEuWrvMW
RqWYUfoWIgjdDAYr5CCjqG7BnYXMFcppTR7NRtGpfgeaIL4ulSZX4JdPz7wwdhZL3HXuPAMFjcF1
YRLS8YpRbqRjERditQii6pH3HDKoq9KkKHEQhEOJbAVLbAgP1u6XOsJ3RPil4pw7vZ1vLu0KOoYm
qCwo09NxETQLtjxukfFiTSmPaWeGD85pNYGraCDnbp6ECk/mdOZKHSDCiuHNmt0JP+WHlnlbxxyy
ziLliflMRBgyTO7BBuxjluZqZYdJkxU1HyOtRIhd9mxURPOVSK8rEx5+fQ87xCFvLPy2lS6I8L0c
FsxwUNN5OETRLMNMuCUUBTeOjIUKzeVooNpa1uX3ImyEM9lN9XKZMEIlSvP0BnYY00oabsyEh0sj
+K5Vx4CLLBCzDyWl0DTdvfo0vxJ7lQ4dlUGftWq7o8jf/+MWWS4HakfZt4zIjiqirbaT/8rfX/2D
tkSb7skUgZBEtFk1tTXfI1POlE4VGpbCQ/mkJglZOrUIU7b0+hRhcee1tbQxrfz+O1eVdxoHePyG
k2wSig2FIDwPQzPGUDx05mUV4+j4ae7FaODFBYaUTBe6JydGFN9xKLQQWirusGGOGNNR/QLgDMf3
eWwzInCZnioMVAMN0G8XZ/NF22ajq7vAU7rQCjvU6C7MvTKk5TlDvDyWuWew2FWw8V/7QkgFBg6y
wzcx55XgBdd5szFZ+Yt2+bJ22oYp15Ds3YLiKwEW67OIhfuN7VLcyMuVAwywfEkoENnpKSIs3/2y
L6QyPlmYmb7+x+sNYae0SxZpRkWlOZsOEtDIuDL22i8JpoDFNR7w1j9hRIwujcYkbiH+Ciq7zfYy
mSb8Y2hoSAjW2hAv+5v/sSsiah8K7Ji4w/INYjrplDfyy90gvWVPnnePcVD7SjAqMLHLwRW7Ma1z
W03/3WFppYu5lQJRaXJ7PSL0i0xdXk8uW8ge8XuwiGUm3trqU8s7R9H93n4bXge3ulVDyQxiNZJT
jKRH38iIEeTae+ie2AyJ33WWDjphCH8KYjeZnpEmTSmtwmP5TNRzVecntVC5VbQM8wFgs5RtSC6G
Vl48AI0dhrZTAtcPx+v982Qg59G+C4kEBOzyoSBrJAEH5A3zGrRSRXvUVQGNERwF8i8+MlYyOkdp
xZwOhqBCmqI2kgoGIm8hppGX1MbW5T/TY54I9uP8J0jm+iyW8laEscjpfuZ6sx0oA5hpeF/lXODQ
RXgY+QqHmC5kzXrhkXgM+XdcrnVEqSaH1BwyUB7F96iObBJjfQgDznIHCD9J4Ydbg4WbdgERl7eH
R852+Ya6E0UoV1qxCt2m0pnPomn4Ulov5vn5vQsI2M6tgG+kYu26RaauA88GJn422tPYKBKa/8uH
aJfs03UMlSgypZ3nOIKhuRhJqQlXgA4IGyD3qJF0sl1z5x9H6Nq4FAzrYYw21JYzNU8ktyz3+a5o
q/DmZgyyyLZYTLRy0Us3OCiP5po6L1rqSNMQrPSTVyJUkWclZMlmmY9UKN+06G8fS6kQ41i7sQNM
94+tfAoKl8M8QHpylkit+LWDXLdhHXkkMvyaDxbvCiDmrviNF+mB0HxtjB5cC40AkJou4BCoyJzk
k5npUBO96wepbOwYr7iDUkK/tHUeKxjLMIUMM91DjeOHX2AT/lKIJuR7AtGHOFKqDBBNTduyruvB
HDNxnJ0Ew9e+1FcG8bkLc7F4aHBPIZv+w9SJVtyiXufJk1FUKd/V0mFyy31AUrvzMANeLZ57qquL
RupNkZwqUxz9kkQqVJI5Q00189MomQAqHfIArD//8YqsIBBpej+NyiC7e322j7cPfmExDuy1aoqX
W4nmJcbpgbPd4r63jlaKTqBZZS4u9erACFjg4ANYFC6vNUQhA3FSfMbfbKvJ8bb+zdGs2p3VKC6K
phTgddZJtKMecl49M78QsMYNM5A9l3HwL4m1hPonStbKt1HyYEUbZZZGua5LKWq7CCanQsHxHGal
7/xG+h7uieJnD3Qb6S74MSl8r9YNM1ddcp5FsPRZWPx0XTgdD7c1luRE0G1o/jp1M/82rNx0uTDq
N+qWh6ltGGtiK7nVY0MBmkgsr44FIT51vUev6nDegvf8poyXk1Nz/vnSz0DKl9s3dB47tIJj+u9y
IaEnQJrO7nvqGFbHMZd+W7lnnnd3EJkPSRLzieESRgNUy9jZJsv/C0szt5gifRvHJRJ/XDgB8kSb
FjJUZps13yP0IWx7B/3rZdpSMiN/T3Jhxj7wfJG7pINdiPoYcl+v6dRj2BuAZBQmGOmiC8kQAhpw
RRqmqlCuZ5JGuCunDoHOfkFhdBrW4qnAn/evLpwcjPkXq9A9LSiGqPaphFtn17UWnDhWyr0s76eP
ex+k2loCZwX3qblrHMvYzcStZgLQlexRTUrMI1DVWenUWnEP6K8SaXc99SX/NQAqKq5zfGqZZDKs
f6+Um5vT1XcrZ7lQZn/8rUPa8plVBK0nktiotuqoJhY9kC0L4ldeev8LFAcpYTN1Hgldn5llFa3S
pRIDIv79cu03lgU9peicqCWo0gzHy+YYktVCjDltpeM4lrQ6x2VWheq42gNMlk+wXrlAORzvOUb8
/yib9xcczUXdwaWeGlPHCalGUIMdhhum49rQ0+HAK2Uuu/Dupzc6lMbuSXtmZyKsyYQ7MvIusEDP
HnlTAanl4a4fWMZU2JoD0U/B2Li8kR62Ah0oYGtA7NGVnNy1SXAIFG50VuMErjfcBrTbClclQvzJ
T0yg9VpTyNwUgPu5QeMq2mrD5mz5Nm3kUXFbOOqa7kqmxHvZ2WkySqT2Gl8OR6weCko7zvV2ttxE
pHT/JIeziDUo/E7ZDPXV198vgc/+NQ/B9ZLdSCxukOZQLgpnBkozw96il86mF/8hVr9Cm4iEnLfc
U2EoamOw2jcbBTY5uWxQZW2yDSM2q0BWiy2e1iAm99M+BsX0YY/JwEkJl7TG/hoIrAaFGKzzOt+c
R/NdYLCOcTuAY4XfJ/o2/5n1vtJ83z6F03MfmKGSwQqTnSEsH92mybtrHAY3w5Jb6yveJX3wDjFa
M5fjNylQTXhcIiaVKIFulSVSAMTTn7IohloK96f++kILh5Dm2EmR0MrcsTwtiWx3Jd70rm/9Nqg9
gcVMV3uZmUUdQji4uTK47FPLQMS3xCOPDOMyAaG2D55tYK77kmCJ5xgjZkasx71ZDjWup2iD1VG4
fap5VWkarl9/81Sa3lugPCfW/4geTWD6A2wj1Fwv+G3/78ZLEroFThd2g0UfNhZqyon9tKuacuUh
pzzOKxiQbyYOveFMhOjqNyjwEFrloE8y2SEwOZTy40/UvfzVshVOuDsMpn3Z422qQu3fcCIOC/tu
+G/nKNXgyw9XQT2Hg81W33Ce0DNKBfMOTYDbgUx5fybmYVJw6HkRkG/S+jVjv/xSbZpzOrP6PQde
kFFPfgOQAULH/r5kmf06u372OVfcx8XlaKqpM9eYwGrCOx5nJ0Cz+UTWxHJpscprbVAVASK+ow89
ntoDqkNYnoDeJ7RDNXWHIcRka5x/ismjhukGoC9dMZfHXmxVYnUXeY4rEWgkAYU9pgms3G8DHITq
g7XqVZzxc8p5Ya7TB2sMce/36laSLmJ95HJXjBJmRV7gbfs7VBwOinl6pq9jUXFK7QmAjsR4fHaa
tRKFt9QQ58pfoow3KHvAi3z0POTeAkRB5WuuHXonIN/pzj2ple3W2kfyQD1cbuksuKXFViWcDf/X
En1ycv0RmgBxowtn6IASjaKJVXSgWtuSY3LpnUzGMU1V/+yMVxjGo5ASq+eHULaUGk0PN+kJeJD9
woNIpab6C++KMCAKDEDf/gjcuno5H1FSk7BQKUV0HdXIqIvj1nG65rpcjkSv+CZ+TVS5TF8cMkNp
grAJfNX3xgVeP2YvGRqksJ9D6/gkkxbCvgNPkaWQlbWrrf5+rQxmqBk1Sane2uEXdG6BW9Wd5Rz+
PXLRoz0JsQknguoVFAC+9bzV6f+4NO18JQTR4Drs8fYgcsDqFBuKwundNcwhb+rsk2sF5lWtE13G
WvN5pMvPBJghh4PPadNT3EZLs4AUXAp7OKllrA2Ac4n1Oc2HYkQzN+1HmLtz07Z8GY7eXtckV2wu
1Cr4/yGUIzoDDttupMATt0oAko2KeYykQGjQDZba2zRdbEpadNz2yL+dnL0479R4Pzbg+HsfM6R6
V3ompm0vMqdVK+MqLe4W6FIHVgZYhuDBpOtXPWCD7FT/FC4LmVBOO/OXbHKkPUUVc6Qb0z0MWGhk
zkF7zkUN/h6tU2DlRsHTdeaKj8ImeqZgfl6qDS+QH4XAdvndX1X8XSG8xXPP7X4gxCDlnZlDVC1C
FSVEyCysR1VBpp3QuC0v61MJfS4a5r6UouxwkBhC03XiQF9NAg/nQSug9woRBzy3pCz3ngfrpf+r
0+KhkmQ2qW8VANZIRmEkopr3RYc8FF/OWc0/EOeflALMBRHXnymAXYbU0piDI9kFl23uQFYRe1I4
xRMO0ry1FrP3xlxk2jgvXoWOkSYZw+RXG6KY2jxIoMHajr2lilXh6OnZBkoCq/I/OspoH5Tx+XlE
Y0OMIb+4nsT54dlclWAL2b2t8ehKp1QJOBh3szch8XTxaUsXLUnzxu8Hyht53o6Aj+8se+KHT2IZ
iwFJkl8l/ZOjKygUW43W4pEQ57OB+D8zcoysIgJzStrGqblMw7DbjDn8fRULt7KdzZnxo0Wx8YhV
5wY6cS9qveqQQltavDnJ0qWEgp6PzqOZsEUynZOSGeOF4c0GB6n5MehkfYbxOiGz7sNWO+Do/zDb
oUvsk/augaFaJEPa1UWXDIlI+ZJs2VnUCUHt0fE+Id1pMu+l1CZieHwnZPLGcbVL41aD776udqm0
cRmsKgMn04Grp6AHlABgYf5O8lO0VCKYCbbr+08s5aULISuzlOSGo9dJbEdnxVJ346ogBdv7N6Ll
eiLOLxqtoImwlN8rsII2kUnwGJMwSbMMgua9b44gsOq1ajqq8oHpx0Ru0aJmo2bzoQcrsk7KZTLB
Pw5BfFDRULiziLDLhn1bTDNPTMXKDaZxdoHfyuXFhvHf3sclEEFJVlJwsT1+/p9760l8BQrwJoRH
7ot0NCffH+iksPR7/ewL2ManX+TrGi0iUQsY+92PnK+vxNMmbkj0l1nOzohHn8I34sy/RO2Ticp+
tToKIkcz/3bi9iCUBvba6kAGmFAExpW7wK571Fqi7TXxTH6SmEOAyWej60ZRt3GTku4eOWmwAL7n
izKxenj7VtY0dJySqdqq9hqIH2/Cp60fGy6xG6HYB/rezCCv6UJzinMgER50dw9Uw7n7dDuKM6YH
4/tBb1uR60LIUib+FPnWi7j/EL0kRvDDW10meobfi5FvUi/XQ0fmLmrn1sgQHJLWVt1D+oxwm6x6
qr10zWp1sUy5FjXaBAmF2Z+9wXHoSzmTaecPOeuVRFXC6L1+4vWMkvi53/DJsqlINxTU6DDM54FT
PNUu6vbelTIMqgswhlb7/B6qnITpxQqW/iDUA9aRYCptxn7Dvy8DC5xWAJl04E/R/eLdFezbICOF
H7SkfvMySuTHZzpoQYUY3AZUuojN6PnjikYIJ28XDLBmy+Q0INUMCENSeIJq9Iq0Ip/O7OLg8el2
NeTZBnI4xW0+CXuNvd2YVBNZGqbNNgKKwZK1rc3h2pRTg49dQoLkopm7caSVpxzZCMg+nwW1bD3f
Mpu5SA1Ih61R1YxNq1/uBaDMYp2NtWcbkw0cc5C1S983IULbT81ZDonzHLaWUYyi4FFzVvymeyej
QHeYzAc6FPXx7Q/vNuh1DPphP7LfEvuCw5y0hTi46Ge5RDqfrybcqT5BD2YxYaihPHDjfZ5aKkBd
/+LoDWqLby7zZZXi2JOYRAQrnlKRS936S06hyK/gsev5Gp4oOq0aRaxMrxzoeBwMdmeMxzyKi1ow
Rclz1j6+79KVPdInRnkyhFQ+ViASLnPCA3i1KG3MPlB3UqsknmD6IUpiccrz8AYXLSEpKLcHNvQR
TVsTaGvBXd5b++v6cCo7SKTcVhytzu8wISKEYSCd/j0U7q9j5OxH0VcERWXeG1EgUmNUACBKI1pr
kgyap5Obak09goj4r8ymYz/l4hZl/qkGRwLUBwepw0FJ3S6ocxoaj7IobKP18iGzAqv/7lyXrWc1
7GDWfhkflcy2IcmnjX6rh/HNVJNkqFYz66HAHjaBsKzqHxbN3AnAr3en5O3cGSxoyifRe+DlSItW
4eINIksd4vp6SnljBr3I5+ySd+KbWYFEyEmF3/qe4hHVz3nWyjESk1IkDh4IFHXA7AD1NU1g095M
tv/RbhNlNeeVf5qecLTcNjea/Zkv7zUGalEieaj1haPv5eleCaouNaZo+/D4SsoQNpLhM/qZJMfy
czLRro5SC1xBQdjQqn46snDMxaAuzgm14b68FxZX4YsiGD3BlyP5/jHUHl1af/4HTldYEGjO8KYG
HAvrPJB8ogzGZTYULqesUlkJgRoQAHEWMPR6vpBSk6orgcEN1eaTgsVNNah4qctrWH1KZZH7PvM8
e2SS52YPuqPFSyAoabvpkFEqaY0JZd4+xvd0XdD/synqP2ESFQOigykqVjATDH3jNOLbRBjrzkyI
YCU5Ru1XXxSnirp7dqEbSS40r1ur6UYPDTa+dc9c61d2xijIfkhtCB7PqqvD0ROR3cGepSLoF+Hf
PfhkJPeCdt+WMLdf+m6jSG4CZMU7iAlkA5FyKIMdr2G8vOz+0jGeE+9ZeiXHS3CZ2JIJTRwliS9U
Qd/bf+Uw4GgQYjObC+mGhLN8gXS4pIYjoPaISY+dMt0V3w2NZq4Ej0EDB/sYLTuba7/K5pIfr/Rh
UE5pAisgHFaNgn3CpvCUwQc3hRhplcLTiitlZIhMz9WD6uwSckIpiRQOIJy+gPAjhy9l40DkBWxi
eBbg0KCa/JEwcg4JslzvkDMcu/dp7Db13H0Ps6WmyD8gncuKrHqL2vpmbYiczFKTjqD5G8pSko6H
zgb5YEgts4eV+yNbPXshsvrlS9LHQoFUvObPIw0Q4WlsciJhCNZUAE+G4Um8a8bV50+VRvqvI5Xf
1ykm7Sv19YE5Ksy15ORHVR8ARNRyAp+wIiXIB0If8lRZ5n/bA/AlCCurMZEwXyw+5u7vITf7PJ4e
qd+zEnXgYibYHFjEzGDyB4ub0IoPBVXprKkCsajYmATQXmJp6X7biHXFPPuJJxaynyYzQqGpn18l
JxfuCtxSbeMlkPQK8o/gBS1jzx5I3kgCsSqOupznj1HFDq1m0z27jJQiNecY2lv7W0Zuno4UsG0u
lVHn/jLAVrJ87g4qsHcPqILNHxhRX5m/EEkcFYqDVREbA3OM7jlforrbS6TETKBO5RJiI8xCIjy7
1THojmQNO0PE9aUaEAOxZ/tg/oBt2QE27jIU+z29zgdgS1KuTyLkDQcBKC3Ht3Wp7TPkBXPM4M1g
6xu0wBGZxCHo/ix2oWachRaPcK3svfDmT7jmNfIWCoCpVXHmyItjSc5FE11pTGcyej8JLMsUZBRu
Ca4o39TPo/dR+cHCpV9z6BZG5s9Vf/YTX/l94wP94a3gDfY6niQEv6ZE4z/bdGhFldt3DbxCVmv1
PhvB1FZyM9T20eYM1bSFRUZXUSqabUtoj0ff09fgSJTs1eQm62QQ469w2KtBKwo/JFdIVf1cCZ0b
xK9n1w5SKpK49c5I8s8TVt8EnzuZ89gQ0NGjuy4k2vrWodW3S8XS3cOPKd9BVNaTm+uNGOxVbpzv
vqniRXG6JofVVbnS1NghT6BluCimkBDJSUKCp0JmZ4u6F4Am8AgbS2ST/GPGgUHUWgx5JFLfCDf3
7kvsTq9AK5M8zxoEeUVM5++bm6Nff6ny9sfPiBHVKPjARZ2VlBLQmcYAecxYnSvS/9ePcHSINMTW
xP1EEM4Yio1WeUWFloMRtRzeDQMZKBXpf/goIYs/OgEEN8WsKCaZDVek6arubKyHKnzC1qI2gp3B
WWZ9cE2q/ljaAYIC1BCb5IPLP8Q5guOzeQ4hR6bfkDwvkf97TO6jP9PRsKIQ0bR3IeU35gg7fnly
jZot6Qq+Rbuf0sPsGPVCwplOlH9mnp2zTVaP9LI4tVXlGAAVb0yKtBQraC/UVPC6dxtZYhhLW3ZJ
kN5Fnb0D1ahjYJhxoIhdzClgCs1TDehCmUiqldtmt6jf1Tz5zMNjzce6ewyl1Lyde7ngdsnF7+B+
+YqYXDVunDZc25Rppqp+k6ttJ9Enek04KqyRQ5+A0imJ9Nyd30VkYc6aBLzeJsuyLfcyImG9cocu
wUkPDxADnVBGKszg2hLBnG6MjGDUjer994KpICffDYd2CiE+UwCE6aNZBqAMWKRAtvk+Fg/2Xvot
QtRARh+j8Kd4WLgm7uXKBQfrg9eRoRU1XmYTbQgwJAzq3WzYXi0/IjPF4UblYV7LLKxdDDMbC/ei
KVw3fDF43okZrMdXJrWBbhGefBJcUXeN4F6p7LJ1e5tt+E/PM765UEAl6Dn2gfNxrSarguncY0F5
6fj/swcTbk1NUxX8pXg6Ewy22fizj/x32sds+9iIPwpsekmASCwzRUHOufy7gGMkWciGy/FyjLRB
fUnjelZqMkuxzCqq3cqJeJco5VcnIHayN8NJe5dTQh7K9PI8BfvIDPkb65DEJ7/PbLAufXqKPCXt
NW6Yy2dUy5cQpPKkSXtHpZGMU/M4HkINMWKF7IGiYlWA52+sYRuhxCI4Mtl0t7lbta6EelAVZxGG
/8h0iKLPdc/9CWnbZYjSzCBtZbKXlkv5D1fuUVUCxIJ6eiTUunlaD+UQOnyWhVdCd6Y2tJ1jY/Si
yFYRDphpFxrVMh5voYM1L++qbaPola2oI02U1/BGm/3R81u3Ndhy6SYdUrUh68yQVLmSQSSK5c+u
dcxHgB/nc29td3V8IyayvZWLd89UCmH4QnhSLmViRe4W/bZODRS4gjUYpkTloOkECrzWFWGxzGFu
7ZTEie6xrvewMHODP5cjddczGJBE0AAOHfrMayC3ZzQfRKh6BP3a4L37G2Y3wtA+K9tLAbyQ/+OT
FwiX9ZCUbCxYfjiTCF5yL5oHBq819jtcRWSfPjVAc4Q6ZTfLkolFJ8uJO+RN3eabzCksnPD7QH0T
KqOHf/ofim32oA2PL4kpJ6GgsmzXpiWbW//K9DAwzSeg7vkjLLKsvX75RGoqYVkmnWdndpO3mQEq
c7IWP6jAKmGU5QQB3bRoPCNQ9WYr5nVbDBLiOK5XP97DJY3ZW6kOdfEb5nk+br2/gjlU7uvvMNOw
eaXYOChJRYTZ84+u1Ap9PTioBiydSs8aIlrN61fMnUaRqsxfe397h7+5XvvlJJEXwxWFC8hb7ixL
sNfmuJCcDQX3QUGzYzNrvOiFEq0t4+jeQxhCgHuiFeCH8g7KrlRfGk+LlvCgpvlhih+/w8+/o6v2
MGKUYLv4rD+IVYVL/FRK882Xr4m2JPSYQSLAQSf2tPCDPgC09DxvQ0iPxQ5G6EViG2fkaTnOE1oQ
hDuX75KN7z0Fr9Y0ZxyKVFCFsf9GVVOcLgrnL18zuntZN82o9E+JjOA+fLRKxbPZbpMivk2DfgaS
lEAajDfPKWu9HzK7Pkf4+eghib9SrMr6biZ7IWJDQxyZ0XzFlJfPIh6i8WNJvcpilTm5Ms2D14Ef
5Y8D+ZrbnV3d0oXYZMOedDtIKvOLWuf+O3fz8aM7ny7rQCJUyQlJU+bm1cX2yF/tKXhsKt7TalW5
NIqBtv8nn8+f9r9zNSBAmAObUTHr27p/Pl7EFLWdaVLpezC4QgiRsr/D95a5kSA3W6uTZV9ZPxZo
RxOm7cwEhVeIru6g1ZJJCegP+PGMcGPAuySj2FilSg6stQrSGMzSwYyuE7xsgkbGFHsdnqbaHRI8
cvj/6bo5ZwzKSWPAfdaJk/6Q6xJW7uP5Oon43GPNdsIiy7g9C0+Rgvj1JmABQnnlJ1jpSzBokdAD
9C5s2PPddnNEm0xfBVRnBHIyadfvX6X15Jvjn5dzLNceU3vV4vzzamebOi0oR6bdaA9+Cztw/Nm6
Dd0Y5fM6lV2/DpzLBttUg89dKWGUGFbLyntvCmCNDf0jK1Am7wTsqNKfmxD5+mTbHckVL/T4pKVX
y9cXxIht2oV49GAFarh85WlhzfmzyP4rBTw/Mar4WDg1ZLrPFSeIsmurWm+7r625ian+DUVj6BrK
ju0rQBLfqSR6DIjsCquq5SoP8onMDar3+giFQAvJM99/tCxHsDksju06qQesrqaSs3ThvEyK155u
kBnuSKyK6HoSDxEEol+2KipvLgeqwzAeFXSGDwmU3zVtXMBQA/Uxd+ITsbDR7Qh+s0ewlNT9s00Z
nFe81MCrKUVJTGnRV4JHHEaGKN5nV6e+gCfe9b1icsLy/7i/Tzc4eMYX1BYEcUCMKUiTuODzWe0l
ev0ej2Z+wROdPbiUwOhcZ2The2WKEJQos3CjKtdqpQ3nELgqrgVaqyHBKFn4ctslm9o3Fs9tGzLK
X8T+Waf/E0FmAS/ycZOvu19vBD3In9UDFtIQFLbL1lki01IhIUN68sQVyQ0GZvvysC0n3+laoiNG
5a4byI9OzpSJXJ/g7jYveIvNoEmme8bXs3TkSKgex6SGXDRu93qYUITxh3CZpgTmdcgXkw2Utbqx
VyIsmc7XQB3ZFfFHlLOGbmtiy+q2AAD/F+XKbxVOhbUSjavMmo/+RJ+WyBUSC0BdnKG9XHpMYTFA
sYFUUEnpjt6w77gGQY4US5Vfsc0gRO21Uk8AWFXZD/jGMMq5hjcotwgc04+JW/DEu9n6BowQO8jr
06odMCkt2H6EAinFRDCHQBhAjF7fQfEOaZ59Jz+FoJStgi2xRM0/5KujQyJCMt4gJfruRaL/3UZL
aoKacdWeXSfFArtzAIbHYHjYn9lCgzBSUdg+PdRkm3edT7UZuj/dDSwWe5Peq9pAesg9RsTrH9jv
QhNzHGP+0jjVU5hjWkOX175IOo8fktVwsdRq9BYs5jLRzwn2/rQxuT7rUlc4wxlGtpO9LLE5nOQK
IhuukAsHnZyCxEMSt2PHgug6vYBRL2xLJp0ZhpMwAt1QAKK3JA3H/90Xk1zMjxUTr/xqDg9yp9v6
OKgjU1louZypSjmK5mQb/4mv2A3a4Ph/XbkQwURid0wQ88kKPa0WQlHH/dmHQtN3zIrB07qTt3/d
vKVxfUtuHOL1bElhqMCQLcfqXX5yqtl+nHFtDZDkNQJv5tZvBuoIN9J8mK55gteHwfIz4wDoEMZQ
r+t0yqNnjgG/PZoxQgcRwBKKJ+Vu4zpuzcwW5n7wFpM7Ne0OLa3g++1B+NLkCLjJd4vNaZKJPhGx
Q9NeIShtxyaXz1g3zMZ1JrFW5mr+ogNOiB3HPNbwGMFS0uPa7UUFwb04p3MTz/TY9XKDq6O53qIc
tiUx+89RzDbpKlgiAiphPou6erK3LwPrlC2z0NInJm3CE4M//XGGACxYFHaGzwJ7mXhhFx8GaqaU
7fnGOXxxKioLxigKgHnAvbIDa/swbfUn9X5N4S2s/9Zg5t/Muj8wh95jaWm7O2nDrzM0piNTleE5
6BBGSMWyqw7otrcZk/gy6rLaLIRO8qcqM6XvT8oC3LkzQv40vDgYogc2aR0zBwYJvM3/ln/p/BMH
bCm8kRL84lvOWuORPF06FBulV1Eqdh7mDcsTYT0UG+wnKNMFf9b3XS0p2wsqhHVjRT8d4OlAeqG/
eZ8RcBX0SJJrD9ebPswSxpcA/lo2Q+586i2i/IaDr1MDmkc4CPEBLh8VEqs+ffrX67b1VebxUWzs
PTVEzt3mn22sGYS2h2087iQXTjGkl5r6fH8vCAiJ78ZTwGx0EI+Fhs6GVURVHLOLHEfS5OcDD6Pm
QzzdVmABWLTr4dXnCPIk00K3PLFIxqfmDAndIow5bDPaFyQzBF+cXPxhpsB2g9PuYW2hc3RX8Cjn
lJQWaqG+hbIK26ph5WbrcjbufNb92SKfKzxVcgQXDRTqB0lF8bTkNvGiWvPwTyMeSJZ3V0Thdc4R
7yjRk5JMuG3TLYWsNLwF4iVa9uSnsp5aSvqlEtsVbRl9aXIhCF4nY+lyvLoSnU5wznBt+oLQsPYO
21UiPg+2kNgOVdFazaa7FxaIUu1pi9lnqWEwJovfsQHG0o8Hk60kn39t10teNeGyCbC+pksufAWf
r8mTCPxt2dEfOTmdt4Nm7NFu+kYUmhC9marlnfPX0GtwZFhrhV/4rxq0tU9b4UzpEG1kVmx0RvuC
kRDLJIGKuC2x2ulXw3qc4Y4V0hbaB0YIkvDbUTh+ZuCxzRDn6uxqc8ZJ6MajE7zOO/Jy/5QoDLBI
oi+B/7fk9Qsijbhd1Cq7FzWdYDJaaHO2T3WiU9FxaNveEma1R5Q7H/BiqJ6aBhRCoRe65dv5m0sM
43jbHAnGqHlVNeOTw43l5RnDojUGVXVrXqxdbbdjYm0SbnEHKnVMqghx3iws6tFQeuWI/WrlQgBX
sgYo7z7cm0ZGcF56kVhCGYECCyz4Y6NdipSyVxFWigv+KhT8RDLDA+kdudAwOnarTkMw+yRacw0J
Liga5DFdQmfIJs87kxKh7/SmtNO3MqteAkc7Cxpd9Eu9bhrX5DYONVySFPjqyLhtbSlIan5e/UjC
RZD1m6KepxBOfG6mBLR2MUSljFcsIygjM4lcg6+/LPS2vVeME+V0f/N4MLw0St4IgIEJVN2fO4Pd
uzyc/OC3FE/wR4B7FVSqORPzif3gRIn85RkST0zhCGZ5qqpG+hYj1qSatDKqnu8VpNcLM9qv7DXH
vcrrPqm5AbKtKVRAoyznYJx3ssdqZcy8U8QFpg+6CLXXy9HPU/vhA00cEgEximofdRSe+v1KfHS7
TzeT1++a/81lDGHpXG9PMGPcQuDuE2S5u65CEgZeY+PDBxh7P9jwOc7GbLtX8YhgQWPalO+gEKWe
0g+xtka/qvmPNL1YBRvhYNfBNPpKDyEfXS+eOCzhINL12YG4bJPWs9vytXf1UJA1TZCrkIUpIfSs
AlwxzIdRIs4gzu/DTzBNzDJX2IPMxkiweUIbhZ7+81h9RELKCG+2QxAzp0OTQv7jBoMBlT7v+c8W
XrqKv2X1+7zfnK0C74PjmjuSxDWXXdx8G6JzujsCpm9GtYXXTXlYNEHQzRAZIKytCLXnm2mUYjA1
rNd7ucqQCfKejgoxBEmRLLCQE63V/Bv4mmuLb9GrVmeZ/JZU3WuK2DYBcMcXnV9imn2K7MZRaQNM
6jQ0t60g1wKh5zauDvZAEBX1tsMXaXwK6/YiQc4QPcm7nkxlrjLY+S4SKmRbdgu8MSNAFrm05VNS
Tui8vhvwSbP0oMzB0EJQ+JAAE+Dg//+/PXaoxRzgjsKPvU7d3tj02L+QsuGKR44Y6Ue02fI0Vn+g
kUjyrPYnFwH1mktMDXBP5Z5lSNQgUcWsZ7yGUUyY8sRib/JdrmmDrqGfSFaQ5yfuuLWSNXwW6koO
Ec+HzzCA9gMdDIggEwdzYmHyYry9gg6kSe7e04F0BGCFktmPWcWVgD9sA4FmDo6UfnB6bxxLLzpu
0Rcp8w9DYeBdDsLQoU9WmHT2XhMJwf6gINRgLP0hpFepT7zJWoEe9psiM3DJUsHz8+Wo4t1NinYB
uFlSZxr2HgKpYJtapioRfxw3XTSphGJWksDqXxfg1Yo9AiEf5NQAYgj2zeNJYX3hQ57GqHKsIqEO
D8ZA0fUKCxPnvsaeu0+eAcvN6lSpNkUE8JImUdJd+N36V2CpKXvSfk62wg6t2IQpXoYcWzjtT3QJ
o6zs/XJSNyH2tXUM8LDSi0utNWx4UUQzI9Nu/Trv69pESCMf9+UkciIrCT2FuoJNxUvUSMcaj3Sn
Qk/ilrou6kLP7XP6Xhj4Fs7t9raW6scKau/7Gai+5cUBAeQ7BMyX0TfqYbtpx5PLZQ3EpFv/+/us
vv3GrJYxaVtUO5jm96JEFKYHN6iTijqBOpXekGvpU4rVQZKvzM0/jxz1JXxKo/wb7DZjXgAN/CzJ
G6EiowNdJ4hTxGlFgXjFF4yJpNfazjX1sSlwZyCr7Qoueyf9NxBzX6yp2xGz3Tq2W/hE/DJiiqQB
CMV+W5ZbD44vZGC7jcG77SRmiZGjpo+oVYRb87HAwDigo9Zw69SV9Rn7sCL87DDRepUAFJQWL73w
iPW+2qLc96hJRR7XE+Ews1dJHmiqQNq/BhFnCx6dC5wIR+C7s8oVmdLqd/uIxOiT6zIiVXHINyjT
2L+keSMo+1U0VFPDGZzIaTtgFx8VCJ8jXMZ0e8xVElB3Mv3Gj/cCbANEMgfi0d61Ro86lXs0HFZ1
ErEpD5+IrPIuCLZgVYqxyrD10ivgzyAWgIXhn9RzfEjeZ/ACvUnBXruaWbJ2w0jAgD1EZZ556t7C
fT4uCkpOiCORZuafIn6QbCq/eQ5sKMC+PWEPy7ekqiPLlnQKen7LsRxUU7rmSEmRyz1lN+bWP3m3
2afNPKaNFMI04DTN8yR3CaqB3ueDkQdmrUcFerhI5LqRhk3WgEo+UAAx5o7wpwInV7aaBSCdsxTJ
ohdsC3iR4UHrWUpke/mV1Dyn4xt7eCiZIfjR+V1bUMgf9F3NrnUM8YoUxdwrwRPRykBzv/S1O9mv
XnWZrEkDcc44eBvenKczPhW3jsS/zHTCnuTQ21iIUevnxTFwMSTVTSr2Kb6+mxpeNZyZZiyU4miG
qeowsFAxvHCPJiymzoCKwWm9UM90MHnKqPd+9g51GJP84+DeVQY+MfRbPlc5lRJtmZi5mfU6cJcg
rWqnRbolQCUsQHsADYSi4MNbNgOCADKove5TUKNu7rcL8wq57m1EVcPIXlOT80/oVZlLb68YqoYB
N0oMVWqPBHbMvsh562wiagsFy6ECBb2A/VOEJrld0R3oPXlyZCYoYAbUDC4Jw7DXYolV5G23jsIi
p5GR/Lp0TakTEGi85fu0eBCQZSxVvk29IDunnp+OcmGYMWRsLVIvKy6zn25sp2BNMO6JAIgZsMcj
xgpI6W+yZlv6SZTDH4Cc+hnD4nnOW/y2XQHaOt7EYMx8NGR+A9BxzBuZtI7KvCSlKO9+hVWQADf3
wMV6EChtB+k7FeQYbQbqU3KP4W4zAKvsiAY8y8nLTJaDdlwvUUPa3ZFoN19dwMmMDJjymf9UesDo
xfTWY+mJdsY/NxrbfWmCZEdJ7MjrNglGhyT87Xd9V6kYIjpxjqwRoOQjSyHdWtCNxiIHMaaliEBw
xygAn21bNjBzl8vL41aRXncIeg5hpe7S22UHe8fwVOI4LVIReyfvJ4XzFMg83q59HFx2joN2ZFvk
3273C6/bPrGxXZZJKSM68rTpQHNx39WjplTYuxOBnafM1+SNqhM75oC8x/3wHQqSNkzP63AEzhRc
v7Hv81Qsr7xlSvzHxyHX6MF8C8FLKsPfNIffxAoHq5/ZlBv42VrS7tKDQfOurCBuznxEkBYcEywg
5VABlp1YakgoWluhnKgYYfpur//TDVSjS0qnj4y31/f4xjklulwWVubDLsTmKdX7XjHcpaoh6fJ+
5FTXlZqpvi6wJh7PP0z4tj5gJ+zUAyv8RRnVTE0Ajd00+l8AJ3PIWhgoANWJ/QEDOKLPgWEEzwua
gPJ5eSfxHaPrPnX/UDoBlBXnWleiu3pxV1YmO2HhLgoViXlL852EPWiVR7stbxcnyDKEKNiANzcJ
RLwgZ9VlqBRlvij7a9G0EMVLnkRNpFXV0hg02cBp8j+jpKilU/1eOYiuqgG8z3L6UZMZPy7vRBve
/IpnxdyanYyTiHKr+YKeSTW4U0ghUmcjA13uWMjGdq0R/N+I2Zja8LR6/EuBL43KnwaznYnsyQJU
GPmUj/iquU88AiLj0NZRtfzdZfzhOaDFN4UBhh9Z4e/yQ+I0+PPdf5ThW41prF6FKIziM8ZdTsw9
xrNXHtY4o+7BexqPXHGWf4jmIHE4qRp62TkCqaVqtVsQnB+uTIE/HsG9q4zRnqf3sz2q/6yU14qP
85/JJSaCKpMSvzQuFYuOSdhtmc1QPer1ShJIj/6iGMh/0MG9rM5MkA4y0FEEPZ5nsDN9rwBuulPj
rexqMSdh44EZ96igiWH4mwv0/5/AwIrRegokS+ju2ROIpao22b0eHddOI61Y4pPEGgZexBLw3W8h
dHXiimA7HYTbYP8GyqEnBuLsGXf7hE+Scyq9ARU6l+KkuQ3jeU/PM6yY5AiaP0D1CwSCefxRamDi
iCUI2uQ9cq3czTkbxpOUXMZSOmtikI3dG/orDEwECfML5bd60VXNN/MR9n19EkHGk0vXUj+j1YMO
gN/8GdCE601wPzBhnyMuryNNp9hAElNs10GTZSPVvDOHVeKrJEa1MrFJjhVRi+2pc7XCp8jegqmk
vUEMQ2J8suWlb5xdoODJMT+fl8uec2ylCbIkHhSU7BDDiaM/mFwns3xomb2kA94h7mhc9qfCJKNd
WzbTPGD2W4iXpYNdiGcJqIjsiIqZinm7rCsvS8qZp0WSYPCj4hy9oaVKXhotCH0yUPAYLj4aTZiM
0Zx6aoenJnV5FLudrB8u4IPEMacHV+cNdpz4LcCFHrRZ2J+7vl/k3P/SI59aPwuH+LdGUI/g735w
hBFgafBQrWyw92EGQv+4EwEEjkwL4C9JNEsLIoYYQnRkCqWHF2Trn0OL2aakNXNZ2yQt+5PxtIm1
HLxot2zxIBt7BvRXTT8ammCHxJu5aS6ibSnSP50VevaSCLokmceGfwCabysBrG7mHL+T5L6hQqwb
s1f7cXKE5h1Ki2o+uIFQXcOyl+QfThYyA9QS0XAX5w15eLyFSchhYCZ9VN6UQb280j8Ps7DE/01q
SIaZ+OQIg88g8z9YzueI25Ux5me6UGFfBmXKYUtPTgG/x9p2Sucs0OHM7EVmPuBVA/IaZaGJjfge
JM0hkhot5FCoCI3cB1V8YNJUHYCeJccH5Dsb5YW3CDEREoCjOug+HTSM8GsN1bw9XOA9dN69opMe
Q0+1KOt1Bdfl8Du6ukqaxMl1cyhKvmD70efP8nQnU77I4uenepyZ0GA3AW54yTNLNr+o0bT4q7uY
iGYTAeXYdI+Pd9NIV+0luST9YQX9hxel/Gj6+NMRmgIhIiHI6yjQmjqZDibofXU6LgwPAzujWjwl
zBaP18Xd/OSWivuDp2CUYP2f59J/bmRSkRSB2Zv9kEP8aps9SV5VfN2h+XVI0hoRVJEsrqPNGeDu
SLZa4ICSBOPkjyElvNxFrmYY51ipNuEI83T4KhBmvdXDYvYsNu49+z+uNmYi8BF3nNHPWcDyJm7w
vNH0zxuEVUZG73avq5XpJAvmzPOx/WbJOlsy7/7nhI+RcU5yATSFDPF65WW6tpBnrMcUIzDTgMgH
h8Z+U6DxWLJEOzKo1iGooVA+Pwshe8gMWZf/EIgFkeZ6eTrelOOemBC+Xhvh0fjBD5mTubnzli/m
eM2CvicbLIdF0wAkPQ7CIamQQ5EmUeNtH7bENqMDma7Ij+CkNXmUwp9HPumRRjJPthOuqGuuqfOA
piDEz2nZ7KgDuYJVUTSnDk2jxrcwQxMR25Kt6C9ZInb8noL+6bQnH7iLuIw+N187rUate2esXt+u
TXGcRcK+FWvYIgDVz+BBVEopbTwm8X2E4e5LVwYGxZCUaVpkx6BX/HPznSb7IV1WPnm5UyLTzBEj
ZNtPFu5cNXBnYUb/R1AmI8k8RjNh8FioTuhArzV3rgh50O46wBJmhPWtKra0pPgLGEiKNUuO9O7r
SJjb/w7W+0MfpMrD8sXOrGnw5itCs8NsgXiUAa/sORlbyswb3OVx1rybukMGF5AREsUvdQrB/QNG
+sF0g3OZmkb2Od56umFepYRna1/ST98oJ8hrgQHI0hh6/WZU10c1/etelKmYnaSfomiOXaTJBTNY
vbyy9jVH6uMgO7RviUo1OGH9VkGSKhYd5qVEbu/WD7X5k1WR0UG7KlfX+/zEZo2D9z+G/adItju2
HtR2QthgayCCqmTyMZ65H7umk0n4xzVv6OHpQhuKtnoz0uUFaFLB26x+31/S1i8gnTesMUN6VpN2
8XsaCqdAXflDSWWCSzrqPSgHFgOyWSJbLz99cRRpTT2KsZ7hFedDKN+JRLaalzWJnvD89WBbKyCH
9pruwUOuRXYgLuTBh5ULx6XooAhjS1unqPrd/gaQs794EIEp+vHsibB6bAfBZCmsVrKI6Zyu99qD
MeE4CvR9dMnNp9ZLsp+junAiDEtY7XOXnDiUDF2KfdVRnVU3IQJPTLVK3srEqUw1gBstFJqU1F88
+L+q/1IFP/+VIB+DpW6LJLhoyC2merq0zWuZTUhQfdvtb9jm5Gs9bfA0EbnjTJeWvgD/vu6gjxO1
bdkXJvZbIEUo2lyZfibAHzATi5o7N/2FpwGBFb/mnc8JHaGCX8f7sqPo2y+iC4nmWXMH7r2HrL+g
/etKSAcrzloEPDzC3TXW/bYAaPjG9H47vK4B4CtdeR6O81lVzCTzmPfVXz+lqLyDppjNNktG0gBC
+YYBpMrwm+P/oTQ9KpOU9u9S5bd8pMCcYrIq1UrxTSjX4YY/sy9fkjgUBvveyjiZLPmCgkOfQhXG
AO3q3Uer6FbGwTLfIR0xp1/bPg4JzYLBSt/NC+eAORdC4eitEUR7dJXbYYUkbKWfkt6k6Q5ptFuF
M7hrNBPbcS8IZieHHKUQe36uDAYx/TfLkm7kpP3IIagr61nEk1XZLfXQVwvHWoHX66lhW8knjECq
a9qjuM8vld+uF3jJQy+6t2erJELMNvrxfTAM+fRgmfIqpc5U81v3zFvzHQwMdMJ8q6+xwPW+5B1T
TW1gQTBBSsivpUpUUALQs5q+Q73V8wVhIoek5Mu3wytG3S1Y+4bh9JOpD3x0VNbPulN0W4QveS1v
F7MXOuX7Vlk06nfPIs/nyrPG+pgzxpasJXAIXxLp550UKaBtCW0aHHHkNqkNni14yUIzXHdtpLZI
ovCeoRGOFs3y4JN+ji2uGiccUF9ju7QNN6YRSud9NpeJDEJaT09kaZ/Sfj62n2bFd91fv5kHqNYk
vNEU1dXyu4T8KH98aKoVgqs83gh5YODIO/EMZixbh/gLUf7G2j2vGc1vokwNPkeTIxtXd2h1psCQ
bHlzPagDMb2M/2hIq3zIy6F3NtF6n5skEYEwIBsNc/Wwz386+xJP8IDJB+0Fmdv6cEM674kwo6O3
2xn5ESizmgdrwqZhB/3x0/AdDPOh6DN7l/gG/gmr/jZEnx3FsT/ns0r3hksygVFvWbbPZdYcM7IG
Y1mF4yGfuXsMSXpiQcB+J4pzDaIbYumnmzrKHxezZ6Z6Up3fYVFEa/7qPMQcwh9NMFfKp1buOBbz
MqvTBQTNpqxtC3xGdkHNV0zNetldeGc8GSWHznZnmwP2zv7VBM1EDSp0PuYNmt9SYXygl1tuxQi4
S0zrPumWbZwAJaucsa1qqkdXBJYsP0J3DZ+/fdSAEDYkveCmFipoxqN1EWaiiwvV/38ApdiKr75K
hd2b4/Deq9+W8A40z82lUS1hGTHGj2OKJ3qiMVpDxKThWOwOesw3JFi7lgW0+8FNfo6ZJwGXQaVF
/W93sGC4byquyyuzIhtNL8L5bCyBBiJtx/DeYeS63o8TunyZlkeD1jSBKORa4kQLqTxKbW+UASDY
a1U7D+mnCMptLus4kf7FP9ABhLS2K9ey6vjJkBbBMWdGtOszRFMsRFcorYGpQNJUP1YCVI559thm
RwWjcyt8VMgOcwyNppCczDkhg5shAN62lOrSy57YYS5Ut/3bGdnFKnSBeIvei01yt/V1eP0Bmd87
QQ/XgbrkZe8xpeC4k6mxBzDegO0dVRFhENO+mUsF+xmvwImPFOHcdTGfi9EuCL2XfuqlD+ODzB0s
JHd3cDSqkUBtt6KHY7YTQ+nMwsvev1MgY/bm5r6N2UfvJB/ySVDAffCWgsD+4yf6uJrm6Cs7IC0O
VoXT293+UNIyb2ge+qNB4fHS6J7Uoo1jdEvCg5haX3ElYK4+xBl93tXrHQh4bPSyD26Ac2S74U9t
6DFiIdFafMd6JTy6IenB/yxCMpgQq+bTmGshBfDc0kVnF9pSkp9NLZ7r5Ph3yyh9Hb9foKTBxQaW
0pWyzbfnBytqJ06GZRCRG6uMRGz3xoE126kN17sFtwDKEz0UhHpXWwecOswlrzQp8VfN3vJUaQRM
Dy2dRGrchPaqYUNemWkT1yfONXIhod1mN+S4sPEoAHiv/nUQb20kMCAvtHvi89t14JkJLjJjsCmX
+KN/bUSUncDiiGpGQtCVS7XVKwvzplMBdCVSi5fyhe/PFMd+HCSJZ8Gp86h72z2/HlshHgzWxx7F
XGaqoNF7WojZvj9dXR1NcbG+/LgLzdHRGZNFZTAd4MojKvfbai+NxAoUEgdh03AYC7qhkUDmfQO0
WUmNrm2FgR8rkZ5jHaG/vpJul1EDgX01lrO36gH3sFECeeoylbIQejKkzJSrvl/1aliCRGvq9nSH
E2WE6zpCCpceKMSZTMIyBG7rNoFZ+SVMjX9xnwZalAW9FNUXRJA99lbiL0Cz2RuUrnPwkOpmijRI
yITca7sHSvdtM3GwX+7jlPIiOupUL213zDY7lqbsyq0pTGEpiED5kD/0UOwetwiNwShgskl+2J9f
nkRNiI6kP2CwgtRDKJAx5Jx8x/7r5udW88xwkflo40j5v8wvu/zyns5Pdr/UXCKIRg0AwMBGqgDs
10K1rtl6s/z5+NYOE3s76olqjWoP0uqwbpS2dVCFbQ2h1pBKWt6FAGx7rV9FgCjVrNb5m7KMxlyl
11HEv+jJ52k5I5WEfyQZwNqcrGcpVPo2JBAFZYgQ51qFAmrBHvO9vqZp2xdWzeJ+QLHdssGylLNu
w13QqBiQtixgKTXOsYzN6/RC/sOJWz/qOYjnRwJQVRY2hWUAxKTEz5wLiNbVJgyWKQGwUkpI1g5Q
lPLthB3k9IJVTMCfNlj1fnZ85PpOzqdMlxwrDXpwrvMA03pLf3AxRgrLR3diBT+IfZLw+5P1Zood
Cg3ngaAlwnSwj+22b1VGwwfn+gyxQXzLKfl3VoREBqmcRro/rEOVcT+TKjNCXxBbrXfXccGsvRY5
K4HT0hDPjxciJVu85jXN6dT8oFN5QJ/O4jmtCCiapG2CFkQRCTKG3ziEwctB+lC+FMd9N+k23Yoy
t9hyaUsMwUi+hwDkeVSq2EAIdBw9jVoptqBLQDB/T/dM8UQxUqM1zuHTIDrhr3e7JTgXqsZPqD8U
axJAg1KW+D56JhfhQ0Gg/zf7N/AeSYxS0tnzdNH7pCRJkqNsp58Nfy7mOn9n/7DhWNWS9ffpDYIT
UaukysxNl/SkFpx64HnIZVngFNsgBU5KOwx/TU08Rb1i9PgbHYDqKSwmQyK/QUwHKzdTIdYM76Wk
Hj8HTD5nSMFMhmuauoeLx94Fn/X8vn2ATSdQa+TSSrcen13TnyCB5036HNG+rcAgv4AUq1qKoX9U
me9WLzogZrUk0WQbOWJi02Zd6+JABnT1oy5oMxT7lNMRJ9y718CrBfCqhA8qf00amm92k+oafEv7
43NTpVgTueVW41afRX8DwpdzRTICYaiuwbol+r1tfYoeQtsyoCVXZPkujwXrllzT27Wts2/MN0cl
fAW4LVER2svG3puboCzGk8H6DD3D917x49O7gG3KuG81ZsmuXlfAJX4NGcaoackyY0heXEIKw0kg
UiIvtDoSnJQQRzZTNbdrAtxeSyp8+1FBoBwotzO163gjSbu8DWz8LEFDpbeOnBBhu9XY4y/WR3Go
2yWvFXaoVo0biV2Fzqz/pn9H/lXvx4V2Ls3S9jvjrBtqUiJX/gR1QshYihnMP5dA4o+snToajTAo
jiL39HnPsZIalA3ZDyylZ+5NC9JvWw2GhqfNdrfWpLxm146kcv+34MKLobCxmvoz+uuxRotbDSBq
N8wl5Bzbu0U4JThJ+p9QrKeh2TUY0HwSdIgPH3oubejAzxAKDq+RlOpfWlgGWg0DE82kvAffJDyw
p/3W9HCiFo4jWqorEhVCHGtrA179a6G7zPq05BBnDwVfVtXx8l3uM7KcWR6ROzvjQwh8nJAa/6K5
gtTeDT5VsQ64wm6KV/aCQp3T456jL6UdardYBl3KLziut0XRquWhiDNszN59vkSYcdTb0rEnS4t4
ezeNngMgDHrph3IB109ZFDy+vc+7k4pzJWxj8vd5wYpj/hykD4tpssgRMPhdTllBeBspQ6VbeWCb
TMigwkmZ63T6RVDpGbPM8j1PVvS4BQ/K9VJ79rsp2YqstFe/vGr/605tGzaVKBRFnOT5xowNCsUD
qgPCnJ30wkQ67Qp7+mL8+R6KIdQGMXaLz/MQqqKFJnf+Sxpzep5ySZSQgEBIQozgoMwF0N1N9cJW
DCqbw0Ewj113gK3IpBceY4AHOy9MNzBbbczyJl8gNBAc2vVSZ6DPLOBICaogqMmfRy3ZTWSzeIDU
C6g1HcLcP1O3PWTaQncKX8g/Z2LBNW+Ba54X988W4L0QvzHxaJTbfDIhpGJvOGLLlg8ZtFs+f81t
XM/nSlIosYMaLGqzxIna0LWbTxPBnOCDAhbF7zRQEBnNFFBGWy+EJXX+2AWqMhrJVlVZS26OkvV6
ka9nUdDVM29Yz2xzeM+Y+xDQ+JGtj501tmp3VTiT8dYhwt0uAc4ggUINLlfpUfI08oVbWXfb2waX
97pGJDzglt+W2WdQwFnjzf3n2f+7ro3sTYf2rfBc7/iVa0F/RqVtLP1ELDyy2LYYKZKqz3HBa2lj
vQPGZBhXAwKdTuWkgNeToSk9q38G9Tyk0gQ5UpdOJcyIIWynUG7+qk4g1YLH6xsaRVIoow8zqSq/
0S4POsr+aGpLWlOPuXNUKeCvTwCdm7Yuj71JnPmktK7hA01baRAJAXTGLRvd0xr1wrm5D0FvTDMq
Z/suEeRgkwWQlidar31QY7q036Tu4gLBxjKHdWPdexeXYajASGq/otil5ajHQ+knaTlAat81dlsc
mS6CKcRtKRhcMuoYueZ1g2RMkiKVLBenDq/V3vRQQxWs5Y0PR39MNwY/FUYXWqKr6jDCBjHyrR7c
sfMQM3Kb4kTPTKrRzTNh6hhKu1Be2OL+0WxleHqjaF9EMM6nu28fxGZgrKClHvvlPQgNfqIRXG9A
S1b9sMce3Pp5go2i+2835efmwULdafJDBYti30wqOx0oN2dP8aFW2IcJYpmyrY+VOUDRjvrqWMxG
XdlYclWvS12EIeGB0MDCQDlZCBttopSKikvOpyKiHBoGKHBTvFAJyxXpOsUqxmunLTKKWhQAWqkh
tGAmjk3E+HJktayI6EjAc50tiNGM5rTkmQSG+RYOrxzuZKC54oOhhE6/BadydrHtehGZrSfHGozQ
1ut5FKjNJeOpNjHYwGSs8upVbU4Ht6XWMFpXc5dJs67TbNHCJW2avL3keT5QOhA8Y6GZp8OzOYiA
ItKm8CicoRXwr0qmeKiuKM5VYLqoS8eLCLljAPwIfRE2YfTONgngadNj5p6EWrxmx/chaTt+GdwQ
R6U9oRho5919aZethXcHJ88JgEmtxfKflmR/pDalEZhrMlqMluP1d4/wTMX09pgDaMUbXcswH/+7
jKckPHzpRcec8urCWFCdGiwsqy0p6dQew7LAijHhi06zsLU+I3XiQgdaPfeGNWuGv2ZJadVjTz3l
7qfEN+TO5Lss4gZeYbIQkHV95/GMk2jARimTzHUfIyWSKIRrgf+NldRv3fg/TtuBnDLYwxPpFZkf
4Gc7f1QZX7oOAbPp5QRFAWPsvRftlIEvuZCTL5nKZZHIhGWrFWVPQPW21y6QmLAPZlcrxJbPEsAU
becZErV6Oizaf99RqwIOgRQECNOqPjUaJm3hLnAcm5giylYIr+V8s/sLrCZUi/dy7kfG1h6QJ7nC
JwMuFZC1hlZ0SBJqOeMTO0Az1aSe83FTDghE1h6jOnM0ayFWl6PG7FBlpPBFAU/8ANIVSSZGxQ83
bmlQxws5SEsgexVrvZGWMz5qWL2U/QLDMLX1000Tg0v6UqtNN8aLsE+4wiQ0ddhSczgs44zp9dQj
seN+9wkFoohxCiS3YX0zSLjTKyjBiKlfbgZxgcWSuaHo0j0X7rWxI2wp1AkoWnotCAclbkOp8NYL
tzrJJ6IXsCVCW6ReJaYrJebK+SCvHPhtff3OInp5DUstHhlIqXHuWC22Jm6Sx1dwlZiOie4ib0y9
f98+YXsiMSJt5AMzOEjNq1qgR9G79MnZwp9rhxVQrtdTU7uWgFrNWIgNg7Ej+Z1p0C2Lba5jnOiv
s6EFGl2xBLwKONMINx6RGPTslukJ6pqti1k9j83oMtTHFm0uJh09iZNg8wEj5Q+c7QIsPnqNYUDz
pDIi0SFezEEJMP8cUNYDsDZ5jFiTxeL7qPSGG6AArPFzL+9USZb5atwAH7Zzk9ZIlXDF5rQzGvEf
YoIfbUcCZnjTq5O2MaFQ96BSUQ6XIER6obLSi8t94qqh9GFMG2SnpxjCO68Rt9saWqEZcHvjaY2B
7aVrZMx1BD6kqplK/MB1eZWua/LTiDitlYvtdKqq8pbwp2snnYMCafQa5+cj6Up9g9BCorcTFz6q
8XKLDEmhYQ32h2gLFcb8Gzong3TkHNRjQqyvXCUye0oU8nhcPtRbTyz2b/Lk2aJtX/npRtIpZCh1
/us8d4Z/LbKjA1wqA1jbBEAOHCmxRL/Z9l/ccagnWqShfH1qpnmIzbdup1Sg55ylslgA1znF03kp
AA3Aj2EzZSax9cqNJi2DG+QIBQFLcgoaCjTgmX14b4+DYW4i4Whj5hVcPfjCtgvp0eydY4mXKDwL
aGmkgXZKR5b4sHz0Vn2VQlqBivm8erpppiFtQh9kAx7LXV6jsyKB/3eM5isZWzeKvDqd/OM2RccM
FHuHiQZBzI106CaGZagslwmuNh4Vkg2gblWCMH21X1FFQWNzxtnW2CWN0TrzrwVel2s4IJKe4i0i
9bA0K5qM9cnoCHnlo9JeXvAlRJbw6zco/73HufxPtGjw3TZLNZ0bo8iDEfiQ5HslWFwUTJUHlO9b
PbWplzUAXrK0SLKs14XHxKi1/H/OKYQt4w56AQWavX7O6aX355gUQTlLWHkGhhTT+ymhwssSaT7S
or7FEHKll4MbttBcrzrRb7qwvRQAWP05vyD6cCjSqSX2IMj54lDSaQtSZzDUYaKoPd9w+wSgN6lF
3svisTVD6YCpdB0GmCOKMIu4V4XRGXNmjXTvA9+EQfiyhaVhzVIYRab0jrol4ZVG5U6PZpxiZt0n
9EOeVK2ocLBJM1Ga93Z0wogaTy63xxZOoJA4h33IdtxGCOTFTPXDG+f1qArAMh7CcUdEP6uNhvHz
MFrgc7iCbzJZaYGGhikgcNGya8Hyoo0qM9gC/CS1Zot3fszx8n7pbOqTzexGD8ZlFwJjLPTYcReG
WzFqJPkIb6MOmTrxH+YeRiHUYth5VQSEP4za0lctBsMtUK+8AL0VhwyvQXFufJw3+kv82N4c3asV
vVjJGdxlmWO3bNyk7d+k3SbBIBpXKD/1jkLShkc16hqIQWDuoz27SJCkPk6JR9g3i+zTnsDAL+LV
NtyehZqYPc6AneXI0eajs/fiml+veVLr1hM3z+fldS1pew1bIWk09b2SkWlZrQ671MRcgTnA7LgE
kzxNp/+CgNQJ2IbnXWy0WT1QURx6k2SvOx+RlOybNgiwCWWZFF2G1f3N5mSOnHvnIAcNeHPYj5BU
/WqA6hyU/Ux1qVVLd/aGb9UFr5ZN7x9V3Bt0vdtQHHSFPQM0hLFUIpXD3o2b+jKlQ61yXWEOiQca
sObBdLblGorcNVogDSIVTpXfAUCVd8sORAF+oTEdDiKc3MpmqLhtwM6h//jp4QreLjdtG0lbBVC8
J5ytDpIvubqpwVBueaHpEkLEjPIutvhLYBZxkBVdCtXXapPkwsq7TmYpYzs3FYdPJC4x+rPkVr2o
AfloujlNh8F94OUhuIPXMA6G8EbVM+iKE4ijLXZNWoxxJv+v48bi+hAThBDcgfNswUuGu4ol0Pw9
lc+nPBgrJY8uogDig+uAuakvr+hVqdxgFVDt/8yMGep4JqBQ0oM8SsOGNO+5eXSudokxyDOu2shy
1lYDtBXBVqueaPpuXhduvcNteS6KrrKs2TS6uK481keeRR0qVvsvWfnr7zBZt/EFhhjJ3zWeRtwW
rUXGAMYo9MApSz5sK8F3lT08/VzC27/y3WVv24dj3S75GO5Q6Le9I2i8Cm/xql8WLHDuO11PjA7t
cLeTSJUGVKRR6a7A8VH3/m7u9IN7uFLGufOukjxfXdPCGFLIyti8Oi9hjLqkVneb8kFYW+0kEiTe
Z1XWaRE5LOsKQ0Flay8oRLV9u/nqa7R/ejLgacNUspN2OtXoPBihj2xx0UejF5sLKHjYNAQYJGQD
vA/AXoFyaGZ2diHnP0w85FD7pLdmxnImVKJWuSBIzQ8VTbv78kVZFoyQoxbwg2ZQLtfcFDTt87Fw
cTSFYmA2iSxeUJR4ooOfQWndsq7RIvBM1rgiZPu1yy89DFBQPZ4wEt/tpbOAREG3lUwd1qq5fYE5
EOJTXxcMRe65HoUbcj3673L0rUvUzWriRKN1HEoUq0JFLgTKv86IiPdj4zl/YoocmQwiLu5c1UgP
Qj5hIs4PIuUjVbopKkxC2H1MwKAmp0XiPh5RMV+uHQSSyJCdTLjmezs8XpJ02Huxz0Vmn1TXlNne
3mXIp/qjbRgrS5Vk6hDLfzldB+WRl5ZFtbzDA4dLS5Fh4S2YgNoPzGEdZlbhMTuL/jMytmH3aVFB
ycWzvtr/Sk5KNyQ33ZLWWApCV0+9Y8Z1wR3ixcddSIBMXXcDk3dHKFlkbS5pwvTBMfzsryIBNOMy
UQrhw4XEX45OqFENQatejZ1N0v1zLaYY+B4Mx7u5aVoh/VU8d4rL0T/yVflSH9aO4hNG8BB+ZFcC
K5UZTwE+QfoPJt2XXhEg0nlTlHyky5Q1+xpMWlB0VARTQBkMcCdc71EtMiNVk52ONldb/JczeZoV
Tl7ZwGMHe+Wpsx4zlK9qL4s6RA8R+F9meiOl2v4eIxQBHevxsSG1K+MDCw2Ix3eUAnHqXokvRVyU
q0GAQ72AwoFlGTfczoawyekk2Om/DiaJD3Z5VbLFJ+xN1Gumch+oYw3/7yT/sJM64DCbd3PiNlNr
Q30mb63e47SfkHCT82s7cCE34aY2+n/NGzOiqwh8zwq3z59aR6WF3DhsdyJPwuNfif3308hnKb4Y
EH6lZha2kQItH1mjXZu+gsmiQHDn9SnV7gQErOqAUjDBm5sNWSRyXks/WNnybfPo9oyPtg3jCWws
gHlUSRnum8dJ+obLznvq/llnWT7ESceq1DR1Lqja/My2+z1e8tvi2D6kHtc9bWRzoFpY6hODhhE1
NRDQn/Fxfw7lEXPzBW74KG3oyxmN4q+ZOzDL5SPOBHVSZeoHKeb4Vn8T34Jq0LuOI5OaDo2tWK3B
Yqwwzg/AjpSxih9/SRdYQC64K4clBfS46LFZgOT6uwghwHJbTsVPBr1X8iqgnqtgWljylJHa8StH
fG72AhfGvkg9ok4fG0eOga0v7wFyH909E5VPzu/TmyKiXvdT+m/4NFANkrFib3Rv++AFhvidjrE+
QAOvmfJZcdxzs/VQN8QaLAnJxB/EVqTF7rwW7aBRcYKnQ0kAlaVaeMS6Fmmb7nhLtNH0UIhsg4ij
0ARYNBsHqP0KxYtbIHk79pvKw71FDLAr3BJwOaysq9lUFNXtbuDnn3Z1a3fMTdOYyMglUI+Bqq9p
xpOZ6aG/t06f7f+L7NSd0B6naMhvgR9V/1qIlItSh0QUSmmSLe4IIFbzwkc+/L/sMPqDSBll8ZcV
wldf0uqFrzRRztz5r0QzRO+TOVNOhgyUxsLRIHVwvgHyPB7Ny27UKTA9AlrbOVv96IC0Pdmb/Tj1
ASYiVL3Saeh5sRiCKaP0f85IW74JQ8xQcRnkrHbUheas5ns0nDz5pXOfclu+dSqbmXJRyl5l+z45
72FLc0x6a0YUZJ6zl1wEN5ZeGxamHE0Tkd26VFUZAZFAkvVX6dQtL0UBYURpEc0ifWN4GI8eY+G9
ra/d/g2DfX4gIc2clIGmkw9oNq3qmUQni4/lmJadiq6TVroHOWjg4KB8hTp59kePnWhX5nRvfDCl
z3SYG8sAsBoodJ0miFdW5aVJQwr+pqUFHxbYWknDqeb5GnkOI8OvZDTHsEC++qaE5gUnU/ohx0An
LGKgqm4gYLXgzb3Q2wSqPLK7DpMFZ7yQcxQIEjOJS7W3XUyZzr66C+fQ7pOglbvru47zS8wczP+q
sqVbxMq4TK2eOlFOFCaL146aLZAv+7vIDFfQsZekCrn9koH8oYCsNGuiIYLqgP4D7qECX59JAv3P
Q8rlS5kox4SfMl89Ok5Zo0xZZsZkfWBnqr6ioMKLDE1cGpfwDXF4n3/dBZh1IUiLy4/Rrv3RlI3v
LZ+/nEfB8E4XJ0Lsh8Vw/Gnh/9hFH2lUw/WwHhEiMZu1EtpWzk9Xy8Z+U9AolQDlJbMCfv3Hb1Od
SC0NNSeVn7mq66J7ObIpkHvKOV18PQF/3cBLuv2+Xm+MylnGvSx15/Ks8rlawA8FuXlVAmt5AjXM
vMJcvedO81O22sn1uS78SqEhlJ92dSPdia+Dc0QikHvhFXDOm2LvNL1rsyBWKHcZK9v8CMkzJW4w
je56Bs2LYQb6DnaynuGtdpazHPEz6O6BRhGxAlIF8wydOICb/naCcDEgjfKv8bgE5nQR6hnXsUsM
avp51DU825aFAm85+x5zLtp4Zi6cZ2McTuyU6+eA1cf1E3Gdqa0yS1TvzXNruXgaKfwRzbQKW98Y
vX3saq5KSNHZS5ySArNq/9qF+C65TkPcrT2W0gbg0rhf827W/LaCJjfjrPNY5QI/zD+J6rEaX6/E
DxAPgG9SWoPBpRskbBXyWgnXMnJCTQZm2xjJLo/6PAbs7bWOsxir2O9rQVJh8f96676IdZcCZZEH
mXQSsKqS/2hvWLCR9QP9OGjPRZbFnp8VSoLh750S2uZNPaUz8kXq0zj1OGsgEYoN3iAKOKGOImGQ
XKY1tmMvc0Z+LPYZFTVrra/k3FWGRhC4ckFNX67jF96fvqi1Q1cBFbC0nHcyXSqVm2RX+/k7c9qg
no4jfFoj2KrajH3tjEM+X0GHHLznM54ttzHV1oYWiMGGqS3VhvBtVmXL+h/zBiqu74jPXNMqf5ES
H21wjN51pkVnxQmjaJlHw7XQ3mayWYj8kcxIfOurYl20OV0JgeZ0+3Rq2J/FFmROLinCLSxGgB4e
tM04ACZ/6OaLKtpG16fzER5I2YRvyT6FQFoQS7K645z6OXk6JtwnfFBoLp5Uu7gXAhuTvFohI5et
FaDN1AkmyWNKemEKXTIwq2osj72FfVOemiL5ERIE42lHoxeOnliqJfrOE5Vl54070OtZQLapXgkx
+XIvb5zZDYtvUnRqQRPoC2nAV/AKV+9CkXZzVAcyARcLq7WuDT7xpNmyyUrkAJg/I+FcA4f1jEWV
Xja+ITWWZ5SC98W6dbPAlhEmSCzKDtBXo6WYaUkH3bOdlCCmcPW/U4p31WLLCKnkROvep+C1OGC+
N+qXzirU9a6+MPDGghB2GTKUoCTr68qhAPYljsyjwe+T00aBrKnMzCE7dRC6Vrp6AOhuSjNr6JXg
RsOtS7XlF8wsZfIL25iyU8cJ/+L7WTgqyIAIiQPhtgNnJWtJlYETS+Ytgu0+YIymQM4CeVm8PX01
TSfo8W9Raty2LmM8UyCtXmbI7hP3Ma+1A19E21IKNa2teVQ2OUQbWhES4BO/8VO3n4EgIlzbdMm1
ysw43QYXrGXLkjD7FT0WY6TTB2poZ063/Mx8bACZw6jpxaYMVGgCze4gymVzKVGN70u0Ya93701e
gtKnb/VIl3izVKhMelf+167Yg5xwmjNdFMuF2AFdFtSOPGq9anebqlz9NHZa5tzrqcYVVullpmQF
+rr/7vtW4BI9VYZy+JYbMEy1wWdPW0tfxh4gQgQr6J3t1NZ97n1z5DzeBKevjlbnppQv7/XErqG6
+FTx4rTReXViSLDEI8q6c4BteRm4rMNdNX47Pk/OCl9uyFaDCs7u85NOqu9nn3/VVyJgPZt4AyZi
n9LnV9+DEq+ZcII1F8OXTzxN/vjhxz+qCd1xNrOq7b9tF+ahxOHfqp7LWdDh78iy7CWCZe8VKrLp
dFBsQP4qof4VkVXgSIIUbMNPX94Xh164KlI2diW8P8BRHGgbOmYlBU4SxBhLIjiLyiqV6SQxJNOd
tSeBB2MBqV9G9DaI5aVE3t4p0N9gEezMr4nfI6ymeXIad+Iof8ESL4VhdEpl2ZNjXFE4Gd5x1NPA
VgOeUzfK2xlFFNLaRvNqYU/8Z8/96j23nvJBhPFG+nLU9Kww2IZB76eipyBJrWNFM6vXAexqqKBs
c8m0OZhEV8oZ+hoPTaCT6mpxqEOQM3ga7TwegmKYBffIYucE2WI4f3Kk5w5QNF2pIN1kr8FlPBk5
adPlVT0mQUROFTyHEbYUYgD1M8v5+qiW0Z4FIMGCVMhGJEVV+VONTeoi5jyjWjZYC5i236LdbSMs
unM3HvCJl9l/EP4FnP5JShxZTYgfu9KcQDUYLi03MyszpCCTpeiN9xuDf5Hm2KsdAyA9AatnEMoh
GW/bpz3VeOJTF/3v8eeTdr95Qu1VBNv+zjUgvWO+LJvfO7xbOZyjam73dFklshN9oN/U8k0YtqYu
GaYjuWslGOqk+9x9Stq65aPQkT01gX9OjyjVQbjSpGjj4ngG2ffI2AfI4IDdKwAcE5FU8O3ErQ41
70YZzQjwMbP5lJvle1XRIHezRb6t2IhNGtzvkzvnHeiyCvPil8Qk3F9sc0MYFslh1ZvyB0CfX5ne
gpIjJ0N6d0MyCEUtxgO4Qrz6CEu8p54uOeX89rLLI+3WhQzGh6uPFaKC8BA8fXKT9czNmGDsIFqA
HIcADku/9UO0l1z1z0tM12+mHexMHrozZB2R2SCQ+R/kHfIH8TTznkZgPbKFiTjiIC2drkYSC0dY
wbpqwUzCpqi91wocYhuApk9XDriUtZz7fHwtcOfNgxjy/M7oIttxUFoKMi81TNqzt/WisCGZdb4x
8PbmJGLHqCCRF5qrvmFRhOEgelEhoUbEc8hHtpo5QU1lofF4Dmssx2DZtD/1PTq8a4jIGKHDQi6Q
YNxOwOZv6zjuH9bF2JPsMxFxC+xFMgPPQVwKJISeTU6Rp4a/RA5NEkJmQxwr/H3IK6A9p6JXNuOA
qEWOnH5IeXm9dAS0z1A/bS+k0figmlwOshbvkDQTlqeWoUEjF/jcWL/eYfRh1FLT79bbMOopwBoK
soCdjvarwHACniMkI1nCXnU+rvFj93Y85L8R7YM8KG+dz4FHYE+fiX1zDQ52n4Beij4SRCKDgJSx
T4ifb4C7CEsT2WcZMnPI/8JnC/tzhq8UQjsATCSYT005dqAlyw1wF9k/1zN/YLGNfHRIXqCHAtIV
l87MyH42EwsnSWvFrEmsUH+KnLTP6V4yoHRrWUG/pOO7bJ111OMxA/cN/W1298o4E//RwkeloP8M
cdrZFio+X5DI3YMg5WXAdl1mQvntAzwoMxWvqfjvj77tM8DdE+3oO7YUU75ciOMfZcZ0ZDIdMd4P
w3Y6hsOqj2LmUC3w+QIhOsUGIXnpCuSv5HMIyVGUxHqA9Mrnx6KC6Qx81YRfMl0xMh+yeeayilvb
69x3k4jzcQ1IJ5tS6fFIvvCQ+9UXqRe8vndJQ2/MiDCUadKLHu9yvcfNDOPC4gV18n+pGmOyZE06
I7DnzzqtW4N7TZC1oR8NEEaWgqacN7NonVD/lbq0S40OEqtRmcrbn3yNorWqTOckPauV2nHKqpxm
1x/LiBhwIsZeLN8R5KarqoDLm2psQ1uiJZMsJWCTRoW5td9sfma5uz15XsaW5myl6WXfcIQvmONF
5YEQ6rEh0Ng1xm+khS2NvqnSST531aV01dqQ5My037F5mdMrT/NPofY8bT5bKQsyTWoBAhzH8mNE
1x9ASfFiElnqcnadFkKnMwqMpBWBQZHxMSh/7j/LZSVYIByqFp2lbVgt6IubXNULO3Reo59BSQNO
ixUE1BnH4cOyYILDDJXbBpgyEHqwAWc5iuSTUoeLy8dn/WLU5x+VNcmumjPI/2RcMp+ZMRvf+4mJ
LeBsDA5gc/tlUrWKapDRjuSLtMzApPR2SWZS/5qXfK9h1Z53qu50JPwCGDO0X9DKwwYHYGNGPiyV
HaWUqisKDrpVu5BwyL2/bFNrP9OnnA9EBaBUQwkO38Ge44aF5pUNh9PRU5/ikPK+KI/YVfXLOjJw
XSTcaTTJPm/Wy5OLe5Kf1AFQSnAQkEJp9hAmz3vktOX6bkmHus41VSviMdhZIDWU5zEBr9X48MYy
zfapS5ucZhjfceH/2IAP9gwVmiawm144XuT9ylPnQ8qflYb5njVWvEgVCgeSSxGCmrXnXlkUSMBk
w+Jm3fuwUjEo2j0pz4KCmztN2X48Jlrriz1jcVJU1DAtn5y8lpG2a9wM2p61aQ29VCRKaRwiTjSP
9c3SNhtOXAboyB9gTtnroh+ORQRcTtLe31sgR2yU3UnMXAHaUUzQ1ReqBoXQa+ixAuOUNWdMNt9n
qYolDURZN3jM5gWypWRsx8X1tiTdX0I2zp5q6eVF34uVLiJTaOCCWhvg99C3fSWPGp0DnKuWxHFV
/z67BezqpjTyIa3+y0UJuDyvGsqsdZu0dqnjzAaKgh1H0s9yIdOTKoHBoJKvtpRUvREs0vVKhnbr
ppMqczx5owevWpYMLwh7NUqtI+yugZ7SsIZ2901Ha4IsZR4uh5gMbHh0EFvfUbUEe3B702p712sP
X3ILna25s9rHiPP+2pIlYYtQYWvLy4BEoUKU+gh6DDIRNFsB/BhGTOo8KT0wZdfwS3WiKZmumKlO
GxEbMNvbeLQgodfSyXsVhv7w344tYusLWxRiXvnrdzf8D+PtuGTZIQlxAhNLp760ej2e49x2fHH9
5dYsRBLcd50eZH6b3U8cEbwsjy9ZJiHXTd4/8zgW8s2bT4S/0MpgbUedd6Bv2V2lMlN2e6SqffX4
UZGIZ/I0aF1YxaXfF7mbAS9W5WY+J72HA37U7V6QGfapSz1xF1qGdMaGbojuPPeHfpBea8ddZKbs
hJhvXXKmtFj4OSW41RLHXkdZpnikbesiDBVmvOmcIr7haXrrDDVHdp3x+f7ucfC5S6E7CS4ZAL0N
ozYP8UZ1IwovAOqGJ8St5G6+zZbcezvVHUR8xbNbXPJOrRjh+AfedZv0z4uvAagzr9HiTdJ/aMAx
HB++z805v071ljfA5G7M2QAdXUC+KL6gLxlgmV1GpulHXPYTc4VO9Wh8GSswx0qd0oHe96uRpxy1
0/roTPxoaMG3U/EIxep6gN9AKPXpDWhVrFzfMCfGhQFLfzE0v8CN/zfPLDMhAIjq2XICdmd+s1wc
g+OgNifPwWwzBPAXkHLBNa8k7nIsBkC4Pos9qsotTkKbnlkEOJ729tq0MeuuF7F8kyVz/bz8B1nI
ghgDhEZztAKShE9GNznCOB6i5NYZ28KUoLKxXWYck4APMjm0fJJ4dN+vvNIxgnj47H6Lkr1r4YYV
khMyDKk1v6wqQSnrdD1F8IAJu7QC3FX2bhIOki4pY6Lypx+97cNOiY3Ew6c2Q1S1ZSpk2Sxa1jJr
9If8vsYFbzKDxc4q6OsVOk32K0Y6nq3eZfgIJAU0xmYv5zINxDZGIVLNuK3jUfdjCGxkWW9ouasP
Z/gwLrbDIOEuhCLDZMtdDtDz7EznpUNP1rFUKFe4huqyHcMR3Ki7NFeYMIB4bbbu+OcUtPrwdWB7
V7+IplWZOtTbnQKKc8QjcZFeygU4lOGMZDPpis4CrKC6vNBNIrCfz/UZ9oUGAlGU5ItMA0JZWmiv
NYY0kJP7n/jWjSfgGQR8M7GlQGtLMgR+htN2gnpvI7bFlbm0biPGqg16WG3StysKmDUvdRMsFY29
flkdPFmvXrANA+oERWA7oj695Ui4urkzjQDzbLK2q8VPXzQzO8lgiSdzoOKKi/+cQ8oF8uMdE4Gf
yMCN+7Me2237kvCJ3wPtIEROs4D02cH1pY2ol1LBL2DUUGsvpVMbfJKoUOEoBRrMt3Uj5ujOGwCp
k0LmSg3jHOpV/IstqWLP/fQW9og7eu+lqtVAnIDgTDt574hMi6a4vOOdMhXRhObxlGKUkFlz1CCm
QPJw8r2d/gfFKr9GH5EwCJCnQGz3QYPrV2VXADcrQU4viEw7qYWHs/mjs8EhTkIDHzPXe5KDZtD3
KHjH+WMWsMe61yDm5n7AMaxNDz0ZUCyL1RSaLlgM3SOxsfeYMj9H8ZQ0NpO7I5/tZEXwWYDN2bRa
wChWV8Qc/LoPuS/sqQoF53c1qs4Umxe+cL03lSum5/nIwUqkd+3mjsi389YTF2QLke34+oboy3k4
LdGN/cQs4sz9ooxmIzIhJGUiZvtoP4QSZ6FgAc4qoLIN9rkFLoOv7jgaZO/GJ+Xd+AGsyBGzes0K
yy4b8ro8YfgYPAzx7zGkZWptSD29y8+70NSO6b2MRrM/KnOfM5z/m3bxfIKB4VR8owRgnpeTzcKz
ba5kvpg5IBBjyITTo0cvTa1ueA0C/F7HE4rENyPLpp6HO1murXTqBjsiJBuQaklEmZ5uNYfKAWa+
ZpdsVqyeS+qQLZC/mFBsIz88zSUlpMEzlravtunFLkbQ8T/2YBCGR1bUxCYhppkHgwEK3M0vrwDP
uF/x3jzmdC6X00c83lDHORmOWzWsi5xvd3XtD6iqNQ4SJlYp5Ec5FcKzO1olVrAGelakGga2yc4E
cYAfaKkK2wUNL8cMrjkIy7HZj2HVuZ87QfnoVTH4BICKe+E9BRX7bBQfAVCVhGC7lTZDDUx458IB
DiOz2M9VnDgNE1vUGMqsQRYjV/MTU11Q2UJETEv/IVjD6rJUXLJ2b8IJXvnfQx1+kX0Qulbkg4A1
Wq2oE4ZQAIvFZ/2zW/6ofprJDBSUjaq9hXDr5xpd+3QP6cMrMs0H8RNwfAIjRL+oUE+PF7uisRXc
YRN3QT8c+ESeTi9olnDpsLPwMCrFZ5U9fQV6MbsEmCfY7mTu4ePsJzuj6jC70pQoeMjYfkRSqrdJ
4u2r9E3915vQAU+c9dTilP5AmrZqxE2xg69+unWr64NOS0bZHHQRlzS6o7QNJZPEnjPTcHEtGGE/
jz1SAmVgLz982+Czrtil1le+A0Gfe5jPI6Dims+7WRHnMqENnvczWLJ3Yv6IkpNxd/MVitZZ2PYp
lgc89VBYJxsQIWc8Vee9PHYKcZCTaJjqkFQSXXSLFkO/boA1l4zXbAtXURrafOYKnnyaVYDyaLEL
gBJfR0xRAe66nX3tYO7t25a9DcD0M3Ed60C2s6h4z+1SqlnJN7EPNsvpkjVBUyg3kVrRfVzD2YAQ
H3KahBbMnBHRTGkW/5Lhx5uCZ6lRaqGoI8PGvqkCnTwUBWe66JFCBDUgpYB+lJPGIjIXIFYMTKK1
xQ4nsWkhHJdL6EmTp6sbv6NCpvRDcLJhZaf6P7XDo3T+U9MwqBNBDG9BGpOvSYYgZK06rtFS8J8d
rEiuG/aOjptpyHIMya3CWbj5fDED0IQNU0smEZVPpBR8bbWj03NTc/PUikHo8x76ewQdDFE/hqTO
Wb9LUF3HmqoBz9Y74A13Q1YfbzLYXrsktWfEf+GIjOPQYXDktOtWZTLq8RCt9cTRqUnz3AMrro8p
tPBdrdBtXQBwKB14obpjDC9mzDBHT63c0L/JcadV2kRbwoWnfo+YHbfDckukcYfcNF4G8h5UlSto
wzycD/26mtdh5PUxXB6gEHpRg5TrRfwIK0X9N5vSbhetwf03A50pOY2hNRKFftBAtuInsLRXbE3+
K33Niq5lLrKvOq/Cw8r4tUqGdJa7up6AmeLktmlMHDpEFXZ7QjWdgotA5KsyNFyLXs5ODfMeezg3
nOiAzw1jtrTjd/oIHMXvqMFoEDp5fbS9HprccUFjr/CkItRTywO/jOfrnU8cdVKsNbit/7FWrrYs
6GiAxh7dPKKGB+pzCIIu82rVtox4CWHllzWVF9ex47eKwsm26Yzjpy12pyi0BI0da1tQP90PWslj
cB8MSbXxOXmglNoSOJMolbTxzpgdRgoTp6/fbtP/cGDdr64CCsE/ciYB5gP8uA8X+VpKZi69aqmp
Y8Om1P0jsSinng31bg7sY9O828JGYxfRhzKmCyoubTrtq7hMstWGB4MfE7UpTu2EVKKvuE539z25
qhv2tHq/jWDX1fZ6ocszkBWEkQ3Gi5Ks2foiIA+L1rQpXOsrZkwQHjYKVaqP2EPG04BNratq8qST
fSNbylb5Trg45kGwAYYFoPF6cIlFPu+IOw7mDoa9zHusq6FboO/kJCjIWwjVgPQRSeizLrftKjVA
CwZq+WK4/wN/UWx6FMB4RgMQJ7x5doC1tVvRsZIgPzf2iscMUAqByJ7kHOs+GRCTLUYK2EIM2iTK
ywGkY+NAim0JBNbfD3tBdqgRAecX4oZ+sK5lUxyAb19foZp15PmeoYan8PiahYxh0ZMGP8AauNWL
BYUWj6ooISzdU41LrOCdxLRjMpwS7XwH7qj4IZ6lOERd2milLexMXS7pP/TPETnfUvPWnrHVTCVf
76EpqLovr4rsaZ1i+MCP2pkLDqv72a17oMxaZYCjLnA3hLNR9YtAzA8Ql7C0HYHxe0dviyLnHfLr
xc1/B4T3IqBZRP7F2qWVg8KdLdWhzLacJQOkcZLWicuiIoGLVjDA6v1L9QKXt0oLyXcniRsvPfE0
5lYZVtT24PJ5Tw2mFZab0OdIn2XaimmIFSPwnRZMjvI9g0ESHgDuZr5PmqZyxvUMNVAsV26uu9+C
rJxxWHWMtV2Gj0uKaIoqbp2N2naFCCBitrhFM3kPIUv+mxMI9K0d9CRciHq3+NthAFLJgss4GPkX
heOkw42slDvI9oAkWRpbnpdQx28SHg8NMQbYiXo8w2W6YSNoFhxx9uSH5NB14kZj1/M8hz79WMSM
tt6AEIXnsip3KVYOTe8Cnzsvvm8nsFbzd3j888/41v1tW6Drg1xgxwpj1//THpRIcN31MHSZCcSc
8kZZsghiETOsWq/HTfrzRVNFTLxvFXrZGHMSvU5w2OdMH5VwzrUup8FSnf6tF4VD+5lhJVxmEzDd
hYKr4UehX0BhW3/+JG+8Ry/DTW0B065PuLvmVhoNs/qgNI1P449clp6DoymvicWZRS0a+o4ROT1Q
oe1DQDfSBpfRCODirFeHdhJrXrreR32hQ6uGnf/5PGUXJXXLe6wmJmyPOwn/jTbGXFjLy8M1CUEi
RjM7XvoXn+6fxmP6wr9/JN6/6SKlorPwL4ntZ5DNkF10f0Gh/WlxREVcspdks/dxOFPPyclpv45O
tt9pzolrCP6MGuJ8tI6H4Qc7IEAU49dt9en+EV/NbF+AQON6BidWfSLxhj3vDA4Ha7Bo9KsOx8Qc
boyq172BOtnIVls29Kwk/aJ0vDWurS0V/hmEpq90OUpxWpTcwzlI1XXfL0IC8J61TKLeWNlUt89A
cawDCOPo5JnHZcuMgEuvbl8R12YPQ0F8HK6lfHy3eNucSmy0lAYicHG2bqKCLVrwuEbJx84DliE/
lOOm7NyKLZVB/YAbHMurvJtE6VuJluP9KegC2YFNStgwYBhhBn60Ei8xpfU7vOp7xtQ2kWP+ll9r
xb8DfdwQRMgqLsHasBBcFd6SPBcUGB8wdNi4r/foYSBFg3hAI8SBRjlAs1V1/MTH8hFzq3xtQte8
F0rb2dyzklL1torEO8T6dDV7VIU8RNSlur99F6p6+QX0Kn/vVkXokS8jVd53pIT0kLqbw6fUXgm1
3SPlAPIC2IGcQ1Mdu3Lobgcsl4Mew89YvK6DZqOQ3KgWC40DaVqW9yckZroCk6qyFocLlNNxUjUy
HP0OALoIIc/H1e4RQ5KHH/prNfXpdi9DzGfjjDJrYudw2ShahSEoJZ8TXQAXyT6hMOFiRN5j3uuN
g/4S3OYK0ziX3ei0J7hBR8SEEIRMKz+j6UbWcNzQ0CdQTGo+sQQRj0ZN+5FLZV8dbsQX+qmUowG0
XTU4hzgSZbNeMUloEbJynPKMwtKAktiubdb2luGeHwmWCR01ZQrZeDp+h3TnzE693dECiE5Kog/1
W+1qiruk5OIJ3O2GH28KeNTVIQG2ff0C7Ps8uPEU5xFwG1d9jxJoYmrhfoZrPavPYATMxnNcLfIR
iHdEow/0l0RVWZEwx82rEg1hVlWsPYa3eBeTZYNN5QV6p35SnnB2PbgPUcVdX/MoqyeeX921r6pT
kgoISOGgBbq7me16Ksa6VrjzqXQpNu4byHi8GC+CQOCZjDTccwJqHrP1vUdnJ7dhySBJy1rYxdsG
F+LGDUv/LUCXVeBBP6Yo33m0tB6wGXXoRIihH6nOAwZISjt/ZiCRtfPkv+UhBPwgH5rWUGZZK6qM
KagL0jqThNQ0inVoo+JQqWPAGjFhFzeJATOr8sxh8XB4Vz8TZt+gLIjRggaqKWpl0/25Bzvbzspm
w1DjdwWGl370HaZ2r8D5jAabprKEZRM0+7YR0M0FxqPhtLfT8phnu9JuuhqQagsMJ7EJ23plSqx0
uM7ySBg1v5i+vSQ1m2x5BZObIVWdZ9oefkUzpIlHlH7O36bdjkIvEue5GtrMYSxMh2XrzaG+OXwb
Htom87C73lxPqe+oskRXBHHW2aZ9CexNubVEV4VN/giCXLOadCGZ7L7DRvSmr34Tm6K/TmGkMT5N
w9j+g8NdoJExOJj2BSXA7ddX4NNnJbbIU8au0rZdwGWgzGDQF7uB2EGjptXRex5epetqXBU7cuty
5RadZgRqz2FHbBINggCncvy379xTTrdpRjJBUHttz77MQAcKoeyb/lKrcHnl/6dRM1jQOb1QgRFd
jlNgg7k4cEv369dpt7QNm0TliS38+rTJHklM2kR1SfeaYBr+tKvBQqIur3z4JCcnEIdqH4S9b9Ej
1bayE62EJCl9PCTC1/lvj2GW5TfhR4vmlPLV7FiLGfaAwd0++k0Zrn5YhNzQPQyTYOAkyjK9IoaH
BOQA0zSb/nq1Yo0o+3v6I4mIHWremvDNOHx5nBjetHu7SgELxWL1kT2M5YDD52iJvGMFBioPVOKW
4VMwML0R6Jx3wHx/IF4JyiwX47ef0ANSionsutWcIqT1yjRygmSX+n0SEE/nk1Jh2CJT0N1IsBpT
M5DfDi50Ew8yXzPxTjRyLr7iC1MoqygThxQ1G4y1tYcV+YkvT/OX7ZcsRhe42MotVzFUiYK8rsoe
SVad8/k6UZw3LZigB5CtoB2UWrF280ozuLnRjuNL26l3R0q6fldTFZaTMs5aTOsywhc1xq4A/AB6
fgE/TNniqs7OEOvfDdpXPPR53pBk9GZTGR5ycyOxAnDshSxWXpews8qmGYq5vGY9aHn/thArOpsw
qmRxwZWokLqotxpdjWnEO85xJx0pJGFH2OJk9UDliB1ZgC6dwbq6kQvlNRDiPD99GKrVBQJws2EF
Rd4MOAL3cUmt7bDDy6EmKKDHyE2KYA3GEh0qjoeQIbnpxKGgxsPQTsFwjzTAe0UHJVuoCrGM/84a
Tp+CrebYdqDLHJwZCIDmGQ2VPWYRF9ycDAp0/OLHvgK5e0XDU97v9MG1T5w29UA2KYY/WHRYO4WH
41NsOGeFaIJaPVrCKWWZ7sR1EumOS1V1rITnP/yUTeGd9jbImhymOPUl/EsF57tVdwfL8sleHRjr
Py5FFMlaTtGKIGKtBylFT8emufKUnealfp2yh7AzzJiIaaAme9nI2JPclMLSLVdKd3ZWxW38agD5
8IyIMgG+zDtStfv4q0zsNn3LECo8xHdfOP41256541tL+toODtlFQWpMHOmAnEDcmusdgdIYdvpl
+QjlfBuzlMoFK2PdtXLYLmWysWFN9dGVSHS+XD+bTrNagvh1UOIYapmDMjS/AClj8V1ZE7/HCC6Z
OWv223fBlFHcRHg2R16en4yZ3QVbZHMgY8h+UjoBxBH4zMSt7dof5kSKppDhgLfR0Ll+fcuw2ZxE
Dh24bv0LX6/DTZRawq8w1Qlj/vTVNALYf6/O7cDr9vlRY4KOeFgCLA0BOxrHsnaffg7MEMe3x8bQ
vlMs6dWjhRreu+aX3cWOwldfpObsHa/tmXVv2KRepgGYfa8J3/YOOETfTpCbFP/F6tQBxDEs5dZ/
77SI2YQkgbqtM2PNBFnK44848VhSdTFPm6cYd87EiuOih7U7Os5ltk8c7+NY8AuaEa6t9yEJPfYb
eIBkxPTwLXlDzVP5chCcWztAyOL7PdhT5KSpLpXapnd0Djt9H/0wcXh79MAIh4byYr63z6uoORGz
wFoxXXCr/kSQ2wX8fV9I9XFF86eE9TC1UQYnMwMBRAUuBwzOHFnxE3zBHmbGZlYB3FZ/PoelsCZk
4uxHQXEHOtZ46BuDUv0Qlp0Y7/gn7EMo4k2d+EijAc1CJWTYvNSDXPqyW5FbSGJI5Btu9sGvispF
CzdF59bntDy2dE3LxBuYfWy+DlyZE3ZKIJqz2bosy85iZlXI1E7NMcobR4WbOqscKqRxalO/tGzs
O2hDskdGbqwc1s1c3FH5vTteqWaPfRnSq3dnpLTcq/nGrAXqA8uWATYytFXRvxPLA2yAQw+brdmN
TZHS+A/Vi5MOA3cmqfHIPfXhpglG4z/Bed7lGZ77tiXZB7U/5gW+wiJdBWgCImHBjpNFlbG4V9hb
ev+BYsxWybhdcJoD5l015OIyLVDVCnMvrG/otgPHr4AZ06on148l7OtG1uHrqyHrnec0VAb3o3Z2
+DBda95rAP8v65IWRyEOxi9mn2qcmBcTXKMatFOeE6cKCweoxwHVrrYwkh4ApBIZEHE2JWdYoxn5
cbCBYLrhGYmUKf+jI3Ks+gRgNfA/YlJDjs0p9eNhKLeGp+9HSd6xOlKsYRsLqC09kfCVaGQZ2Hbr
2J+QU35dlVQ4PD+LBf0tTf4o4aNbWxrKo64c6nbIKBeqBRmskXJOox6qdk7/KSq7cr+oSz41g+9W
DT0qftGaJPTZw2B0q/wun0nT+aOoiZX+yZlGo9wWu7vK3lONYaHmDBfABXGvFKZRrxqdHoj6thEG
jwiaO0Dpr/UI0D3vzoHaCoHKQ7seZMbsIOJkXhdLE9BeCN32FrzvIEOgdJWMFhL0DDUjPKVOz3RS
S1oEbo1FyTIqL/oAMa3ll3+cotiuvmxVL5Q4Jk7A+rQuzr7iMK3OCeWgZ5U4k3ttrrMKIwYXBEZ8
WLezp9DDdaoZTcwa2AWGzyT3nQceqx0FS9bpSzCwo5qTz16bWk0VQKrfFVK0dK9LchRipATvwzHM
PY5FPdxqoz8lyMmvEg5DddZTSYRrdFnjSBJ0CRfl5i1x1w5sVd1wAoJ+4K+Ee1oMJ7lJmNXPHFW8
FP58aBH4H54pkfDu9yf0IYZ1CvD+q++1wqaPY7redaYOSc5crUPTgj3p9i0pTS9Ud9v+ioVZ3/sq
LFhJ3LDPZTk/RRsMsAHzU1rhwlcFbob/cnyTQRZZZgzAC24rSkD3SvAcmZs1bgThO8uAumg9Fz9Y
f5MkIufP1z7IbIjrBDZc7TBAaA+PEJII4ZRtbNtU50w7/y7oULSvhEjHbVhHUnYiLZCm6NFq4/MV
IcOX4oskuQIImfJ/sMM0UNGGpv9sqsl5CusJG4Yx+FgwYvfScArAORWt0677nMhN5Saf2RJ7EAm3
ezVRUSJq63Pj2mjzL5uRqNOpuFy0NvCvgB81XT8l9HIqNvAcqAADr6hGaDjd295eoz/SrhDAfa44
X4xzdgVQDajvNIuic2dEX3jxQurFTagR9tStpoc/nPz8seDd5eXN995+oBcWzXG7gWCKxAC9gSZK
nRBKn7omz1fLMI/sdwsuXGKareh9YAlOmAQQolGk5gztlKJh/N8WANOJQFnTeqVgn3kYP1Nx5+zm
NsYuvXWs48+p3sZySqUZRCmw6lUDqSzriuxORK9D93Q6UU6IwI0d4/qWj2nlLN/df08x85MrK8ld
DW1OWfQBhoUe8uukzmvLRcBzOmLXM2s0K9JfXAY9UKd7QbNVJf9Cqv2yuqoNL4AizAEJDhAKI6Zs
FNsnQc6OSnVE2CZuatN+bzsyFS0NokzKCuPZg5sphaLx5DQ9Aj2yoEI4qDPsqHfcNfnczJYYGwHQ
F2PmLUWb1yOHU5DpHCpNKLSb4mZ2/+DxUJsX5OnuCkVnHs6E6LyJVdnnwx0oDd57qgq32+9nIkl4
9HHQG3b18vICaAz6+c6mkbL7JkAc6kNvjUh3P2ZtvwgdTOXmE2LG085UHF8hbtSYTmffcnt7wNF3
tyooQ82YIAoOarARFi4MpBGMKG1EbK0PZPIPkeiKkqMhriP0H7gbGePXTkhg8P87FVrfArtOFTAd
Eg+gUl1P2K6atZrWz8c01CWdE9ARZOOPCv8h/D+YLfSLz0RlyPFIu5UNkBlW2jN8/Th8g9LZUMvp
yOcpIglb9eVl6Ck5/GkqkJ9fXptLxhqnUIF66anEeK/TG6wzGWyxeHnhbz36WRlJ1pj6rNEBwmq6
jx9DOjw8LyTbu4uhoU0mOhH744HDj3K7uLrxuRwScQ5w/E03zSp6qRqnmrAKcjEz82dpXHUStjev
HAg/vs9fFE5ilm6cyPWV/LUBF5ofN4mHglJdH/jku4If6qnjlljC0lQfY1Mg/qHwe9IeHIdZ+Icb
sQB71W7org6q8dCVRKPdEY+1C8JZb5bgz8RR1FRCz6bQbx0VDdEA8Vv1Ba77qpfLO27p088pgYNC
70uGGx5jshvIkXetjnp6AL8LAAKpg6ygMD2aWodGOmHRLqD/U0B10MIjszqgdADlCmdkATC6mUkK
VAv7l833E5fG5Aw3LGSabBjlKczqwKOP7t+bfMZOmBcYsyrzZ8m1esB/jowxva5TAYtZF9li2mNZ
FlvHvvUoiOCpF7hapPIKMtgw6tpO4SFHho/gTmVg8EvaWDfE8tMrw762iEStT3T70zATO11Eu/uY
2w58hhpXl2UOiLc0zNr12LtlOHzUvyP8IgFzTWj4F5agX7ib/S7XWgJ/KB+gbhEePtXPCXHuT6Ap
98CYLIHwaksP36vMW8G9HFM4hPyYOhwXYVv2yEpFHZOFwMMtc/uoTk1GAaH/7Q0+ODaSboRe6B2b
1xDbo5cj6K3XU0eyn+yMNme+gNF80xYzYz1Uv61Tr302foucsnUGO2U8ydXdEcC73NPOmTSCBiXx
ZV6xI24oRgO7+EtekXcY3Vre7xjCFowCQRCkzrz5oPZ9Ljrbjnhc1j31Ruv63qrvnLVXkFBad/Hl
IsA0ZOKT1d3Yn5pw07f+TOlP6KQ8LTN7dOTOE90NE16RbnF8DH82L8/Nby5Rwxq/ijdDJ0bdDKW+
adVlR+ukFgSRDyEUdmjroZKaKHAkLn8BtfL6H5j5LMhXdp2i3+jZsHN9v33RWxXWDELHiSwmh2l7
pNTZdNRgl+bziTtPfwbCRsLmQEvvDUbzgnPiUXq2xHtyu8fXCIm0d0nx730eo7PyZJOYrNoMS8D0
Fz2Pm4lhxG6Irh/+PTWbL9sI8NcyRYWjV//1qEQcsPDoNiJnKgFWbQXd6ZpedhNQS1lsgr1WBAYt
Do+0dgSlJA6can1TGYHrO/yJU4BvCxHS292ng1Fd9KRY+CmIp2NFjxuWm4QhfxDUQH7Ajs3yg9yw
fzkm08PeGZyBBWbFKNaKYnUNbER3CO95Qvs/AU39ySMgwWsT3VSlL7cihPUqJ4HJCFaw0dXr9i5h
ByM7WF5ZHicv1f3ceKxKPco9QlhAmz5ATkSRMLuw+JYXrYM1tyeD/TN0ky+tmp1xO4PFr3fEVD4U
3rQR3ZUZIorVaaddqqHJgy5nU3bNXvgCKzyIYSkw6VCr74eEmV1uBqSEAHZnmrDSJ3X++rz4NI6g
ST/A/pkX7bA0vIK0w0qi7Qchb3HvrL+ERyw6kd18HP+OXkGcfqaGTmkidl76gWTzeAW1TDtpwL0R
IFpl/dvWq/5zk3q1trTjMilaybRahtUuxGI9TUpbAobyjBh6tHuymU/HO9fDnMtLdpag07R8jfLU
vaEuVpxDp0JIL6YIMhwFMq/pZxGbK8xPLk+6PiO3rRgiuC3md5bXu1TXGHaYoocU6ggbsTlkQmCn
5UrtnWuQSGV4SY+GMGqeXUSieKc6Ki2FxR0bWKhtlDSW3CgNS6D9UH5ScI7ES/euyfeppMaaCS5X
YCz/WHFc3f8JAWM8QILqc8Q84TjW7G36xuoca9ZKrmDBs5moo0TMtyLV4JKqvGikNMBO9Iw/Hlw4
05IeFm/IJFevAJVwh9wLv2WzoZsE5Iv2vonSaBR1ryLzUicQ5B0Gq62SbKSz+uG8MfJ8tPi4tYeG
Ja1DjlGF9xCx/6/Xvz9vQw0zknAyp1cmWkWZXcJFM5dMw5r96fouGtP72uOa6z88EbTlfCFIjVrv
2DrhSJyPHTklATjs4/VLYboh6jz5Q/bcKxdNDwyzFwC5LyGU4I6Q3WmdnrG2S7gRs4eEfCaXh+IY
3mdg80QqG2J3H7vKOhXUL2EnKrOgQdxs+7Hv1D2MNZGL/X4qq7P8dZoxUGfGPAvfSO2pN/uPWvo8
KhbDQ2rgzZJYli9hm3IiMQn+Pbgp1J4ofz6bD/lUUmXFejQtMEW3yH3+9px37a/8XQ1HRhndjWzb
EpK6ibmdrRDNmKH3f27PfZtGo5/rJf8CPO+1iwbZP1O+3t2VjNZah1gDwvHvlJoZhC2T92rZV/az
tptFkyUBxHQYW3UDoYym+TAaayqLO/O7Th/jDNm+7H1B+KwKYejsytdpSpLCi5aVVj45BdCHolUw
2BR2ckilg558EjYByxomel2yNR+BXySBUk7qzyEegldELazbHmGxLOxDgLgz5WAMmcrPd/lOMa8O
B43qqK33ZIout1hAaqp7oVT4w9bG/C2c/hAQ6N2Tq+L3d/EqAQcllFStG5HUO+1JSZtJdSxc5kdF
gFW+bjnxulYkp3BOuxek57IvCmkoLUytNxApLe5XwnhvtpXfr8Kl2CYVf5prnyWYn8UUPMOGe9Ok
mShyQo/lc/Ci1v4JEQH4/BxO3sN3m8+/dnmBPfrfhqP+hG8sv9hFAXPhBEyr2Adyx5Gg1aEXO4Rw
MNAmvVsb8voPHBsuc57jGf7fgeChnrHWEtL9awrbSoKDmZ5KMUyRS2vDR1TCfU4+tTrUeFHjpseg
fnFoJExf/u4bnpjmLF2xLvK5GcOzEbXsd3Lk1tzy8ipXYiaIfAeworxRhbGwe47f04gA4UPENrKw
Wx8Eel0XzWBLAdCB7hBl8Gegbt6r/1BBiS38CC/5+ferZCAYHLxyGQZNapNfsbALwGTHn8niMF+Y
Bu/lOWnRxaLbblSh98Gsv1scEA5+k+aChWm+HxcmMvI8u27lrstbZM2hAFbD8M6mRRofvBdUz67T
ADJPlquKv5itNeSeQUtOg/0CeP6cc+LmT2kqT4u9jPKeDIeW9j55ftbpU3bgYm5zRsVbyRORpd/n
tpM9DK5umrWu+YtUxyMX7oHvfbq3rCUZRsrY6ndx6gx3qbP5YZN2CSLl5LzoMUSE/aA2e3qjttGb
ZxP2480aiyXaVLHhUHdMLxSeOJrH+5vjypJ93s9xaWpIdX/IANWpyn9iPXZSRTDHGfFM/AY0iHxy
MKAzpYh9l8plLutdYZI7VWoLlcqhROUQjjsui3mX+WTirYg9abdZ3wPxDZT+OUZsvL5DJB/tls1M
guV15XQqdE68D2JVlIHZdBYvN/006xZdafV2Y3YXXg1sMC4OhQERIVo7jEcZqrZzrRzO7P2v0mPU
X0uJVNsxdfoyRIJROe4acFnC7fLmahWW85RF5fr1Knypv+7ToXgW5GCefUxFmFZ1t8SrNnNLTZOa
jdeCUzZQgDFOBFKTuijZuGYBqjdhjS1J+jFnsaLm3jr4Qkk2PSEmeDchcrbRyQ5FZPajUdysU2qC
yRONfVJH+CMa577rsfi3qFQ2dBFD2iRiPYMXmxHNGrb9BmPEkGK86uFHFiR/qSCQdwxfC0n1YEqJ
jSMhbsohmD6W0dQYZUqbQG6fYVBhUhl4Am7ATzEkNW62cp4Gj9iVJ5I01+Lx4rvv5wq+UuHPKdiC
iUpV/+uMx5KvFVOarX+fRzDOUeDbAt0RIdlBcTUV5PG4E/v4m2GHuvN50NkmFIoAJ4gErXPGAW96
ZPoRMsJD3EwTNF2/kuRfC/zcl44em1VyWnJRhNTuVQHpbfVVbIi15w1nb1I4WtQrf71TKdbk3gjK
pFQ5iBY2Szzv7foMBRNWzuHFOlCgrje2ZktRlrfBNBXNPPo4hivuwO/ZfW5dfEHo3hSV/1wbr05e
ZMNABi+BkSRIFz6f/DBY9z87SzRqUeynFZJl/C5EXhmRKlZSRf/fTakcJ9E09iSu40F9ujTdkMyp
IwVaq4n+6xkPChVTQhWbifzI0wjZulodddrUItKE9GeoOUTgeP232uAnkPeqHWzCmU1Bl5DbFXK3
ByHsdkMEW72DTDZWCtbSC8Kp6BgsJ3BRVPEJzjOd2SzYtvmmGGFjr6haiaeqzWAbkEGnTw82B5gl
i4EH2tKdwPCpTvx8GhTBBYCSsOEk8v/30A0J6jgPkljcX4iiDo6k+OuoxkDDMGOdq2gNW1lneVVP
+BAbUWZ5ud66Owlda7oI0e0gWVGv/XaRRm1SnYnuCR4n/d9FGPPlEsEEgpf1k4exqffFiyVaY2iK
BOV3mrCDWX5hWZG2eVNUD3fZe3ElmwmVEVCnIwLXxEjykglCaRJcwWHXkRH85gjccmendXfpdUu0
3kwYVvRlBcSvYW87hmheAm7WuhINNLLSDiGFHiOtphDGj3RSu0UWiX3zmaAxfmKMld4H3uNFD57L
pMzkAzaXCSV9RmJcTnHvFpzyQ/zd0eOSeev1YfSKRb0f0xFHERMK+oS9H+akBReQHn2CSFZJdqbS
PqXi8l0eLXqGvZE3Frhv5BaZP8gvFNmsoTQOPjpNe5QqPxlIyA6rmj7uj6RM0knoSFnGjZg/cxms
Nvm5uuXNTNz9p6c7JVJ7D2U8zgpV7Y+2Ms0NgeWY/YL/S3NZTZDFwIUGt5ufSzw3ZWkYEsIs42uX
iAJUlWzc5g4xUE1a23yRkyteUvnbOFQqQJJoqeGTvyYYaFcViq44s5wFnEUMEkLlX16rkgun2qRo
gGJ/AQX1+AK2g5W8ebqXmjwYIyIqJBI8Q0cxXlPWHcUw/MXaLpkTtctC8Hgre8pyqId6YmdnqOHn
dbT8JNua0kgKv8uRCwkBr+xQFPTOhZwjwNaBeA7orpbDvPmgJRclICoqBt0uQgobAIFjwREaTu9W
43ZBzEq10mQyMcH9HFDe5J1OlVkIl8K/A9ez1X5qK0/u9Fsv3tJETGsgwqeTcQ4ffMPjEAbhUFkd
5xEXch8QC/fc+iASKGnPClCCkEqgogItYbFZrUSxWathWdw2scAKWDdAbl0EotC9wo/AE5AXuun0
dTBBV+cwHWp0yH2HZzi3c5w5D2/J3JLxglaE2UYAZZA6Q2zGdNoAnwob00aQkq6y7WttiedE04m2
2C7ypdslVoIwyjbV8dOxxGSNYtlwB1DIc63hYsy0yRSIjimR2YM1sZHO/2IznyLUo5O+CO1TWZID
M8809JeTXzLrEMkQ+rXcbD92cDlHdfeJ7c9DLdc/JEhbgRdEUVhXl3fTwdSb+OulzWeKw3A7mlMY
eGUXnMnCp/BBt3upYweVYGfCw88cNjngcmuE+8iTSgq9aCF0/+g14G3Bz6LqYqbHWuAZKGdEU/5Q
/koDmiICshP9XRdqq6cK1XAEEtdyadF1meAHlhLeFmMEtmt1EkAkZvmUinQzmyqn4FUl4I4EYSey
vOXCe8UlvBpCDdCEUMwMu/eG6dnKET56jtNX86fjn14VZo9d4ocSGvptVramb2RNEqUfwjkD6KEO
O0SnKJTyCUbweMPfgCBGk8FIDDz/0YP8qqMprTvs68dEUQEYgK9JhfsAlMRvZ4EQ7SUeCY6VSAap
tq9HHfocEkJfKKJ0jyTo84ckCypPVQOu65gee+7MmwmFHISdOzE+NuxfaNZWmLtVtQ3VjM9Xd/8U
lgpGQThI6I0P1dmb3/hJ5gd26BT8vuHipUmQ8dS86s/kTxNh4azTal8gKhivIpJPht5DcP/Yirkm
RUOc0EVeRq4sZfMmf6wMV4yhc2Q5HsKG0ocSvfNak2+PMJwtzLi5V+BCFnzaSzMtySMjRBPvii01
+xcqN5SfSKoTi1/lGCc+QYs2HfS59VoUQfGmP62SO1NZVDB6UKXnLbouyytdQdiRcr6gB2sH5qKL
oDIIp89q1Jhfr6UYQw03rXdkG1bIGcuUpXy3vG30JY6uxKT2LQWgoCSIPOHK5CweqMaV3D9KBSSM
ZdKA3oq4pDHoH2v+k9WN9Oux6fH4f63ENA59NH7YSQHk/HTEnORpFa4sh6z4+LaHKvRoH8x7qMEy
M+Xs/cmf2SsPsPMw8s4JvtK+cbVxdxKwVOEtO3oYx3PdgZ73ChU0Eugt2uLkWGNxBA70Nomto+wT
hVMnhmfetRrjekbfnJny9eyh+q+FXsVU22mZGonKW49XnU69U/dJ/bmRKH82P1+scYFj3ZOqOt+a
QMfPRlv+ODLEeDpSAIDkTSoiLQ5RxX6zAS3OZKNj2CCQR1zX9LF8gtWBzvGufX6pNusDr3mEhipO
ZQoEvXj5CtPACNIi56edFc+4VLxNl8liGei0brh+iZI+wuPxNCIGARFoUSNp1VeSgl3G9W4skcLl
DnZl2Vh250jXrlQETcoSpcBHsW1nzRuZIhHkK2RcxLGrGbIFJZbEJvnl0d22s9Iq300GjH4I56M9
XFb7hARev8+UxQRZwZqoE2YxB4C8w35cBAaCgBPPEHhUuXGvTgGqCqjQM6JVV5crm3DfthTtC67S
Q5qnr9crQ7xF1YS2OPvT4DkUUrfyM0IvL0J5ndHvTRSqFe3S4OJwir2+g0pM+VW6bkXU1k6W9+Iq
87KbaM6x0YY3GFT/smqS0rG9uY0NARmcLKQAfuH/4dW1iq1zXeCHn9FUkxwAciJU+6N7WTe3kPyc
sNct1scQVCxmpn9Un6xafECwn6BsMPJGYPgCVoxcDbP7eRuY3/KPQY8xwSG0kgz1wzhROb29PZzt
7XNoACcMPotpqYG6nE8WlYrCOPXUB+4tfdBQwzLd6r92Wa5PTH4Y3RRwSYHOxtSoW1p8oUUICCWs
5NpnoJKbH6iiOnXe7xbLHW3C0Mtm00woNBo2p+8mXm3zl9f3ZxBaqvixWPMz/rAkUw32wReqQC+G
TjCJngjzR3sVEF5XjS4T9W/wyv4ZGEERBbKZI97Q2Lw7iC1CGUmsepqFgQ2fGPFnkqqLljkjdXRm
s8zmUPWWU/lG49ipsPspWXHqs7aoimZLADQtXBFonqw2WZdnkinVFC33EBiwJoo0VtXje2H7TM7J
d/R/fJFwGXdaX8eistP8KZLtYMXmihIddM72zRPei4Fg/LaW5JLsbb82n+x/Iw5rOrpAZIJCHVzm
eaG2zIGxcmdmwIl1obpklTVkkkDQTd7bhu/vkRprZrSJnal8s7LdlmgbWOzhFHOSDTaTS5heLyO7
EMD21W2oUWzHP30pgX2q6SJJWA175R4tXadBh5lAaXx0oRq4CgBLU8X3k6KbFoUw+5l/f+rG+rRu
GfMKT0JwYJwoHRT7D8D+s5WviZyQZ3bE13yAzV2KlTmkkk/KUNpJCticcKtycmS2URX6Awl4RAx3
FGMVxWa9+PA8FYahc61uwVGkS4Dp9mfT0OTaZ9wAqf6pKMTvgJTfs8amHNNnx3MpOh/pvafryCia
JjxauU7M9SW+ip5FZkYcQPRvfZviYzknStXU+IxHNIW0NUoKFTrUU15sHfPzBcLDAQxjrCceTFAW
ZrfkeIDg9VXGcoY6b1drtixzxwfutJwUuow/CRuIDFjN14+aLA5M72tARBcJkD+jb6caCJaAAE4s
13WqQKaFzfPLCNYLj/cjo0GVQhZsa5k9ORxN1X0sXZyzYotvkwTR6RpTnIavHPHpOZ4m/27UUU9G
YfAin2fBK7BbPJlRvOeIrtWzyFw4x+DZYytDofa8dSOK/C7KZF4ljfR53ipHNr3lo9al/tavJMay
vtekiHIb/57bUKmmcVMYlKW3ZbEL5VcnbaizK6E2ArkPZ0i2wOkbx0/j6fgVCQLzShfrqkAjf/Xb
kTGonGP1A7Jv23pSeHSPTQZJ4F8Za4zminQyx60DqhAjLF0XAskiEYIHLtgKu+ZxeSPYeQm8tuBG
1EL6aSNG+aU/aa+/GUndx7LeyInASOkbGXhiHhsbq8vttf9lqhB8ly9ylxrg3PPkxcOagTwS9FEn
WOc0duE71p/ENNH2wp6PbH3KtqVAkS7LPyr47D0Rj2Ha81yHafebxgugmOAWXdyZLBkpxY762j8Y
Y1Nnm01UQUipwwkugXVhtY4ggTAEhAqsGsskPZ5zL85W9HVs1S8AWIiEm5bljn6fadt1I9/0E9Lo
Wx0okdrToNIAHgKnt0MlOB8cfxBF5VMbwqu+aURK421II/Kw6dJWXo+W0Wj5vHh2xO28NwiqE4Xa
PLJTCG9ITPrRD/cbf9Qlq9FFLkCpMT6ETJMeLX4tkmPpwv4C3eqJXKDPprlH+gW8xS0rGnXpr8py
Kur6RGgQwH/PMbynpS0c4uh4c3G2cLFgNaFM1OAWDvyHQxw8TbiYrgOqFCuh3AgGD70V45mW2vFK
d7j70oLxhKBJBpguqOWxGwZ6urhlJSpigDDP31LI2Xx2I4F/ZvPGszZ0plhoVGwV1Abi/m4fPAn5
C5PFbWU+Tp3aUELx0xbPbmtnDHuCiZbzQY0P56ub5dAVx2pt3vTtpZDCXF8ZIan19ea4WB5YUtZQ
E9joDPXoml5y07mP6KUKI/Lzg3CjZZf+BfU1m0PoIKiFae/GgrtVSHf7mbf3HdrRl1Re/P+zfE2Z
MSoOKHltoSPfQVZh6xyLUfjVok9gMa5fQPj9DfsKsEPvIkG3hkeZqwGeMEk91Lf2NbQSrP72eY4L
d71GRnCo/8HOFYgQSXmHCHIKZqIPIkFBLuh3NedCETIsQzlOAeliQ6gfnGk0M+1mMuUuUuLjcpom
UeLDcFt3fvBtIo7qNT5bEzIx+o3doGe2VgxKZAiB2xHVBNA8Ln49/kNUF2/qwSHZQrXXpBfRnhIZ
iGqFkDWOn6DAMsPbApIlF79TeYIhzqoCw9oTOZ1mJx385ZkagfqvQ3tcs9VIYTN8GWOvvZwkSjDH
K1tA8P0Mua8kZt3YH55rytkAAckd3iEPa9M2AoLKS44Id23yfeGWQlJnZiOraQd9kS1SRyZDq3Q0
ZGX8mVKTeGjRHnCHYFdy4Vy53y41GpKCabHEMgtuuoPNhUoSBqzvHUQx72nF4h46yR/DLy0z11VY
9OjGEiyPyFPFghffeiAe72IXfHC/KSTGeMLhUGNeSeWNoSI2ManAoS0yvoEehBMU3rbhrp36WnTj
7sKFQugv66uQelejKnhbp5CY1J4lk5dspGx77wK8TM4xe/BjYz6UFgf5BzMyyuY/w1IkAV50z+9W
gJc6JTbpOnWIRIfwyutHB1q6CNQexQoakAGzjT24Z2D8r4c1fn30/pE7wMXc8KyKn6t2Y+TBRwyy
nt6KLB3t3GQ222Nc726m5w55uz9PZtN5JvQIg6C/NjW5N0EiSWc7XyjNBEt+/K6aHB7qt3FaEnbE
gyafg2EDf34hNbdm9SChJ89l0l5RN8JdLYg9NyCAOPDNVUVay5dSI9xu088aafYfx19Sp14f/yC5
XHxllEB05IFaYgy0h7/t3Z3uopLFACCI+v0ZmkDgbIprBZq0Ca1aMWDyfc4MS8SvXQ128m5OEGb9
b4aMeojKoB49ykSGukv2DNylX32a4ej6ZYcbWrmPMKc84ZPXGf0xY4gJluLkXIqyZVCT6E+3opgT
w0Hh1VF72XM/1thdmZNQ/pl1AtRQyCSXC41hJZz3yKUOUFgArZqtay54xhvK3yCTsw4fq1kWN7qg
uOnBEuJmmwHiSI8VmiwJX6KJNC/8a6hHeCkrnxVhL0CONonkk6U2lFCFPi5HJosKaSNvZHcAIKEU
1DzwjvkUI2PaJB0pVmpiVIMTz9ho58pfj/Q/K2vmcUDA4uW5kOWDpMqhfhmJZfRcTMQ3qC1Ns8Re
Ilf496Te2ekya87NNKaWf1/PpVo7gcD236iQe8BMidYzIxofHhLTh3q+oTeoeAbTn27PMRCFpcvN
mqFaiY+M/l8Yy4M+xND4Tl7d+uUILagYKuxuWSwJA7bNjhKZVLyRQGnPuOY3nfsc7HrRQanPlWHC
Ykh2rR98RUNOamePhEvZiWdSw7g2YsRmG7m7W6sVskCZl3Mj2KN2JV38HgJuaMLsENQOcvrfaRvV
3+knWuemk/iYtUmL7i+XvXjtOjwZuRUZiArSZIBkiEm7dkgLWgYp4hsnpTpc0K9nbbAkCZUaltII
QA3sBv4oHgE9EXR2gTjtWd8xJ2coQ1BQa64sEJuesP6hq25075BjeRTdQrivgnZxlLj4RHm2EWgY
Gb4vLIVK/p1kSAp4nCXYn3KEV6wRis/4Hg9OdGGw9VP2V+rt7wml5p75Wd8Td/w43qeQrTm/H09T
ig6MN/leBg2Ij9X8XSTAIyxv4XvEEQG+QTzK8nUVK/a1Vp+ZBIAQF98rUvhSTfFfQvaiGjV9AZw8
dZpmx7WP7xTZFFtaxRyO1yuTWgI+JjYfA4V4II+/50FwGh5UBLwVn9qsE64bE1aIj5d0qIkwcLBC
tqS6JmTnR3WAryldiFsYGyIgfJFxzegP0obiW+Au5OJ9AOUa82oMzcYrPd/jfalYYJCItgxVPd1j
6BJRlZgauJYY+tHIsJk+r5y+Gjitx5B+iLdt8Fe2ruwh7LxOyB1dBlCOlvvvU/gB4T+hWeQb6790
EncGB79muQRZ7NkL4wDlpTl44IqTWvMpZJutVgfCbjFExGzHRgpjKEz7djvgwH9hmd+wpZMSRFan
VsWO48jqb/yTZVPWQH5qQXp6WWPl9/HAD/qCLV4oFbsoME0LVtIrhYG30kC16HpyoizAzEIZecyh
MzF5ebHs2E2+b3TzCxl9DZrJXxVjue7KPtYvE5gQY6cKheJCuIZMOpbkZrgL7WLUMvBt4hRtkiQP
/qIulp20ctQwFT7CP1wzSwaXN1aLmlohUDK3YVHpQvj51D5juOHK3XetSS4QaIyoPDuvT1P3Xw+9
4uxCzHtsFab8MG+sRIllgmCalPwPNJonERLABA2MGgU+NVeeJNXsQytngC/2n0+adPLsK3jsiuQI
1CP/qWh5LEf6VUDGi0AobIaCb6M5T9PD3i66AhYEJqrqRSuDpYYRuO/zu6j6tJmsqh91GwOWL89a
uR0pXCy6ey4jX3KXuLWjS4tb641MWcyLp+J06mnoUa8GEuSkwCW9dnjp999o5e/VMDYtVaE/VrQ2
XX63AvDTDzIC7gJ5I3/aOFu71hyGQSk6G/odMLYRVEUJ3vJGcqkD8j6U1SSr5g9gHaGLX3rub3vc
BwxesgDoyd/EEAaW8HQDjo1REZhoCcAjbV0L62RZLlL5f/FAxoA4jxQOoxmLUaQfjXGSFsIC41mP
59e4vRbTQLg5ttcsyM2BCEwCvtvSPOFZFgnLpRIm/SDJmnAJ/n0euiFaCBRQJbcAOkOlq6aOPODP
7SRF7PRBe4fvxOs4XG2GBr6Qyx8OYWb3DRU0NmkgcVGhc9kh50PBcqyHi2WeeftZfNKySUP13XHr
VgnTWREdZa5TT07REfrZ9doLTVmGPNsZ4w2FfBQWQ4UuRhQEcumVPs9WMw95BJh+Nc+V086zbwL1
YLw18x9tNoLSARzUIZ0jHTNDDavQ7Htyf6MECMd46m6QGChAarbfbnAdpl/3gEGu19iZjHodlSj9
n+c/VgR69V2Su/HpddtqXnc5kYM/jGafQu2W/VLSt8UHFxAYVu97LBFCvJQ1BEkVrnnbyd9Zi2Tg
ecmM3/+lZBi0cX0D5NLWnyhcWJdjDxLQ2pDDuEWbYpnv4QvDfZG1KLcYdjGk0sNM/lcvLW6grk79
bSzavTqvov+FA0FDF4VPawYrO889c40CRrGjDxZV/l1Bg3SxrXp8idVTUQcxP2114iO8Ao1YYjdV
O8H4onJtuwX1/rpkDZViBS/zrKSFm1Jl9INE+fuU3i/UN+1pzOKDKlTWqDHgdo3Bx/oyWHMJdd45
S9EnIxMVDgTIzyD7BEsDir2crMXTAozdpANAE6cGU1mmneE7qmNbDHl/yBdz+w9Znsk7PUldqLjo
br3ijx7nZBezflJHAhKUQCMAsIPga00RXf0aptnVrMShntilcmUn8tqEF0av4qQm/ZMPaiDEYBbc
H7ImO46T5ZPI8Hb2+ORatF85vNVeO832nBEa3gGPa+Cb6dW9mZnXObo/awyDGUxPm7JI1yq9YY5o
lUuq0/0FlyVh2aJ0ZFZJ58TT2RwM5bq+oh00WmNyLrGJLxBbMHF7yywzmIpOjiC+olXJz5M/itsc
FH/ZC8BlYzgcBT6IMyW4ZZOAY1WfZHA5tkECG2oANWUu43LqDmM0clhKr4VgEaeUB3YbWOGfE3Z4
PYfomkHwgz2EW6+TQcTgSOMOTG61mLNS2T+jA05A5LV7GoTxQwGwsvMn6BWbDAjqnNE8I+TcuGJt
WU5ovCH1to6+HQNB24sbdkovooy+EyroPHGPFpoqmyf1vVOWVqBcvQJLJtO+ydYLdLsQQ8jFtPgD
IDgdkN1tPMW62se7XovnG7UWlYxxfZECHkRmnBzqyXf4/Rdm5LQhA6iJEOAoWTIlO1gqOgK9Atkd
ISGP1MrX+KpM1h2Vi6gLvZUh/gvucz8ztm9069ufr9MMuX4rWhxtJdfvE8Ics1eRrXG95sYfG+6O
yPvznbHsZmcn0mg7GzlQIEmCwmLJGNJ4HN/yOZ7mNuSkkWpwHcaA6RWO5pbmYKg3dxNhECkGVljv
knARJtwWXnwFrLUMGugiil1n1A3XEk5HWXGvp3Fk/PL73oFsbbvOUU97+cQohpv6gVEtp5yMx17h
gI0x9elUoMZiXOlVU95MqaqnZRAz53dQ7q/6zfWj3L8ES4Xdep05NBnJYaZizB6hTzutwiViuxpj
V8SuKlczHNaC5EK0Kqb8kMAi8HM4EW4vFG/RKU5dELZqPu0HmwRx/+6N48WQyZJt0BTfN87WuVr0
9DNZp76MzQpT8y3z/vuN7doZPNDky9eHbaK3Xm2HIPcvKpJvzWQNIDh814i/Fm+W3KKcM5oVuQ6H
Ht6oyAEiwGHOi0jAI88UJZrOQ3EZU60rlIAAox6a43R/n0cNWjFgBZkxiNyYb5Yg2otNSA8g4MnK
08wWHJY1elfzmR0sEAmrLEJpP+UjnG5N9b9sMbnTp5b3q8Z3GKUUHcXW8gFz7tRFAwh6kzTP4++j
adzYgJWU7QaXktzO2OQJGXi3RAYZuJ6d3nYq50LugT4xXOCvyv9vxVAROqnKeTKheIkFRJhPmgSE
jSOEYxXEwVQC8s9gv4vNry59796Va/nRNZVMM2uSHwdBRsjk7jtAiNaR2ShfgvtJSc9Qrk4jv6EY
FgTh9R4llroTUsveauSQMihHAaYdcYvSlfUWx13a46m+ignBebjjYSor0tdWbtAXDlitkxitGtd5
lo4lfAjp7Fs6GIXEIPmTilhUaII+EjuHzy0cm1WyQ6JUf19xxdbsGL4mddJlYYSOspFJQSPGtReo
QlVPSD84ZYEwC9Vfagi/W7Y6BW5u942ude7nF6z5s2Kk4mffOvSfgsv1tnsmnz2qeTdfhQvF+a3X
xJYFFpBIO4Sn7GeOftHtoOfP1PJPTc40Y5q60oIoldFkFC7Twd0EmoroykhVsKmo6KgVm4+mUGEp
b4bwtO6bqR+Gtc4IIP9gPrthLIAZRu/wG0TIA2GjyBRUvukwJ3WHt+DrxB+VxbyWgT67en7OqUQt
juok7inXHOoyP9mESblB0JyUG0NPRpXWHvFf9H9+E4a3hvbmskuEDex/uyVCsI45TotvU8dD5LWe
GMB8qQSWDmEwC+6phP/NDuMBW3XvuVmG1hUNAW2kq5Wut6DWqvTLu/mc4ARgNAKpP/U5UBV+ewFH
s3iVjE2ku7MU4cRWubE3Pien+sOBMvQce0b30ZnwAJe+Q+Iawm0QrUp0zZMabaJVIMORvbcQDIuj
IVcFJabW9LPXAxGX8QIhFbDaeWyCzvYmDvnpA2pd4a7FpMaAQmkL7XUVp6FI7ftw2IQ0BrTz8TDc
y8wpqHG/T1DilxusRkEFm5h+nkeWeF2P/laKCEuLKDgavyeAUvEd7lBCEfYhs9sb007gtQGOisna
TwoZ7gFBT0NkCJe02jFMCYWD3UOxKRZ4516Pa9HExDmjsh9PL26fnbZ9QpnatB7axubcNtGFyBxR
UWSjopdG2bByLgTZrkl0I2nEcRYlcxxHjPJk9Iknb/KWRnPoefO4Vx9rUVmN6NFmjVVRgVgkbJyM
o/oKka8jtyW0sSaQNJ5Ap0IGZsovF64HD2bDMxoA2rKp1pwK08deGy26E88yD6dKGj4DvHeZci+p
i3Wf0cJB8rJKepruafSglqBGH6VT5+9HaWF85PmQQqvOGlrUBdjI3ZeuCcBFiCPCtlLujrNvboqZ
VIo3Eth1QShGesTHYZ5JXwOsVd2TTXnV5fjjhbkBUBDrGG9hxV1QQgdMiyUMsvp5cWDJZgZNwUvp
hWY54eYHJMAbqkVtR3RW1aZP7Vl6374s8tdFyuxH56C+pWti8ODQw8vWDtrl1b4LxoZUyJHl4xcG
YB2jevKrVm6+FOW1RKT33soBzy2csZ0O2bmXk/iAj79tpqPMAh2LZmCAVYVCCCJOA1cBSmdYaQ2f
DZyHpzz1KPjsokojXnFRGYBg31rTQMD3N0Cuzdu2ROl5yQMXJo5aS5837M8dU7bnvwJdxCl1KCET
/SZt+fe4k/rDUCUw8bWGGoUU01oKAe+iYTdET36spUmgTB4uzAPIsiKsPiIi3tGTUgiRzJmmeEMh
9Ep9GkUrKHesDQDoD9pRyj/kVaGcHj0O+fZ5Re/8CsMMsqFaR+iK6d3VXJcJVJVatii/2nYiRkLp
iZaktVgjwhbjIeDhT7BhkyK5RuA9At6P9QiRBBBoWo5FJ+jT64hfpYQBguxrGmbnDm1Vh6TLHzjB
0WxNSqxKbPWx46j2Nw0rZuwCquTNB2NulOj35eGl4Cyp1nPINv/4q/izpNhmuNAKCE72u9bf6vSo
BPUuWVlxmlPVXdXXnEPPtf86Luuvwp9FQRDfOv0t9jx5FTKSaqvMHylCrb3txDxsvxLe/4wp8w1v
XeLPa4lsKwZdzR/JOXehUoEKBFGeWxIWhx5nW5K5aYPT5mnJvbqP1wT9p3ZpFcnAZNxCiXOgSwb7
7jNXu31i/aGcfsm3eOad7Ps7xbiq8mfKzT/edVzjmlvMSvj7l/9kfbl3QnzhoPCIqJkmAYzL3pvv
QW0QgmzDBdW6oPdCfoiGi9Hu2xUc22Hmv0HDwXBi3p3eYmMKce8lve5xV9YVnAEls5LuKONb9aPj
HtNrK2C2hlkhozwgxjuJRKeJArYi7r011hW5tlsgqU2PDjMR/Ql7eFLqfNPp+H6UXFw7PNzAsyX5
awcA0NWC9MclcvvHPTDE5fBRF8mEAsAGKv54QviC7JD7ZhxRnYo+SyNmjg9lJ9r7dMwbzWisSnKF
PoZd/lQLe/LmvNi1WlnITqwh1XGKYTQzoAEawFZ0f7/cD6CAm7pP4bk3mfWDA1WjLWXZsw6EJjzv
0rwBhvLuXfWuzGMA+N01gxjy2lrDZ4uRilGrBicQpyfKEHTp4Rp5fg2GRGmWkOtVATY93KnFkZb9
Zr7oGcqN7CMvMxYi22QWSSAK5NssKZrzRQ/AM4JyuX4bLBUpiCcgBHzXpLqEmtXhORl/U/YLP7dC
Q/FwT7lQvZ8Bf+QI1StZSOV1/TaoOi877Qn8CXLd8kKlPf66Mm6q6ApjBHbfw8Uma/kUaqZZCDOb
vWK6HgdF6pziWPKpBqjet+qfgQT1HMXZTq/bmoRldqkDWXLwLcpYw1x6iQAma/AnP/InnnOLtC4/
+X5xc+59lDkcEETD3eOg4NsRGEjKXNMBvrlkyK/m8mmUKd2LA8bqPyrIXObnwb03SoY5ZlDN6XtO
NCmZA7EdOTnOECU6a5mla/ejo0jxItMzRaVpw6I/BUNhL7WDh5m/UseqTRmwMIXi7JotpMKOR1F2
fBCarFIVTyoDd40MfXnVqFxnPOafACQJR+rsG5+Ry1uy7VI/0hdW1XwrWieP7q1kU8a+Zsry+O/E
NWozeBjQfpefLNQ/k//ARNjWbik5KWZRhwbLRPjGoYhGweT7938OZHfj0Me5seoRVlwpT643Z8zK
sqvGXdBPD+iqi3H7PiSGTWTh3sEHlX5LanZTi799JbukQICyaXcwcwGfncbNmuA6/RHfHO4IJJGh
Zx6YDMJgJ6NNbnHxI4ZgzvGvqnxbEISsEGnIb/0V5apcE0JgLa9g08iBz6Q5cgYNIuHBOltZBoGC
Rsufx6mHLP3yCM5TynKG4JrEBDIlivKxTNbd1DAGCSCxSTpPAJdT/kEFJ5NfVSC/f7Il2UEWUZRC
E8rLqYJUWUq80Mhj41ST5T3ZyRmuXHj4A4VhQsA/bwFKdde235h19W90E853bCnpNyliFGr+uGsR
W27ylbnSF0RFelyXgp3uNN0LOYjNtK+OGJSRtzG6pM+EFfA6rFiRXQ/09C6I5juUQYeXxtKHbTgX
zs04Wp2SIHhwlU5oVsxvPzjxTpQJzB8h+ucnplvq/L8OiREtW2qCA0kRywJ1H0QEQzl7T7tgGPju
EF6gS/C2dCFqgHB3qkLRknxnc/dRoVvrJ6ghYOk90dTV4f/rO6GaIu2lmbgY/Pzhw6W5otBU8C3l
H8AkNMjTDCxKwKyi5mHaXTykmKB2iwmp7xoB+bfOhAt/KhVDfnvm83YLxSnGxdo10pcE3j2Uxr/Q
qmD1HKgsPsVOO0Df4+5zy9FfKCrrz/Gv0Nl7zHQSqraZ0MjxGVcFC4rr7VVVzA1uhVDVZWzgPtI3
hsIO29DCn35VYU2hhSdGgxncbsrp5Yj4AXkWYt7m3xLlorEsr0U0kNz5ZWsWNPVSNCZ8R2tcJ/mH
92LOpIHzbOT48QnLnfWuGRnLp8hVAQVHGfg76SZdx8zyrfLM9iyPav84KCcnj6LMaEWtprQi5MsU
Xqsbn/uSGEqNCVKBQV+IOmwHZ08OkY5WtbNznBmQY7GfUZeTQeSEGXzREFJMAE3LjEMErmDgcaXG
teBakGTJCoYj/q4wZeEfhj6JzhtSD1OGRDRjNsMEzZC+q1lhqQBO51V+5d9iOn1c2ddbMQEP2f5j
rOfk/qGrH4WK4WDT6pxj+45o+62kLM3gSIi0LjC3U6mmi7v8zemYZ7TpORf7thrKH9UPIQakbvvd
IGqFSOo5tGA9/SFjH2ZJ6S9YqsFEqdh4dvegGgtdbuSHjJlY1F7WNJlaoXN3sezlzL1AujS2GlGg
bbvsQum1Ld10fqJasYaaImDESJbAJv7W3thHG6fd4PXXTds7DqHjK2ODDJHNasS3puabCK7GZxsy
PJf+Xw8jdIW0XuaCcCOyzNwGg5z3EaYWdwr7NVVJe/dKnyvIe0bukUKV2C7kkoQ6lfpwRQDIRBV/
PF235Qr7vgpVjQMjAe8kQVjvvjpFoBJqjeyhEHbgGX2a4xdOfCG320DhfICrsyn5j8bxp2Cb8ufc
iRd1OD0Ntnmc81h/hhVwXfaiJw3H7KvtbM5oqY/ICQFSpCugg4AdR2J7imOYro3ZXT55gh3dtpXB
NRDwCktXfhdOnMLce4xgCS1EmW7CzSI9888/z4gaSQdyp92Ekulb6yaztzvqZeIcAmrZnMcMY4Lq
6zFbiXLr8PUGnGId3nO5CtGPoQzZen22a3/lW4gVn8bhO9TcXspry8Y2zU1TpgcSgF4x1Rv1iUk0
ylsk3UQNdknjd8OZtXLWw58+9mbIRFxOHMa+PJcCqYa8PT76o6SSXIlEjujb+/BJCm1kkg4gkcbH
rl3XJoUpuI5H6Sz30J6kyoOfKK7AHdVPScLCcRDp5wFuzZYVpOzVe4CcjHDR7t0yS20qP7Bcis1s
7C2ZNTuG2YaCWcqBUGmyVX7JagDREtGpxLKTbGXrXRA92dMeNlAdi4VtKAbwmX/pb52KweAd6qCr
xsbWkH0xlWC+WxYOAf91BtahHdzAjbz9WkIg9voDM8zEt1yangQFfndV+CObmzkuCz9ghLH0z81g
+FpsjHmI2Dk9c/HZ65WSOSXZuvo2o4ymo1A/tJjopux+4JsImK5hCDRYxMlUKQbKY+P0qDjgTqff
LND2Qa1k2RSi1F8OhyQfgTKQLa0lZcAEOsdHgybh2eUcoQk7xWKVmRiC5oau6Sg1FPOE4BYniPw3
6rTTlx3GWN6K6Dbc1QAr+lxlvP1UoVjOjBUKpI7BcZ0vGq+GtGrWOjgCN0IQPZsP6DeK+ZeXIOOZ
lWHnkWcuplIk8xu564YWIemxlCrlS5nTg6ewQgA8NnQ58sgR0BHSZqHYLXQVYdbX9+nKkwTiWsLG
x+DDERbdw8gmk4DtQCZWIpXTNsnvnwAEC0ryiPZPtmCTrpwTU6g/RUn4O5IY3Os2DrmZtJS/LrCq
ZTpw8mQvyO8+yduCIIWLLYKJOY6626fFWDGnbTjgdbNVpzjF2CAiXp/WsFnio3SNr8p3v1+aHVQr
5CiqFdIEMbRhd5jk0SSMsl5Ot2sJuBVDk8CAnXUU7E1zyil//s7VJ9T5WJzRaDh1xD0EUBJPjbsK
KuAFoRR7iirSqrBXd88Y6NOUnaihQcG0GIYfGzvZxV4FgtkqEg/mfIneZ2h4i66rWvtUfvJQinnV
R/NCUyaTRypVT2LQ8n73pF9GhFwmATd2ww2oSXsc21VRE93dEdpsNO8lAhD9PIMTz1T0sOXw9hM9
I8FurK+2rUN8w0OU6HKHQLoLYRTRSfyGe/m/9si2e2X5mvmKoONgg+WRIqWklyUKu1eV6XDMGjF5
/t36Iy8GT2iHPwz+8hpmwNGZC4wfy8rDS/1TppYZlUTX1jFewWvfRtp12wnpQ3zIN6LZgQDAxSGb
r6LEVndBctvkF1/im2Uh31nmCetAhXT+ZtwN8PLlgVp3ShPp0L8qhfR5vj/OKjxaswhQRa2zm1Up
KVHygQPsn0ClIsl4WnctdHZwxvaOLt19gYoaSytD/xjZTPV4PhWqI1uIik4M/yjUCvYWO+gUI0yu
4Js0s3qW1DdV8OR3Idr9hpn2iXeb946m6vgC4KLpOb8RHoB/yjsPRhLCOm+brKHSunYfK3QzYUAe
VzKe5Fi/nsbn82OtqtXHsOft0zlTKVLcEAo2Syw0soqMYswk3YT55PXRfyPeScXFJOqJAeFREIno
l/QmlbNs99WHKtKeaW3vtxMvSbch7miOLYVETxmjLrOuouL5kD2zihDyedEzp80L8biSXEAzGVaU
rsO0g07SAb+jXz6XyFnDnZKn3kggGQWyewuTiQXJaub09Jq3XXOHSmldKqQLGq0UZpJlX1Q0PI+x
6Sv3Cv7kRhEXccBZUmJWewQwBN4uDGpiYfmtPXI0kHkQLOc2TJbrLrgNPD3J7yETzGeIQPv+Vv1/
EBU8/2usbnHaG20EKCnDkE1gqQ/kId1BbW6lCtuGkqK/HHnSJZpCpmlq9XyV7w8Q5raiqRmxUL2Y
eMAjGPDtGpjexXc13j2lNCOUNDGc5/xB3HocA8ILlFskYXthzyUQgSe1nILam/8JXAYeRWO+STNo
48Wdlum3YyL4bZ+4i94qrWUA1nx3HmCyfG7s3AQKAExf0UItTGD5SUGgJ73cV260oq48B1NN9iwi
ktC3I3bBb+AwpC/p6A3pgoW0KPKd8mNbmE8I/AmDHALrLKQZgO0NeL76wBpaxutOtT/bjtRx37l3
M82Hqt6hVEdLYTM92+zZ+kh4sg5DPxAbGEz04hpJ5UVfw9CxjQLtqo3REnu5EoLmWayO7mVXVhGj
zdeqcRSs2/6wXX40Ro2l6gnBR9WV+XxKu+gpCPcyo7u7gSq0SoBdgDnbIh+Uhocf06KxQ7nXqdpQ
zOasgBxbY5U4PIYZ7BdsyWPCtHn9MISXaD+xhYXpNJxfiUyO600bLaVk+kAaLO7JCaPblV36wvot
CItZX6/FBfWOQUf6kF3KFbq0i1VrR0rLOh4PmFDhAk6W+mp8vveCHyxoZb5Hs8Yr1G7PU73jZJtq
zGWl5g/C3kkGqFKe4BCZNXVihqret3SgXxVwWzeC3eRzPSXwXEdqPIMq41m5+qwMjJoeTPeFGMTU
rjy28TkFRudhPjIJUlm3GCD7gV2JnZrHe6cQXiUdUdwq/NXVlcw0NuumxT3IYEq9xhURJBfjRP6n
CZJ7xPGTJsma6q85of1COhMU1dK6/tNAg6ApIjr/ou1GVXdfeQEHMHVRzjZEouVvOD5NI8WutDrs
WNqfpy77sU1qyDevjA1523gqgkTIGQLjJ7BbHPOLOkmcNqQxpI5fU2sI1/2FNRTwRcGqGCjykhdB
gw48h2pJWqahPl8vnmpi2YUvjByWDW4jsSVBV5qYJVfYcQc8F02Ax0YmonXsJJiHFQULZTW/asSJ
1bu9QyzXjGsXV5HETdGOJ8vYmQM4gYFT+ADoWivJpmS3BDfN/ihqz9xtwL2WdIumNFu21Gw1EENf
dxvz0cLGQyFp2w4AMEKfnLsSOQjGGk965dnakdwr780OcEcM85T3L0+8fgo2kjWRc3VA8KdyaYCJ
o1gXbypczgGglkBkSaavxS1YEBT+ohecBFcB9aVLFzgBjExMnhpm5c7pKYZwgny+oVyCVLiRFeNw
m18geupGFMH/OUDLkTXrkZjqHkvv0JHL1NwEUbHyw3Tel/4YM1Buslr5delBe+1fN9zzPNtm6btX
57GGJjg3wpnlklxMcLSFFobq3EMDSM0i/om/Vjv0mw/ME5JRCSkhuQLvUSEYMtkF9HDvmgtOKOql
cMHvrF3NlgrkIje0aMJjfzHBZfFuWmFWhmrGhVJtRrcPp3eeH0PUZ/9tAFduVT7+uY/MXoSamFeL
O6jo14hLeDtjz7sdFtr1cBZtjtYLeulMfNgRD1AmUaDEIyVq1rr04NuV826EU1l68YF2BJ6p+edl
YcSE7fE8NyzCPZ5bnG2AvK4IG0b303PLaLUtvsDT7Fu/jS8qdZScZ1VYvTZ87q8bTNduLrQI5mte
AgRwFskGfS5jiSvTEqNtGKHqZ6b4tmhdXRjGwxz3eYEEDfLTO2NluOLDGPpTktYDx+A9dokqIlxt
uEPK2ESf4pAbMI6B3X7WAs+szt67S1UZ4h9Y4W5aRGxFOZGhfEQxMpCWO+bh1rNn4OqQPjXeqI7F
jWN7IfFbgtJh1LqlJZRbsRyFWrNkPEzdjI9BXiB+oKPpi0AzvneNdoemcZmqzzRWLPTkHf30S4J6
eS5x723VIROjcBI8goYPvPKqtJcOxd1Qgq723kHiGULhPJos+HsMrs5Mm5C71i1tCy90H1yHccIJ
wIokPBzgS3pBKIzwg/tExu8jatLUOJv7ZL42KVdQfowSkpxWIBD6FpXqXOSFBOfluKgern0mpEml
nkBo0JuiGqo0k4tvRiZV7fwu2chEUyVWtcxN4Lu2JhRmDuACHpy260jTBOhNsMNZXroitCeiBLbU
bT27KowkDUHSBgsBIMOt5J3Z/VLZwL21Vj1Wfzi5hWSQtjB4lAI83FT/sQKMm/mDMC7aQkdbaqnL
3Ps1F+BfYbi1vQizpHg02DAhWjmlFILyhnwQuPmaCWSwRJbFBuViB3V6UEmQEg0KIyA4Y6uyC4pS
N5KHe9wLW5FYCamhDWHhSnoJCfgLUo7mRWAdUi0HbQl/Gb5TnlDtJGTBvhx7E2PQcWXWLvxsZaeH
axuyIWRvx8e51Adl5VWw8+M6hIDD7bLys9gEq1hnvs5wLhhSQVmrTQdDTaINXGZs59H6gQHkfpP8
mka7Qmb8HCURXpYHfwN/2Y1NPyOE7Gb2RPHpHd/RblG5HoZ/NUwop1JRbxe+e/Rvv1kwFM6ps1sO
8TIuEGVtK8U7N8XsSLL7627UuHnHSj3aNA5PXy9xDQvTje4i9WuWqoH4SvWpCW0/AHbuuKYDkoPV
70m9m876SNotYt0SyHeVxevFAoD7ocJnyRW20zLvQF7/x7BiRehUOiPRJCCRzhJZzIwlaW1CPirg
1zK8H7uJ3e9e0oBKUIuAhwZvSFOwBozcA/LnFY14XPGV0Vaq/wrhofA5TClnEL9gyNeQKMHp9zHS
4Yi0/UWrO/fIVx1qUt2N2faIbiR7GnJgCMCCiCHmMAgL97iu01xqg90Uu5m7aaePJx4rg7dZBs5n
piW5ADYGVLXXGSrq8SSsObWjSBPe41Tinj9rC5iB8kAlM6E5ySkeytCj3dUc3tSIR+9QKAnS2iyi
mlDwnatuDwrVIi7TjSwx7FXMqLAdPRYV1v25qlDRhEcajvAXcLrIbkmxn6My2npBqGAjYrZJHCWA
BCYVV2CXplF01EC8R89VYQphIXVsH1Sq5hLu0oRZtvqJ9GgeY/GCRbXFaW2wPg0LjzZId5k8gCBD
J2usZC6RSTJauKh/Xonm8JhBdiRy5qZoZNLNwMyOMN1uj4hP44ACsKI0y7+tr+pJCiyA3XV/mesP
qny0+ZUufADBQOCCoFn0gxWq2dhCYisXIwFd9/i9TH+b5gdi9TjLOyuXJwRSPQo1HriKzvLmzU/8
gf+NAbUzfVhmPutUho6qEqUVrj/elf6uESP/giWe4HAHtEGuqlQUkMM1Zf88sRhIk+T83+0RmWTw
5szJElE9XsGmIVg5sT4S0YWUE3TDqpSwtuzr2wyNVsoMk10JPa0E7sXpwkIMchyRm08mt8FPcbXq
9T5rhTCd2v2YC46VGCWwY1pcVFRQBGiQAYUwMxHxsXYc15xFzEz1PmnXKUMcVf5GNwg19fHYjkbZ
JafOhKUMFjXZI3qqvpSLTOdwoWKSyOyZ17ro6B/5GeVhRosZLF65q15Dvoz20c0xunIcbPO9RpVg
EGS1I+XaTWWaqPcPkT+vil7YS7sy4Q5JqQ5CGD28baYZQKFPkkE1O3zu/+/yg2eiKe4wtE8nz2WV
QuA8AeyMHJ7bPow5yedUdmcY+5ycOztgmrwNYWNCVzl5mBejl9IXzN+0fJPz1TJvaUL13ndlEwzS
sMBkpp1RoKAR4rMJcs5SPF2S45f7mSWYnFlV5IySAoNHm3k5ARIjPwk4Al1XW0oSYn8PusjFCXgC
I0Il2xxcjfEOfumQs2Nmoj3nFGEYi1etXs/tk497SrUo0fjoZ4ewKOF2vyWrerTZEUfDcAur9G4m
ugsjvq3PAPER2H/IS30bUZ8f8u/uho/mndtIvTYvRfEimKAyNO5+bqk9AFu/wZzkz/LUDydYcjOW
29iwMvHCRaUVp7xyqjPWlx1wc3DTFTDS3+1NzckRGDk7RZAuvPabAPRCYDfauW5qoZJ/9JDFJSVS
Wb1ZhjAdFQ9GULNpCkw1GldMVh99YrypK7pwCKfp7P5Kfq5gtpdLdcbfbbE26iyuQ/TiuZS58hAb
8oO3z8Sd153N98zC2vy471DGhtTuwkqsq+hwgXOHeIRPgceJnwM3/Dvgr542ZqzAm8RbTjT8kMaD
uhRuUKUWOkF2twoIgjnTWbX3SrKKMJMuA5nEpfADQj30uYQN3YoAijdnegPabNz5xplWrTYmvLcA
cDLNwqSW37QXfxcTNTo0erwA8gsCHz3WBmwRjprtt4rqr/C+n7RteMtRhqSqIoD5fj6uVqskgP+u
0b7gr66hhRu2UUgZnQ1UgEpXnDUPBnI7vz99luii41PKGGHfviY8FdA56qGI6I1OGARvgO/FFkw1
wleKeuBHmkGRQ52EA3JFKUiBgbSZGwBhnESNpEJPkokJXZT7WduvVnWTgdOh7hd6kO3k62CKVaYF
xVp4/gGzwVkqtw8LW9k+sR1X9heD9/ZSPS+82bQQOhnpf7HXkrfXXPyzMYwku9zAlT1EIHsagNZe
G4t//a/mLshUVIo9ad0GAMNuUgzxEFamxhNI5SUNw7zN9Jw6cApyFspc5o8CE5Fytt5lCJHCfcDv
nJ6hj0yeiv2S3p6lrPm2YpwBcZXm4Po/AxgXLzkvIHSmNV+xTXQZPfr1sjL1g0gwohFpcnBzYkFW
sDrt95ffDq7RpoDsf4FjM29YbK84d/8LuYpyQjRQaSnyn0xMP4qw7n9Ky4zBlVnLWNnrmUdB59TX
cUaNdPOBHJkv6H9DCzo5vB8NluyunRZOx1l8HjT+nZ4YMP34U3XaFja7ErO83/bG+Lr9jKSpFP2E
62irwD1iG9D6GsoLcIsbnEUiudJ7c4gPVQV7yWtCp330Bb5dLUy2ak3k1ZgriRkvjNcXa7WyAO/P
DjUW9LKhf4o5gd+hjWemgUZLcwPUrBuDn9F8nh6/0C3vZ+eP3yMedpbEhNvYPmcCdkWDxF/EJx/8
9Bl2yRUC9MnmvFqwbCB97MmzL4pt0vFwwsab17qezmWUUlBrmNLzzctMm3Zmt4/T64toSKfRkNyx
9kq66o5XXotJ4nzvisiy9ANLrtBwAdiMdeZ67DMAMhuxM7EHdZoLbZBGM1uzCyqpB8MpLPen3R2/
zhHzw2ProhUWqiP09qt3BgRj22HszklY7QVzioxNVtI9amQzFY2L9IpzzNbQWty0IWezRf+H33wW
uZg6Jc6/WjEK/URNlCew1pLjNNRjMLS5l4ExSKmbel9dIdmWU0wNm9V4USGyASw/G8jj/z5ys9yQ
yCIoENRuiIXZ5bFygcrLFJF21rUXT9inZ0gIArjzPXuCk1mnEWgYOeSNYGaxq0iaueGP7HT4ipns
vPJNW60GH47ai0PG4ceUdjFAkmFBLXK2L5QzoFxgTXM0Dxh3YlxG06nHmcqMpYtpgCoFwoWAH3rf
6bIBCbs0CsMeJTnZbIVWO4HltcAxtINs4NkUIjRIynIHNWfYoTrxPoT3yNHb5rYWCmfB8u4KynZ/
S2syiS8NrM3t5FcsuRgSd0yAexRMV4NazLspc9/R7gNQdsUTkjWcxX+gtZYWilGwI1VWmm4Cg+0l
jfI3KrK9QXHMjIb8EY2xJktsv1oazxrIpnE1fphRO57eNWVX22cGYrS6BWqgO5cKdgt4GvKLPiPn
2VXH88dt5bsCDEFC2t+KXmnMgnUAGk+FeP+qorP4nYhnxuqMeLsjPJNpNuFqTb2TlT5tM+OBnKWV
V7QExaMA027/tDda4ihH5n8X/ONa0SmFl//0yPfFyk6gQyHbERt40qZTARYUCgn6KDiKcVf6mE4c
VZLZ3V+FZtvhbsxydd7h+UY0TRVCyXgD3MDQVJyApRRQIPuW/sl4McSzd1jWHe0p4t5qIZbU+IEn
EKhrMMMbEbzfWYyuhPuVUeCeX91N24IuUGef/VsbcJX9B61JSCIhPy0sw3EEW8quxmEqU4As42Ly
LU7kneJUvbP+CCgq5tdMyrhuNrJj24TFcyN/pRhYTQDO4zUM2C6Kn4mL8KF9BiGJvPyH+suxflTN
8BpKjkcR8evzWXHQ0QC1e/BKpqhNUtGf07IWPq1NeSxrRIoISY7EMKZLTX1bPJUVMzZPFjEJcsHR
J01984ME0iAzH2awbccH7Yc9qBBA663vgrueG5HuzM1NhJQqrEVmxZ+fLU2OzpUX5k/TDBwD+ZfQ
ibhOS+kpJy68P3Kd9kQgm4FcvazKbD4L9I98GNuXW87BQQ+kbUQpOxczGDh0UZuJKJRVtxrGEsDO
KTLZPtBnsVAttPIbOiRPyl74NHKIXz+DTGsCEitB7yvNBGw7CPsLAIAGMx54tbZVFl6pkgdMZzEI
zesa8eGHc80Z1/KPAYzQHlCqVwVnGfvneRcBdmvmDXM7E7UNqDvP6YG2xot3S8kQxmOWe8vU2xRi
kjjbqvNkXeSOF0G1lI/pOkOpysEfdy4I1iEmm1hiVH6SthfcYcQXL56gaIjubetRMx2sTVOiH1uN
t3iQv0WglRQAdgial2zPQpBQtQz7YTiRu+WMBwEZAPe2rL4Aitt5cO8r4uRnZVDIHq6Haf6UzTn0
I7TOQKaEviU1SKnM2xg3/WnzJ0kAe/+CeoSKhYxQlFXlHOAI2NB2w3hl3742sJq1XCQ1+dC23KpL
LxXOuWtPMI8GJ6iXiJ+e95AjUXSxSMGTj58R8tea7PAl5uBYrW/xHDnJOhwLy4C78HyDCKKR0sMe
zJ4bGTiiKYh1kxRm6PRxNqx+LukGuAnvwb+fMcMnsivppkszgjMelF7QA9/JxrmfmlySt7AMIcQi
oPR+yvk91ZqKJaph/fn/Ju6NZ3VwQJ4RQG8SnaSIYFtEmMttkOH5a4Rad1gFL5hoLz0RJQNv4kRU
cgXaipzVra8Tp4eENnjAw+z8gEfj0oHtbHIg5NrptkZEiNClqYG6dwxILX6U9wefMl0sr9CYEG+y
X4MeFUUW3wl+QarAEkUc1EnklEut67pvT0gZH0rqJoZ/ktZIm9NnssRihD/joWH8GyDNkSsU2zDq
I+1b77NtEhzYR/Mu9K22zSp1Es/Ft41uuD1yyjyo2WPSaewkJmv6qWedZgatDe9s5cEjoKdUXNSP
SrY7Ted8tYLdEarTMZs4NOv3T/dMbqkrBN3kIFGTtKC4odZwuP7l6tO+tnMttQ6A5++kQBBh3bb2
9LhGPGgGLcfEQazYeSeMlpOBVhvyFvJM2Ja2cIc6v9B49dZL5G63BtrPrIvk8xoVhTQuPkBxyJtA
Rc6T1wMMVxqPww93DWdzKIgDvzgAVoxj2Hz1n6OidF4bh94v+GTALBt8SBfhm7HErGpXlAOfqP5s
uZIXEvCL5Cp7x+vrSevbt1BK/SMFdkn5Bv3RCHtyNHrPJR+rQeS3FHcy6xoMnYG+MjrL8D6Qph2V
iZp109lXrDVSjMNo7FBeD3+lw5wqgVLow0LFFKGY0zCN2X1ljlPlMwfz1n2hNkS6NYXmP5PhW4nN
jSTodDJmTxsiFhAuzTgWuVtq83OHdlVhNoCOUUNo8vTbYqIQvlLES1ZLjzoncDNS6n7HpzApd6IY
3dTOzAr1ryuEKxWzZgAWU3haRdq+HAM5nqUKFr17X6ESybP+oJJ4UDSkUg272MH9/GpfBfPRQBfl
kbUI8oq47+o0jnSwbyjjCrO7OsUsU+7+RxIwQhMIvnibRYqXkLKNC8n4G+FZZbdg86vbeyCTHM4G
cCkGft0m6qVJ7i69KldpaYPRf9i96C1BOa0GcEV1tjokDclu8/E2MJO8ingmjra37FKgAeibVklZ
4zZbDo1t1wfQA3H4jSq4B91YAFG7UC88WlMnaG9naMy/AUTu5Y49qtjWNk6htd3sLpMIV9DJr/Gj
V6acN2Ho8ZEnzszeCxzvV9QpNDk4XKtUv4zQRJZ+p/is9j7/ayQ9PnQHufKFFUsyRmzDw7f40f68
yXGIPM2tL3s/GA7NWpNwWhLwlhp/qCpYMwMpSntsBrH6lk3xWC9M/kCxhxWRFJ5nVheJDNORaC7N
rYmPPDf4L3kgWL90zJv7SN3i6AE3aVpo+K3NvMdB/M4KZ2KHI6o/I9IPhCACuI5fxauh/o8C3e9i
ggTczckKmFOCVYJ/ZJQU36Y/sEF7OQ1PaktdZHCJViM3mpnnNXld/Pxf4YOIHuyvD+uiLTJb63fA
RGokzbPQHffxgeTObU4pHmM5jy4WyV+QCnJrfb8L0piKwS6SNyQfEnFIhkTzAeZhbbJWeHaoi8CL
e5TYnnhC4BnA/bLTg8N+Hzz/5GrZ4DZVRD8EvIyVUWOXuGFZXiHV2PR2Iy7SS1xWfg08jFTw4gfN
jt9p7E4GKa3JvFD8bdWgoLDuaUYegYC3oeV957t8jbmRlFbBz6fa17qNg3E0pdid3mcD3nmP5Al7
8LVIYARXzo5/ff47p6BvMmWctq94O/rMGISRUlybxx59dgyHv/6a2tlnkmf5QFXJGIHr1yMz541y
o5a4KgEYU+htdk5Qnp992Re6TbccgVeFmVmMyP7J4M3XSlsYwLEKCcoEY9vkqMEUgMXgx210raeT
6r50mp6HFJ2YBX7/W9x6pwLTVlwroIg+vuVZ9IH8ETMZ/evmqAAYJFRjlXi3SFopxCNVnIU/6Q+L
6iTNkPleEyldxwv8VuDFwASXlIoQyTtJS7gH7AlzLQYj21KTaGyV+6J8qjbXrXIeHIuuTnJb+p2M
zwv5FrG2mXc8lQdseGd57wLGTp6liyQfETgZaFVb7bm50pJ19/Qm+UeVqzeLoTnXbLbArP7kxsT8
dtOV6nKYVma8YSheB1n2b5LTHuLSz4HDJlsjbsvJlcGnR3609D6qOV6zg4tyEsOLWifIrlzptOvA
D6nSaRsN9oCF8WvpiENF4uDHXq+Ixcp5FlSr3BilVU6B48DcucOzJUQ8lva6OE/1h2iiFsIEzgNG
Or4SS3yYMm0+K0TkZnMSTxEetc/XANZcBQnJ7qH43b3MYs3lFXb3CLGW7hOXMqwtwCe3yZl38+PZ
giyUTXeHpR3Ksxp5y9tpitH70akWRl7Vr7ZyCisOZjEzBIjx77L75QV/sF3wCjGfbbdODPhFvDA4
FeMPbUU9qwlyTfK23wntaaQnr4nTXv0RzJuZdSHMpTT5TFeup97QfBneK3KRbIi4SPhbTp153gGs
L2+qN0AWjdY46lwOMIlIgi9hPT8bajcm7r1Vix06HLf7R7x2jFvTgj+VIQURZnEGkRqVyX2SNl+Q
0VWJ25N7vYBkT39ZdzCsuAQOi92mdbwzddpt+PAyD274hCt2/C3E7HFdpZ6aBaTn2KCrwR6d51tT
ZQGSEGCpZNX+w3Nc5cagl1ObyLJjSZAqmGg7bMKVIlVgD7Kc+hMUdBVhxHEfpXapEMLXZjBRKFwt
Mx9FZ7x0d9d9EcUra67HI9LIhX34+mtprMgLUTtd02YsfNGBI3mb1auS8wo7R3GaDNR/yiNFl/+c
8XHu/LELT4y3bCp4GyWJ3vHqbbCtHnK2IL00763F23AWwp4uxUnbkTBgUGr+H46kE7Le8qP/yVee
HQhB0/+behh64UKsmmmIg4Z9E3qlW6Ah/aI3aVmfPMu/nkfvHC0rjcXvgoKxuG6b5n+41hQU6Uaq
YvLSR4qiSiWjy2lgz0F1NjTbVbALp0AtZSopfd0N0yGPWjMmhUALXRqKOKlTcGS9RclY+5D02LDs
AYOjLmL0FD37hccZn6v+0DWrrzHv1sW/UY14jno0xeHIThRo9SM9TaWTj+ZwdkV3iHjXfDGuz7B6
NNMEYVUdalN13ZcIZ7vpqGxddC4SVQVBNVCovQsc5QB3dIvfOBHf7HCuCxgrVn0AXa+xP6gl9E5I
Jrf4m1mMkpMLTTGV4aXPpX/JyHjHZW5LTuzhCH1bAT6dtPYlQQQjWZmYMkEiLWFh8LDj7MS8ZmkG
hfr37sMi0osOOO/b1oG2o7oslNHunKINkc+AnhTP2Afth2bcn7qDA6k5n8nsTsNGMzxEYd7eY0r4
NDKdAs+87omjlE/HOgOMjftIUbohIR0XNSBW/8IkNK1ZZl4+E8PLPdqPzj3IuNzRx+D1mojeuoKH
0pScin6WivAnJUwgc/67gc0AhTqr6aX4TQpSmrCrE0vOO/OF/nfAk+rwYFJ+8Z1HL+un1FU9sjfY
uU1gG5TdrC35AENq6WISWbVrzx9HHEoD1Ht4iIufj9PeVZDTqPny6G7a23aeQHGTU7ZRZzDxKVMM
c6rLDUi/7t1LSumC2DPBWvfOG8f3lj5kvXIcOIAP0N2kBZ69561JVSgrUfyiR6nt9PKSE4atVA3b
BQmyIstnNs5xQlNjB1kZwUhD0wStB0aj6h090qHcgXcboObgC3OLI+eRC9YpHA7Y4MmpTi5W+qnq
0sUhLJ5wHoS/mhTXmT9xSn9arGO/k1AWD5Kp/SCQjQr6W+qPpoj889gFDAe2aXC6Pp/EKiWysk2v
16QKqnKIMTif+dw/o52gHx9Ch/f9FVroBot+9RGObQkeXic1loxPO6TRSSB5W3EAa2sk0qZYFgIt
MzZTViC/n5RLKh4JpJ4MfzBTyFGY1Vgn5FxssReSAxpjSsAm0KluLemGxEOMU0yilzSHKuoPNiLz
2q7k+ry4jK1WJvufzizWK58vrcpetewPYDYL0f6dV6OaX+vdVK7GnyIbZWzpNjugQgUaUSdFphF1
ETgMqzssGEfPu89+50A08O/CRfPuFheaGlfmFFc/H6fkviqxUDr03IqAYP/W/Gk0qTk8lE9X4K+r
REq5Y4SYwWJsrVQEwWe6mW8HkNC+ZicgeW4kedt2Gj04ZQJ501UjRj7NBmta7Pnb41O17Os8500F
E/geHdbleEY89i4bNQMpfa53Iespd8DpL5IPfleSyTE6zAd20ds5khxJlVqkgQvaWG0HioLL4Mmu
cTvZjkvPTqptDCw2y1DZAqL+snRgTu3ICkc17gxX3VC/GN1N0q9FgwvJRgFj1HA9KyTprLj6YLLv
EeBb8H1yZJhHw3Tf9JxZ8o2Cn63QxdIs+egNAqAU8VHdk/asjY0yLJxKFjV9R0+ET+Y3UZOSunKF
o1jS5kyhl2ngE5RQ3m3YZDUTA5LKbHkbDX2C0oPdc7fWwxd3o/R2qFN2WR3/ilVTAEXAPtfwdfqd
vOZIlM4SSX4HhEjuGGC203MuState6ukajKGGvhgalCJxFt8fGNQRlccXi0ubnNsM0yDFPkEGVjA
WFp0ZPFHve1Ag0ExdwLuSAYyMJzpgNdUTuymMbAVHTWgSHqN7Z4GdRLitKsedbnxzQGb0SErQWj9
UhpybGeCQRO9Mnueu7wIbZmX5xg1IMJ17yNb7m2HP/re2Q5QUG8ygw8OSOOSnVgG5+nSRCR2U/eX
79OVYCAliaHTZtDM/7Yf7h5thryi6r56A1inIYDzWE8ubpDI8YmHcxFgsxBPdnoM7AfmvGWQM4tg
tAz/y8S+d4YINqpjSf55XHUBFwgTOVgeBd7Mvj7FfMbIBIQ8CUlQD6QtKs1Xft00d9R51YTbQumb
iN3fytyn0UOA4CSYRogKZ2FC+PjO68vW8++OZ28SZTU59s70G5QPxCRmR+I2lG9suh/8lL2LIM5K
hlR+bwvxnnS4GvFeAyu2E0RrZtvmzFHNfLHErZ73YxYHCTUQdfEZ3m0GMzgNNrP7HF2B+CnE1Rix
2ZCabqatjLT+IwUO933oPQoX/mXG6PcELPDFksO+fNZmwHLlY/G1rOgM9SqKvloeedFBJEpPW2T0
yqXXCfa5IeZBvtaiY/4cRn1GGeQC+ezKdNdnDWCAZt5rtLX8rsfXKsdCquylgWfT7aA0LRiT4jvi
O/9m4CpPvMfg2DH41Mq6HGYomXGlywzveuVdPQyJ6pDHtnZBKg5Cwbk01eoA5ZwAv7JxAaSlS1aL
tT3UOFDZ0OuzgYqzeUhV92w2ArRGP5PvRRB4jGd61dV5l0u94YIlyNOt6ConOJaB08Dv/QVqBQVk
Otw+4N7zUel+C1ZPHXgBohx91GSaSZw19CTXsu8qZFBnAR1IvXc2mXRdkq28zuUxbdqn8c5EnVcv
JoEQKrUwSr0y2Cloil9EYO/6oY13URbXyFbKlH2dzerC7mmYHkloWlTOUAKLBoQwOWUb0I/cAbfO
4YUoOlESC3i7HVF+oF89VVwBQhHBWqnQ1IIfr67I3IJApvnn00ZX1n4nayY5P9+NpWte8JAEsH7O
F3rkun879YqsmQt44bbvqnYMH2+f5CuycdN+GEWi6lJusLTky2ls37iyWIMhSb7iO5/IjBZ2THWl
eQve11IN+d4fmskFK3Ts4j8g/eTF6ZJXpOOPWfGX+5Bv2+NvNr8NEsWaHU7CO4E12sqyH3FwZgZe
XEyG7slCnTbNR1qyMr2Xb2Gtsu3JSZ3GO2+Xw99j9qpPCWjdstpRb6pWKQRIhfNy5kuBqo5IH24u
iMZfhAwssnFlSmk9d+QYqPnu1VNQhR46BPxMt9Gx27mobOMNqE2f/tEVNwB2MlmvXBnUsio2Eb0L
Q52llCumP5nsF7q1cWl/l+pLetcS8S/QAU+j04O1U4H2IvE1PS5CMTl/zo2KS9/jxIuw8yD5jLQ3
vnC3SkHGPm/wOlsqjBb9usVZ5fyYr7SPoBII8O+9OwHwHBQnHoWzaOvcosdmvlWJxHtUuWeotXY8
9ZAZTNBqlviwL//8xnCkY1MbLKJWU6N+lfipCJuB2Sg+6FOMsprDFdL5IbXqlzqF8EpWtewOsM8h
TGke5epjGRzE3p9ZDZDFM/0XRUjo5KM+/AM4f4wHJeXHslOJxoR3X5fr+gLt5P1ZJj6bQZ7A4FJu
+Kt98dqXHibC2kKiy8f79KMzlvJIOJr8YrIthvL+Jr/9m/cmofDbaC9+9w1gJ5AAMkE0hqHwdFfG
4dsDJXM09xeBp3jjNrNqkjQ5zh9s0NEPi90YNlK4GaqOT7404fFxYhtxkV7ApJxg8KZhiSfaBz5u
2DY5A5wfexQmozrJKhYBZB6PkNvbMYiKALYa6te0lzXOsJeH9OtPlTT4RRRn2g5WPRByl1pSHlI5
N/X+flUiKbvsm5kYCJuiymNFmRAiTLhznkV2/0UyipCswctS/EtmkKKUrshYhEWTL/MIExVXXIwA
3zHOmC6wFnXUEsnpOqWRpFQRm1Si+C7yPKa0H/FJkpS2WgFBdvx8jNebqx9L+KGk7dPJXKTol/zl
qGum2nlKa28UOY4I5kMUOnMnP/Y3FxS3N2PMA4Ot5/Gm9FIoW7eLt2AKIbdo0qLsKyAEnIXp/RC4
3QJ69GC0XsGrdOTYqdhqfhUcnWHOycXeETCreJ4PTncLPiDg1Ey70d65CjXYX32HMoUSySzvXbas
2DBFxj0bru8fhrei4FDPcwJmzHH8GQD5fd2UPvwjQt2ybhgO2SdQMlvbnlz5CGpy7k9lJmFgtZKH
VG9rZ9beAnWv+ELbG5o4t5+usoJ11NMtIxcRoLHWjS0zHSdvd0fSl24heq2VCaflb7f/UxM4HH3O
2H1R1iGq/53jR/4/QAAjoNVspG+p9xXCJ1kpAFWdTpjlWqR34wxT6hKaqwMunC1Qjvft57g3IWuu
/lKxEqJbBewt5n79k/fLrqJipBRFnXGYT5GkvPPzhPHOFR+Kmj6RnDutQjmUHJ6E0jeT2f8Z0H1f
l2N+4469x2JOsw/7u1ZWYU3Luwv4T0N81it19zN5joWseEmiylrCN4oyvT6qk6q3oU6CqE7f1e5c
/FSdSJj3bxq32sKePVcZwVwmj/VDwkMk7GmpAeHCZqF0eblF/1qziiuXvX4cGMfCOwi+aJ8pmsih
ZO0AZLvEEQwz1RhwvlvZpJQ2Uo7fWvjR64vV1WCCCC84AO4ejsiC4EEiQvr/aNbtRKxA+8VFCHI3
uNzdkhLimLPWzYZCWo75IgC8XT7WKe2ndgdTJRBUuEYbVnA8SN7daB26aZxbqrLXNJkmV6hyxdCg
a7HTpzQiyXaYvTtRy08yO+roGH+w+PWMjf0bGHc/9uPEzNLwjB8q98ptTgxtfcbomfVpquetP4Yi
Xp55yPDxP5U9G1S5RZT8GZi/KcOrdLc15qsYOxGIYfKuydCdil+3ojX7aemuwiAAJ/KhpnQtzR6B
d3iDJlP7xREV8cNNFbGiTPRR9cNzeiKjB050jFJ9XnNWJ1DbdJKOknKpkpb0ZfuPwgTwXClJ2qFS
52r4cPBgnT2Iz18g2v8sp6SGJBVViTcTbypQ+HlzAJsNyEy/EQUFv0hKhROtrSReKFs1AIZIoX7l
EME2N+B4qG7i50N1MKfEcZ2qk2HVjOmixog4GJdiPZIokvZFebbX/0zw/zbNgZrVnmMztCLj4qGv
Pzu1GhjxW7pZ336MQ69AYSRQyvScLW/+LoU+sEAjYaDWval846XDkkBAx/7oMIDP7QsHHuKl9MI/
BgtGLDwhofYjPx4EXBwoZ3WkabY80uH0mQmjqSo+JtWD1/zetk4ag6oqVifMnVVz9bN/s94qRkRg
K3rxHKDbfDGo99zID1eAUR8conaFNZiA1bdOv8jue6SE605l1kCclx665a80We5Wxxz7iABb8vcD
VUrJvz1rz3AI4ABVX8yxxaIiH8S6uGBfIMqYaunMC0LBWlIheg1GErjZabsv2YOJkDGJq8XikDjj
4eYGs1eKUmFlhc+ct+5xMlUiEBRNkwhUCskFFiMsz38M+9EbQoVvl1D3AJcngMJayPXmo5PLQXC0
JOzknbUQF0hMFx2AoyCVJKJkW8PfL4zjSIUv5qGXfuBQw/z9Zcmueqnid8d4qrVPnv7ivaTdg8LI
fex22pC9OIGLt5R8pZja87Ocp0PwgM0kgkpw7kDCnVXG/Iwz4hz2LWaCPhXqVtY6v1MDqPvBy10d
Xv2/cphZ8SVmPR3O5iICijJ8wCC81TqUpktYn3/UYEHMHG59sjv8HRbRly6J6k4ou+3jSDr1vfoZ
JHdKnF3h0m+JHgY3Fmh0szQ16NPE/Q/bJ7Olt+luP+A3poXwg2IyxSb/LJgVSYU3FLwWvwYz4/cV
RWbkc/vmrLyPcJDs01WLX5SRonzN/tUMnnFdPJVqF+xbmsBUp+E47/uXCA/gx/Ulw/b/kZhAY86/
1kgxkj/m/wC6VZ8dUz9aBz48YKw6WHYJFbWZ3fFlwy4t5NMQEMnPvuRtaBfrv1ALPLxQmg6cTIjF
ljycAxgeoCeQxjSGhjIa0iWPEki5AfzM+snyzBiBzDGCJJS685H76RqhB6bxwIMjfXBoKkANheDg
Dh43G2JwhI56EfTKAI3VxntDesXtD0EanUXkB0qU13JSx183ff0KkFhpT38kORWO8pYAyJIhIkuD
ygFq9jo2Z+/lPIXTsFGX39J0iNoJs4hXArLDO2ps/BMK7UsyflYdQfIp7eGE3I+xriR3BkcDo8Ti
XTI4JOfdD+SXu7YFueTeuDNii2xuii7mym+BVyo6H+yrae8DuendNZu+G3kYwJVXsrd4P8jDOFkK
t6ilu+agrMTKGyjAiGl9XbLPAuffkfEDIPI6sRVhI2YIDYfS6xN/p4skV3S/iPaOWvudcMiKdaWR
HE6RvUDRKawRvQ9y/xxdnei62amCQaqU6oSt7xd0BW2lJcdepx5BLtObMyIIIC+F3/mGCcn4yE9U
mI5zFCX+TXNeQ+m+GDabAs0NQ8FlZL8iojqCYSJZkRJ/2mS5C1syHsGb71l9Qf8C5yLJ1vpApvIB
KMQ6JwJsdoGb1TIjnWVeI8MqtwiumUxD5JgA+6JdDjiBfQITSepG/Ew9p64tYwwT0eNf1TWsqK6L
2wTE9lbCK1pZop1uZNXCUaGbqA0UPC0KXTJXvkhxmziU6tgwhpbankLF+qPnuIKZPBFxVSKjFtCr
S33kysaHPusW4HJcvB0peR12Xyb84/wP0w1Rrgju7157kuotTHo+BaGrqbqDb1hwX0wXHExgqQTb
8yUojwI8H0LDFWgllAQXAD2AMmySce6gu/Uy/ve/wrLX/xV3rXtbfVGRqSZH+wxqg9PJ4IF2Bwze
RoG6JbWDqt5r/Z9lYa7/B8RcQ/mIaz4PjoncFi5abNA/7/mp46OBaPfkw9nSftcud6j7C66o9agI
djJIc0RlorWqjxn/tcUbq8wwMMYCu56eYENgQCAaVDZQVuorFUYmvvQqFkDQZytf42gdVRD0is+D
hmIdR8Y6RiSI4ZSWJAOcPYLVZ8zTGbfOFR/4VobuvthmxwHMoKDwshgDHJEQ9OxtqOSJC6S3g00T
5ZKON2sQ+d7eoqrTQNkm9uRk8zZRVX75I6Os6luS98/9jkHaFv7CnLaHvfBTosrrjh91Oy8YMYRT
zILLg+3ESZsd0Kx5gTCbJoxUZeEEWJ05p5yvv/QWc7tLwbytkBgP0vZ8XyQU6AXU5OH4WvujROSl
SQdeim8bEi5zzXUAZtfKicV2cOudo6kkJ7Vvu9qxCBA0PUfCwJDaHR02Hb6xR2pLX7/OcPgJq4tw
CAYiOxzjPhfAiKH9MT/zcY+Uco4Rn49ZKh94G4tN+qyXTkeqcG8HvNMFaeZit4LVVfV4NH0L94iQ
m/xoACWUza00mELSIaXO0MWYRrCq2MoVH+igJB3lmA4gt98jftQQ55K7DI2x1HkQgCvixs47m9q4
xFPZ0rnBVxCCsa94RMNNOMIOTqwQaCMG93JEceJiUUYb6ByofK++LrDivJ59lVEzMeJBjhXpPbvM
Xhl9lx747qPhvf1bkrBdkiDWCRlFYWXtinmxrOdnMWkJnFa4O+miKrjlxmm6jWhEUmnEiZxmRf66
onleQv8jIJaMFSmg08E5xx5V0ZsqbYy0feO11ixRQ608t/mCfix4VecKnYXBfz3WVV+uTrxYGc95
5EE8QEqVvroRwTeZtCyuSZtX3Gpkkpz/bXm31FY4243iQiC/q5uRFL9mNosR1SIcDor2JaRJ7wXH
LCa0ml1ffG7Ry7oLihCHjudK8jEpqjBR6RYYNqym5ktblaexWABlROj3thANYXxy7p+3CkZ5i4Yq
Ue1/UHFUTEUQVxgw/y7BmNfXZDiX3z6EnILlY7T71uhNcprtceD9/MA9r3FfR6ZZ5ur4GhfjwPlS
B+gmKYJ7z5RLtmTA3tLof+W1OlTuCZBDyz3gqqjKay1hcdmg+hUeNG+zOgjUfmNw0LjvKkgBdOkM
xnFtxl43fKl8HBZpfq8fLks84/u7n8UEjghOLcIpzhqDvV5Eogw02DRRgMe7Vztp/cf6vZekYEvm
LZBFA/NQVsSFya8PK7iz1KKoeM6oK7TQja24xAI8Xs7S3/i4b7y/WGy2hj2uRFmRDhVdAMAKsmiT
QroZ3HPhvlTHEbXFSdtH1lHX3jLfhlXAelGqY0OC06IA/W4bQmonxRl9yOFKNN6EsVQ51+vqqG8b
mxJalD3VbOc7USWzazFJ21aj3TdFAri/KQNd9RCpnBub2RcYHr3WEJIF/55eQPt5eNohiIluktII
97NN7hj/+cSNm9r+ARgnuqiaH3d9gZL/b1ZANMydjZOV/vVMtBPJBXBqKSfJUp3ceyaHSyB3Y+ud
qL9JPu1ROkrnmeyi2SPDV257UB90h0Wa938/vWos+7ADh0ql7Hb0G3TNQq5QC8mscmtN7peRZ65f
tmFJpJujCmAsCovXMXbATvFW3nUazslI7h1OIsb81FlBbacT8LwNCHn035htWzLadIiaFn6b573F
4xDr0tspE27f7JcCLUG137R9ewptq6I95OhG2ffpIDuQlyFrgJoZR9xkZ/Z48O0zd1rnKXIJ87hk
H08feW2i8LiHwo4igV20TLTeHXFIghOWWyoj/H9L29ed+t3woOrpmKkY8iN3CtEKniX+tXwGvnSA
Yfj+/DVu5L/wyA781kU6PADs7kkSWicSCcwyBDXwaA+4Qvvz+X//SPUsXxMIzQDjlsw40kLuWuDC
QtSJoAX3uc1jxOqZQ1rAl1ljEfDSQk2KeIORlcFPLs6azLraRi7WYFBMLssVmjYzxvitUNVMNzef
achHpVUpfrKIouiDYObSUu8wF6mqxWRFDGn8Phjy9aRYSwikpY81liwy7USplsURjtysoylsIe5C
VzBo8titoZG130NahNYMgp1zifRsWTN/thi0Ww3FRSGXIF/ChO7acc8zoJGZdLEVUwfkvFPaJvoK
hovD5o8eSk+cieuVtHddf6bsq4y39aJABQr4AxzReMVgIktwaJn5QQNr4gIEJ3GqPJV93QlYEfqI
AD/Wga8e92vm/8HpIeCb2vwTnH4bJoD1NgUYKXJoZaiaf9jueUQDD7FBfpDwdUQOnlGFT6FU26Lp
xkp+P0bsVj/ZNj14H4a7CVIx9LNO/RFe4tX1RmjKtMnfe0/EKFtMhIBkJLe6+Xg6JYZLthg12Qaa
rCOh8pegDHBD7OiXxXSAH2744vDjBYca0bxS5J1TkFdUq+gJM0ftH5Dc089apz8w6DmOAEo5imJ2
3ua4ikigllZI4E0L52Xby3Hum6Ha7Q6Tf6fRa5c0m4f/zEAZB1O3zKVie4+MC8ArCSF4Z6feNk6f
VoxGHAROw9WwWww9AChYJLYkpZ0bSgDFATG0ezne7WTQCaLtX+K5I4bVv71rj6+GGXCxtrJfCuKB
8cZhSbjSGNZgjqIjYufTAhhrHD1NXHHQtIlvemIGmCL/WEQhA3r+gr3eLCUKilrwr0pyu0Praeu4
G5Jx9uc/eyJYX0lozAOiB0ndPWukrsglS6NWupfFw7K8RENLcU36QudQmT3f+euOhXNMYdqno4ZT
TcfjI9wskGMvU/KhBoqw6QnecWB7AkM7rUgenwL89zDS0ubwkhJ5Q4WyvTfMV0iPWq5ihYSaSGPD
+/aO2MgHHXEi4CVcskxmtPbOCXYuIv/syFe65XpuFDAcDXdkEe2/XbO5dZ6NJk+/hqKZiWOk9uSS
hBfJnSg/6fmquyYIhXHwUnS6QqhvLG+FJ7iWPeOtaFdghxlhLHtMVgOwXDfEUaStqLIaIIoToxDQ
iAQNoSws5k86qCRIgbCVE73otqu1if0zMZkt3dLGifyD6pawMxigTgDBct92fOKYzCdeoLRj8PyV
GDgtX8kHcJ74K2zQcN21KCxVZnhUcFn6hHwRy6RqEvArCuB5BzrZNwALPp7m5Fm6TL52jxoFUrGW
lR2KLNCgeOXXKgJ+2kwXpsH0rFk2r7aOqUd3qAGvp9ghT/wtNuwZltFVliXqwTUlwYktlNhAC7mP
sP4xodTAyGeT5hv+HIWawuF6F58ICz1odCWul/xGXtL0CgW8upbi7wOlnaMCVnuBdksAHY8QXw/H
bCnst0RW+tVO9CMkJ9O7/xcwGjGJCwR+y4PsmEjhebR9DJ/4DGQne96X5ZzELb0IFmJX5xe+QqyV
ZDIDnVPMoRJfjR8qWrnRTUdiGhoAau/g5SxNA3oZN63rzS7tKSYJ/nFGLWxIQzG05LmJPOegEkyz
6uHFsaeuTofK1/XmRS43XvS9YM8/J7S4LLv+r+RNyfnbbs6g+4Yrf6H8p/5OEw+eI4JZspEtt7QX
BRLOVyAG1UxpPVrzCeK/WcK/Y1taDtc/BJ4cJtDqzccDAm3+7zMcyZGZY5Szji/sPHIcDaP44G9S
wxSZT1pTwqgZpLuRB97BDH5jzDvVgV1x2W4GEV4naCM++mpIcAv3PTWc1iKR74Ed+Gi7/60gNXhn
aaytYQYx/aAS0sWTBwZ8N23QoiAadqfhVx9f8aTY3arDispwB24cAfD6oi6awkwYm+S4J/tajKkM
w/G8zOQMiW7EEqTjw9SH1JVGEFODudHUIyLqwH/W9LZV+Pq87wdY8KRIEWM89oU9ghxs8CSemW/3
p8b5nbhTbCQframeNHe/vGfqlo2xyBTqQoSK4IlWQutFUosnHZ9i4/v+H8aE6eImLQ2JemVuyzil
f3PJDBq2bsVvIK9pFSjyfgc5IBSEVnexxaAUW54v2AYAZXAh0y3Ghoj0CTDV8tR47Q0/xCwQkhUi
w9w2a7eV8g8pqWHvdxhP4dcCDp+IM6kAqZEted4LseK5ZOuNArqk49QVjMn9OzaRrSwOA4QAW2CF
IvGBz/1EL/M1PJA0QwB8BEUvV1tcy+xMTu308P1vvCZV4A9h3NOp6EOZGZBL0E2Wud03Nvlyd1cW
d+s23RxbKYx2RXeWhUWMbhInlgCG2BcTbIvHxl3c1jHP39C7zInjY5nG2FKrxLcSEOcIeif/z1NN
IWq0OLOrG8DYwVjpClo6bTPnIXpOZt0zEYyARLxLFTzbrbK3jry3rQKZQa1bsR/fzKJUm6QArZTm
Go4cgoiQjOqm/DbDNVr0ExD3yA2Sxp9zVTmfNKJx3tx3p2IZL7yg+1iTanSgGUm5mBT07etyddyE
yLitz36/JxQYTEHhD9rN6lIIO4vr4hHQ/ZneaTzjgzZcSIZ2V88ScN9Z4Ing8BxXAlTeX7mNbZ2F
QI5dtl5kCcWc/lhX93gicsmfC9EpP8DHgM0MyJCZbKD4md/f3pFx8a+dZzWYTZ997TNVv/Ixo2H4
fKS7j+VdI16o6lJAYxQu34rEhRfEr8e/ZMWoZ1Ih3XO7p31PSCr7NkD73vbMT0CB3p9cmc2/xBV9
+yBGzCEnh/OEnFpVwAt2J8ucIEPtayipEmOc0nG8xOxsVc9/YQZ0u0gceDdYzL9Hx+IB2OpNS5Gm
0RAFTnC5uWJa8I4xM4Y50eVzs0ks1Sz/5hEtyMOR36MvJqxQdmcgexM5PVIuLKFYKS/t5Zj0aih7
Go4wHq8t0ZHrq54Cccn2RI/RWnTTzdWak7OSQCvC1Sfu/LfC04Y7bSXDZe8TH5ksS5e4XPhVUMTj
NsRP98/PX8MuyMTxztP5v9UMbSwTN8174ZlJa6A5sCwPmMc+7NBBRQzwvKAqF/20G+zKpoajVQvV
Fk9rUdXCDyXWKNE8mGik0DjC2eOKYh6K2nbzCiMi8sdoGuTNlMx7twdblbmpJzXucSeDekW61QZP
XBBpb7Sn8z9C/vUmJIq5yVA/DF/sRcBUEnMLvWLEMiLNGZH4GF8+pmB8/cuxLWNM3H9s7fJTHtqu
BPgGRk65kjFNHwS845gK7IhubnXAWm1nXanOsj96Rd3aroScCp6zPCsaFPnpgZVSHtVNkrBEdHiy
vCaO6cGWwxxoNoeXgP3ubdsgKMW1CuWJnS5EpscDR1M/trQe7geCPDjr359KQhq1AwrxhYqRce8X
cOFeZMfEuDatu4V3/O4EHZ1v3PLjwxPVKvoJJEylzlDGWx4a/ugBd4LcERvE1EtrwyjKAPiKrmbp
VQPuj9V0YmKmf5nwZoB3ccerVkFgxSit2ejaifzAHZREuTYaOXwoRo4DGSl8Ud1hK19YZVxcnG52
LymdHK6rlbJNrmqjfY7tUZDxa37bucxWbAoVK9+lmO+JjlRb1N1egyKyh7wf+gYJM10LbcVz6KDR
xTfD3VucOnQqG9lYrDByg+DohOB2OdkYV88tb9LwHMXgoJC+LdwvkAjspM86KcH7L2n6F6rfvzIX
/bEEeXHZ0TqZUDZTDvKKI0N85hSm3jrX8rNJsWOm6YMrtfXtdjotwJ3ekvK+9Kc2EOwiwqdwdQBl
dxgUyoItXQHBiRgpQ/4dP2phhqcCwOqM84/g59fodVib72Ihm+GqlfkNniXvomS7kLZo3eGNWA8a
27TukHOHwx0SQ8ZBu2x38+ZCRGjGmigqGLKXchO1V1raHD30gy3i/g85C3cHnDnIH+WATUFkTZRv
BMHbxVK493swCjdUl6izZEhR6cBIdbxsvtBlEMXcjExX7mgqQ+iSYAoRbG8DK97exxyFf8C9bJ/e
0FfOgV4tFiGgJrF3GlsyShu1PyhzTFkIewaVZA6HEszTDi49zf0mzdyi91ZhJ6ODngIf299p6PtB
cStceIpee54ydKbJEWrlZPDnJtXSCzH9wKgCtnW+MvhMfAJXUhdy3dCzoNtBFsYIp1zL05MUelyx
eqIT67C8UY828xWELbBz/sbhkSKSAu3LN3qZfysnri1oxljoxDQOnbhbOnqCJTTQB84QGPMNeSqq
mdozmNesoXkTQiJTiDXaqyW+tMNti+iuvL9qqm10CnPIlVMsPbu/QAqRzLTo+t+ckekBIYNJRerZ
CaUJJNWJpvfKNOnssgeFAmSLf3elhb6uCMw1dtXf6HrHm5jaPQNW3jkTBH0unCZleYQTPYJEvMaq
frOuPPh6M5jFueXXasL5yRw6j8qigBlGXQnQEC5KOFq24oRfG2w24eul7Ol1vYmekMLb7p4PEYo2
a+wEaJQ0jzqYXd4XvHPcWa1rL0ZmQCkhdMgVAmvn0gVCbQO2p/GYiw3x+zrW8CwEevkPtbi87tVu
tuPaxqbrT5BfpX8hiu8GUcD2TeHJ079qJxWgL/FC28JRiOzvAzWif36Nuy1qMsQH1D0sutIe5OKw
I7z+5sO5wdZWSG9lQj3TZ/V45OkCNU4Vw9eH9COmv42vohfQss9MGB5cr/7XhC/TTZOJOBgHjq6e
Z8vdAvNMmx1JfxsXvQOGhk/jM7fHp/I/DMGhtHCI8A21ZBYP7WLOmzFFf3AihvGz4Jx1aGGc3GWK
aw3s3COwdjHXQPUc7zJlFNvuk7Vt4XKkOL3WdoSTwTy4KGjWY7016pCMdhF4h0sP9/GO+K64D5ZQ
Ji8QgkOmxd8y9hsF31QXlitK+2Acz8hHUg1QETygwOj8YNPXvgRb7fWzha5EaTvzWffsevYh6dRC
UBJWek0lwaiy6RteHVFkSP2cdJRPADbBbbaiLhx2lwrBmTpUbk9GbJwGKlm07EcGNaxllj/I5hsP
OhkOSDaB7jsBjzpL9S2VMeLD21XcOJLoCjy5Zv3XdRSOHwWlc9tXm1TTJ6qQYG3/tnoK9bYQu57T
4w9nqJ8KC8N1exockoSbxh0YWWTjeHw4Gq1MSOFJGZPBvKou2a4JH00vZwHBWLZsYKqO6QlVn8XT
FP5XHsJXDNNWhhc3ZRr+Cly6oCFIsnd4JMEAdRPqYttK/xY+zMsO5fPT4j6BiEDRa/WXFLeD/IyN
SqmbllAmJ9KfVRSEKfXbwUGXV1eITqPUSXFJ61d3yQ553YSSU68W1FaaEmjxhUJwC2CXbkrYMonE
yjAn4EdEtOGTlqTHr9ELN0/PuIapB4o4QCCo3bum2vnRGZOWzGFOjjr5CF7D1QniN1t/8zN1HsIS
66P7YjR1TosArU2jrRZ4LYZPHeHv21xpxpnBG+k3umrYwevpDgamMQCgiAA3w3qxRaxGSmfyyfVD
TyPTquWlx3TFGQbVLf43h1dUtXPOpFvW+cYWexU/ikgEPo0DkMvjQ7H8JJdhMObKrPm4pHnX6n7l
/U1Ro1WZN/A2ydD16g3k+F1kHAFRe2TBQ0PowbbfLMuWmRF+/YGVxwsFXrj+AjOGmBoOyQmPzpWU
5Ut1hESQ26ZdcqD2AGzkzCec+tuxepFh/xTkitnOZn3kS1kvornhr4XlKcRe4bcTHQnB4X1BYTUj
GqzeTkaVuSQwHbNfVGDGcRLUznG0Q6Df6L0uBFlyM3jbd8gpO60WDZ85JyNn8sdE53NGjumoHfdw
mxw5YQcGwCT25fLtPltbFrUVobjyhF8tdjJeDIykoMSxh18K+dGgfU8VeycDxGw6cw/h0RqeThST
fhZaAsrPFJBx5j9eXmY1eSZMdVlffOPQFSChTsA/Al4Z3ABwvo3FNN5DN95gRb/fN6VE0e9vOFfR
QbS3IeEVx0z+PTipvOBnTjFEgyb0lDczK8GrTYg/GrFLKdTtyWzSjTU4aoI+a/BOiP4AQJKLY38G
erVbQVAIjqofSCw2xVDVOdIbs8Gnws3ozE528lozRdoMUZCywuOd9gtEebo0ULz4Bmi2GiTalpK9
eNEZ7iQcCvsKb+GfRYuBXJkGqAlihrfOobJrOYpmXxGL3jlWKxZraMQb5dEqZK63noFsoFuxucaj
wcaHjk1m8KrHjOyPHOPPHljUSbq5/KvVew84QkrePJ0KTUcouNddz6jFWN2OPTGGHwNXssGKNWHz
QXZzChZlEZ8IcmR566fE8BxQrnPKa2Z7Jp5klNjK8wyOspnTaKggBBn9END7hLThMgUSsu7mxs5o
rX16EKauEpn2l+LPtd80sZ0PZNfsdIZjM3Y5JrReAv65TMTlpdQ5id9irzkN+ewId4DTBlCMblFO
o5cfp619mbfsCN/YwkQRQ3IfQJ8IQiT4/f7+reaDHVy/B42k3Lm2sGT0wipkQ39GO6O+TVC6uxZM
JIRzEnLN8kvWNyGZ/roKsPIPGfPYIC3hG5aJ1acBMf4KCFyYoVHM6JcvR9p2m+O4Wg3km3uHr1wf
2+VvdzdctZyxALx9wProjCK2HWNKMlhs2l6KQgXJsV+FiBAoSHIThoL8ZgwL0MXa2NyP93ZO9QlH
LLxNNzh2I8EDR10H59dOMMsNcA016I3X9SywEWv3tXGro6q1xnTr0n36G9j+jyOBw3ivgQHCfW7w
JDP+4tmrKRCDxqE+9UIYTTjACu7dB0g+5EHrnjWWfmUOhvvTP9gp4ce0MdtLeQB/1CQ2rIB7BSD9
mc8LNImc2/JFUZAVEId1ntwciXU7fXqf2+kc+Jl9yV1lqyVcOn+tXnM61alCEc0zM//S4p+9+WPe
MsO1d7mJkS+Ug378Vxdh6T4QZ34XrVkVyd6QIARBhghbkOEe8RtWwy+qPwciOV2X9xQQhJOgy6xw
tKTaPdxPfYdG0ixNqK4MFyVKLNnXxGd7mzFkYDSMILmPHPcxcy+6ZAiQQjvFKVkU20Q0bkUY+91z
fnvccFBUHkZvICk6lDnbOiiozgJx6VYrR93L1WAdabH7+9y9E906gpOPWd2hO0lm0kmka3vrmck+
lRAa96tfBmCntaQURYVwpCquPchW+P5aOmNsZJmSHlLtLLnc7yyp8wYMWkLSKaNcIbrv00G8cOHY
8/ZlnS+ZBQ+KaoJfok4qbSD/v+xgkGRLFFdAIjk9nMa4MVq0dKiWKxO/okaaWDsfwblE9zAqMA7M
M5+RAPSVI+q8YmBFN33rZ4T1x89+QvOTaszTj8nFH/EOuSo/REF2YStNyB6c8ToE+0dVnkB2VxXI
5DmEAWQlrEtk0lLJoBZ4aWDsavg7zeMP6OpsFwoqIG8wdq0DqlMK7Q6y8R8F1IPW2DSrHFSk2I+9
djuPubynMLJLEYvhigHJfl7mjvBUp2f9V+rAgatLv2e+yfSFouyjdGF7uTICQYCiRe0Dd5sBBT69
USGCPxCxam7scpB8sGOH2LfdpuHkHBSK2qFrcxMcyMmPix4wVwal0pzx190GT/JD5o1Fr/pb1mTl
4GE8j99vT5+MwKhLdH86EcKRRR74MRefVrDzRCh5UlgZR3BcA8FcQ6bzGHyjHSvg0/pwxRWWLehj
Z+t/LXdJSNSeNhRW/pVj9PzclnQ90ewfk1wa+H6gnce4UJ7mUz2HzC79lzGJYyvvJxzbp0MTgIFi
WLRaRV2KQ6VBbaHdRLDbS5PQkejyG0Jlg6JoVJTi7gRm+86Qm5alyxuGvDafhFyCu+YT6qhnMb3I
3hX7Xo9N7FUWfcEkJdi8OzZi+U0s0R7oyqI921QdBF7tKLHEOmIJOvtoy699O/cEJhnf8qx2CSjn
9jqSjmQ+BrVckH5c8jvW3RafChEQh9eWmS/uufcnf9qiRB/fUaWSTcJenZ+CqV6paCMQ6EJEXnSs
i+nWalL78/uMTvUETrRpGqsLfQ+51iZ7yP6GTsuXH9iqY1cpzp/0JLQtG/idDkmgS5CHRjcws1t8
rrMzEfu50thbe3/o6QZQyCQO+caWUcfKAesKZUJnzvsWPXtSjaJ8f3dNI/KeyxN1Dm3eeL+Yyusp
Wxod2/WBhxuQZZYKHFp9TmVnxLB37jgtHq+d9UBSsD39YGh9DGgUgQpbdAnD/lEc1+jOYdh1rRuJ
nwtfsXQ1lBGQYCUdun4udjNv8yo11q0ZISm4ypNzwD6HFRuYv6dLlcJKltLrALwne2XyZjpXrAGF
a3ZmbV8BtmeAC5MGQYuYNpOC+6psA6+zNd2yrE8gWZl//sj4Bu0pltMAj00spSD3Vb9HaBNhPcpg
hqOpRmVKnJM40KedWIXwEoeC0euUN1Jvbt62sza6djf6tlt4QCte2b7h/a/EE152LMUf73MX9pMi
w2GonGMNNAPyqvE/RMDAYb7himNXQVGFqlqY9wh3OIrug4aRMP6FyJQwAet9cS008N1ikW4GLCgY
2lKd1Hx19okYmfXZT/71Tj0JGSXaEoatJvLS+WG9Jnbo0dMqJzh0IrGZQtiDzu/PIPdiTwclfheX
oxv1oElwDaK8aVTYtaHE1+UK5ert+MdD6kqWghIwUb+A8JYVxVBmDExpwu2inFg+7icVpz96Bgrw
g+Un7gLRmEPr2Nr0PKDjuMliYNj4Ub8Gogk0OgckONZxSdB7TO+mTljfVfP/OpYiuXybvauIFyqB
JVIa0OVNb2biXOfDDkuuT56i/mWaDBkU4+3AaTq4n+eRV1hRO5BrcNvaRCW1G2LuL5OptV1h+XW0
myQJHna/+2WV0DcMqz8Og5Fqxm5zbeKblNozhiuQu3sij9WJsWTiv1fDd74CkYpDRnjaFGxdSOVs
wZFhhbjAWtwzHmPI95UhxVM7pu7I2imgE75+jJAi+2gRBlp4OZt0+EH25l71hgcHZsE4ziLYsyCN
LA4kNzG3NehLpxWpaG5KhdBdxbI7X8tdQLW6GBajE5bisarzJ2FTMdd0n8ysbXqeHYYjkGeBuyXV
ThAn4Y4m6h932ZP2cBTtD6qYqBEq2Ri9SyWGG3L+QuQVg0C1bzd8kIaHlDPLK1xkkhZqkgzGdOjB
UOnyBi3GV8TEET5yLUtmGcGNQU8QiuIGtJgsHeo90WX+h1lybRI5sFDgXKVwHx3KGcJNAVlSNiTL
0NRs2dRjJeU7H7CTtdMTwZ2GkLRGFahunMC/WWPriMJeUJvKuY2z24wRI4OREX8BdoTdNSpAB52/
s2P41/DGTx3iCao6mZJQGulTUc4y2hb43Cbco7Nm3VIVTEG6V/pfNp7yCdBKj0zkm1Qp4k2027l0
tyA2wgP+P4jfBy0VAi5UVhoAbLQm/T8P9iWCSlMBqaLMkJU3PR3qfmVMky63QAEDX8ci86bZ4deI
7Uu9w+03UbYb+/scSwCi651QNeI5JwusN/X14bJZ/My5Qe30rV5ceWkzxeWwj20cwV0B+XdzuiQi
xO/6F81yOjAbUsl4WKFe5CnyM9hTLxXA9nfhdUjDWgAUJeLteFOjjf4v9manSDEW0HXDa4aVLrl3
WzBj8AnRtrXlrTSGBdqBpu/bTt4emFfJWHDhjL0Alnp6XG4MaxScosqfPfnrm8OynJW9DUinULNd
hppf33uIt46PiUQONSesi5lEkF0l+8Lp5wRv+5lShhPCbnnBPDQJZLmLvfWxCGEkeF3+xf1nhwCq
2cQ5c5y97m4kPhB+9M969+4Su8YoGFp6qVWLxirT1Raknv8x/O8zUXdNBoIEA18wQYHBGiDkrzGO
Q9G0Q4SVCCxAxjE8ZSOEgMAXBbV7B5gb/y8YKBbkmQ8OwhYlMhQqgShFxafeI+ux/5k3hvGt9/3j
gjVvXCMe4QvDFGdce8Ly688XIH7/q0PfBYmh1DmF66BxQ3SfkXT6V2Enwqs7mSvf3OOG9Y9oxDXG
73VUkgn+JrWiH8a16+04i+ZqQTqjTL02bWb7jaeJe5xxjL3WBKExqQqtz/M/o1lFDXi5SGGxpzqj
dYXRNeRdwWQTHWIcP5zEpPCzkVWVkDer6h4kOxcEHDFKdVJ53e5porbHVFpflFwDXq2B/OAw/JZP
KB1kfnROTi/yH3usfdEGSht+zXZ0bCNl2ebfMp5pw75qnkrLASeD3Rt8/ncI/0dpbGzXW9/DxW1T
IBqbipajtmHLDdrcPiZ/FXvdKCNFV9lrk3ipXKXxRGE1UVTkM8azD6M9Fg1nMvq4r5kWVDzcreKw
uZU9P9WRI3inFfBfQo9jWMNzoBiXIh3snM0FHR8DYB/aAB/zwXAKh6RxOkw7I09naGDyRbhS2FmE
gWt6+5MTXCo5naptDeO3Z8WHXL5RReosMZeLH3sM3XX5zRGpy0S8cYoAlYMQd8NVssOdlyyb7ScK
vxFmJTU+npVnOgRtd5dCRoFOkyvza0cMN6+r3xREeE2+C6m7PSgb3gZ/n2dl3y6nI53icXpt72fR
lJ/zllKOeyr2Amdkr40UajK5C/7jdoe0i1xzTVetXfbhX3fA9XRncf9ad9lyZAM7/VeeMhU7egfN
e23rxOO2CWVmoba4PNwUTX5ifXkCKrNCLtUZbXERMgsneBSVSPUymvPq+BbNUpT/TZafowyLihsB
y1V2Oozxp9/JiaQbH7JrE+hsg9eIKppgs09BFSoU4WGXG6mFHAQEwSX9UMGueGeEIJStURPTXkMf
cJcpsQtQePKj6YSodyogZQDRrjG4nH3ESoP0Mc+jaixLrFXzx2IbPLzg+I5bwnf8XYrjkwrwW1cW
KBRGSXbeEbtkKD3/JfXQVOUCqhPqPcwqSIBOnNyeAO0Sk39TiWj+e8fz6pOo793m4neu8D7uJuEs
NYC+tz3J0BN/KHp7KeNJfTJIO2uWygGhNcE61/5IFQYtzPxKHdbf2i6QxLfRWydHl82NeadNxVTh
/EYYeoD/Gqs9D/GQb2ZXjmX15pp8ydGrw717DdxBMhkFYd3AdkMsGFbN+UaYW4Y51JVCCVIjDz9d
LReS5xoP/oU3wB6Rh3ROaefGZNvQXm5QzK0vvD29nClEdMevVTOxI7JaWqSqcHnH/YWQT8DKJorf
8kr8EJNCtbSOWGMumnsA9uoigb/wY6j1m00sds7Auc6B58Yyn47HQEMIP5M/0/vPk0omZUA8w0XO
PVfsmEMurjtSaGdzzwzPxubp61+wqoVBR9UDtJdYB0U4SlMgYLp0+7A6LA0lRAPBpBArsIniN+tn
zKrqT1BWVXAh7XhYIrfx/0z2BAzOTNEmjGIn1oSECznP3wrB1gZ4tsANNXCeaXDsvGjHfi4rJ462
C+Smoe7uJ9n6p1T0UESbvjI69VtucwpoJhu6NGCU86ILkk56gSQviNKdk1tFTKEujZ9yOECsvAPY
u3VH/byPYwOnsMDsabx5X4NW9USoT1ssPdREuHNwtHWGpNFstKYPns9JEz9hdMbVvbXQVMCqCU8c
Kileo7+j6ZqE3GKDucOOwrFxJOXiHugQ4ZmuGJFE1FOgt/ukVIslSf2WvGrod0NbufYe4TZ+aYox
DrIngMxgImAu+i8tQ3oWmiXc0MKwkCEX5Ti4wjMIrWTA1DsH555+pgwnPKlOU8NI3TFyDObzoUL9
bfH5LDKhlXsB2ZbgOAUBmBdE2TOQlUUC+dS9Ho/a0lSbchSN9hJWYNf8KuCLKSccbr0Dg4gqiNv8
3r2nvMjiKNylD/b6fmXb/i6f7fZpaRxSCQqWJXk0EEjXtMlmgtp76RR+epg/zuodNTvUjUvnwwSF
n556vOBk7pbDNsjMko88pbcxXgu192pvj4NSe+hQaylVoCSIsXHqOs/gyu1yHfSOvIz8B+3yN8lF
dYXEWIDN0JRrfVrOH9GdwDhXwHYX5d93VCiynH2odZFKOav5FDSRdGFtOYDOu3h3WTztP4+argut
QXjMQr8uIAhYimsvPL5Gs5swVvq4OY2XCVZvvCdW2qU5wjStuVFpXL32CCJrsMMdkOsjRUJcB1w8
fwynRAez118wZoFUMp6CPmc/aa3H2cFBI5f2xbb2pPv0sp5kLy3KxBLrO9zUMro9H/sv9fVc9A6U
A6slK9AK/FsgFHJgIOfhkFDDwDZNVQpbVyJkcDnif0hPD7eIrEiXSIL+NUN54e6f0zEhs3rR+JWa
SGd5S4VJS5cQMVxQ5lHzbxPI2VXlj47HaFE0dvJ3+HgIT0jS9R7pMj0lj1sKTSGe3FtR/RRaBxlW
kx4Q3g/NnQHfIsUBGOAg+eNgf4Epmkqi0HJ02sRaVd/QeXMGn8KKoOqlDqtzkUxp5Fqe2TXe88vD
tteUOsO529E/cSbRL8g/KIsdMzaU3F1JusVcut5DDRi3iYQ2vVnkv7QsBFImN3mgbYn3u6UnjLuW
UPWxjWTUBzii8VJKs5IpDDpbt4XiV539poht8Z4W1MtZW6j0eYekktWo4NZYmqTwXzCzBSCsmAPr
/uuHijWi21ojBu/6Ni+I9AUe8KWb1dfU9C+a/svXeJsAcNycgWbWjedaTa6dWcPP8PhsSvyx6yVk
9gwL3svLvMyvcV8BvEa4eoi8VxtPlhndRgcK6SBlfpXlQH+s1ohitLMZSuWUNMKk7yBH0D0Df1Yf
Irp+3DUHUDEECRZOF56CZltqsg0wRSCaq98AbPdN2pol2s+SN3GTeM+c/KUdjsw5k5uyAqDt80lj
/k0/VZnG5lBk6u3BJLa7T80Vd+JNExYmKNvLBVVVyv31XQc1vIhYqQHWoJaORD/kCPwObk4AL63i
bv3+6tyWn6rChEdEe1ka5GJ7GkBnygcOafs3ln71gPaGr6CCTxxSOTzoJzTMkRtaZO2qsMxR61uZ
/K+b2BAQ6OMHV1kaBNYkfmKiIpzpOOGCMhM/ID6DwTT61H4G5UQSByGOwpRGo8q3ROXkUMIj2IlF
BMw73c5v6XjLZ8gP65rx0ahxOSbyOXhnH9wCKrL6O7/Rxk61GhOx1hqUwiF9ich86t+1+NGqrjXM
qBZkOhd0ai5VnLEMGyzddV8Ps7qXbFaJydHL9lBS3ARh6XnMyZRBFTqbbTMLTPKGme9fC1OoFkC9
0UZeiV9PgoXk20XWTqJ8Wl3f5rHIwV8t1d22rMNLVS7UeFb82B10CwXP0K2yt86Zv/1fDcots4CJ
3PFCk8nB3/bEWuOUwLo2LNWr1SZTt1pSH8wbYXQ1Yfc5M64V7zv9BeMmVD0Ayym78VOHqclZzEdt
HsqkWz90A/6+SuJ0npqlNL7iTUubuNpuApLJVbstVonDfqVLKK3mn3bJ3yFnn7UF3mzgryMPGsOh
laxtHYVI8CqcRG2b2bmFovq4ceqrXBg48QvVTc3wU0PPydFSimn0NrKZMfnoW3EhLxNiRdMJsF6y
EzLHJhLM4OMhcz/Wo3KNCYz0HjRe/yKyvat+tO4zfXhAsfu01VKhdWhOhNKR/va2w+DDi69R/u+K
k/Bq49gBJo9KqJFrO9idBE3garrA1pIJfapUAQpsoN3SDvhp8X1n0V/mZbXKS4i2ZayMNNiUycFR
jBATvoRfpYpxFb5PkqK5nA01pi0cIUEc23C6/bL0brxmasXfItJEByaq5l+OiNipzAjoWIZ1BFWq
RiP6Cmd017YJ1BGrmgnZQ9hIkEHs3Bv+fjy3TnoZSXjXOv1clPvfZteOzevG8Abi3UwyoIbc6TTV
IH2CTG1aPfnFdCpXgaRNl6uZPPRg2OKNUGrYGWN+WEN5iN6iJAo6GjerCbLQnpBWU3sEy1fp4zB3
XFEX6KBJN62Gth6FtieSj840aC6P8Pc0et1MYkWBsCClaQDb454noevopri3mcOXURxg50Ivpd0e
ORwPfMto+MBOflXpqUCJtUDBAb79JDR4GTsEbSb/h5Pg5jNZDEviaQaE0UbPFOSj7JOVPIdc2Pr5
iAlqqX/Gj8Fd10RIPz/o4U8CXuLGqX82UOft/3jcE7POQnvJcfv7FqqJUNMjdVhsWV4OWq9BBhZ2
oBuiCdXD+ODVR9k2SK3eKZvaI2RQP6frnX0Ras8gwnKFKbyWNfg9dhMjB2WHlCjEChyJAg5V1BT+
6t51nCCkBF66E82ED4L3aORe6/Y52FjxTbeTn7IJpzWDTBbRqJ8HMLdKzucKSGweneiAUgy9sB4U
cdSsyF0K5FR/ymXZpaDTNonHosF7BGo5M2OTPTu2s9FjTGP0CYUuJVSDy0MbLGKW6IBcgIWfKpgM
NLNVWYVrmOJBe1S6m0WJHO05zQOLv9TTClQUpoPoURJbpq6dknODK7+XFWUgi/9hvf036WXB+Ue/
yuatuC9b5eA/SEkpqXCoZuy7ndNTHvfEvHxPsc0QAYmo2aIn3QyCmUUVGqlWRpWtD7MxgW3GOGJJ
aQudIK9u/NfPoSNQ4rv3X1B4AEq5uugr3uaR1L1I7PYuWTMIJQwMgzTjHklXRai0DjkVRzK1ah2R
m3a3WJpOp9ajMem54Hykp/Jel5hzvqs5bf5roRR2TS5gFXjjmJAnaz8diA617D3yfaf2li4BqsTw
vqdKlrqpQqJfnX5qjhWmBef2X4Xnsf90zzi2yKpIJ5NHuI1DUx7lK0jCTV66v4Qjmmqp8an67KYk
9UsOlcJhDWYTkSwBTqDCS3NtTA4ovYe8mhAWAxnZSk+47e7SRC9ullGJYpJ7m19T8WjcGcV8WYqJ
O7oGuwE2/vkDUN/3DFH4anNCFfa3QYXWEnrslii7Nlvmqk3OGqVuS7HH1j0UVTrHygvEQr7okmjF
REdLw7PAULh1IZ/U6ON1zCFLirZjbV4kr7qby8rU95IQ9+un2RTYFzm9uK1ACcOGCrSuKv7YhDdQ
TjV1B44LsQdT5iO0jhR7TU6B8glOagAH6aG2SHxRXP8RzN4MuSdyDJdlQm/SxA0HWVd1p2/c8HQ0
8JtAmP/9aGWZaFe0jfy32Z0BHnkbdvovk21HL9CTGS3+K0y9RmXWyTxTw7b82M/EbMD6YdROgfxF
OJHxVzFZvcATzNDmeJ/sy4nuow5quycblCorijEekc9RkI4zDwej1SDa+7bwHg30rrxJywwstgq/
XrnW7dtI573IXYtRUKl0o+s+mx9lreSnYTFGON37KTht8U5ZomdFssFYyRly7mkyfVIFdMAPOesc
71fCGYdM1ThaDMQzGTc7GjPhErfLh8OF9xTL8ZoZ4s2/IsHVIO0onUhHb33mEyDpdtGClPRTEIxj
Hh6f3V6wEThvp50YVAXgDenuri5eHeB4kQK8Py6PkTIAHd7/eFB+1AqXXkeEeXX+Oyo+p3slK46O
pvvZjTnMzIJX0CkiKd8hwisD65iRJfReGpawLFp5OY1vXGuMt1cgLih6nPdcrfI5H1DXTVGiyaTp
BYBiYbOmPgQSu4DBr5l36a5gfXAF0lq2GyvoIA5IDXHHKrM1b9w5MFa/88/40OtJ/rBvgCiYOn0A
WHYmiPqIZMtBT/scZtlKSDoa6qodq6czO8KvjKDfZyIVTylrFmyRdD0FEH8lBaOSSo+F47TA/AFv
FntII7im8RjA4q9MpW3pG6h7X7oBzhS/I6ajAzZPpLxc2mDdmm5+qQb/C4H9++tO+baIEMXs27vf
Ea/yZu49ZS3GB4ixC0WOwqzgi8q4l6WHJsSIjS1TWdcJ9y6bx7EKC+BAPfItkrQ6aof3wFYFEm35
FGX9xZbpYAULNR/tc81Mr0sbwkDer/yzHJb0H0uE9/wGJsLvyFGEpdd+PgfMutpImkz3gs7u5rlX
qyUm19Mng5hNNT2LvJlqP5zEc1Bvv20a43/cQQhODhXfa91lCP/jhjhLEHDLa8puZkSl2ViDXUlR
but2OTnbm0qlsv8nGLPPQDE0jwKHvSnTo2+1F1LnonkrAERdrCq5VRyl4B7/Usjgb7l1NT1UzgEV
IjegHe/ZEtA0WB7tKwzU3q2wFyX/EqyFBmqjPMCt2A//IASgChbylaODod3ttWvY/8aVQW+ryIOR
W2Ilh/JHCbA4r8Qwl2RZ35aV8DueMsM3s0j3Zw5FcDPmF6EqhZsdLQfzEe7B7o6A2sjNa1nCJhJ3
Ex+hGOg03qmOtlitulu+oRhpBY+y0qB4Hj503jpHCOcduR0D5e9IEkppoVYsKHmZVxgfvyYjXYyc
d/ibhSHL/x+D4Zvi33ldHXHYW0ivrOIj/t+LC9nXUakOdhlRBvkld0nmD+oGwqLpip4vcnnrnW5B
/h97szwM4oXXnlVBpvUYTFwwkMQ0TIAP0thycMW9EKO0d7deQksSAaNtpzjJ4OBJBJN61M1CcaQz
VX0GqnZuMUsu8GlWArW9G9soEf+7KtJBamDErPDHT4HeDYIBM+pipSxwJbMgFEQTu+EaMgpPv1Wi
LA48H0x38D2ITRmsY77LCZJXUASYvIcTFM3A++FG/mS6tynjKqdB/13Zdx1RzAg3B9TyF13HaWe1
HRGkUg2nvKDofl1gU2xzZb3Oh034WiALyLmWrywqvDtvSDLzl4dbo84dRcIgHum8Sayy2pPZqbFA
uzQN7dAWX6fqOd1cPfqaWYk5VAtMgpTYowtFLfUBDNG69uaLslHXsYgA7OWzgM5JdbEBlNYyGVqe
P6Bd4B/lakFwmd6lh/pvDhZ+yjceZ8byTyqHxhmRxZ1WKPCvH+uIlh5Jm6fq5wiSvzB4lZLzoJra
CjhrtxNIzVChN8MIZHi3xjSUdIJh8h6QGyJdi3D60cK+Gf3uEmTcdvyDn2Q4j3OjrLNhczR3c4fA
CnJgTp4+3zCtSVDfTEK2rrIAKmTmE7K2/V2CYfMECTrmBD1JFM3UQURdg6kEE2Ab5of3KOQLvaRI
rN+2ShYgEI+Wr6TFdUzll1IC0Z9tgRkLym58M+hbDBgAQ19DEcqwuEokvRo5Jr7oV9Otn2Kgb4li
X3s9bpOsNHYBCOAi8wZya8HtQQPs7Yiu3bvbY/gQhJAS1swSu/5472THDge5UtQq2AbHGhWD3V1r
ZY1TvhXpzaylDpxb27pS0xb6OLK8agSN9WzUNirWo9v/VDC5s1ktNhjyH5W0pO4HKpQd02SRtOGV
EjsMaqX2Z61bz9pt/v8zOuPT46JNQNlsyuMuD1QsG2jGD2QwK74IqZlwUV4lidPbletKqUs3zrWa
fVqgST81mgT49lxfo4ZPB+lljtpB9NYcfk/pBdvCAZBOSPA3JrrMdfuu0PaMMmvfeIhLSp6a5NLQ
WUmK1To2VxxIcyqmR8XM96cqSO8nygXD+2GNAQ4K8zgEqMulwuDpexYNsTnRI83O/Up/23YH3f20
+KvoHG5ho7yN4aZiwROudBXXTA7DeVAKQM9ioK1IealG9Qu4B/vQhT8InJr+E1N33puRSu7NepEN
0VdCn+UfPU6Zqd+dDzuzvb7t3tbz1CuPQrmsX0/Nv0ZReDHcud2zHnQtJpwacMBSlOZcnzpERrPa
ufAWTvujHkzq6g6nLheQ+pPm6sQCYtr9vhziuQwLiP3OKwTXNok8/qDkAFX23I0/cR71QTp4lXut
3lXabXo1dZ8Lb1Jb5y/C1kUmsw3B54DilxJSo15JtYm9xnx5z0OFA7nGw+F50rBugHOy1eO9BB0u
/AoMgK5lSCZzsI8YarrgiQh7ATyw2c3vJWU+sYY9x1L/v0QdhZi5TFd6u+/7IKYkkEgcXwPkjMrK
rdX0qAthUidB8b/NudUCLgxKCsdY18aUjUZeny+0WZ6QuMAo15yglf03Mf0DJele7DJUzp1dCBtQ
OG9sVWnoNZgUYmJ7Vw1paqptSW32WsbI9Ec/0jh0v8CY275T6sjtwb79MG/3OISjHzkGa4B34k9v
ZYqeRVHceVixNA8pjuT3K10M1bNEMaiYwqBsxBJUdeeNKUIYX8bFr52Bo4d8aY9kYkdASYHMCnsv
lfc7I5yNynsK/mFCVg2XJroAMvr44NAxtmifu+SCPb2P6gf1kLV3QVzbi4LS4Cs8/GFCvriP1caP
wngTSUGw3rb0DPUyzWfr/AM1YkhcxQUJGcC21XIMCE+xmKE8a0WKjRoPr3FBF+8QN0qFBGJd8qgk
N83sI7vUDqSAD8hW/tVAlzlP1oIta2LWjKhISJXDhrzp0Mpin1HRL7jEXMxl9+dEp1sJNI/sSJXO
d1DN0tet6Jzl7S/6JPuGAblPgqAKYqtIkRhNLggNPSKWlbUM2ojWXHj+cs3TEqgxytPRzcJOdQYK
WX4mYBDXgH0ktYbQpUkus0Mf9YrqBpD107AFRSvUpHlOhEF5t/KbZETBThJwX23IkKtDFYagfFC0
E7iD47yDIdfz9iGSdcY03g00HAI1EKSLyFbGQZzuci8Vju81q+afn/ed7ABJhEz+ElaVWEWqAsUv
1B6WVfvoLDYzI/h1On1P7cOM7LIFF0SXRCXIJGT8V0gqvo2zO/XlryXNvhu+YLHkQ0fcA1mqGyHY
t0cekcbozDZVQmx/BKcnMCzizXCna2fJrCxZSVPczibY18qACsGoyupPlXGww9EUfcJZywzLH3/y
2KoS/SQC/+Rd3GbwtZY1JnNFNGnvBptsoV11+FMEY0LGgtKOcNvXeVifjgvEAXexGIKGu2iDA0Z+
+2M9ca9/srw4yEoVuWU0hpiLgvZzj9b0QvsXVHbLxbQSfAZzTODWKWzVNXuLWzzsp4Hiu9wF3mND
SrXCeyF1+VOyjDnx2LQseHWZXHc8EvJMQl34Oiiq/vDIJ8bpPkch9h1QHUFseXycDn25o+rXBq+a
RfDGLrUpqixsu7BhVjfqoMAt7rDnl2jJlACru7jqN4Lork/oXLWDj/IGjCnvt+GjNw4nt6JaXB9k
caa7FX9lBCO/shlymHUhe5WPwp9k7K0YwxKELjtG4F8rNybfErtXmvem/GB3AwIkUCzWGPt1EbYx
0k4KvQXRZBN8whw0UedfHMzPec1p3qq2ogckKW75i4A/C/hatJ00W35B2376d2tDRbYIFcODORK5
Nb0fRRSs/ffP2wM8s4zTq+w9HDLQbqGsuiYpEJFG4QACjNFDO6TWKT96k4DTZuNPbT0//Fyazp5u
PaEfnzXBoWO5QUZEoKyz1tHvRD7t8N4qeNQkH09pQoK3R2AxjRVGRq+ftED3yYF5/qEBsrorJyu3
xEc7enr+5b2g0PBTSPhM5RBoahPtttfghEjqJmgE7vltqLqcpSLZEWfTZe/O+QqImKsRsSnP63EB
CT3E+BmiPRm8zpz6Ru1wsp/G3zFudaxEebgzqtLZ0TtGzGWqGKScaY56mGkCegRypicSXHNPPoi1
b4UgeGziH0Ql3Pi4HeO0wGU2hY92IxnEPctPbRDfy2eWpTjXMrM53ANyERrZsNqbmTMtNn4leYS+
aoaMhcgc1AmpJ5XxAupQSBnb2ENFdeQb6NTk6syd22RLHoOX3KVFlvmN6hINdvbQEj31C5jJcswZ
FVyBgk0kKaLZwhbcC6BZHOutbN4dxg8SdWpZ3hi1qHbvDpQA6fBsFT2YY/MLqsEf1M4pq+MphTs6
IB4rnrZlplrmnOi3KYzKNzL/uJwFPwl917lBXYgQV6DfhepbNZcnyUqArCO72ICs4LJFPAffRAIs
+nk4E8rkjtdTvj1gPyo5mBl4AVwvJZn4GjEsXFI7ee95cruQiw0Zf/5kHqy7JRwukDX9OO9oMvXf
6M9pDOFX9Pc43nRfFjoQGEgNVzHto5PxvXhGxMKIo2fZPfgzT+0CZC40yiAa1uvwLf+J55UOiaPe
PAdat+149/6FiglkaDXbIsVlYW31alP9VB5EDiPQLDDshNF9mtfPxAU+Tuwekt+gYoNntBXnL/aF
T2E7hSRId4LjwXQJKUk1NzS7L+fNUzEhpbsW9JwqCcejWRICFGo4Egmb2vnFZ9Uc4RmnKjk4Cbx7
752ra6lLZtJzf4W/sVNFIKrB5maiUM2n0V/sVooSCbsVYdk0H9HF9PWytf7W3vX7TGln/K8F/sga
r9ALeIDNIJ8oB0LNj0xuucQpdn/fdCAjhaExHuaD9/FWFmuSUKcpjBkLzaSFfLhoVRLWOReJ4VnD
5sFv2OiE5nvjOke1ujb34SMnkKw0h31lzIcLFkLmja0cVc9dRjW4TJFIe1RYMZbbgmvoyqRZdbII
d3q7WZ1wa2O+BV9XIHgTmLQq2aprMkSJ6OFkSvMYAAjG2IlYb1CX3Ou24smJpCgj264TWB5JAmb9
4W4z3D93CW0HzmC22TfHJYk7pDSg7N1pkAxjPWxG3PKQhqyi0ymneOkCZkNO1jppiWF/XmhZkTXR
Rg3OkCyCVxCWjIlJKTdv2VJJ2Q+5nhCBuoNhNEsljALmF3c5NlPD/ahF3cZOX466RwXOrY5mOLx+
Gcc9TrPiyy6ZTOYrxLrRG1/7XdUijc3C5+GZHobACDPVmnPHxs7tJHd8zAA/iqk0A5hqAnnY55pr
6VhH9V6ApjK/DEMEBN+IUEQpbSfHO2TtgLkwUZPikUv28PsHoTmpr3/VXSGixK0lmnKBsgqfeu4T
chZGyHjsgHJs3eN+NvhrqV2imJLp8NgbjKEtJgVmdBYH49TT6nm+NHW8CWspQX3i2YXbyPbsjgzI
ceayotPobiGb3WehwnQ/yM/b/i+MC3jsku/C3iWBFYHi0GIzrHFf9jwA6P64MoMQJbvhRNN9dhMs
3WhTtHUYo+skmYV3Dx/y/AwyMiDJX8QHWAsghuSic6XH6ibdlQrp/tmkz7TCTwl+S4GXe5cCUqmC
WN+9pNBZZtQQhlyOjOe+PdxCNV75SpXeZKeF9WueVfpfshU+OXvEJpJveA/H4yYVr9SjV1QlukAZ
qKpbK/NmYQ4pGdcvaHVWX2FCJ45/I5qPJMtx5W9hECLWL3tA5M/E4+Bnt9/mO/anIOENiqMxPsyM
eveuPls0Md0xaMwyQJZmeoYsxgd62+65mN8aMklXCXH64hLsE/4DMIlGk2BhOEJDNL+PVkeRUy3C
XJRhixE8B4QuvPD+9scDQVVZ4sEwE/FRZmAlP+IjVoopf/QkgQq+lCvNFM0Ze2T6uJhnLzynzy4W
yztvjdDU+SaPaJXkyBfPyzyk3RkonONebi9UrBNqqFGkHPefy4kfB/34dcosxNs7cP/xUe0eUG+4
AYjMDm37QViQyapKIfAszhuA5qC+WsoikfXuiLX6UZbbCjyOTOjgZi3L2V+kZAB+XwYnspCeVP9X
N03KSZoF3xsIIb7R4YNctYGOIAX8nOENiDpiblw9Xuw14hqFEO3XwQ4SB8uLeGEIEEEQMVfDULKA
xGNKl6TDLwiqFK4hDZCpEI+43CnDWfCNMQWnfCcPtYVriLxuEFstFUlp4dRBeGtrexytoVHN1BbP
K07BCYmDltNVs+/g5MMXHsbw3VicR5rUxiXBQjXL8xoH1nolpSFetp/ILyjARutN083Mbe2AAhG2
o0Y9HescMT4ZEtRPfVsjb14Fi6GxfpCrZsQzPCTnW06BH7vDsyWkvFS554jUwQfgDVK7n9RFpEFd
9OcxzWwLXnI4SN7tcs0zFA4yhnNZ3tkn5cuFEEa7b+SQjXoI1jbg5c+fTJDhr3s4JihmFuwpPkQf
qlSW4AHjh6L14Xflbnnu6yhaAcExUUjRtnCDJvMNp3UwYv488MazY0u6T9lMUBmVAouSEYWYBpsY
1IgRdJcng7LjSL6uJbFAstDvo3iAzdBBytKxL1jlVdEy+0TES/asR+dv2MHNYgyudb5UCg2Lhry3
m+ZKhVdPViJunC83dl/MBFxiTPduuO8xBW/Jh/xXSsRuYfW9qigvQLng5kj4kq3jN7i40j3tJ2Pe
tmdJcLgBlO2Sz5eZ8gMK0Vpf+NXSqYzPuZ+1xHapLwH6W+9bd5AuhcO+Q0RXYrI0JoffCFjI6ejx
oDz2fKq2s4TZvDZWb3t/tFripaKffwHmYrskCBY1XssRjggOEPD4xWFY0CoCpgMZHi5Ytvl/I8ML
+DM/yfSLkzp6eynBodKJ8MLSrv0HX6TZtEpzD1AJ+47WXnZXcWZfiB4yGbVgnDoOB/UWEr7o/mxo
Uh9yNsCTFS8WHtv8qcfuygEI/fINN3xP5HKpvAgryOWve+a0mwQ1WBCby0QqgDtbKAJSe6iLOjTB
3GEbKJc9v/XWfi6H4uY0k7y0MEAXOCHe72uWsU3fF3oa2Be2cfJVL1fGgCcE21mBxQ053ZzyPzWX
/mIhgWss153o+m/Udi2a+LeEVGP5k5XhJ7dTovVYk1SDV4XqgLagW4TPNi3UyWXBsdYGblxPRlva
LFT7AyrHqFmYyDo0GCRWj4AO2CfQX8gfq9Z1TTmzmfNSo9qgMzckKX+Ql4h0s93AmXE4l8E57Qf9
D4gwRQGTnryOuPYeoKRYWnN2njiR/YG+kCFHyqBsv2Ygn86auRD6ro7bCgcMqzz+ZLcdSY3OKDxn
YGKCOJa9hnrJb4QzvApXVEQalPJMILtA25DeDi2tKKxcaMRSZIGneJNtAevgNZ5daPq3/6Bdisbg
PXeGA6Rlan536ROQkhBE1Gh2WR6zPjAgFPFVEIcgM7wVIHeirpnWKrbyhLhaFHnyKmRlPmW8L/9E
Ms85OmnyQd0/FXk321WQdGGvSklp9OQF5/4AsjcJLdrgtahNr4n0moupfJsGyhkh2l7XltxV0kML
JC9YcUnCpazYbGGRWoMkaK5Gw0KcVqp8RpZAiM5c/o+n9Cn7BK2Upcj4lRaewnBdy8oJxmgkt+sU
9PfrMJJQ7RWXd4cJQA1KoKb66iUYxbioyel3RxDSY12kao83phvHgD1KU0XIbwCJOYOgDIsKhhtK
km3SubxwPp5/9rASt7lCIMirJWxzsPdjc5ktyBnjrs9U+8wfFpRYidg6wvYICcIoUIz2LD8c6DDr
kcLOwE64noB7CnXOb78vu/seSXWkMuh8ljRAAExHE/nryJQ5UxYG56YdwYLmtCmsKqBzIChAp18R
jATPuXRhrQYp19PJftAxV53UVesYHSAW+Fj3Fvx3XTVj1CzEcCRwqwVwoI7RQiTAIB8FNR9kdoCw
1GuNc1tzXPeDAgDm6X2DVrSIkhN+8d+qAYGLqfN9NBWa1qrj716rCTVxcT1ABcZRpUpUNsygYUnq
9u7dwfuWJc6jrRVcBmcBBUTbgOS31BImMKtRD8n3MhjJ3koHYBv6EWwZbp7apVwZE3GLYNPWjMca
BKAkaToGwVcexqSRNpwXrPuHB9ym5Ofh1bvxWPfpzp49HofyTeStCNBXLLaETbvRrcVEflTY2IfW
nycosFn8jHtngo6qA//TUCyDSUQVkcbLaG7UL6zq+c+WF4+sr7aPjcoUC6r8K7Jhsgc+Tn+q7PVD
WQWLu9bflYbFRcTaj4MSAC+AHC5SbhjUvj/dBBT+hccwpRONzHlSiyUiAImdJmEpmdoG22x2Lm1A
6v8kLbxMgwmTxpuO1/nW6Trs9gk1v6t137lR2GysKEN7nHS5xDKsCLZYtDIDUuBza62pWj36Nyds
LFprvtwnuixtPVgq15IxREQXzQC/F0VR/z78GFEuZsTg4asz+lkQRD1yile3QwL+dp8Y8NUhWHEH
E7sofgB5uctUdPX6VuqWHgTrqhunF7ZVQ9tOU4W61nMhq9it+eoBReDCQqkex5IERJqjUrqfmyDD
tHqwed8s4piU5EXs66XAoVa7WPvB6ToqQGFPd3wIO5KMTQm72tKWhxbXpzuqYKItESIMd/bSKREB
RRfPJBzUMKtRoTEiomcMFn23Nwmp6nsjt/oTz8niO4Cdk56KbGrXbIxV4Qe0vxf/5cvPTgm+tRJA
+FJafIEtqMIb2LpBAMHNUqDadhUWr8+4Q4fP6Bg28TeaBZI2iO4pu39kN/3LlYFYtrFm/z5q253a
3ezu32qTVBFnMSMi9FPp25R21U4OE8nHFaA5LWEFNB72cbEGHYdioPUxEPZPXoF/drdQ2HjdatNF
HiGpSkvYjfnaS5duHTkSovyzhBb0RPdoMXmgY7aS0hB3tjzcBS7IPYYYyn7W+bzgPLPSBVpq8ZX3
vr9n4SqETx9QmFORc8f6pZTTGWmU6DRhRKBcR1GrJJf5h/pquSra85wYwQCB6l7ik8FUqEGNj5De
zcoZ80TaXYjZSL1WO09VPOSKR2cG629Yc6B3q7Bj+zH8R0qhZPu9MyM6eSvGdqA98/x7/sQKS5Wr
U0/egrXd97UFKpvnn3zaHXFGyIGQXDymdGqdg0vZ3mf/rQIII8b/RtBVBYA4kRhDflmaI1UaJEJr
W5D7QgCVeiAGsKrwWaV0YUbSfoysBu6xrt8xaXAwBJGlCPods7ILnXnUXjsAYy9l0vKFEZykGrzS
QE4yqqEkaYpIxFFMLssZGD6O/G5N/MBqrsobdo7qVHQyu/FX2cAaRNM5dW57LdVymBOcVC/kLv2z
uuvlSZx95eV6myetmt8mNXfjta04GzDwbqPKmyppO+Ut4LOOG3eaa6Vgm6MpHezm1z30zFVZpl8i
fb61oRluSRmsdVC0MU5eppm4BPWesg1E1ny+U/faP3StNiPICFyaYfa/xK2av1sD/TIa10ppNGCz
QR8gro/jIVOwR0WQXodYqgPZzsqMuL/Xz2k1Tl326X55WxrDMRZGL8irrbO3K1oQaTpBCX1nHDa9
ByTYsqTslcjTFhoO1Ttrynpd082D1qfm45iohAJP9gF533oEHB+5sxY7a22GiC11q0Wtoo3AJ3jD
8TQuz9ylVsRcSGw2b0pVXzsoz9NUeQ/4rm+2YzjJAff9e+yzz2eQ99Gf97gn5VdhEjc0d2ygAjWh
XuRvl5jfMRZ50dZKumdhq1hdTXCZ3XHtKNL4+TpAaMn3Rfb+YxNziAWntZu3jQW3mCe7g7toaX2N
/SNk7nFJHBTL/7QjnSXVoegEp4A/4HbiyT4jtYe8hW9lbmYSCP/UFRNC7zdJa04w1wpRweBIEKL7
CYNMRW6VfjyfyL95C2GL6WseQpbEmUU73wVIabNosuPOI0t+H4bgXQtpsjKKjhBaiQlJQxuUrfgY
SjF78YDe9C2o2dK+Z5eqOH4YGGT52Pbs/qv5EArBNxWMWFCM54UOQkK+hdMUOOXDI0TVlZjW04sl
WoI7pHB3ruFwKo0kfCaZbzufNSGGl1wdYnvkLlA9+47impqEnPje3W08FNHI8DvOZFQdmGEYtIKD
TJ+2iyYGfrgqJWMD6fMVEPHuK5PJCErrSuVTLZUMAe1GcRd+JThlk5zWY9tsHoOkNxMwRH/JPF38
/+96YJ7t2th/wGOSQvfkrGlHznSRVQGLZGN+2tksD3EKjRWV4iZNGPAlLgfbY0APhT2qLc8sVlbT
ce8OOJlXKEc4v1DuNsDiyA6DCFoMIGjeF7QccjLAVakP3savIBXDdqhbbIBentRfTlLwYPfaYfwy
L7G3lW8jDwqyawNcrHRtVVPktZDPNK9YZCXRtdPrZ4mGcLY9PobailPq975s1NtTt3XFujOxgM9q
77qbCLC5RNAuUfLoPvIpKCkmnCKqaNQh1jxggRbmk20rT1zSspRM2TX3VOXthVsnxyUdI6NNINnL
4qWr+eMH0OgQGAjUrgKCtuzII8R5pBiQ3lKNLuaGhh9ZTxmpSjHuiT+UJ5pJHz+uNLENIVJAEutk
IEvS7kZjko316qY+ZHkpB5/M65RivHvSB4egZFNvrpsaOJDJuL7EWd4aI9aMlL4UUC6rQMRTCwmG
66jaQo3ST2VonRapzqOl0CJDJRRALe+Ulbll7ZsHyv1mDLmlPCrLDI+67nfx5w4URh//jwE9LDoR
VHQEFloflFtrjIs1OhfHfqudir42haGUN29BMPx8T0CrWkB6eDp2FfFxiOGIWE9Y5349eF3h3fCH
d7TwzBH3wVkQrwM5kMcn62d+uiXE0TB5BSojbM7p6rSR93NF600ROF1isNNiZd+1fzvcf4AuFGMt
JZ6A3bfmhl4p9JDKA1nWaYjx1k5tjCRtG0Az/Ir7uYoTRxAP/sOxhGNE+Vi7x2NGjElutgttrj0U
1+Rj8PR7x3WSn0YXx7Z3+Yp+btunVmJa4GSWNozglklPCPlef0SKhlWj/ZhmxFfHjzEZoZPTPhA+
bRJaZAaMDDR/PJ3uUqNAcu3hY0UFw2Pe1vznUlXca5LlnrkfGNwDEiykJlitqhpsg/7LqizNCUfp
6gew1JKXDf6/9YBLbrz34w3rH04fUNNfatqFVofGQyPJSrHh/aVuMlPsyyJcQpIOkuVF8sqZUDhC
ABUP98EEotLmK77mEtjVWvVW9DB56KxA8Our0q9KXM9TS92Wayfxxn79p7fxH0K+qOV/+wnOWVvg
DwA8EQGrSCl+hK42MSZTnRVWO6PUdcQn7iDYNewQNGZ/P85bP600N4IFX66nWwE/+E3bXqgkqbzq
pnW/xmcTvmW70EOhtnQ2oqQyQhh3XdLjG2SxQC9dZRFQBIhG3ITzBiCAqsYCxxrMqxKY3/1XMACH
ViqdtxUBpm4ryEfAdmZdLsLIamfAVtiJB629Eq4XSVQJFWBIUXOMz7nbCY/RN/CcLSInOLoq48Su
cvH5ZS+uRx0tUw248VzWNdtbNdfi5B9VXUCgcaUiWyGLlsq9DybDURFFGQ+1FTyehWJZ1ewWitGF
EXJ5ZUDLIYWs8+GHFwjrIJuaB9jD/Nr3ua9yjHEAcJ/X88LP18yZk2UeSEAunb8D1GhqBRfidKqH
K+KqAxhMf35HSdaJD7TiD3q213gPF/KG23nuQJJ2BDEXQ0qTtwQSVwj2jFpAqa2G8/aVjEtMueRA
6QNq6UgYrfd3j0qzmtTsbAnfbpM+Fs/qcbv/Z3iTBCinO5uD1Zb7EhoCJr59pOwCknWEmq3GAjeM
WHUD1S2i3xcomEv+hX8qkuU0303COdYGIX0pZZCp2txsKsOQq3KblT88TQaQvKNa0188ZGMGZ0wY
Crs8F/HIGCcJM1YEpE5k5DaOd08V5q2UHvF8z0bWnt2jViM1YlOT0V6JoaM+HCw4ItTHvQOduHBa
R0dUPdD8e3WLoJoWamrkTXxfP9d1KW4kKWx9/NGK5JeyHDquS0e6kgwMjP71kjTwAo5SDKWa7iVA
1cw2wyn3v0N3mPXh/2cvaJNA9ZgoHB30eQiGwawzsgr8h7VONcn7R5yWRBWBEhJLuvnnVOtC4sWC
0iN4Ti3bLF4Kyz7K4QGteiwPdh8TWbUMXU6Jhw2O9WgfjYkoaOyw+iHtIWye+FwsZK9XaUYkL/rD
VGZ8ckgY3Dyfq/osv6ZvFcDW1h0ps2qedbG4qfnhW5ZNnGmVUeIk3NdLIea6TTfGRHVF45m7QqLC
g9jkmuGw7HvBZ3e6lUaesXZXnXP2xIyxEN0aFlZHTJhY6GjblFhT/23CdEA5eFpfV4wDqNBRjv37
hGztcCoLyAOnFbBBR95x6V3cU0jlbs5oB7UmUI57Chx7rmjxJzVAngPQARWVNefSoe/g9i73ogLG
WZLco1EvjffMrX/yDx9cAr/VG/xbVWNz2HQXy2Zr7gmHyq+fgcDxApb9HtLcXjPzzIsXLTtKH+xY
hV92CMlVrihGoBjl5fLbVhMyXFsLXiY5WmM8nVTPBhV7Q3xHheZVOAna1tVyg90lGkBP+/HIVMl9
+Z8GSorCr7Ycp1YcTVTWlLfMkAm3fhIEzH9dbkccmdzggNIVP6KoynMJZWbCFH8JXZ7wrJNexjnN
TP3T31ISmXCVASKQCFQ07twlUkz4BqkElZ7DY0dYWr4Ge3PvIgffiKCauP00sKHzsEDo6PfKHbs/
3/yVByLV1EYsMM5Dt80Jj7lULJpQ5+SIArepaU4do/0w6YfFc7BCXRjHhhHZkDiMYaQK+wh+AZ/5
a6lTjTD879u/E3XQFMaAOPdb1WI3lOo/fmwua6uJwORMlhRn1ZPELawtaxMBF9arR9daQh4lnsbA
8I3Ygb9baaxC4evYyWDLW2gpbKDl4Rhdj/6LCBLDT2k+JITdMXNy/Oz58rsJcsapos2MFP2627H0
b+Rz2WcSS9UdDlgDNH8Zp+lUojO/2ADmJjrjLaQx3Ys1cB6G3JSjRWs+aMgdLkM8Zk/kxQd97qVv
YHHgSH4T5W/tVYM2OGW/fcGEzCKlO1tqTCboozGwKTXxghWqgap8JpOj57pz6YPYOmGAL+mh8tHk
81PSpDeWvVKVlrbfxTMhK3DqCcn/Bi2bo8/KpG4L+yydRzF7wyMWSdEb0CsYqVNuwCklCCiV2PrC
+3TwRfP9GMHHJ4fCaSJgu536ENzYmOL7r8v0x5wDQNL2X3wr3uOqI/HWzD3VPU4V32mw5oEgHUUg
iTCgLiazUh0J01dGbdRk063hcQqEy7Bklr+b6EQ1QDkc2RsVThr57t339vQn90k9tnRmlTQHcwAi
7gE6wZSBlh9exEh9tJjtiocGSNV0yR0mMkgg4Qmpx8IHFvjEu/2TIuDKEr6d4znoHKaJA1bGDWbB
2NfeBUPHQE77vYlyOPvSYZlraixYsxj5SE3OZWw6WXmpwhNBppHK96wQuJTki+C4TWkysSeBa2/t
mmXdO/wou9VV6lgK28BKXvm6T0jodyZ/0iDm77mNh4rgPyL4xqka/sxBbrybo8hdPayc1ChYl7n0
EVfHmWiPbyyhXg0CwoMmmvXb1y3iu+MQXIBy5HWZ0quk1GqQg47Q/h9b2fjRPKDSAhDOTeMLyqbs
V2kgjB6M1pODTO6XMKGtDxfmIaT5SjSDz8JWoLgJ+Z3OfwqwVD8yBGasZO+ex1JIChNU8o0CY09U
OTwCnpxaPsUkcp1vR9i4Tns+LAk3ugFoiZ4N5J6lTW4HAj3ul8+r5SWtiFoCBO9zGjSFTUnuOtfu
ih0Q7+EXlDdNkhK85OWUz2OsRuwwG3roKEXKeNfVrr2FkVXS80aYB7lL89NJhXIGgaXP/rslheKb
Dpn9RyYf1n/kR1KzfyisvOxtjLPJR+rYbefuNQ3lk0t4Vjd+mqC8qAnt68BFglPVO/UcewPHgzCH
2QWVh6grPdX4XojNT05IpY1a+QmKmqFTIZMbHYxn3OwT/Q+JMfVUyzgNKLpTn8TJMf8pz85HAvp0
z4txKtGtDzDPsOIHrrLUMeE0TQ8xk4rgsg1IQf3i6N6ZVF0HQKTKj+qupR6v5BFBNmoQLaBfyIXu
7uB1dAEcRmXgWs2wdnq/fwnS7VseIrW4WUO+n1GsvrP+KAm5j2uHLRdxDXvyJT9iGDF+QUrLfkLR
R0OxNHnvs3zUxEgKBdBAhsQhOxEE2VF0vnRXRo4Gs+kEJNtI7TRH9LqubwC7lryi9AwHNT3KqYhB
FvOGRM8XvenEEOItpSI95MUJnh0pW4AmoOw92FQvfAq5idoFXNg51tNtk9t+F6Q/21nRVajk8YV1
VJag1UV+K65B6AzjRZTPQoRR0/aWCv/QxQFbqsw1D9QQKlOsIWHVpqIvF8oEKMgO/SJtjeIazYVU
LUNgCM93nJ2qK/bH4m0GgC2nxeZUfkQwGWqICEuvy7pprQawJUnibyfonWElZPATAJRoQBr1CTSQ
lFkwFWEFJh2hV9V2yGHZc8/AjsqxuF/uEc8UWkIqrFweSJLu05YS9cr3e+K6zNC8MTzxun9Suhbj
GOCUPQpyHZ9c3ToaVekyakbye2A874Q7zCqqayIqKZFrC4LtrXBhXBqApFETVl9ovIr3lBzloi43
ip+Z2+wdJvlx9cd/BdECOydoB4iPukVnDbsW2b9HzB6w10TFxKq5iYPUKo65WPo3QFFAxKD2YO94
ZrYFbHDioyvHtOK/IP7dUeWDuElnfZAVj2+7vaa4al1omUDlD6SeW8iveYBTREv8ShOEZn400oWP
m0/KtxVuVnHwbOqTDFQ69z2Jz6FQlyQ5uhbVbqAdez58ZO+MaxEk4tbPnBjgaiE3fKfnZay8Xvpc
9ePjerqkSjAEa5ihzqiMQw74Wh5sfjz+AH4mlhIdEWufXrbW/e13mAusSGTWH/v5R/LaQi/SR65q
q2dMzyh89vks29EprrCw4MIWdDjObLsZw3A7pMwb0hE3q7M951WpZcW6UFv7KwDbXF9Rj4BSjbo9
QXc2ctbpKednL3a/iPQqSNdz7b9J32QHv9eaAcTjhmgmR/KPBefhcHIQ0sHnXuD2W17snBoUaCBH
wlDTwb4TayARairwh9/Ajd0yesmnSNSWe4MnSBELA8qLjdK6LojUnTRnDo6UtKKPbQIQHQ7SUMTQ
1s14Y4OzKfc0bTSn1Dziq5L0fb5cLayDMHDuwnpbGXHfucRL136FBQbUnXb06q28XdBBEcB5jl6w
/zRymrXlKUIUFGNOpe9GcaQljHZuMI2YOi/359MGfPlnvn04G8uogszlXAe6AQb7XmWijGrZinq3
+ZwNy+uiwWCQtsUT4HAVvBa0y2gtnnIfI5HedWTFOMI/3Y7cedwLKU3WB9SdF9VyVB/gw6HV6xN3
HE5N/klaavJoUXZySHsmONDpAktYoguy//Nf3vaeIof14dz0iea590BLKMBPsxqRWzTUWTwYMXQj
pCtLhxv3KvUkfCJ+e/u9SWmJQBe010BSwR5WYPJsWcKHp1orPfjrNg+KayZcr0fv1VUktHOBDmzy
5DIaF9k4tP8UM64P4+Ys97G94LgtrPIEW6YGV8K1lUmrBjpikc3BAO7KpuNIXWN0dbEGABCkIFNW
ZKlPCuNAqEqbfZEZOFk3f0ONnX7ziWMC+1SDEFTyEC30vEXbyeqpm8Y9yJGe+dlbnv4stDL94Fxk
u6FnOq+iso65ECAxDIr8rHvqlMigH2TVbdrRBzv0NVyefgeVOwc5xrlHaGr9A7f0WyArWLSFSgSc
LPdqtnbPWoemgh7/KQzKYcGGDfZjsWf37WFhKiyc4VYHV1yVgFdSb5CCcxkJjkpAZTi8rAgVBEx8
IYIgojPKo3BTmp642fJssBz1jg6beqIZkRsxiw3GNUgyeJUzxns86El36zMDUKsFH/zlb0v8Brxr
juYhlVWy60X2v6e1kUwBSvW8Q/WFIlkGXE5UGGmVknkVj/tQdZdjN+UOlOWB72dsOa3Trv6RJ7Ns
YALpq4X47Zg9FOvE5KWMciIw97C9xxGHcZ1A+4vR8GfMi00G4NAJdcuCVX+ihiEHxBu2sX002U8t
mOPbvODuNGU5YQqVk18eeusQq1JhzPgOiHVx6yuycpixq58hM5DIa5nPkKTbcmLmnZsPcCt/niUN
0+qW6NpoahM4C6LyvAhq/bP61z5yj0UE3dMQaLIHNN5Rd96xx+ylAJ0gKFrVLjDosLS+t8gXlTJz
3IyP81RkrNgVp0p5AlTxuYDLWoPfuNOW71CEn8bHlM7LwPhj25pL3NyAZTCfAD9mkd9A8ofJp908
glii8EI1KhN+nTkNVjYcCXzqKJ2tF4WWrfsyRakyvg7VgCMZifdkhwDdRwVhPXU64WAqyEPgJuuE
sm0yRZlnVTqbmsbo2TEDOi2SimjDF/o9xjK5kl9EIC/kRqkVIFXpaItsWvCJUVTycPBrEFU56mr5
pnp8UJHxWU5QycQHKOxTNTUD913yJOK0r05ueh9Wr5sotho1Rnodxzk5tnYfOijz05V1641yH6YU
5DpFDKqe43jmXpe3Fj1DFWczZYDWTZ4ebBT2cDf9ASJVz5G4txeQ4uroX585mc8MHTPdGQdQMU54
+VKKzL2ngM0VOpO6NWYiqMaZ4L2qFU36DakqKVj662mdlj77sji1iyPJOXv41bvigDvzcAv8h01z
LzSh0rQzq7UV8t+mUdBh6ehcupSInO1punQnmWxV43XIasodKTgDxRhQew6Gqf8FPfg6O+tNcr7k
ECxHxJ2DPyWr8IbftUrAArXyAUqMkwfW8L09d9dW7fpou2UclHZlPEA8x8emzcxbiZi4RUrBUlkS
7dVRvtoCHGOoTsw0OBKSl6IQu7YGwWvLK9MuNf9v5hy0Yyfy+qJ0Gj7oIL5cRbYMLv3gEL3F9Q+W
AJ7rgvb2uAtVgNd8Y9zpuEDsknQImguTxyzIf7TW1u0XNJ0GCZu0+412uM8DVh1t9nVhnjX8JNjF
aZxQ+qqOETzh3ZIHToACil8qZM13ERkHfoch6700UJxowCtRWWa0GdSb+1Se1IdVaAioF4xCSBz1
Dar+PjoXUyXbXIWPcLcJ2NY+yn2mApymm28foAF0LiGbIdNF+J0jurFhv/6DCeWigiGaXwVINWsI
JDdDwitR3Krx3fPEajXAsDhnjWhI6lZl2z7oK8ZYhZ958CAeBeD3SXPlTeuhAE0wBr9tFs9spusb
zaODGjpvJvL11LW8Z32iRv2YkaaH8SJioi7ZpOhtRZwfKN+itD1iFQJFlHlXVo2L6lPLykD51rNG
Rea4MR5nO6O1MELCfXQ6i4CD28LaxCEPREARMZs22ZoFdW7mWtq3d9XNTbTg8+zRVYezMdmhs9Wf
e/nu9/+VfRqHioKuAED4YazxJzBkcuBCLxr+eBsjQx760/VOu78rr3/qRry23R7xJr0GDjie5xHv
E4JcmQUlCM0X1BALQxp+jclyJCxeO8wb02EOc2lIqfp43s/X9cD9R9wWRGk9xRUDWGnQbUkeYsEY
/sbhCQ7j6o9Wi1eXJw+1Sd0hH37rd5ZuD+J4p+xim8MNJ3ymAkxCgO0GtRekhSclelVSQqeSKskt
OxtXrcYtsTpvSfi73R0kJ2XoA3riBQnlIocMve33LkAZ0rCrAPSFVkJCROCdZalv0N1nXfy0bDNO
rmJ8p0tx7DGRNMSlruVMI7EsLvDPJgxyEfjg1pcsHR7JFU7L3PJbh5EzUrQGfANS/L4nv8lDkZ66
gQJuAw2chs2I1jxAi+u5l+benOIF1LIEOoURaJoKtQY542rU094MR2ewWA+KrTrB/OZkWV1mrXZp
4K+U+8d+IfYgWy0UpQSDOvD2RgYHms1kQW6utquMMk6r4JJ0GRrjqDh2dHZro7SfgH0PWSBu3Dqk
YYobPjyUMgqNeBPrmLs6L0QgBHzNdoz8Lrb+P/5keDp4WkN7MoTu/Y78LfjLayGhWPNHVz5m7fXs
yFD0cUdGubwFcnp7I4ULwYjvIAUjV6Qe7vsh0i5Tu/2v7hQd+ZzLKYOHAd2Yp3wv49l6xiXrCK69
nDzMEpewwZHCG6JIbDvtVyQXUrOVagxZvSuUzgHaymbuh2gcnpVFGovY2ncjf5LQ3pdDIkfo6nyK
5c4/xaDXvfnwdzsFxnWi+7crLPMvQl3EtWI+Bs3O7NwjWwmb0IDlXINlbgY27H4R9LUu3a+K3dGX
pBnCxT2GRjbIT9cJA/r0Rhpw2THZhRl0US3K2X+fBovRG76a6xE/EABc3YQC0h+q4HlJfTcXZCcF
FMTCKz+n6037qBbIjycFfEG8XDpd48qEJK7cYAUC2cN9qsV1yfpUooHtmcumFq50wgEdMKC/m+VE
NCV0kQYvBwxoVSdzOw4sVm6GXPqQtqRpgHuUCPo6nBWhaOK4tyorIhcF8ZU+IbPTEPuxWLBd7rLw
0N2T2pxDHIgb//FrTttG4gByQMZFrzrJx3TuhEhXc1QeHV31K3uq+qxfaCs9MulBfSCJ5u3W0gLg
hlYgkAPBMaEXQey/+FbJ11GHFj2kdwJIMCW/Im+WEYnmvfDX2GHSNDbMDCjGYhZr2QF7KtFpENq5
zXBXIUL9vb2hDxanTlrQpSNflzy26mdpn93T4LSGIldw1n7ymrlz0i55Gg8rDY4U6z6qM7ZU3VKb
k32ve8D3czwmMEgg5kbdxn8VbdsUkn7xBc0Zy58BWmk0Gb9IaqX28rkSoI7PxVlPTDG9jZ/Yjwb5
pv9wGU4mZzK5Oo3lcJXJnhBYWRRB/5f5+D2wthCHioD84JnprOSL/YDU2CDlZNohOeMCKqiUEzbT
ZfNJtN5QTvcKwGa0DJVasp22BNJwLXlJ96W2Y4SjtIA9R6SVwCr5zsGgEgU8ieSw+7i1cGnUMqj3
8zPHHj6iaKjYaQNLAvRfpja3Sd6NvD1qgjNcBmmGM9xIHLsAxI67/TErnXrkdHReyC5r/KxW+/dH
NSGaC1Is0Eb7Y7bJD8pxRiXwOcWmGjuT/tin8UdQ+jVOJaPFCUuCwaOYbj9ESakITNTOcXX0mtEe
L/rUZHag+jE80s1iGDnUP9VRIceOUeFTvp8MHclZurtFsjbdOomaYHiWMZKerDEeC5xJIaa9x2RV
AWyzPVyqRJCn/I+/N2YJsqEQLOx8yXmpVb9uJTlbH26F/ld5TA8Twuhq9AySmaYyrNLScR/KMG5C
HNEfvDmvOuCwlEj2E8DhjCpzTKBXzxTahowhlphYM9HvqkpNOVVxml3ggJBhT/gzpNEXoe5duKD1
49zwk0nvIhm1LHeJXFpDDSnKzJkmKT8/aY8ARViQ9wcx5vZX+Jy4jqO0go+AQZCPQ/FYhUw3g/y+
Kf44BBMfczSba9QZzQABu+HLuzoA71tAYISxhq7KYTBh7ON8V+4NetVpYFfBCJ7lXXLW7eE/Krsf
7oyK6VrY0Qhm6SB07jk7lGI9CR0UNijWxhjwVNZh1nIMwons3RBYuZH08bubIJtAJ441xL5d4TLp
7RX5qAbpgVPBBXnlz6hSIyro6F3vD4XEWjvOHKcXmuwSSRZOphWc8dULutZRaFcS4mrGSH221vnb
YA3R3vEf4tFJWvEkKG1NNlmnNaPLx2i/6i9pJuD9vd8eaZFCly339v4gCMO/V9EU9ogGh7s6t8gT
RzjKS5i1dDO12XuUn8LgKRRXb6Jkhch0eOORL7iajTTuhz5qwZSRzA0VZpFRRmbLAz3s6b4eIaGH
eJ3/S3459pnBW/XN2YxFj3msV1kqwNmt0QX+mbkoscY5tGtX67ZiQXmqv3k+r+hEjSuCBmhNAQvS
ufeLG0DEu5MKFY3p95YVGPA1RANoipw2T3UoyQ8GhYz2kgXo1iIKZ7koS4cfkgf5ThdBST2/Ujof
INaV3WZYVp6b1ZjQ//NYmaDZLjdw4TkhSf57h1MEpnIil/3vG6eiccaL2eACJ8MwQRHqMOg9i3Lz
YlHu1Je76Uj1+5dtnl8bFdrS4fRgi01Q6qG98TDH7QQ8rC47zkUub0r1z7UbEBrj5iOqWbP7kvMc
VAODYzejYasZUXfWrCSp3JxgKLWzoe0ticnolcjHyk17nGyPtBHX2n9lAwRrEbN8KfV4FNta4jiS
WhWdc0VIVODdyjFfMW1BmAyR7MhM/s4SqIYltbjXUscs2ZzrVCE+UF3UIOi/1yiYYJBuYx6W9+Cq
R3QFoykitwmZy73z+OAdaMqupj0i0/7Jbaw55eQRSx8aHN/Dr5c/gO1zZW7/W78680mppDgDxQqE
9QVsNltOc2bI29pI6Tl6P+qlXv13h0Addf8nyn6t243+24A4bYzy6ODIfMq/PoTEwN/ruKlbUeNU
nkO0bjwyF83DWrXYbvlJZYZhEYD9RciGC2OJ7SgoOU7zViJU1o9413oRGq13idS6ZMW/xwFlxtd5
lEvxei4sRlYZKLaLwUO3/r33gNQ0m+Ia8lpPn5WCgYH4p2aqhB56+AP7uIxXCxM4TSM7T32uQbTO
LkFZxSFhwTHyc7es8DytIqDHGV1MHn9GTgOXcBlbuG/1ypenifS7+6Ua3twY3G/KH+hIyLOfxUwT
wa8f18+RPO8YE/rp/0YekNaXo7Un3x0axnFeQ0GzD/LXjVks5lUElnL+opk8/0kg4uYHmHi1HsLT
r733+SIIKklPNWeP6vARHNPohugJVg7jwSKRx00Q13bugjdcdO9uQ9xDNkMQGOUU8XpXKO1xiZVO
kvp6z2Zcew3XSSDtFXu5gZKk0D3EFtmbQ+PstUiwBP8pO3rroiS4pGEpjLlwpFOJxneLq4KjRrWG
fvvo+C0ub+2yXxpuCQkTlcbK0HQoHPjoPYtnwgA7sXUI+D7dJ4VkT9+BM+4nVJuc/gp2ooU6kwAh
qQfbv4/r1kq1o8McurvlvWAiBwz54k/zGmqbKAi2L/8zXkvXKj5GVp2y953ynu24LLjn2w23p2LB
sCorrmHfNe40g2Lm+z0IKxwAt7LGlfsxKIZ9HI+sBcqq7h7E6XgF3ykbtohGKnFVoM5vy1auTFSP
NY3QeYsxUR3B0g4WIDO47Pq3MQ+qWPkdvxgrZCJpJPUmwYPmm4B9PFBHUUzwdZW3VoRyT9qeUMHJ
12eLrrjWjyLO9xNkcr1PZ7rwYV/0v0XMHOi2Y8CKgvyR0Bnke9A1wA44PxTNNE1en6gE2xe9XIvG
wGD9z0XGRqDbDy1TcYtFHqiYdq2R9wStMDk67FqPrr+DUTeHFSOk0SycTSPVLDZKO21qN4wS6vMe
FzAaMFZNMtWUWcLqxigYh1u7ZjYdjd2Dw11HI3BSadzgBV69idKH1rPXl2Q3Q4IBIHAppSJOCdwO
11I0F9lq3rqoNRz7mOLklSZ28iSvjKPqMGSQL3XT2tSDN2BMySsoJjNDQKttuSwB3f2NJDCH54m1
I1Xmg5QExxqoHlP04DUfvU1WmYLmrKNc0Zf4zpF29KpeRl58bthOCynssOLabDqgcSOelR15KAXy
mXRrrpt5CZTX5McaK1RS+zHhL4QF+vsttnT70VtN8TUNRk5DiYzo2bkVPUffcK+hrq3uc/1PoZeg
tL+3fjaHA+0Fyb8kB3+Xsx7Y5S/TIZvrKucXwl/tYtj0kDC5xDdTAT5yGTPGb7VG/9cGHvWMq7Bo
jGryMpmIyVaUFwkjKwpiBBA0cDVEtWOeOxUiQsj/QAh7RUNyaSTQOG9/thzsC3UFfUannxgkCTjM
FceSYnkfTV4lMHDdAUf+0zvafFKGWjljJ2Bnv7FADI1uvVPyphC6NsHxRhAE9jODJg2l/B7GbNGH
YNoL06ctweMvVhMvN9zmrabBa6bjhB2aznfmQUPxFgHNr90dhFKU/p12hDEhNrRE9i3DGGPKlxgN
QGGNWLD8OXpMsDFX2TTPMVbNnLCj4DV2w0zJbfb3QBs8v5S7HqQ7j67cceR2e7YBGEQb0PVHm4ZB
EhlVkVdi8d4l9fDC1q3QNISqh4Lhfth/YQN0h7Uo3hnzsC7qOiKVxtC0gnoHMF1RYgCERLJzQ8BX
SPj4QqVBUeebEvP1WasmfmwhbPifttuM2jdHFxlhRTNthlqjhgVaRYelQQjKBjVuEBw2s5lpwQ34
a28GbgIHoRIxbyvObOEigb25Ck+2CFy9W2cNDOxl1kY/06aA81TnaJcY9R/ooI+6xG6r2z+hsXMO
UMxpDUftxOGMi+W63EZygevcVQzHCDPrTWsOYt3hLUkiKnbfgAAc4SYXeaagntqQUVgmLc52galY
ZpXHLH+suA8sP3o2ct8MstVaPIzXU/++Jk6RklVTD0bwiQb6N7t5q7Kzg6U4j54xUwjxNlg7r9lB
5y0gx+e5UJmfHL6sswchx02ImQPunW0YCJ9ww2F1Q4HhA9w+NeiAHUlM2aHjeKryr28eeyv8lhH9
AoqwvaD1TF6lo5LT7PKej6bkF5jKijpzssF6VbPKxag4vuNkVTGa00gJzArG+nEG+5IE20kmqEWE
HZCG0+x/FLkd76yboWTyWeYAoL0sYwB0nSb/nL1OWWODqV1NGtAxlYJT3RdJzyYiVKrhlRz9BZx9
/PhwxIa0NL310ajfbReoTquUxvZ3scx2Esa0j8z59aR6x8vhLSYHTHbSzu3C1JpdNkTPjpbiBEjy
ZVWltvGwuJ8EmmoHmMSCIz5R+muFaW7JCIAjvzJ7KQv5V7xKeHOf8x6l444Ib2cnN2vjGSFHPqaw
7gORRnXZqNJBROrobAWP2wh9n8JkFoXBHKNB7B2yydWpF2WW6i3sBhsqQqpx/asvaZgvQ1w6KQIF
YFacmzvStplTCEfmiZ43QlsFF7T5pNYeQDXpTISxjs3RU3/ofGUQzoGzB9il2kYQtHitKL5YV2Uj
9QN4FleWq2iu07TfPr3K6+F/YKIdYy38cWPnnUNgmOe09HhDLJRoGIsFQoQvgF9+MzKbYeILzHY7
Wg0c/Z6oAUdORe1CsgahHnw7sFQuj/VjSOCX7VTp523Ffi6YeTfJr22KVLTSuhbkxOLXi6TOhe1o
5UlTw2g3oW44AIOBLM877RqqWt7S2umOT+xLkBhBTWd7SKVx5puhIAWI6hZ+xNZ7NGz7c6mFZL6A
ti7HV5R1FxWWOvIv2r4lC2BJDaicVzeiiSQXiWh1+H/qYv6KOTxZxpZwwfViR2V5yxAWqbDK6lax
uv8+j9c+/91QVWhR7bLdM0ycFKY21I/HuB3fuxGs+Dtjm22uwRXiA/KxiIzzn0IlF2F85RvDJJ9G
gON+rIIXSg9eMjLVg+ulis9td8Z8ZpRVdpAiKKUDKWkx/7lToDs5vU00AKlteyqYGhib3Z48Qn7A
Lq3ptt74CRawR+o0rc0rS/8oUwenp8JKdxhRAREnKR/6zBEaUH21c9fuyDZui+BhGaaTc3BHuK3V
9Bn2qH+M/sT5hITM3UzuLwO+NRsUGFOJM+JusVI9Cep717LtuG1HV06jia7VgiirGqEg6vbTVOt+
HAsxGmzJUlV7Bww4oN0KQejLG3DnQWtyZvekFnRD/QgpCpYyRqKdm+lML86t4fa2MsqROtVEO1Aa
d6Qu7sLKHoY2Q8tqoKol6U4r+C+I2+mC3EPHFTgcltfZGpogFZ7PhOvX0GY+7zqKwpK2ThjWyk80
v5gOgH88vxv8KaKAk5jmGJ7K2ZzRpl0TIqJ9n56mYtBLIX9uVkqxX6lK9MJOmUWT5NoCmycHz0E5
0e47yAOhpdLh/BSFj1owKKHGRtpB8NZ5sgAFsztvxfSl6FENgh+eoClJMnZAG7zjoRJmJUUdgTqS
qdWaK7/gZWxuXNZNZ/mz+6MT5gUllfjJggW/fXtYTz5Df2V+TgtWl98XgbQxaEc7iaxxJsEHRfBC
+NiqRd0LJExfNkEImIrE82C7hV9eYzLd8jnWMD2qRghxhnNMxHEV5rWbiE0vFM9ZX/2aBbkbgiqj
FNF3d3FUkZMVJmptandIZPSQBwQzgMmpEUARIsivpdjmm+0bFAjqa6Kdw8DYLai0/jeESMy7LfhV
0f88cnbUtsD27WZp7oB3QnYn/+uzqPltAgAhXECm3315ajGIfH2tzx69RUIZdHlpIDTk+DRe9Ok5
x6/drOrfYCh443fG9ozP/u183mtKq/sXYY3rPttVoscpQbFsOqum3Qa4ctBmq2lwVBMNqsMTMrCr
OKW1OghIPTg/JFOGGCgHdN2YYbvuOjEHWEWMmGHca9Up65Sjj/8gNlmG2fOwWb3u/hFnZGBcIMYc
Y95wl2mRyCZFd9iAIRTSUhoiJf2RieZk1UX5JR0+XfmfAu6MeKTHHJf69/uDeuQecTrKQG92K2RG
4TpwcO6eBfm4WImsc8cYXbwj6/6357sZHZ7P+VwvUEln3GoqSsXDp494XerPjyO2G2zNSlr8+/aC
z8G55aO+bbU9uPre7E3Fy+3vg/xNmv+YlbIKNxFb+XTh2ntOlJA/xNM65yPr9IekL85hYNHVX297
DpkNg402afIK/YCj2UV+uNXDj7Px4u2DLwUHRcgtbFfVK1cw1fybmTmKpjj6ieGbav3kFlBiNGfu
foiFjRI8Ab+Ry80PtOdtAH1tE3vsCHJ/LxDBvjwHmeUTQzNdRnNeRGwHN/dT0vzELWfF7nZYqdbo
gfwhxD8Xvzb6F2P34Zmgpl0yilbQGqLo6ztTgN46Bsy5YT3S7SV4WpcDlYvWfz99AG/cZPgAEEUL
VNgp2ai5yyVKXCVCxpbsxft0vMWcbTWH5JKxnb7xCxCpnWNbMzIoQuA3Yw9yHqpT/vsGerpM+x9M
Pvh02Lp+vhULnM0WY8Ct/PFpKfcFQfx1Ld2xM3JjyDfmXE/lLyhiRGf6Gfs3l7slrskUT3eRqbA2
yMNBAxkzgPVbP0NOWTDTZOtLEgui8t7drIMbxO3HrdqAJ/FFXxrLOv0CA+yo3n/7TfLWJrX0Yf7x
h8C0hZGoO+sDTi2P6gPD/UVLRqfoSIlrvGR0Kqz/tSNsTOm4gTPhaHRzhv/MK582CvJEXj/ZzYYn
V1VXVJ/rPexbC+SlvEmlrJBOffL0KEq8X8yQzCdqo4D/aJU9NbiI1p6bGEaayqFAUWjPdVgUdsJD
SGC5q5op8ZNsxSFunmMqS3R1cy4SZgNdPhopl39DSeTX4lRuZi9c/GQTkTPCu5VWaQyXNt3w5Gwr
QQkoNe2GSNgmFPv8wM2AIrLfVCTWJadDz72XNlIebjowAQZ29RCdj2m/vMRgzTC2R3Ggrc9LynLa
YkOQJSeiFEMOn1DJvgD+2GQnVjo9wt0R2CcmdKy1r+GGhsVBavQ7mqBfTynujgNFptUEdtUQD/Mx
lccavHPjZi96IoZ3VhIf3iWQ5i9j2nTcYIuabVfHyHDjdGHzDyZd2yDiTxbLGgcrL5YKRRFGuVxS
XRSDLNwBHUTbIdXzMZwYY/CEsaP3s01FYyrrsfVJ3McMrjz5x42TeTjbCXr4g+APvZfdo8SunJZX
dkgJi9EsqarG2DZcg3996DXRnB8rrmTjTRpwGzGSpLhgH5Iwhpwb7sgJWpGBSGxTVPkW/7lezgWU
/A3eVhiOzd1EjYVuoIzVvJ+imTAcZvh+9Jf8D3luPuSQDuPI4ep/S8ZbOLC8kbYCprMSfbNTVNlX
oJ/8T+/rcrjVWLWSTWXa+VAfVpuSlOZmZOtfZRv/jbmfZ2WazcopvrEH32RZGy4FoqdFvWYA5plc
MuS6hsdl2L3vCfuATtYPgGgeIKL9ZSg/8SVLv1g1xgoQFzb2o8Y5v3CyAFT0Km2kbg9iGjxoGvYb
X0S6eKEQyPkjDZUVJmc+Z8lUHjr+G5g3ugxwhrpX396L/u3uuocrL/GgnkYNvxN8Ytsh+tQZNkKi
qov3i0r08JxYrQ31ujTnoaudOBbtXinRtn1RACfPrvUwuMakAZ3D6H7Bn8spSezSlqMyiCnhI3mx
qHzQMOFqtCRlfSAMOThR6fWlrZmVhcgufTsHV9g3CCMPpI9tAIl5CaJEe67X5wmwd851F0LQjxrt
XEgO2QIgacQ9Azhruh2wYQoKQu2zSjFI+YplwfTazAFJf9f5UurSSZYhbb2h0r4qe/R1Wy0Cw01/
Qu5CepK6Jer50CuKou1FERxM9sk6qRb6jDvRpYo5Qe37b36txPkHhHuetf0YV/NYG3eF60lR0QMw
xbfOegxdoCswO6YMp4w+mt3FwFLAAxx3ZxVN46YIVdduHfA7iI3JUyTA5N8uZ/BzV1s0N1InIDPJ
avWdUK85Hsp0QKcMdFT+YoS1Z7YT4nj0+D7pqmGf26+pOzIK80cPvW/9IQ74J5nGB95fF5F75hLg
F1Hu7jN8o2DGtNEGUlg9zo3KZ06gsELBOpIlGewejUJle5K+7rvUt7kM9P01V1JnYrCc0xiR1OeV
w+uldAsCtnD/hhGrJ8xaMNtzFx8n1Rf+hQiJ/A7HBHqJwqFD8dK5ab2OIz7An1qL9tZ4zIMhp1rn
ZxQ0FUF5zEDaT3fPMxTlQR1bCy4dWxaVPzXiMseWiCCSb+8MzeeRO3c4oBME9qzzLO3f73QFXuRn
IFHeHE4NC5DJcjPGkns2T6NcigiOMu7Gol4azj9+8MEh1N9V6hKMmImE3Ippqp9ggSkLYmvLgLu4
148zNkJKjZLpKHq+DR1x01i22tRKDzOKHpc7zP2gE8+dE+1RVB59o7BtAQHT0atN8hN1q88keuwG
AYVlhLHJkagNNN2KZcWLpHcgp17aEJ+pv0oDmnF3nhT7CJ/BPnMfFq1Fusr6Ogx6pMdLVDFczuw+
4YNMlhE3IsTlA6d+PXmrC4S8MhUSJL7kJWoaWnMjtcIqNb4+mr5VNOVOBAvTj91A0CMXNwGtOHlw
Uz/B6hn/1+JUpGwF7qCoo+Vwlc76QEgrsPK0jGTTG1jl7tukZkjIqqTefH35ihzt+3TAm6GqCIs0
e6NwSStqPpHm0O4p5ZdG6+pBfjIPSzT+TaG+d7GEGOARphU2WsK5+XctOQjyz2ZmLmRq3vPC/PQG
ysx5bptuI0w9VJ+Pl7AYi/pG/cRjdtLJAkThl+g2F/je/iqUESxpqWi5C/tUELw8kZjXQsiud69L
wYAFDEfqsnzpPF9wgD++wcOB/KAk4KS+gyu+aYRos63FjVP3pH2a6BSG1YmI4FTqoVPZu/S7M0Ls
eo9LMIHPYHfi8tbuFJ5hCheqdTEgT4MfoqzBqCQJcKttt3w2dho58r59w3dxvWhJ2vby3fGy66AO
uJ/zpkeLREq15j02XHnnzoaKIAY5xi9HQ6iccGYNniOt+3gjANzT1xA6Pk3LdrkWfr5aKrIbob/p
Kimo5RcCZKC6AE1qSAXfu6XmJbZ/5GFNf7PFJ62z2Mmctwfb3LQOLhl8IGS2/XV0PvWnnUOcBkDY
Q3w3+LpQlJ7vaFdpKMH7R416Pdi+w85CrzM+rwFS3Pj7HvW3WxyxnTJuwjxVZDEN6xDwwwJ4rxBf
TQra+4BH4ZlclbuqZFK7vwjEmey7rQ1P3srSLb82jAYU6l/Hen8cJcJweVgom2jQli9bbMbdkXhR
eYJD4m36L7F2NHxXtAUZVzr5kTkpYLpXlccYXuu275goRdlHdJ32wO3CE4tZ4nCOntY8467X8Urr
/9Hn/e7MNUKi2Yr8B1CtLHPbKMxEniTM4hS+mRxqlQjRBLxM9GRec+JVNUkV5HbyS2Ye/zgBVP3f
lkFZE0Av1Wa6LwUc2dT3JKTLy/KY6nJGWqPsN4F9U2BceoxIKNGcCj6yTa3FGZbQJyaYvLe0I8TI
0+93EDc4py1nLxWGPOJRsEDIC0w+7OMd5PIRWN727zTWTL2RcxGRJu0gJJlYQpz1E8IU7ThFMNgq
H1TgxkAMOyqESRKCpr6mcKQutsbQmr408BSMXTnazWq6+O+me3DhuEdBwYjUXu4vW8KZByCUVL8l
9OwsNxh6Kwx26FQUOHMoGVN3HsDk7cNeLmZMvahRM18dfqDY7nezJxlQ72/PExnI5y0P3QMJE9zz
yZTvo3vPW03hk7gHy6Al6Zu2LlNn8xTiOwabxwKGW/nFgmXnp7+4AuXknkhPX8/Wx0J7f3pgZKux
SzBE9/V8nN8l/TCLSZ8Hy84hb9WCuaVVOtM0yKTeOyGntG+Ji49VAAZO4yKIEsC6sJMZqgCmYuhu
DQZpUESLZyFJMev+Z8y8ZaAqLzop16Ukyh/ufl9UslTh48C4QgT3ilFck3EcrvDfhbQRm2hV3mzq
WytLYroC11OC4eOGiU4Y5vjzL3c5yIi+66nJtcpBKHl6QExIC7Y8BWTLy2wSthWTdc2eI8HjD//m
g0eCNdjb79FBpbDf2boMcqjIYAjoYwJhsslagvOxeiswghtkWejo6+imFM3jiyzmIrSgAUssTUjo
hbLbIJcLXECdxD1Lqe9bQ9cyfHyVIH5Ve4dPdgtXGQPL4GycmEFYMYUxQi6vYPI5bnM/R8Kikqub
VqbZrVd/T+L8utTahofbhwMmIgVsX8nflDnMO34LE9lNVpxXFkxgRoa48Aix50aMv3USu/8riQmg
/QOHq3jAfkuH18SiIJxJndoZG09m/I8+kTF8PodSQ52DhXHkQOcdsctlYG+Cc2uUrXEl+gxzrCHl
AzXQP9a3VtQhedKvx7QTrbyl92GeRdGeBCYx5UQL4WeIpvst2bP0Uj5UXnfxCd+cLQAUiVbu1N5d
4L1Tu2v4YRGab2ATrj2kvgz8aGotL0t4lShNqGslMHtm4U4yLzv4AFANfCpCSWcFh/lC80AYQd7V
rlJ65M85PYKiWNFP633QlEVh1iMNW0qHwJuwJSYYczxxdu0pMp4tMKR4HxOpBDRAOIaotx2AQ4Xx
rQ1nRqd+AraMfCGd9ckpXxG/6QY/EJy+1vUccwqwaR+CVMxDhSkWcwPZXHEdx7pRt/ZsPCwlj271
w0ubFBDJ45BA7WXasZWQfo5vZyghUHtFZhisER3dkAf2uDOAUPQTImqnVmzMTC1UD/nIQxGdDTCM
0q4r21vHVV/S6yIEwWsXsjqZapKuvf1f9NmX3Gim18LHNLWS6bjae0mZEJkBDCAp61zLtKlsgAK8
m5W9KKzeyiHqPxY40i0dnzyE+bmENtxwNW45DxYrnfMctVV4PJnhCqxjBDb4itkL3u5izsyRVs/S
CGgjbqrxL8957B9CGt+Xf8MKlGC9bzlZrkRw+yHuxDZLc5yDVjN1QYDU5BXZ5+OwEuPHlPX6nl85
hgoaPV3GWMOiJ2fYjTivcvK59KliEIc4wdAWn4URHZPZSt5G1e5M0iCuL9C15Ucn5vF01ZHOzss8
/1z7B9DmB7A5503r0mx6DnCVZjtOlBinjcEST6kEhWNsviL3lW8WlzYC6Ecd+zmfvWdVQXq12iQz
bxAkA6avCmto8VQtdpmWmth184eNRf9PvmOvDG8YREWqE8p6KJeQB9I3HYwKRH5KsrbR8H5no/HN
WtuESaSdN+rOmVptLkUmhTZ46i9QqS3G9/b3Q0LgFVIsF+KfAIb+1fPdCzVA1YJljw2vVvQO/6mu
NQKADbPMgIHc4/9e30qbJXPD7MI2JrGaIgHI3TGKArHZLuBWJnMTHEu0twWA61i2tzcU+gQDSsan
exw2h9MeyDU0D5E+d5qkDmPO0AJPL5DR5kh7Vj/9fhdEGHSpWb/QpUe6sIv6CQKyH7Jt7ykh5M+o
ZZJAQNqw0siM5AVp1q/EhOoKRoAH5WiA8bBH6ALlbtk9SGJudweWur40ti/jclTyzhUzBTLuJTHy
VmYJqVpu/hszf4LfMz2Pj2pREhId7lcIOv3Jvh/syJqzqVrJe4vJ+6unl2y49llcCtESOZXFi5Rv
TZLyBCL/j4pQCBpPXR4Yf78V3rtmCTp4wwoN0+UzifG4x9mUhVHtOS0AziUc5D1sUDwdLllDwMwn
5pMxnOsP3lrye7IjeG0Cwc8KQsEG00Vzpz2jkHBUy3xqh9zxhJv8/I+tVkG9aZEQuX5ZCcwhsCjL
iyXo7w1IKNoDkvl96NxWZPcu/o5PxJ2RAo5+DnrjTgFppG0IYLE6xXaiUu6hx3TdNXkaipEnfjFb
4D7oKR503cir/arYwtPe46oPswYAF5JYZkZXXj7zUC2ZCTyxUdS0J8YmdcSMpKfqs/g+luTNjrmn
WxQEkSPK9QH9E6dEBFMHNPqkIXcMU9S8MlpBDnx/4LrQ8BIWhNOxNEb+JwbHudmWcAQEp9DkR9OI
jRfKbWtnFahMGaSR1ZVcI6vsCSD9k7ZHLCrUjxz5poCAo92T6HaRjy5mrCMNvXSZlN2PxdkHSrOB
wH5IJMU86u/kXGnu0VO4YPyXHVwXSyfdSfuYG/73XAqM3rpAcC8GkwF0Eb3aFjq6hTA0xt8Knt9h
w8YuYOwU5CKnwc184Eb6do4XnDIpq8L7B0mzo8ExYoWYc1iAarFsuJGi3Din+kmtui61XT+Ns16G
m1IoaGdn8WA7/vl/82ix1mvJtAgRL2XbJmDNBUCwbyxC/1+AMFC0hgYMQ653FA7geUm77ljZu2yB
62dRhx8C/W+wLWqOIeA36LgjHr4o/3wmwKGmnSQoXSu108lJYIeuNIJzQ2ouMntlHHYCwxW/NGql
KGX1D2VzXCr9reB3Wt1/1V6MUPDmN2bv8mqqCwlrtPTCfCHLd4hD71MFNzJO54FqflebakoZZ0X9
reZI3yYfjDVI/ME4z7p7UOhwxX+wYxN8hhV95aOZIOscKX6RAfvb6STaQDuOmI6U4QStISx7Cjyt
FN966IHQbRQhBb9sJooVb9vIUg4hgDIY0Z+HfDJ0SVlBe0nxIWEjfz19BJhhqS0VjjL4FwvJACJN
AiAkZKiI72FN6pvbXedeG0NUrWrW+zCstoGAI0Cf/xi7vPgQfi8FV9SHW09LttAAqzDa505ga7+o
y52FWLJwPSdXA4mpzESPUAATk0vBxYdFdK9uvAJ1jjTr2MqjbFFTnLIneC2C7zrocS2/vSIpr7eF
KCo8AxbMqjY9GSwij+TyRb+fG6ymXxnMY6V6ESZx7ge0rxclgmm8W+TQpmfCyKZE/IPh9i0RYlyz
Zru6YB6V+UyZhYk5I7aA53I5+J8OlNXRHTDnLhogp/gMIzs6B/3SMl8q94ZwnrZJnOJA0Nh5Ho5L
nbeOMNCGMQaNHbmWLZiqrs9x+PoR20EDEeCgOj4g2B5hJmhVCcblHc30+krmj5JxZh4jVMomlXNp
v1J1d8hghLoXpXvyzGVR1oPpRB/eMoEOlMcEAXLqENDdhOyklDrvR9dir97eDmWdG6TrW8IF/eWG
pL9TeQwIMuEM2L9K1m+dS4hGh9SG2RI/CRCf3K4O4d7/bcx1aaosveR5XmScbnBUXmR6YgZBqI0q
fGzHliLbBaZ1GKRN3nYbr0TQhmJE1Rrburau5a/gTHRnMH0cJk2RX/MQTaFFi4wWwJylsrditCg6
Tg/9Zw2cSwxs/YXvU1IlVJPy2Grl+tBxKYXfUClFEyUyBnbqz17m9gUR/PwnGhoeAgHfzdhjPejW
m/Y2Omv5PZ6IDBWL+z+ET89RWazkzT6O4XJ8S2hykp0/vcdQtpVXasVdm7+jO9a12of+xtOPKBIZ
c63NwskJi8EmltKANAYJJkJsktqM4ThyxwF8mOSN4ZecSvMOGlfQdLQ5ttftMxYGVqRsRcnsHoDq
8lBvSc4CdD2qH4RrMy6GWlgjXZ0lhy0f+9UghXtPm1y6gn0okEFI1HcuudiKFldJ4b8uzbBMn/lV
xFpbhPg7hh+uLNyV9cVLi/qfklhfzWGEZuWLXPjPa7Rd4l6xZrxqULZotbCjfetNVNM1iDUT6hSd
0F5Pd7NFO1WaSw/JOAxBcSQ2UY676ukbpSM3YldPmg3cnYd6wmI23NORR7t3Kv4DUTFtzhbC8iPN
AzTiiX0iOCETcfzYRzp8lwH4o+nAWv2wIDvN6oad4XYdlvUpJ7XYGd/cCPAqC6VTNCS0Xv3qDrDf
bS4W2ogTBOBD2W5l8yeZNasBDFDTMkeRveRMT2O+sV22t8gQ8YtwTmAZ1sjR87TG626qe4y7NU3x
HmMCQ7cywFjdBWdxAD98vv8dsz0e8mliyLxdEyZJp0H5v7kzeB5C6MIlp40jA5GYxkEGxrDJWU9J
D95+zJ45uQJDS9JhhA05G8rmniGvBA//78GgaiI9/1jSFiDojRaR9C9F1nvUe7zLkCKMiImNg+5H
rbUldZnGkcemZNiE9cMlNJxZN7+IHjn+kzNN9NwuPvFv1CN9tHCxDnaG0ieAxJOklKafBWjWlcoH
wmmmt26uvGRifV8nVg/dB3rXCef/YVb4JGTHWSdrW9tvyfuLO44d2A7itCoKaFdQ7V478guX/V8Z
ujqwK2nK+ao0BBhHmZiWdwe89ssEi6jDa9gVo2Obdj8pRbu9KE3WdIdrLg/4RYWgrjb550O1zPVK
/a/YO1ah2IjI/+erGJnqc7X48X+E+xHcLKIY21oNCgyqBtCRsrL3d5L0+PdZjzdj2LZuE08mo7m5
dR6EQRjFWcWd4UMrHjDbyrANy8nrwd7eTAk3nf3d0eJZoFJYo2KawMFUJ1lBUXrLuDXzTSXQ3QL4
8R3mCX2+xs6vaUAdXlsFsbaWr99tSU9/dHELcnJbgRsqSOYGdub0UWVZV3wElNbpuJYwzRMcqp+M
ecLgkBCmxRs8VyoF6fnf/I069KCPEY+1RcXypocEZjqAY1h4jYF7LGX2/8QSwcT8cG/CQmgQouqN
Po80J5fN32D+W1yVNU8vnvV/BtRG/IrvmeNJ8WP+TDbmk1sqXgTfkydJkRCY2wFHZjPGpyyVaoeD
GN2Fg3bCQudepIpE0HiS68XKKJJAigd7WJzkTWCecT11b9NEV5WOhG+778CAqrzVGlVpN40PbJHx
bDmn+guZs0HmDMswldvm6hZ2sHUyESIZMZ1nGYLjLTaxomjHzpU3CNRLcJ0XtfSzwgK5xaEhB2zk
Hu1PbzAauPsq17rEOEa6rS2027F+NEye5EyEkvs8DDZVJxI4GU5QMOFcKjoB7ufu+9ji8vPhsXt2
pRWiPaxYLKDGCU8rGMkT9KH1aWTRFkwjXQNm/93s54m2TMw/P26msD3rgfx5Jg+QDdmiWIzKFkqK
4Iag0UmU32yJmyYLFuCVbRw3IQjR0it51H+O48j7woAwfiMZNOsZGf60uXW8AZAnKHfQNbSiIRy9
TX6Hp90sdiDRL6OJzviZ7WHK8SQWjgICYu8agt8SPuS/v8RYVy4TSK58M3bizZ3cA5p7HHpv9zd2
cu1n8+yumof+moqXBQwEU8HLH3zrryTZ3fYmCX0Gkxet78d/0LGuHmgA0ID7yw1mKhVW9QFzO9lH
kD0HpP0lphthqE29uyqsN9950l7ViBw8yW/ijaWjLYtx/r2dvrc0Kf6JxZLcFqXjTlVJXAHz71kd
w5hwhpjifPq7i18vXM80T6gkuzr8Pgpc22mhzubO3O4E4MHaFEJoDKYazOMIDd6Lx5beDjnPNLJD
SEoyQrwvFkbnTeKNQV9dxvohItBUGgsRfJ/zbcx8PdBJWCWlwfJwUC9Fa29R/8oTGb8mK7ZKbonf
4BN5I7Ui3tqBkErJp6fX+Jdax/R3LVuvaCSnoBE5sjDS0yzHInoLI+7nBNMv7taNw8KmfRmqfHIk
w/QUz48lnKCjRY/AZtwlmHvxbGH533zg3v+rMKiv/jfuulK6hgyT5mjYTOgrZmxp2TChBtvbbjMD
zW4FFnlY/+8tx+Pqi60/1t+8Ew07Sz2m6KupiqusmQqsg1hlcAjpn5vKeLoW55rrc6jw08Re4j3E
dkd/mDOFuPk4M5SPA2/UwMPkjnZ70Yc4cXMvJbVQf1PFpzn6xINas/7qGtJZ+qoO8TKCobWMJIx3
p90xKNr9NFRwPUe+hfo9kS6aAugLO71Nluoz4b88J4ESROEN5mCxn0iKvrwlt6XwXdyKtIfA/3Te
z6miYZR18UpF1ADoOwqk+jcbh5oMjGjpJCGekY5FxG2ZLFaIr0/xvHAkV+QifzfUkAZajjdTxYMB
m/Xtz5DV7Co6EqzXO0Y9r5wQDzK/LfcwiTiN47FOGdPLGQNeyMPeuCD0/qq2chO3r7114K84nq5T
/EzV7cRCAjioPQ9Q/h5cnkp8AisjTyVp9cADFI6lfPf2uF/Z6YcWjdrV2NxQvQj1xvFcW9i8EBZb
n7qoU4a1xn5ZXFzsQJ7pXHqQT2gNKOTGNIeQHSmq1NcW+LJaB7W4MEw138RYLyG0+ZNTYvdjkE6d
8fwwQy5nd5Ho6/oHxsgbnhMjH/g5M9K0Ga6v9GHz4oVyYBDpScU85a8DaM2UlI/i2HQGCayLZAE8
yDyQNo/5KMrHWtPMnQAB3HCE9sXQAdpkdYepa3FLon4z64/Y4oNpzjey5b+GkBGfx4Y27kgysGMd
RMRlZ5WkF2eBhd76qkENU552NZMqiUGuPtwt3aeew9r3/8uTbgghmm4L8weer3xIdkv7wYaqAgzQ
X7RFLC+k6y6pehd5m1EyV8mxAMRIOXw6d4ZKp5biUscvpjRRP7BvWtP7W5WKYLbBQNODFHfiO+ax
ElqrX4aBAh2hApUtvyLOg7mBPQMSyjmQqmmAjSsqpYkC2Qu5hwZDpJ7DgscZU4sQGS7WKC1BcBjm
tpVhLeWgJ5STdzE2fu801rIirXmMmvooMm0wYO2kr9zxrsdfecSdrVa24zxlzcvh88nDzac69lvS
bJV5iCUqeEaSiBIHF0THzrqGGcw7LZKH8J4wgW1ZIqriS6oGE+yWPXFlkxRsV5bkwbHFaEnU7CW/
kCDGU25NZmSs7OsPYrA16nkdU0JB4DCqJWaF8rPHWflQIwjn0gkFP/APWWaY6kdyHtaZ/U276ZkV
u7IDRKSMlIgpZctugJcK45dpFPhZbiYAfZSdbHPWpfi3F7iOc3dVx1n8Yw/punERTzKtK3zic7Nu
cJSnFLTpPeHwzJMSXHrc9vC8hmuYYkkMT8stGavyVJxKo/Lqk0vBVe3bSB3wY2TZ8nHDuHSzo6lK
X2ttuSd+Y/DbuOa8/AjhRYvDLuB2OF5GP4XP235wZiWViGm0k5GCeCMAQRFBKQ+H2WojRW/jr+vj
jmEcAVD9580IdBBbV63XG739Pk1ks8d1ZRPO+JUEp6myxgrl4HwSK5pogjRj7YCnVGIEH8rm8cnS
we0MlKd9Gz1303K3rnMxDHTfg+HhuUCsh6Mj4va4floyDiLhTTjcDSmrYZOmVzTNVkTuhmWtur8+
m5FyPttG+X99kaHlwJZ2GKgfcWQIPYNegNqOL0GAFO7QcWjKz5r8uJGifh97TX43qlePz2K/No5t
LyEzBhWXQOfxwEYe0u3OgKElNLAKWG2qRXZ69J6Wnq0M4qLjqCc3r0DymN8q9g5aESiIkxJnnTG8
HXpP6xjmjaUi9OSH0LIKq2mNl4ZsuJW0wwjmPnRVwc+56V2D2LxQtNqOwYKjFia2jAHoPzMH6MRI
0XzXyJjqCswucVkuCQb++eZQHWd1sn7ryzHCnxQE2u5IIddsso/qPy9cbEqYkWZGmIkuOeo6e/8X
8dja+cPJuuRdA8NYcjLliQ/FwB3Rxfr+mvMyfDejUbQsqR0naUoABHh5VQZTJZlGXxxl5rWUwNGJ
KGEmiqW7ZxOAryMDAbqY5zpuj47/zX5NN2/kGBiC8QpjsG5YHn55Nut1DkciUVwOpFww0BA/9iru
rLamLDwc0PPD5P+ZXg8KAPlfG92GnnjqxrCDiFN/8u6g/f+3WDRZbR4tGK5fSCeZG8XOO1r9utTc
5M8YRpLZrkUaWClDyyX3rGMZ5XslXCYIX0eiPWqYovXhCXeoC0RMoVavglVaPSr/Rx3NWUqEdg4q
jlMWacYbo0Z1XErsRLfwTYwsORlbGd/6Yy/8X6cZE0y8j7Je6BWuT/e2rfeQGbF5CpG5sF6sUP9N
QhWyKoGOWAiyOFMIwsoK9+oPXsTk4bewMyn/f1p6LNJr17+7nJpUALYNUe3WZWFt8K+mtLxxA/uz
+JmBytslIT0Uu5FVHnOWNwWqGrLE8K1NH4/O4GFHBH7SOFMcLEkzEYVvuya8+KpIwhzxuRkEV7fs
Gc+pUxwfmQ7YIuX8s7670n0OrWuDsEvwAgwY7HRZnQPeBbuTivUALuTSu4uhaUMBxFPI6j2WK3vc
50Vh7zqWsOl7NavRW6j2gacf8mCXFtS8m+/yUg2p/tiiHzaIeNrPHKrGC33qn4wIqhycOBmCRctq
TCn7dJVpV1J0R+xAVk4Cb3IQqfpShndsOv/RuyQySvfAiJqB0+AbZuUvNcojVt6Ji9GBPMEMKX4f
GZ3JSQEPk1q8Vq7n53xiexr6iONgEhqnDtj6GQV/epBB+BKS0Czkol7zkC2oeeA6s7y9KfHX1Bmj
soVte3uuEjFkGvk1xECDXsuQGb+Fa6Vpu6QlrX3K1aEdVA9GgpWdotnOrIXChgQYXa5V4wgEhX31
USLlopMEjASp3OXYPcsnmu9iA5r/FrtorgTY6JsC1+bTqSSN45UEPvEvAK7DGjdfPjsT03PMmsIM
tYnx0kVhJbtcBRkzzUpUXTx1ttj+BlxltZzJgxQptreQ19x8PZr1uXusmpJwu8e4BTO4Q35kPW6e
A6W3VOBa3OM8Ue2eU+uQ7JJQ+KbXwXdkG9w1EOietnknf2tE2mqNHeHP6Cvvnad4zIf/TgaAWnqW
M9kCmF8NJyAzMM/JAKT5VWynlnFd+rClu5ZgjAaujSSTW+MT5BN0O9ZS4eabK3xeTefYseDcXlZp
mCaqLVa44BMvUY3cTMIAsX+Y5E5cjHUJMSlX65p+s8wlr54lSay5b7RNht3dhmm4xfF3gXf363Mm
XnDJFyqtOd5ff4R3cSMMLn8mAFr5TwwisCcfD0/fpRqnosni+9QWObtf048gcmyvt/P+R9xbwW5d
EF4TeMpbZPQruQD8GzuPDbx9LRlWXShmwxBAkm2i8nqfvn4OtKuN3/7ZYQdgC0OVrc5jgWeCbuEp
0szbfJYw9d0hP3kSNNU50/Yxf4S7X2eG/3Vm3Kxi5jgeA7nQYSVJfI3Sa8X8t6dB64FeOzh8ZX9v
ZyYBMuorfHZDacP3izTnKbjMRMX1RfUF/1i4EpF69jlVDvk6w0/cwEAkFQIX3DqrBOmxeI/0lidu
oniLPDLX7b/oPIgDRIDLf26jxNuQFNVJUMl8vOL1KpKxk8Vk10QiFt1G7cNRjvv+Aar7rRztj+uh
XpPg2qZBRc2ef1rO4H2J0Q7fYT/fxFZm6D8jgGbdSl087XvVQnP2ByQMPkaSg4NiCWFBTaqe67cL
coa3cyzwluDX1emg3xpE35eOulKV+cy9uI4kshKBIfEGeaUmNqPbTvib2mPwMr4GlXcpzGA9/bxq
4XjFQlMNFttR5Z6wL79g10+m0/pZe4NA7ok6uMc266qq6URUQ48qixD+44xHZPYENbdkhN7aTfT4
/BSN9WnDyiFa4MBfyTwJaJ6gl5Z/solKNRAY38wT493vgB5RmS8+sLfTWIkHpU2JlUL0PrAz8h/D
dCDcAmZ/VPz7js/lxRBnRwdE5bJvqllJfBwOONxzLPtsHpM8NnZspbKgro61SSb0AUKQVzBUITV4
LnqZIbBRTKCy/fksW5+hq++NSYHWYH044XPkJdmIGYVWIifOTp+iApoKcBdBRg0m5ue7XiiFq1O1
NdHQKtiS+YzUJEEw9fg/rKyvHe11cn0x9H/2nAli0BS+4KLVcrowd3eRCG+KtPydA0wKG37MQmcc
3kjHJ8lSYHNZa9bnJ6WAXxbTsAttUGD8LurgmQGmPOIGUioJOqfs1KybKNeQWU3nOPIZ5hPcboxs
GMVImgOhKqogpKwZU5t+hOOPK4/yTIAKR3Hd/cHuNVLwdNsGdYKGu3+z8NkoZeIYyqquZvfsyVMX
VVfQDG25HA83LsF2J5iIDiHs/T6H6O7WNZPWlrFkkDRPX8RRGfkF8/7AcV7hZB2rQRDdpNzBDsh0
DR00S6NnZuygPqmI4eHPK0Pgi1UJj9hU0JW0YhL3LuVfwkWnkonQJH/7R5uJPNRrrc2f//ErmBIF
A06yGnggefaw7hGWGCQM8u9eMQrTRdVQF+vd1IlgWJRYY8NJJGW+yaMTa903ccMpjrCa+NKB3gYc
DaQCPR+Z21SmkOBBLH6CHMBFbvRrVbOUCtaP1c9QEwFdjp3bfxewRCXoKqQcLwChSH7FlvQQelRm
GWtMdpz9Me1qHK0K04Njlwo7p2vCjVY7w1sX2Rg613+jH5donK7SGZi+207mzjnVFrQRVmH463Dk
0uWorFv9Q20GBBpitTogL7hW30Feat8Ju9hKsfDE1COkhe/OaHAOSo9Ua05NGwi1/5BqHV/JXsIS
sZFtWjbOeqEQ4EA9DHZZcDDSUYo83yevquTTYgB3nHxLHVpYvr/T7Z6el3HybaTLWnIgOtVYKmf4
H29DIY00PRNzrcChaLpKCDtoE/amPfrumrQXyBq1E+MK1UoE9gUcE3k8o8wUSiQr3Yrt9n34xjgr
ErXArJvV6DfH8fNQiqbhwAd1axDbjnPuOezNA9+9yyMALPZGZKzsw6GAjMk/EhF4sZ0FlK5PQG7O
MqpLoR6rj07WtmD+jT+78SFTXap8Ut4fI9cvKOyjAqAOp0tnvfUyJ8KH37eXmYyw7U1dOfJX5LO1
eoUho0HMIWhTK6JiKBJuYQlXcug89e2SHgb9YaeHKP+QSkmKu17Cg4MURz6lYG3xAMuFF9b35n5O
A/ljhLDb9inBhkkm/oAIJiYSNCjSXK1mz/cyn8bo6RGQNlnUZvD9OgJjWc+pTnXrfVKPaaKQPckK
8FAiiOy6oQqXhDseZqh3BjkG+RWosFDj7AmK3sN5dRfAWpwWXwN3tBKJi0xJK3eFWYTaivYijZCw
4bFzDgiD8XyTFHILNDxGLHW+cg2TDWmogE/T2l5/lFoETJXRijZ7lNWBW6scULuckiljsjEfbHq+
JwwfNJ7NjFC/rxhIYxAxIzVJnQFaNV80sFJ6OlM3f2c5PcaZQ0OOAPzgiSlGIoSj9WcAJqsC/0RP
SSEeafYK5FytYCMUzC/V3IPjDMwXkqkGR3HF0nHdG40V7geQDsKGoFIZ8kCFf8J4D9Axy/FNiBdI
BfmXy/d/g4cxJU2tZ186LMkV24HrQWaR4noT8/YQ5Dibkrlrud77iGXuc7RxKnHkiHEkU9Pvpcyf
zOK0bK2XIYOqZohTEPXODLgmuW+gcZQTsBn5ILlPTJPJnmxBbnHVQhZiJP1Reesq1x4Lj+RPw32z
9DmSMB6FZVMJinZk+sg+bFbMTJZe8E7fktXeUzGgZyLUvVD4JM3zHYkmlXlAuVK4nO4LDqm7wpE4
KAuVlJ8VU0pTNFRaqjPG0ivjL/2L+RzvhKyB1SjCxQu9x/eS79hxFbNMcwM3rK0bRPyjFiuHTMdA
2eIzY3rWXDioZxHVGpgoU5TfJUlnTv84Lp1qIpigsmaH67QsvhQHCYkNT6GszTBwWhzLva8lGsU7
aMcoor+wDacUFsQE2AbzvZZCqYmfAzt547naOOj1avHI9sLUZjDNSB/zRT5ipOCdEQEYFPbzZbQi
e+UgeEWHoXXhuF2AFB6quL5Ne2pYHSgruvIo0YqA3E7A0cENhG/bE+t40fwX+AMmGcA91Jogc07r
6siV+Vbg1TFo4KDvFQsvTs80rzJESKo0K95qZewP5Udr6HRTmaTuR5Kp/TAYbmpEMOWw4/U++v5Y
BQ9VXJQHW32DU2eAcKsQMkWGHsv0Oxil6mKxtCZzriM7ux2KmSqW0VT9UqyxVkfcGZ80G5a5dAkY
ZW8+yyginI1JExVmSpX3VyTn/Ioe4HIzj1p4/D3CpPDdYmXTwHnRGLMb7L0rcOm8RVVlqt7DvA/f
XHpPzK1jmwVXvBethADI7miBoygkSn+d4zGSop3gq028P3ObCOh5Qz4DJ9M3KuQIOT3LFd7fCiQr
1Di6W11jV7ekO4XqCAPZs6NzWvvFE7DM9A3+KtCMfpb0UldHBYloI+/DCL/hA8fkWZ0/QsNYjcs4
Crdyr8yOi11r7noZnTpHzK9YwvHEJDBsNY1Q0gLKXyx34W0dALZ69hSIigMuwwjMemh+k5Rf3hcv
iUtGopffI2vu9cVXpLH5zYGJojwA2nbKgYrlNVXG2Iz14EWdhxvD8W1a8KRugogl96IWZzI7bKqD
1z/xRlwOG/ujdhCeo9hOxzOVLJe7l8jmURPk4Qg54SXWv/mEo4E576TZIlQ5T4K6yq2NCf20Atmr
5NRhxJrWl+WAPS3uZXLMMLMXW7bxQZ2YD3fszSfiFLnVT/5Pg3z6EiMdNZ7qa7LvclkxxuOVVz0w
W/33Pzdx47729gxDQQcGYx2ALMeKeAAFN00G5a5d75ewv7GSVgMJyMTYKd8Fxk9RyZw2OD6I/TGt
e/UCezexG+ExV+OqqLdqMaed46SK1gCMFGgXDFtbCi4gqDzLnQWYg5lepMljhts82YhodQQeopB2
35CT7+ZXa8RqlAz+xdXGDX2RhkQqn7+4eHfVxAqBHsJC085GnGluK1456rI3shJyZhYMzZNXo+Ke
zDzLeqrlwSOYrNNDuLb3MmMF8S+J1waAVXk4KIwruBl8Dvi6djN0FQsUDqfpoqoG8Pgc6237JnKv
ZpP4t4CaOiGCjRvetdghnihjW8wbndqDj/DXSs0OU0lbxLFg3pMTkYHHu2Q6YtT++4ssufLY5HNV
8+uUTD1mve9RXgmrROtO4r7j2d9YMS18fqodL6XSUQK6/5hI3ZpUuQuFagMhqnPNs+L9SITpJujy
qIreZwo/QUPSFwaiOZPbBac7Bxi0aRXkKgSIcKtXg/+4e+x3sQYsC2ZjmifbQmtfiz2aQCOrzW73
urY8SL6ZpvR3J/mMZDLqeXJwBNJxVkQwj7EBOAp1NbXh16+lZahV/apXzbcIuFNhdDAT54cydVI3
Sh8QqkNIGJ4W+uOHzNmPesL0EDSWSva6SdaGnDS8vfNkxplG4YUZbP138YUnVkYZfSquw0+wGY6W
JbNdzQRJMjOnh63J1ZBxNG0irRypxIKhcyRL9sXJwEnB9dB7TRQ5e8/ZZKUIzDNYSx7LGIiKfH4Y
LIbKrMTXto0Esi5YgzO0MKGeZUrc9kgQbVpz3pq+fRRPalmtAU6VdB925fn4CrCUfa37PS0gS8NW
76LwIU3eKb2VR+Y+Qx3x+6HiXzl6E3FVfZ/vvpsPsUI701io4dJwOZkIT72svmAEyNBGY3KRheKj
hqTezpWDuuXUR286hiby3eUTWJSVB2Xo1esbgBtVW7hhPxaOJhAgsNyhag2JlB6SSG2DG9bnhnZr
hpxNelFiKPSrL25yMmLUbqGWmz2hJbzqDp1gBUJJGed9cToj9YteBEs0u21vV51Eyh7NGPWFjtB8
1OPEUmKjmW/p2tw4vthxoMdfwdjqrfxcRKvP4XCldsVtLfrsXIvUfzH6G8misU2trNTH10Gbvsl1
SC2I1rthvu8sUj9L7lmT/l9PYZdcebZ1nz1RrtENQuDpVQLyVolq0ugr3fC99thbotWjfMAB8kq6
FNdYWEasW5Ed5h/N7CFJ0P3SrYJUjBPSXw5Cw7dJlUIarYSOuLxZLMetEhi2WSXE30WeiIwL92DF
LzqNl8EVNfXjitPLs/+m398w7LsvBFKwIb0tXzCaOdXgFinwhoKeqXvthATjU0+7sWm1pyJnwmpw
BWAbvAgY1QbuaixeCEV+nIX0AW4AtFEvQ4xzsTg8YCOFna/r8aBLpkj2McQuVbGA5emkuHHHEifM
Li4HVtWIZvpx6qFIKBg+gwcyAO5kYoIq3LFaud+r8hX+JyRjTcC/4VE8gwdwtamqMzYzEwGfeAIp
fn/DItxg5/PiFt0hyiTyDFUbMLvQ/qNd2uDHWrAUk5q1aMTfq5Tn8HLyTbSsbzdGpMxGqabJUutR
v8Ulsp5QkbjMK3HpDO39MCr460Hxiff1Ux5pqHhOqjDfENj9a9Pujv69mJyygyo06ySRHY9KRHWq
rD/y3MF6gkmmt0YOxtMRUS2JDezlYomZlHsn28IIO1QdnQvL3yv78UJwAseS1eIFbsdITj35q+R7
vZx1+LJFn9qrAi0rB0C9xQPCMXbsoPBXFcHQ8H0pcbKs7x86kOVtYAGEYzjrijeKA4/0SKEhuyUI
kssIZ7rWPTHBsulxnoJQzdFZpc/4xnISkoWZEmGPPT3Q9HsLHOC/i2L6Rbj3Ah9XfUB+AkEg5BgZ
YOOQboLm+y5lTW1Cu2Hdjr1Rz9qPWWQew+t/eEyhru5Hw1DV/xY8tAKh1wOZCLqjkNE18+Oym9eh
92fX18q+KC2HY78rOFAbDQtVP3VNttDarazF+Brmwqtma3OVFvriVnnRvvBQBD4J1yqRK5xZxIOV
Fq4ekLtUjkSLOz3VkbyCLYTp/RseXpiuyDCH8JYDfqG1/aIfMQElh80n020rjUkgfOZQdSddljF4
sUP9avmLMLKrpXEfsiXct7ejaIQJtlruR+NcGNRtrQupmq+bvE06d7YScGM8wRjwDdQC7awoGqpG
CO3hONLclN1/G7n2v+1QMsubylfUu5nQWJJob2VuKcgWOMOC1tId4pHwxCDgA8Aor/m28+P5r43d
ioO0AtkeD1jEJEI62JO2m/3H8kNfF4jt6fVfAq/YL96ZlTy3BEs36Vb3tnOLbfusWzHUf9xoGvJC
wRmMuDL0j3w0YbCXOF7spqU9yYU3fOqm5PEkfasbOEWHwl9SPs+F0Y+8RUIIINaUPIklswI6o1ix
EWnlTutFoCreECsKOY+8r+neVvfYWZQPagcePVXyEmw2xwzqHsB6Rs911dCHeCBQoYLOZzFyIe9Q
5r0DwGl7uTvv9RoVi/Gh2EWz2dAB91rnXg1QkqzrVnrwYuEQgE0LP2jqiU5IJKSfRS7dVZc6klBO
xsx3kmizOnmFHfyIIyI4bApiT2qNwSfRwhiPT6jfOsmFDgtGN0x/wYYZPwsJSfED4fMd6ZbI9uW2
/bcBiVoYf2zsHbesFiz1Whg+8aCRXPBKxy/hwJmMQO4gFLJeLLvGMdXWqprx7eLWAhGrmHujh8M7
sEe8Ls4nETLRQovDw62jcHGiwMvNPH8Ua5pRH0zPVQgc6+jwuKN4m94k61rfVhOGFxueu3KOnToV
085g+XcblFxwSb27UPr3OcVgBD1uy8va+wCtJd7QaiKl/qG2NhSoPMCAXQGa7JJKa9x5z/n6rnAa
A08bdHHklvb8R4qmIQPzxGyD5a5i5dcdz4m9GPKpEHfZCT9x+8/EyCWBRkWjFeV13m9MPt3x03AE
96gReNajJQw+vRY/auLa0zpZXqmHU8A/AOQsEYqUy8UjU3M9YKImQ54lQ+wve34al04Omv+25OAG
Klgniv2CcSD38AO66vdTbzQLc8Rn8xXMxSj61qGnw6WNdU8jiByELAyJkzTPo4IS/kmfmK85VyNd
eqYGZMe3rbScTkbrDucP6txSjQ2yC2QAsYMDFGSPsUjep4hYl2XBwbFTHKLfkTjPaq9VQtaof587
F9aEhMfZsQZLl5oKH/KOMozTuAACmeDcC18nK/SicoWtJstsHQaxNvsTUTme9Daw4pWvG/HHxOyr
N0R69hOMhBJV1gOyz6/iOiiw0WPTAGcZ5YjpkVvbbhu0VP4DQMXqr+JrNta1+sI8paHYzCEluUkN
HRe22VsNOctANVMqokehyTSrBDw11mx1edrybyRVseABZ6CaywM9ke0/w5VcEBct/lJ3VM/1wM3s
sW4k0aM8PVXxEzea5TprhNGBkdDEWplO1ULJPiqRweEaeS+q6ugkIF7QA9zH8ZZv8pyQ0et9FE7i
ePCJrxGFdeIob7XBA5/cwvdEdVUo1aFFFPxqOGV2lFmfQJvE2BFj80jsAlAcbnKWqUqhwDYFs46z
fayCKGhq/mVoLNk3Vw/JGX0glWETuYhW2VnaldqvANT56R+OsxwxgX5EqokJ9OyzecoHNuhXMfh7
2G8Qfkyf4g4BVnS/g9z9gIqpigjQTOS9KpDlP3K7d1LkQNI4CjQbPq+37k9ei0YZ7+GoS1MQVjxa
lgTUQCp8yIrakxy1qnknEN7DWDps7JywUU5E78+24RfnMoOks536ukzM5ZkAaZDLhoRcQmAYfA9P
Uvej2Sjj7lQ0kPh4KsRRGyA0150oRFhzQLHHgxHtcxNwfktK4RUVustiw9yu/TPz2LvSW+oBbsBy
kF4TwCt/5GXFCX7BAyraJc4I6VOlwGkYAZkeVed3f5r4H83mO4Kf5lqIxjaKE7VUoamCRsyIRI04
b1XwoSVARCKOmTLEwFZuECE017ZBTZhtwL/7WjFx+2NRCIvvd+Y2ej0gc2LTPfL2XPvsDn57XhLD
oUtl/2yrZnAg+bTvgTB+DwAma6rshi1xqRaMvjZzLvPMNY62lF5WLP4UXkUidUZ+lGbNjSN0MtME
H+oIqWb+iWPdiAwnM3WIULAhF0qFLYldWZZJ3bt+Oou82vTeuCgRkZslFcy75SNk9v9xZ3yhTwN6
Ew6mNdFamsFg1jhUo6BsWG/NaAbFB2tGi2+nQf+/Tt0dAHJJ/oNaNmkHj/+b5ATgOuZJ8m/nlok2
OaU/BYb7iK4fSeMCSNba7zc5L+xTXIhKYYfuSKnN6V6eFPUUWoUGaFNyzh7A1wkfvxvUj4Po/fON
mihmUaAiiWb19+K7Xms2teS7zIrboHjcj2Ag/Kdy/eZ7YLyjq3Cp2b/DAU65UKdoaSfCGiM1REGQ
KzqUqOnp0iJpHPY3ziyia+6rfNdlZqQVigVVf42SdkF3eLu0yQmkUHxGC7HNgBxIiZqNTRKuF/uL
wf4Jv53Zoi7Sgw6BaOR7bdQvcqn3Zy+HM1DpNwsABHEp15vXg3j5DlrYPPfN3vLrxbMRKG4MS5IV
SnhYzaLP6Do+AqDgDDsTMrc1zXlM5rs0vYtP3FeqxE84iO/j+IJj1yxXcvkELwCRLflVxpjxdAWp
ZUeal2YdsWIo6C5RLPQHPAv2pgg/RlyYXWJvQot+L6JTSq88xM1pxz1Js7FDDDFeUD2jBOziyrjo
S6zyxaNitShqi8z98hmjE/biuePK1MCL+JYEntKdTG+vc955TgBybkQDnJiExYvlj6+NOzqVP7oA
tC0/ghtANdn60nfX6VeXJyg42quc8bxTUO4STYcOPE848jDQxRLPHEw6MUkyJXDmTOKiC2HWhQZB
fAlVNz7ExlQxTTdusfk6w/wczxoTZeSmZnVTMKZcEdH/N4T3sIfx0uqIOGWinsa9viztPJt1Ap+0
RfNwcFBWAftgCrVzVy+o0MsOdPjhXlf8Rwu3RXRF9aUA4BkVgMY/oQu+xd7a95r3qfNZLV65vFy4
/nSLAd6FZFP9dJaera5NHowlmbxX4X2jW/HmpZeF3IOfsF97lDsn1h7Xb+eJqyf4FIpZBrmF7vOQ
zLZcMpLS93rkmeqXkjmkud6VE5i19v/AmFZ+MkZZRTiViqZAdxGFJRFpywv+E1V8bEYYMPpwWaIh
txK8V3algCwtH6JHSyOqpI3E+JR90Ck5s1oxIXQfWKIGObYwPpTimp7biZJueuZfayiXzARd4DzM
lXWpEcvqa/947V2KYWB3SyLzYlZs9fh/mlWEtCIaR0Ylqs/JA/heLCW+mgTzxH3ns1430IOAY87T
gvKd7uYSzLpzNWhzUajZ/H/cOKPPBL6vXQ8fRCn6AKBQTIo8xvo55zxHGgWgZAMJukYgKJ/AfpdC
5v/TnS2b85qYDQTaLyxRH1bKU4QY2/sm1yRGDW4FHEAJswGbZjVkFZiSzqS53NHq6ta2R/XuolNn
6CcE+6DBTGp+97VK2HcarI0PhBwSRa9vsdqlU8LsP9sQowhZ6bvH7PReu5qzfKyVJVdSD4FwQ5RC
1fovcX7qbhh0fr6WqfyfQesVmWM/Zi0DYsuR+g9McQD8YSEs677CiS1Ju3dMeSM8NLRRB2rpfSwk
8+jWfwD45YnQsnNIaXe68zF/Rfr6LuE7OYT8vqcnFQH+xcRhkm713jdRzXPcoyqlrHRtVlGb1skj
zcISYkrz4GeS2YINmnHXCpXXryAFLWi9VWTkUG81l+w9JHWwFWIW9JuyztURrNtFk9rU7o7M3KiN
kR0ds9V7U217xTSPOfg9zOV9g0zoRUN7yzt6l3gGTImStsAuVEvgeDbcA0kXpbxzcDPUX44QLD6U
l0V9ih3B0EcOR8RZeJtkutjfIM3C4g1GyZub6324WXizgAfhnG/QejquT6ajqU4EzphS47opwp7o
PcvP1XCI4qpD6lPHkU6XvLpIdFcqKZ+z39hGOVi7w4i15kM1S/IFQAVDSo6AAiahD+aiXvUJTOyn
ZaxqRTUtdgt4YdRJmc4ZEKdNvPuthkUNMaBWLZ5ihJ5uocMGlukh4idtLfflLsJr9x+Tb4EmuAC5
Sl6qmNfvGnCwge/jUcClCv71X1z1R/lz0I9V5UkCwZSwVfwMBQ0nUybPbJPwMOo49ecC8ffQI/rU
qqbb1K1cVfLiDx8pFNyWvPWGBw2GnxP4Utw/xCSeoUBtdnPO4hdO9Jl45sUJpcNljTBXPyhr1FTg
axSeulTXQnEjktwXq8sw+LCWmn0rQ9cZUiLNNLvjL80pNgSX3SG+1sFbP4/z/5jVHrqe3YQdsM61
EAr/nks74WTr6TiubAvzollz4ZsfP5p3iB7qqY41GQWK5HnWlGqXYU451c0CWaT5rYHMLqmqWOT+
XI0+j/APnFu0DZoPuGZAU37RmamVJHtUfXhRE21E5cNyn4BzwoGLabNZ9aUCBdTwyZzHmQOp0/JN
+/nhEhuJlGVP54bSqbkQ6jRM8ZHUEgmNvIXO72nCLtjscw7BwQ/lD9ifx1VjF45tdJv/WQFG8V8P
6QNR7xtxZnHf78I97LCCNQljUGtynkIur6/476tKMyS2CYZkn+ulwgEa0rqP0SLv3npJbe3sOruQ
KWjxJQiycP2MapMMKiTDt92MM9iNe1ZFdwBuihAaiQeRKTAhS+qRMVfNcrGrGP/hTawdVb45K3y5
/c3dg/Jb4E+4msFOKGGh6jqZnTWzwHZChqwelOap5/uo36RWlpVhcTd0WoHls7+B9hYwQP/Sgf/U
K5Ka+SRIlbiSPlj7jWUp8mp4n3CP/E0Yy1PA6dnHVNLLaz89aCE1BQqntGf1ya2N0RmvAfbYynf9
ptkaur3qvQFhZ8uozq/JfWQZyAMcM3HvtrwGuAni/xal/n6ZO64NdhMMVm5JKmU74c77f2Q8T1zu
FTM5cU0hWt1iKY6rl+eyW62olKOc83Ti1aYVZF7E40p+VILg6vPC/FFowg0IAfcQHBkpC/dteM4Q
oWN/ypXSYJYumv2OppbMr14QM2TZbngjRsf+1X5RK0T3hZeKVjcVOiAlur/rDZ/Z51Hf0KgKlkrO
kk2KY9F/tECEszQQ+FOZhIdJYPDSSqlkLAka0q18onA4rROg6SWAqt3OSoE6xlRyB+IyGlCSk9jR
mNeF5LALZ0zwQRi9KaDeo6i/Lvc0tXbxWNrPMqi/kcqrA3DxURs1slbEeW2FfyhxesigtN8qfrn9
hZQWfBmMcErVhyCxrrDp3coVa4x8nOAe3Djdv8JiLz6pViYkM2qLD1QGVKHi2Yy9yAHqD0c+NNra
s6vs6AADUcAcEnHFtUSVJKpEh19wqRPLcbA9WbBYiZ9VzFt5pU0N/ATaWdW/PHZa6GRPlNNhkwSr
SNLtvwXVkawmAGJnguYHgiF4hrIi5C54wmp0WKHHIkpthWRaXc2SODd3hXjMtvr0ma0KlKwDuyzX
IZROLkTEskCQmPKDx51XW3SBvXiDVCISAcTceZSVRMModR71Vz7DGAfAb0hTuJR9wWi5L15efe4U
5FdEFlAg43d0eRrBBj8VSzgO3yTvL0QdZGs8a0TAaC9IShra4ZxBR+OtVnjY3yavQGhDfhVjZuAy
xlYjU3Sj61ucbK+ZvCWa0Y3kzPoqYFFA7KkGwH5nnPQVEycGAr224IoL94oL649+KaMQ9MQJg89E
tcxrx5+05sDaj5UQyhYX1ZSS5EEZrhghJ2f4LUQz0qDPI8YJVXWdkTCCuGuY6DnUtMcjfug+bPjp
MMNYTL9HDjVnrRVXjRi7bbeQ40uKhevvtJsazZAP+7j0xvqIHXWdRf7rqvw8Eta6dTZtErsMcrEZ
OdWBmycs44P5KkyIqeroilUz5JU1z9Uta+NePA3F1oK0rE4RlgIOdQAteV8XHy55w/8i9dq3mjP3
HZ9ckcLa7xrnyeI0Sck8/zRob1XhvkyoNn9FkJUafBL0vQJeWbfFpcSmNqoluYMWCsz16VhN1UMe
ofGYAPdyNkMNUWOJMDWesiB/DlFM/expzetkn+2JGM6RaiZSjzTe1ZXLKrdQj23GdxT2KZv/fB5D
paGVUi+/RREyfULI6zFWpIcRq2mrilgTxW+WMdAulyT/2o4RTCxqm7QxY9kGZolDCzQtxOjjiGQ0
AyjYDC68jADQvEjmwlac7yHOzwXDSyH/gyXmlLMPDs4IQ5l2HwJkoO1VeJgSzM6239/b3qI07Wre
csVOPw1D7EpzxEbFaRytoDtu9+2m3Q+gRcViJS0Yg7t99ZsBvddS7dnWMCeg6s8UPSeebthbNSUm
mslQ/Jy0M3QyD4hxmXk8GQv/nQA5ZEEIhczBaD9H6RfgjaHOMzzouDgluLncuXp8dLk5hAz8PdKC
GxPUhLGsLrqZN+0yONylzATJ4isUJ3zUa/sK8kW4D3TWhfqC7U57X/dEfAhCLzGdcLrJrn+w4u7s
rNwE+jj667cyx8pZEHfi0vCwuWBJvlT1KKU8ZoiiDYm3ZXtMkSTooX1i9d2np3BtcxfMcp0jNmCb
0jEFnqvjGIEuqB1Czri7165VY/IQ/NZYjwSI4qZA8CFs1XBbv0V6sggnz5gu3iqWuyLptsOijrkG
Q+lsmKgLe36VDJWY3FeDaxY5AdTWGOBUpdwS9bmEoAzfUefY/WDJWIq+P34p8Jksyr5fVrW8r3nc
ObSMemPYN3BDyuhWpRoasoTpptb6rg7ppt5ylhAecaZ7P8WEMUEGcE56ktKuBI7DCN3w5Pi5lw0M
Qra8Yrh4so+UJ39T1Hi/cf7TeH9ZhZ5pJrv+nGLxQqHbqVqjY26uMYa0kP4EG5Ewr9XwUQJBty80
PnjBJ/FdV03DF+dokir2MM//LVcr4FcaD6r6brkXX5llDuHwbmKrztjUzZsJT7wZo3NUij3Us1OC
ExFqHlFxfbjPCY38M2EoV5vd/0ChjdhwNlUwzPy64k4Brlt2EVkBiYuE1gRkbJbJgNGGzzY+d2bQ
/7WCvpSi+ANnaSKTXZ4N9ebjyrLXIL3UE0pQy/mmDN9tKeSaTsDVrzqz62jXogd2yULNQ+xRONvn
+Q4bi0liLMNSrbxjGyWDckMjHIkFHeNTRRKRUxVJo8CX8spkFNXrf+CL7kKo5G1hy5gJlNP9x2PM
9vNBgrSuMuhfA+vtBO8mJojhXdP0+FyVEwE1U4clOoQ9CGhamiQDqTKGvcP+khs7ZJLV/bpH8M8E
6B5PEj8VLXtgWyVBeIq+cgsGN7+Z00E60SpWd1jdoN6WGJsggh3tGDJigUHaE5db544mwhDr8fF7
h4I4RyXYEB3wlYKgtODdMD+7YWnwW7Xv905VpzuphJubn0YF1H8Gv5Mx1W9b/tTouWVZ+XZZzomW
qIYC+AbfEHFHPCuHCY9WppncwSVNOj9OU4p8BhdL/PFxmtH1Cq2jLps6KLfS1Jvm7ByfTHlFQIxE
PSF+3mg+adxAXv+LLrYUzpovs6sf4vs+DKl+7tBcq5wIWdLtSkPlUn/ZvQ8zbCBC9jZT9KCo19qe
kUw2jAaBo+/iWXdTx7wVYk2wT7hxf1XBzSgzNHynT45D/vWyH8ZlZYG18mW2z7ZOfe2+HvnOJTei
NuXE9wfPRCvr90b2VDI9PLfnF9mp3i7VhoW62eHbKyRaiqivGUBg6peuW1NNWlxQDQLnX+sCwRZl
QFQIroVESC0mkjy41PCTWeZc+oY3ZircXRdCK3/fDiWs4WFi1YiroieZtj0OCFXu8O6GZSqX/4gg
hnEiNmctcweIlb06rc9nzKN62/jx6eMXnA6EjiNmvS7GxZ2Pd3I++Cibk1v07NwFoDsbnWeC5zcq
sikiLtrsxWBBgwBddc6aOldgE+yYr1V/EnM6ues4Mko/4hSiJGtpsHIB1VfI6RIex1bqOtjz0+x4
USzmWuVHoY0m10MNEkRFn/CwMmpu0L+RaLaHLAlYQEjVC4/ng0n/3uTTIUHlQfn4njaY24RbP8Hy
zz/kz/fE8nhP6QsdKVw+ZalxJ918T7/J7bAVqC2XQi5EU6osQta9PFLdcRjzS/L1v7DMPNjsNwD9
6jNgnDi69prZUgMqgBSRMNQke6H81x4Vp0usAJFP1I+AAaIFgvTkpeV2bKskb9ihN9nzWez/jI1E
w8kfLQshvGDyCZFK88gkuqcH4cU0yHcToaoqsxawh9A8/MCChP2i/QResb3MxPpX27Erusm8H5kh
GMNj5JiuAlqWdhR6DBVQhfTGGkhIMrHk1d3qdP0sEOyF9wgi9h0sHo9bXAXNEX0tY/k8mGRMYBqc
wcsbkT+WikA2ktZAv2am+ZVrZ3AwwJkhQiUdVI33noL5sWe9s7dXuMVJf3rZJEK+5RWemJS3WAMw
KUGM1Uf18o8xdkaS3Gswm1ZW4eCePUI5oH0FIgiRUZn3oIulhL8haQ0KNRRwcwyVlZaUE8lwQLdx
jufToIxaQoULHPCbdzHIKYM7xMSGiPZvZv5tGGfZNpqjEDQFksPYjjLFuJze8KhAubVs2iGskN3z
5JA/XT7i8ZOLgWIHO+21dyQUXPDSChr/7ivlT6gXxEUJ+Nlht+7hbhqp4gdmnRy6rE/A4gUPwnPl
Kf53N25f8CH9M+HWvtuil9Alh+mx6nhOrTyiCRcmwAP/DqWwyCZkXoT8bijsw8NjriKH+YK0I2L2
MyAm9I4QoELKAaMjfHHyqiSHR+UKufv2ZTLXJ2cKN8hWjWlC+24X4vJQuTxOkbRY2Wc9jF7RK5hQ
C68CEWbuJPq4vDrjWyWoOkcZk/ndJ2TGUqBDFsW5GkmwDaIe7FZEEivQTOp2SQemFKTjXB+NH/8W
8XpapcRLmA4za+f3T8gfis+Ul0ivOC1YtVmRf9BkBMMPpiK3eQUQXQQAY1EgdfaRn4aCZ8w3eooI
ujH4vpdb7cicIbl5o3LBWp/DMlmU1+tewzJID8hmhPMx28srgju3njXbc0Q5C3Nv8ONwdB8uzIvI
ZlVguKBoYFGiMRQkXXyCP4YAStEn2hzvarfvFI1QlECexP4UO2TtIu21X3+vh5DgcHpXnMC8yiom
0XjCz1DLgYBuWxqDwfRjLJZf40drV+wuDMKThRccXLTHbe9wD4QvsTDcobwfX5V8UgUKOQr5MKPT
nLAoYrO+ukVaaoD1YQ7q2MB54CBQQXPoBWlKw9DAcF+etjdhsc70O7d/AfczwF6bOzJVG1qMdkps
z+zvYX0eCl3PIjgPMTd9mbbNAxdN81ZUqCJIkYLaAFDd3DjNB57BTr57YHpOWx9RbgQ7lZSQlyd7
yTnsYluLhvtEIQc0u2PRTa+RF39FTPhqnqOZE+woCLXI2w5JTJAHeIwNvzmnFGqsQR0md3IPEjJr
Lprpjqyw9Q5vCtQpCExWOBCIfeVNKmHiwxED/AnSp5URqh3wNqZ36gNuovYXW2dEqdLKRXZNwlED
wyDjepIlVR/Z5sW9xAkQ2X9YgZkS0c6grQ8FmsNchf9t/uyatIAYG+jkvis+jj07jJx9BU+m5VV+
6PODIdlehuhTKPlXgh7A+GIfj5GMxqmcMc5qxM4cfCebvQckUJGorBB0LhFDBcf5jAWKx+qem1ah
dQ3gs8ffKg3NNUAu5U2qLg6dqhMPb1TBnJ8vefBwPnDsYj1vch3dd28DsCa+jyazCLP0TftqG+eE
l0J/oHC2I9SAvPmm03nXS7ImdEqwKus+/jB0PFj9Vlp/lKDJFEEEq62t+13A3LQGWKpppR5xC3gZ
Xmwd9V8GIQ/tiAZwUHcQdpwVki1YnoZkByFmvjmVeTxg26PSdjlFuZ7D5Do/MTkx0N4vpe4o2UxH
cGuQyyOEp58u0cOP7wyUxfW2mUl98NBWt87HNbBVvCpNfRwnyh4fi51PWwWs0lPSMDzf28e3m46y
OYyNaKk6tvsek2XQej8WYYJ2XJF1esUed0hZrqjM1XZ2vnSigKl7vRzip/Ft6ToUUrYMSUxj1Mq5
pyfTYhZRYiBYxl/BxeYNX4Ypxxd2r1TE7XzmfuHcI+rGW2ZN2/x1ba+Ul0Xo/8/dN7q6+0q6jdks
Z4ksrU7K5coamXkFJU9h8RdiDUc+wIMcmmDfIkMDJ1V2cY88ASIbJWynfnSL6X66LiVBa1YQpE8S
9GMagql0RMWYnfxtYNOeoMotrnI82SYTaomrofaMBzNHXfn6YFrHbHbYeqaXsHXgq1mzEsL/nPXm
TN+3v1lk6XFhKC90/u45E9l1q8HDXzs2luet7tNMZ0UqxvmrM4ICDn/GYrWKsHTK5n+jc+ENoyv4
0feh5wXuCeuANK+w7sx78NYMdTpXZQnq86wqDGuMB2rOYGIxOHl8jOIQmQ3lqTU84kpr8Pk8rXjd
v24eN/1ZZbmrkmDs8nn5/+i4SYaR3bzTmYYGikFs6Ct27NngzCl/bSKU+M9GzE6iX1KccKlixJw+
mnZV4HoIJnzhdUXw1QdpUwupQsqUQ528/99Cr2dI0kgJQ/RuLLpbsTls5vl1jZEkbLd0vrnctbGA
uqoXhFs9r8Q2AoyOhQ8azxhfKE2AXWmdPlq+mG+7CElNHtxYW4ubmLD5Fhy9nD7svxbwBoqnybhx
yIp37C8t3zznTnj7vwhTCMxUNlCwtZgJC9tDOorPC8MO0WBHAlo1FqgTLIObSdc0t5DlBYC0qWIc
H23mXuEyYIiMghBCTcs8txSiDGP6bHBmd9J25UFhqoA35Dc3hR3wsRwLm+PrxJBqsFYVI9PcC/4U
qr81vbTaWo9OLSXYxmTBxy8D5XsbQ3l2e9aGOkNsH1xSs3UZd27oitS8jSnLXl+YTkjsCV3YgNa3
lNtiqvkmb6FJ0vN3RRL1IoOSQyD40NcNDDEZla1WazHX7KP9bJbmG/0FcELdsJPk+LZe1CKt1VgU
8bTym5suOLNDmBH/Rvzdmn8LeNoQc9/wyMnheAucIyfx2GoU0wy0IduPgyMsyJUNiqBR4sPyR6XU
PVTWsZQ3RtVzxDhoUTEF266hwTiu6ivioXDDEQS2bMeIFIZQOJMfmCUA+QrRMjqKdYmOrzToh9MR
D3OCAOhk09WnNEkgF8ngdxxPXFLkVeJYklmhANUB3z1RjKxnJKjuD/pMfVMPGTKm5/RSnj1FzRi7
52Edo3zndb4+rB5rvNFSyKO60tlSo7w1K9MsHTIPC6tl20cP2lsVdk7V/Q7T5A+DumpiheRCKLb4
J/9QATivaRitnJWLbbSchwJNK8ZjIhA1dZ+JjM+qb1u1b9bxo/QiSC+mEZNJbp7vGK/RuN3elrb2
vN7VZT7FkKW04a3QG1Pbg5LksuCGv+pBDno/Evjfu1uxRYn43r8jBQEDIWpPHcE77fTBVP/2JD7u
ZA3PMcOp7nWF5SZGzTxrbVN2tZ6IXo/XzO+GQz+iFqTjOZlAWKzPjyOy47M7ss9296nmjEuGhrXM
4wXSDORwZ52fJTJaVqI4NRidLzcgOCZbg0Id+s6SzRg4RIIs49K02H6+QNoHEd2uC1uf0j0B/qpL
o5Z/sL6bmw1XXMQKQzJliWsEt4lFYMrDn76bNSDaBmy0nN4MFkldwUOGKlrucfxZ9PkX7V10UhXm
UdDxSG+RWYoMRGITXc6qodAl/xuwCMv2WzY2viwew6TL8769cIJigqrHTaBevRDi89mY1+/QZna/
eOExmYdgPPJfjhaZwpzd5M82lmNJ/n7EZugIRtEAZOacdc7vC2LtKiRG74OAn0oY127dUFQWYHrz
JdBt+IBvvp8uPOMY8SEGiSMEcbCF5H8fcGhNPgzT92vhRJeEXRdYsmQ4xNSp7FwDRqrdjMJnYq5u
WjBLOHdooRsH2NW2tU1g+Dy+XSoqWmbVHj7Wj6KEYE+cQREFbfPwEI0lEgC3KAddCn3Bi7IthRud
S7CAQVeT/8DeDToyWE7cT2lHtttHQ9m7zMT2V6Fix69sanElJMSOeo6HAvEOgKFAnTGCtrRSGBoP
RXAmnF4etj71i8eikNsZiZOhYu8ijwsmeSZqjnzaUlNRks36sRGiQuWY0n+jNheYaXwg1rW4Qfq+
YvxYCR7royFODYAQ27nyc/sYnmVf8YoqTYgk8ULnRmghte1Q4xmgtHehRJXl9C2D9JdE/hVSg8Jp
508x2u/vp9KaCANQH8G9bJLBYzFNgEkxjgPdsEim7Yrq9JOZEHi9rJNuDGxQ1jk+6RTX4ViwLuXY
L7xnoBs1wFn7sAyA7jMEOpFiEhJrSLncMgGM9NchzFpZJ6BxS8ISsjMGC8iokEcE3aDLFQoNkNuP
WOXld0KcX/jva5espftiwmGmj0AlC44fv3hyo0cEIr1vKYode8NEXkZC7plBnQRBIop8ds5YY3YD
tf+8WOwFdFBZV2djJLdCYQFy7r4vBZxB+syJ+QxNUIcdm4zcJFEljn4CDI2OrZC1cdae9/GjHEaq
4K0XpJrHeqMJt9rgm7DjwBTa4rVC4xJYQvOAsaq6FYeXEjjV+sP5l9AswbnDuj0IlaxMeYosReC5
xPjHDv67H3FsveK7ai5bPAI1Pa9FfflXB1l4fD4D2B5uxou73fGHT0Ezs/dsEQf9b2bLnLPt1EOm
oRbpwl7n7nQOhAOLKDEUotjopybmgzO/AOO2t0+QIhUBKE5rqsLOf/2mv0Gfe2O2JgDdBonm9YoX
MQMW9U4jSYtWeAU6bFhKhdTaHrX2w05RfgZqngn9BWubw3Kal91LSJCGWbHILooB03f+Ysni+wlR
GppBANX+4TSTBKpxLL2Ai2dShwePdbne2tAutulDZ6qpCTTOmQHx0mqPNgAyz0jcBM15N/0GdLRi
cZuXBHyNk5B5/qNibvFTOP1Ys+Q672MhWZ7X0Ui7+XO2hjQn6aMsARF5nHYfxtYSl0uI2H6xLjSO
Pz2xcV+gNYeGKTvBDtl5v6pmiPQwBNYJKdt0ZkjVJSIup2I9QkFoYGNSe3Ul4HNaNbn3JU2dI9sp
0gSD6NVIdj81T/EDTIPWObSbQCZRMnATA20bvxs/MBSaCa+rMHkEqrmmvsSNRYvmX4/h5KlyOnHk
O8wilQO3i3xf8S1EyeFkYcFPyCFWsLLFgfYXO8dZrs33z4Oe36sxUpZDJn0eNjnwXCuGTJz9L8Bp
ppsVQMi+YYq9IcxZNB4Goyen+gBifXkX4qJicziHcjr+MZ2Ft5fCkvKwfcX6Jl3UneD3wNNYLkLZ
vG/5G0Dx8Z1g5OrdwtbgI7hTePj/VchYWBjvS/pncp8fFlR/tVI5+qlyM33ZYMR6xc6F4Xw8XSmy
HIdmSWN+m1CkeI9awHVrhBqERmRm8UpxJOpSeMP5bl42+JmhUI0DYCh5HhpitX4elrDwRBvtXQ3A
kcKYZhe5v3rIuEogQRRp3fRcypERItounf1Ai+pI7iSAND3kt4nzNpg6+nKVcSX4uL66zlkQlQLF
WCfXicJgC8oSlbiongJ7loF7ZE5tMsFyN3sktKC881BBiOTIfMjmcoSQIZo9JNsJ4jUo0wYmvfi8
AxKC5HhliPLHCiWh4iE6o/GdPYgjPC700SLXLR4rYId+FkndDGNn9kNEFHls3oxSoF8Y6NE+Ectw
2okIFMN8YRHp/5lXvOB0TDH8XwBFjO0ulvM1ADtB5QY44WLwX66BLRu8COIN8s1QapbTsn5OODph
Xv7m+wVJaBoQgcGhE1rknbQpN+KG/dcOuaiJDKNtexNiZ3Gbk2H9Q5smMkRYvtXepes5emfhfH1D
H8jpbk2JrgxptZvHE8bLQqZgMQM0xo/2Zan2ZNHhG5QXpK6BPRkj2rXKXIfzpE71o4AWKZnhLTil
xbZzBEaxdYJP/CcVAusEyzFWH0g47Cfn6pXkUu79bwEj/lfCB0h3B6GtXl3Tdcp2DLFxx5g5yBdm
6H2IDsU2PePBjl2w1LKGPxg1Va0aJoLiNkR3CehBLSst6J1GTjbZ1i1A+KAGEh73NEBGT4gpnukH
J+qi6pj0kWyGpWwXM9YJWfNloCyG29R3oEIslPEMLM4pi0wIqzSZPM9MC6EzVk4+70tigPMCZrEM
lzvL7VWzZai1EYgTF30q1WquoTs/BLP13KqmUWvGfYYDfua5VNiIEytWrMer0ef1oZMXlxCU2NTa
1ivNJKxq0lRybAzdudUI9HYlCQ/aXnP0KX7DyTLFGw1G5r3fuEMnFTTrVZGFI6oT2orcrrAuuQm/
AnnJtCgwzX+bE3o5yRtidOSI4DwvSKH3lsKfr0x/tYTSqhU83p+lkuDDUz9DO2sgPNZdYYt98WfK
lvAZty3dmrJ77ocOvjNr8l5mPFnoKs9vK6WAiAhA9z/ZSq3MDR7VMa6ys5rEqqhckIdvRubYbdqB
QkNlkyu/9oT/0IgTN1byhuexe1C5LKDO2oy/aSmU9xqNxmAzX4Ri1bxr+4vt3HAIG/nzcL+9yceI
Dy+E8XHPK5O8E4OmRJiZJf9GaY142UqukYLH2G+THeMaW4u9dHsjx06OdDK+grItEdWRe4GzYTCt
WNBL99CBqQhq84dgXmAjHymL1naAqBI/hdEQ4ioy/cehVGu4a281oRZ68B5Y1rgcOdLjT2chhR2w
gsKE0acQsVaLGDcGgOJl+wZX7QypOUrL8u4Qdvhhpe7zTItvOyRUQ6cK0xriXVA/QZKqH3V/zLYq
5nSOyNAgWxNAeP9z34sWpkZch/O6JBq6/5V2fJDFTotNG1kzZyCPfX5PiYpxS2w6H7xllSkIFwIf
TSxI094gEHlLCZkgA9+8isE7aocnjm/m/La4XtBA6CkXSDt4m1aFUZII6Qey0Vzs+Rus/RyrkLnX
aFJl//aEqTFqsFYMCky+evwZs7Xeo/1SwACYTELdlVCi+ZqCAR7sngI0xn0FynfCoXq+FGicxfCr
xK8F3HfwsNjiKusOaFbWH3v1dfe6sK+mDHaMM+f8Kq0vzX/9M/L9pqI1DL4HuIMOwYgkXt02L/ZI
J95Jxqp3bK6Hy3nYgF/0sAttSjlbFGO9wCc/ORdg/YoAi1cde/INNlg4iQH5a107C+a9DRqyPUJW
rSpH7IiKdu+qUjfl0SJWSHGSlOw/pvgBn16ItSOWyo8whbraP0io+GvLqgmaTabr25+qfuoXp5UK
PTHfJQ71wX6YlGAiFFYlnXGrpln7nz8o762cI3+JghCInOWC+PNUglUeHKwT11mqeki9sK4crRvj
yaX7xzjUP3Nux8GXwd0SBQlB2/2sakefyfJwUNPuzHvF5Ho5Xn28V3PcU/asD/IKeyRtURmc+tUC
L92G2lrX4/C9m8KMMS2fB9emSxh8D+dB1EpPRaseby11IYp+wZZ9qQX/ggU74dwD19hsoBV+kxtQ
VQASrVICc3buTRYD/aX/FYaeIKzpPDVoAYIusn61HJYNVCxtFWnun8OhN6t2EC3VR1Pv6zZyQMkr
rpEG68gfmfrBB8yhgl+OIK9xCv7XX3BRyXOBrAZg1iMxbsVjTgV9i0ABCf7kp89Lhq2GGfN5rat5
J95NWYynEqk1Zzcds0IXi0E+vd9vxRXARAgvGhHFt7iEmZTEiv2cuImMJkgNBRMWxfYvrU6nqkOa
46nIrNcWAFI0353nYc+adyWv4M9GSaE/ohqrYTxZ/3oCMm26fmUW8O1YiGizTloq/ISpp/htOmif
HjNjP3osIyfwOZaGZQGl9vR0JVY/+FjL8i986GlRM2+IstAoRK4oKdBH6FbdKlYj0yKeUsVMPvWY
5oSpaBdRBMG8xcKYa6j2Aa5XS3nuGikDB/0/2ozBJ/f+B+R40wtIZ3IGHHmXK6u03n2a2leoPPzw
lNzfkEC1E/+jxCnc3V2KZnnmxNYBoCJ7JPw4tvgZNUA/IZTloTbZXdjTvTazwG+WHIQ3ULBancfc
hIJrKnD49XsmLx+VIRaUh8+wTjg6h1HkzUy2SaqvPzyrahpt/2lxrANn+bBvGoo/r48g4ea5y7tQ
H3tnRp23p3WQ5FspRKaoK/aLPQ9ncGoBVR1qpYK4uwOQpxyMe7R2mAfS0AQtnEVev9NeYF/9JKOj
dwlA+rWSHYJAq5XAfANqjOKr4lwG1bdtQu+uvAoXm5/nKI0fOiKvau2q9fCVqyiwb3T9K82Sd7os
oeRabiICXSKoI4qof/32IZxuIXN6rUigmR7q8NIWyhq10tR615neOEZwoTsNHDx61kRi6QgZenID
0eMSWQL0iuqUmf5RP0s6PfVEVGcgj0d4npFiv2nfiycQEqSbyahXDuIZ4XQnJwXsgdagf+fhtnsi
emFAE5+NK/ovXiiq/6fqQceKAIE0mPYAVCYsjW9y7WVWLn4+emtoivDJ9n0SsJeAxcNhKtToj0+u
AA8fGgvs0CVi0Of1/4ICIHP7gH1STR+rCXKdWLgB8PTa2NnbPK0BM2w/hGcXkR7Oys51qRW4r3/E
Hhh2NBDNHIN73x5JLGJLJSYkt3MLsMCluvGlfqh4FQ1AySAOFB0PK+Eh8m0OWJZZSt1jqkDsyCuu
lZkv22CFkLBJ8CyyuhihcKzIK+8hL3h96PIx+98Q9wvXSLbvLE9qX4p311fLBOsfzcZvHShHwC1O
K3s5YMIsKnOQsJCRM5YAcI83+4WRJbVww8zLEMfyu8Wj6/bqzdTbN6TfyUlQqOo/4ThM4yjYjw6h
SRULBSXH/lKvmNP74JO/lPhMmCMZOU6aads0OY++Pvscjn8lv7OAyxb/yn06QZbhFGPMCTYiyQIZ
o5Lw4pvTNDp0mu7gZDvmICEcFnGaUVQ9wtzRXSuy0/X4W1j67GjyYh7koHDFWLEm4KLWA6B7xNRy
KNCcwcdeRSc705Jmgx1JyS+XAPC3soifRHr3e2FLkwyAgnjSwaH5RPBHMtRRfcyjLmaCmAIFN7H1
NnBuVspMTijsf39lpOQi7/3Py30NtVs34vcVIDKgrQzXFJsJy8YeBWHQltJpzLxpJ3+528+T7Ums
ZV2F/48LN8+CyiUiYUocwWEp/b0s7m5Lo6++JYGrRw6IkSao4wNzvrogPzZz35ktoaqW8gJgDM1B
DNNVWC5R2zHOBDVSgPxmOKQH25Ml8bmrItH41xAMPYhQS3UMO5Fn7Di7++9xIRh38PR1ijRJvXYR
9qr3bqNa3bq4GYVuLgBbJ83vb9Gx+d1HUJb2WKoTDnF3QVFBeiYz/h0sojoSj46Bmt1IGgpNoTK8
82rDklEzrD0SuyJzCp8isvaIJNQrQrXSjpGigPBamtNt2zgaMjnK907/Eefwx469oEQ4P1jgDIcg
Q4bZw6sOEr2qZtuRzEpSd7j1yRl0qhU0s9341oxXr4M3FTH7hrVfrx2XeT/2AfIHUPpUx0xxSL7x
AcfH6OmEokoWJPDEu3CbGwx1buPHBV2DskdmCDcDJJZ3zmIMEGWAMVqwZ3iMSkKrKOrekdbKrNzN
/uf42trtR4Ef2qVoprkZTnLWcofl32ra9Afwpq710GFkH+uWVRw8+3ig/1S6trBzU5CUrxUeUF8b
prv59eJu7YkpAyaoYHQ3f6dZGHxpp1CK8b81Am5ZaPTRBLbYajHvBIymaWnnAz2q7yelT4hG4xur
ItUy5UqVVGdU40oePQq6Fol4IVVvrWVnZqYD41SjQWCA+eSBIxe5fGM1S5EaZpC9zjc3Bi3vAwNa
aFQWRlgHydFbJHa4ZeqcxRqVsWEX/8BjU1QQDW9jR+els4xI04ucNDiIRYXATXCH7uIhqsWlh6Q9
H7JbF3TtBZpuY3uxq9lbwnC22DedwyL6l6HX5cor/5HJ7TgWss89sgF+a3z+UzOc/JlPYFr1lTl7
4MKKiHYBvEP0PuGMPGXKDpHuxFS8efK2dQpgGkE7wLXRf1zketfkdbdzmbgMNEDV6yfol9Gni1iK
9rZ9tlK6wVw5IEjYD63WKCEt/7WbwdOUmduFH6HhcDln8Jf5y5GYuXC+MWQj1PvaqXwJb7YbPzc3
l0KYalmIG6MU1bfkAHGYoxcQXEq/4xXPszG8tBwPFGFUOcVBO0PFNmAFyXQG6ypv2Uabw5Eb9BTn
3zyMsi/+/F/mAsIz1pA+wWYPFJsn5eDyHANR9Hd2JbCUEC0S2eVZYzrkuu+mnqhwXuI5VIknKzXg
vK5ctV35CBp2lSPUJ1QxCYO6dP5Zmi01FX2j4Ou/rOMyhlogFI/UofU1r7eIRXQDxzu43tlSwiO6
eOqpopiB9IYffzbrtPHo/DDmhD32AavDbnr/Rr3Lh5Aa4YEFffn+ctU8Ox/25kPKjkzeEH4Mbi35
Fn+b+CQKIWr+3Bk46qbWZh9hYMyovIaQPqdHd4jOsPXS6xsIankAKix6TPGv+lVgNwY81Qep3Jpq
jVvYRmiURZWDyohjROPSqkel0uYhu41kOEIjK5yGb3OgJZRPRgAovCuKG/AfQ4HG89UskiDLnvhb
9c4lXk5InUMOI2XQnmde3gEX8Q337PGO0l0mD0zyH3BxNFLNu8nC4l8AqfULrQOIEKlpPzc2EHqu
ioXnebjqgku3fMUHAkTuMCgCQKLvd4MkI9qM7ToZPTgnWWNoq13JAbPI0ATqa65G4XHuVQvmQ3Hf
K5xl5TTcnrqyrpv4KWyRkA47sZBgsPv+EHYbkZezedOhxjO+s1qSKzQ0K2kFHfPe6Y5Tpn6ARRBR
BYtMlySxjPQUgd2KSo/w8pEHxX/eVXzws8SCHh6Fe2shYErSL3o5hJlrukH3VHLNnHmlqKAmtpcB
0KOQ5CvuR7L7csUcNYWVcoMHZGO49bWL0Mp493mcUxl+mm8uOASWGCteqGpaQMhhVbrukpKQnpno
Tqj5+gEpt6zAOF80xNDfhUjvkoPqEYNTwzFafgLhgjaoqTBfLR338Q3EwNq5/VE5+s1uz56q9dyC
j4I5kko6MAkDLP3GWY6RhmxFZiTUjd7nOiem/rVhUjQcl9KToqyouAvQVU+aGbe2k/eg0bbObstw
BBzpNH8B3KFHKeX1nKyS4YX8F0256ZbXVVwJNYNNiqM2159uqbpDHYgFv3J9DkhcGyMxkS4wxSdR
0z138oH7IvqMFAFsnxahoHYbzUx+JSiUYCZAKWD+hKyzGrghOH7mH2bP4pgNE8+QPhirVXcbXcft
jwRmxYw9VAp41P1c4+pOAt1tvF8ZiZ+uGkoS0WO/5rRWy+6aZrczIvpoYltosP6PKe802TvdipIN
H1Bssqdx/HyoMNqH7T3fZYvLqNubKKVSF4CmsCFBl2uAsJf3Cfew/S0HLJ7kP2SQiKP1299lTzMA
LWWnvceRdpb0L6oHj/dtOgHYU/AP355z+nuJci/YFyWNftdF9zZHfy+MklGrXqnabQfRDWoqgL9x
V136d76xzaeD02AZ5WzBjNbLk0rs8xI+iIZm5zkTbFRQGiRLN19SkOFy29UFxIkSqikfa3vsCs42
Ws07WRupqoPCl6gI5iHrLeAn8GaqxL5YYT6ZO1JujnzLKYYxpkoGKyMCMSOPpsMMI1ej9kY6EFAi
3Yzx9/xVryy3m9//bJ5IhDJ5hUAHueOSfnCQn6w9dF4A1LxZYu3Y+/Luun7AZHwuA2lnaV0GPvIq
L9PNQMJHVAm3LqTkclQQImkYIIbO28Rq2Zcv0EFzwKkTXqaykY7SQLsBkUeOlBr3/36f+faQ96/c
US6FXLefUkYp9XaCz8O9HZTqGN2gN/ptpQtynBGYYP3zwnuTVs28G9t10GKaIeVrzGAeKCT8Cn9p
rE21MQ6D3hLG/Uj1IY7GYhEs3GDVcf8u/JKEFlrz5Mf9o2s3pEjozeAzGg5hmmxGKgTvxOjRUXP2
4J3K4QbcQ6RTkYESHfW4Hld2ofjNMTgDIXsJkN7eFq+6ggdADFAbPfAxTn7M7a5M3hZUIZFF82rG
s6seaQUd2wLB64OV3tZSQsmyCXXmGF2zOV2j+uL6+ugJpyzpuE7MaTCwmoRS96hFNrmB8DluI8H3
q+y5wLfwU+4+qunoWTfqf/6bT+LGZIFq9RjYPHTofKdhIhTV0h0VoLnGCcTCuim/e+280jjmuBO+
XVGP0u95azHOLiC6F54hRqRfd4m2SZdnraP77klzU+FwOU6O34H5k+6aUFle4ynSmxcBi37N1wPN
3Pi8jRe5FWQrG4ellQ/SSLgX9QwhUrrwnu9LjShFBU53WxeicMURa7c5Z4N+K/pcgu5ZPcGA50tm
xEozocsEEbPX5qitfi7Z0FPgr0FaAfujFBLP22MU16AgX171pSVEK90bZknlC9REcMQmvxojejyO
OQ6csu4yRrhTn5EXahLKqXs8XgEIb4EkzIq25o5g3oSPe9eDOnCr39/TFbuf8gF2ATv1P59KjS68
QOfi8rDhrPBllhw3EM4i8B67UDUmlEmSluOFsz2vMAPQW1QpPpjG2rwV83ZWX7JZi2ituwFuZ8pd
QSJ7T0nae46phhMh1sTOb1S63FrRAoWDPmGB07j7Y/8tpdhQ4LSG38OHMNiNohvHUGGWfV81/Q6/
a0myW8GUTcp2/jlzOiCmmsre+9c3iSrqxsbOj/jdZSRw7dca99P0JQ+GShFoImtr8rUHdyKW+dWY
TJdImCboa3vIrBkHM7B/tC/H652ni7vpAZhQDmwcpdjKQiDcfIvDBnoLQExM9kP66rjIdw+GbS0p
GaI6uWlxLuWAbjSEVTF0wkp0yZ+jejVR7xy7LLwGh7Teip0p05K2ZSFX2dQunOv4vOHi53jF05e+
+yG367Iw+AQdxaBetNh5RjvE/SAFZeTvpvQF9Dd/PpCKAsyhD/R9c/tgEmfNjQRrHd6dkMjSfAec
RHg6g1uaVONDwgVInr14bEMcCWxBijBYts5swcA/7xllgfan/vftYRehaz6ZMXcCjQzztDFlK3+A
yoATidPEbbaBXPnGxbEdETqHJllRmY03EtwYy0AiXRHND0rOf4MoAVrNWCn2WCJInHvHs5hFqDMF
/USNx/rz4OoDiEeWdik++LnR7UyW1VpZnr+5QjPTPXBO9eOIY5y129bG42Jfo4It6qYoPit1DLT/
RWSeQZaLU2yJ2mmPhn/040JrQ9c1oOMC5tZf3jm66aKWDZNg0hMCLqnz5DmXSTtFTYbvotItexfx
Qi9oG2VD5eFRM0nm9NIZhnx6OjJ/TodLggKMUIBvnJqwAeIUDKtgh+2UTsgfMVCTc3lxevXUvOwd
G0/qCF3u+KSs8/I8anN5a0gC7SKJyWgPyUEbq+TiZMIcHPwL7CaVwS8Aezqlf47Xv35NI4OS5Zyz
3ZelRcfvevIckNmHyR8GghMLoD4/dNyn/QMMHwr0EnfIbiKSGohVyIXGbnt/CdFlI9pVApjOeJjP
A5I1m5g96SLY8n38yWpwmTNlWrUNHEOouXJZdKUYCz+T1kzusLlqLmoDLJYFcxKm5nxP1njemwOl
G7kRn5aAJCuRERhKgS5cKzja8NY8PCD8dC1sSHuInHlhek+b+TeVPVDEnrm8ndCWWwSIP6E3gphO
6GMAtzZynxUfCxLtVR1D/+P0fJetbUUJillCr0/pVxKzKORhsbHIWcDgD/ZxXoYiJ2Vzk2hiY8lm
LLOSqFkHiBhGkWfFfCbk9eLEAkvk+gW6ZMBwgtccgc7390DiSFc9dMq6aIQWPBgwvLURtIVogM7W
yuLYVCAkmCIF+eQME3QR7HFbZEiO7PTM01FCj2+nyBIHBe4QQSQWXXmDvc6FeZ4lq4uVLzmmuWdl
SZaEcmu5eDFseOu0DJ8xi2KK6OBv/P9aeT54towmGtyQonLtdoVGDrUmfe7QhoHqtlPAwXC4/8Wf
SmNC9vcs0cdGmDepWzNEmgffhsSE5vrv3k0zqsqCl9ckbUGtgnM+YNzqv2rKUKIk6u5z3AiGgRS5
2lw0jxmK6JxKOqr84VxBBCD1wOF/kwKzF9QJNLBcnJ0bkssUp2mmEbUtlN4tIUFE/H84+jnQyPaF
R31UQ+iYgVpyMlwoWz7CVPFI+2F/FeLce3quZdZd93/qtRRXBk5vs6saQepUsfIIAH6CT6bx5hHI
Rp7n6LAbqVQNX9JQlRUy7i74AYeTbzJ+wnfXJDhMFTFwh21kXg4cGSk0YmFwkvRQjiGmLIC9Qxjr
1YGyfrWp94fcZFkC39qnADqTLITvFUTvW6KaQdaPTlD9DiHe3HhKO9Do6vn7TpRYPIoCJ24V4Gdu
bE07GghxQ4BC8ZrGXVMI0MW9YoY3YDcn0CM7+DxYypbGvxI+AGafkGJq96MrP/unzPj+Qy+n6QI4
IBj2N6rJvJBGazogRG7NbnFcTTLKtifnNxy3CaoxrmYaV7O2JxHfQBlpeiQo9cd4mFL36kTu8v5G
tFulf6lfQRDqxhxEdfXy9wPnrQqeE7PuoSCC34qYVjG815oBsBD8CBeoFVJgDd1HQLfEMWt3BY7H
JB8s97uqIaMtcd3rUiPYuEyD6Aao/VB8+5xoNPoZlsffbqgEwIzL6e9TK+d2pGEB3U3jLe0qK/6M
YVtGqvFMJZO0T8ZmMKAHnnQFnZqP+/IDaISI8zXOpwYYwHshSwHFf85LCSjPi1SFr6XzqzDIBQ9A
7jtwgE22JOBaT0Ls3RyRHt1L8FpqyGAwddpn+V8L/fQo+789J4SClxGMOd1iYEyrI/18edzH9O10
cLlFBXqJqgwySvvZoW6TjuJtR7QTHzXvWpTgwddMgMF1UOP5V2jWznTn1M9cc/jVpKeBxPFdGN1N
tB0myYI9ScaCxw2yvyd7odgHXDeCJ8maub7eZF6W3k00akmdR1dzcFkE14P/IPfgnQY+swu9kyaT
EZS/YDMDtMIn5RZ9ZzeQLvBV8URk8AX/y04CHR7HlFSYb5WH2wXBpwORqkG6hm8oG1KsVyiLLAQx
+ZHf+t5sr27grWHS7eLHyl6nxBHG13CqbdN92M6yzAkobsVIKp6da2DBBLO4YwzZJVUAYDoyci3s
yTApPqCYvsyvEyxEaAFjTniowAjsbRRjBJrW+aUL0CPcYXKRfGJPuX709BnzXgyyZeAn2updr/lX
h0E2XHKKPo3jV7ZCDl+6teKZV2RoDogV56sOL995jrDc78xO+Iitylj1kdIgq9Rr1Oq/XrC7N+G2
wjlrNFgm/AUtcc4dDJeQ+w4FL18XUwISJzUNwyLkqH8HNLs/M6acZgCpa4FDy3xjTdEomfr8bgnv
ZICpDYbBHRMnXu4Klbwoduz/OA6IbXjaP4JmjKmiCQ+q7ka62FZGgvIB44UnB7qy7cPxBt68IdJ6
9LbjAc8OlavVcUOa0cPb2OcM/1vG+P1jXvRVLr+K1oxtCaCAxCaGdgV1thlukZm8LzMC0PS5wxvv
y9S4npLma8zHw3yvVQPgPtXBvcYd1aEBsvmqNH0F3w3qusybC90Nin1+q3to8kjrQPHQ3e6+5HoE
XlyCHVAvOUA6zgLf3YkMaKFC6o+S0Oc0YQyLIHbFg6vaFioirZlhAbU0gBeq/dDYPNvo/ieolg2j
yxGzG7tUs9RRJYfB6fEx8Xn08Y7giy3zP/EaBmQ7s1kPY0RsZECZma67yd3KnafjPAVSSm2cNv8q
3h5WLxXW/007+n9CCv9oF+jypG/A3BRQ7d1mIRLeJze2cKTaVYAVKHUo01uKf4lBd3a0eLybWjOI
zUlLX4X73/whK9RxSdv2sICFbp7GZN/2IclUwVziLskz259t0HTCPT/hpCMTZpGCALSqGcpAILRI
U/IBwH6cM9alXKGvTyM0v1chBsQaY1cBcslqzkiJhWJzM0KyEqQz8gU95AB9RDgSJTI1QD0iartw
7UghEl6D7/76neUsFhKVReoS1hgBSmx40AhyjRt7n43bEExu1jqVqD2F06cdF2QuJYo57d2sjDCZ
JtPp6um7zKZ7PO9v10HgQ1lhBKGtNti0hy4OTRGBKfuVz6Th1Ca2RkOCQCw964EhUnLOa+4MLHdj
ndyxONqttfmotkugoME5MN/SX6KZbtoAEu7cgdrhJyiVMpujKVPfndMfx+QifC19kE0pvb6VjZ2n
2+5g6tmnRJyLlm3kTr8EYtmIiSJDBu0g+atTJRMcJC91SVcqB2HUpikdcP3nq0iRy0wA84nSdU+E
9ufoeVphxjjv8PhgG/TUX3umB51Nr8o+yVdGLRxgaxp0Lr+nUhjy8QNdcGgYS3olslu6B1gujGAE
BuY5uNDn436UxjE0Hd37rWCtXmDh3WeekxXaMgx+mEZxi2UaJZ8ZLGmW4z6347dnQ9sEaDaAnr9t
m/7jK8bwCrAdou8PgM7M+qL+fkwKtc1c6cM1j6fzUyHwfe2+PNX4DSilfqiW2HWaEq0FSOZ2zgX7
S2vk+BUL0zvdNRs0WiKx4rX0xa9GNVAskidU90Np0bQkoGCq68GZ5YQtuKjIhqyYzdEr/23Nbotg
Nkx1LO3Wxnn/3aXU0DzCMmrJHc5nRHU5gzhzMDX4THb6W6c5cgc6OC8YrneR8mX384ObRKHNMV/S
VryA6ADQ3yosPlO63fQJ4vFuvK1MT6sBvhx+NBW5aZRxjcldByNUq2frpwi+vnc5J28w9kCBqVcY
BCMdcO7j6/9t8OUJkeWpSDfYfSu9OXM9h97dQkLePdlGM4JlOPH6lK8cyu8+VgVSl9vpyKtt81nE
XscrAOC6oe7S//L5nVJwCAgb68H7eUzOckenhvu/NvTzHenEeDysy92PlZ5WeU1qa4x9J3pdNe6+
RChb/Rb6ed8cGxWa4VpamvLMHAzfC8qOx4GlXAe/3UR5bTtb/xrfenzM29El2wCtoB7fXJun6Xac
3mqtLzX1ZfZa1b5KZUp71G4HNcY8Kxsn1pNPWGHUokJWEpc2F0XfgNev5TMFQzVJstPuY4VtYNUi
sli95YYbOEXFGYONTRm1lNJdLOn9XNGO5c9/WUgtEJ1Y0kRMr2pilRp/G0MMpD3z1CgR37pEGepv
Pgz0bT9eEAkLTPKvTT3YKA6JFt9FDh4rQB82nv/1vB52pmNeCx5dIfHZb3nQUpFHjL4VvmwPGHqs
Vm80rUOtbhxmJvbneoiJoGZlc30Bu56EGm5vUYP7FiRAz1H8utx1NHAhiOxW7aU6ROk6ytYZkzuW
1Bfye+Fvy6Km7LivVdt2RQaqBgigSwiIrWWa1axQHt8cfPV1fATXLriVJSqA6kdYOaK7talZMjFF
8SpEDvI9gbmfVSLP9Bj1ZHc/WWyEjIi6NXugnpyOHDBGXY6De+2kKQq4DJw3b5ljhyxKtVyxkuyP
B7gcLinz1/gSAc0YaGJZFN0d5z6Eqi4EdPl0jXCaqp+bsAxgVQwsJscNoPOLXqzrKNTY4/q6i4tA
eUkwS78qYlCcwUBaCs6SIIcXwy1tySQtWhoL/yvprde/BokGkZtp2+JqU6u/Mo2K2ualM9yl3o9f
xHawFNaexlCAX9+1dJuSw6ro+I3mG+Tw3udFLtJ5MUNphLc1eYoUs84H3JyYdolBZNCktkix9zMZ
dY1zD8rnSMRTp+uaewjbiLJLqud8LKsl9FWxlfmlOh2wtI88QUC+SI0Byut/IxIhIeK6XY3Oer5O
gZOJJ+mhS4KOfEHqEtGDjcav/uSRENO6Lw0xvnir0eoZZFf6GIitJB6A3ekcLiDbXTt9htcWogfo
XhH2i3j8NwepsZrEyXqyCYmgee+J8kx0qspUZ3kx/idZy4a1VyuGPS7vuloSKK8Aa48DOsTq9Eqw
Isp+bJLDhf2SNOe1P4Fh65+69tbqHvqBnva3Ssem8qspttW/FjXoZ3VXStfv0IZP3AedNEmAOEbO
T0+yFy08H1Wmv0s3jIHlPkAHot0xWKNBzqsijIz9wrcE5wQ6/zRWxQskHkriDPtzzy01Hw30fUuh
1QbUtUO7Sqp/eCqLB8R/9owW9m3B9cnptibjS2WVLTLB+ier7cfL0XQc3tEykkLd1geZJjMM/PVL
k5v+ws7O3Bwh4DBpV2gAoJPbDDY3KmgXVmNP+9mDHESwBU8Tnj7eXDCq8OKRQP0vpuYCU/AoOdUL
J0wsfjO6Lz40rT6Zltl60e8s1ADkS1H+781rxHFzWY0m2zoHzqJBpidVUJhBXSOcDXZbY2ryR+KK
qbYuMLUZ8mtKDngEwUjQCId/BvhCxcZAN+43xHLFogGRbRriZUpSaq6Pefg7uiZraudUKF/iC+HN
qowW5J8RjOyktM4E0x8YWvA5sokCpaEkDuOvMs9KWHpvv1EvBdrrs3kQohr/jGTsJgloggJAORCS
jmjPG7SOKEAMJoCMcUnuYNRLxD/3z2PxJcKN2r4zto+LEdR34587Fczz57/uvfhdfaajnn8PLfsw
WS13YfYUzRyBRvdu6sraBCjTl+Z1dttv2HAfms+ZlbFGhw0Q7hcpxqdYYlhevAnXuxnqGJqj7IYT
OiZXTWYvP//W32JlKv0vM6sYTnUkjHxjjZ7bJWqbeEvOiwN1M0OYOOPtoAhAu10P7+/P87Avcljf
0FoPnA9IOAOp2v8wfLdT6XpyyBhOQIVPSZRefPbMor9/XQ+4aaIpo1RCETxWWoDN+yZy5bH9ald5
nORPEZLxSGLd3Tp7cuSAPVzjkD4ZL3TEGgibPL6u77QYZw0ahwOeXW6qX/wQ8Hk/Ptlr4bpbCy1A
JamDA+oQR3eBI8tscskHMU7M4CDJlyPe8b2ct6yow3fSqPgj1a4cTPt7zJAFYmnTo/agO/2C9Zcb
HQ5vQiJet7LP1Q+pqjJqvrMOSxKYcawwzg//CtLFeFGiA/qV8TPC0nhz+hhg5QbNmfYwJF4DP10U
xjfTder3iIyPvyyGJbp/P1bcY2yup6op1d0vrfY7KAgLmLyGfWT/GGNLoUYldRYgD8bPKZlJsqKy
TAiqc6D9wsl5olbOM0PBtwCuk5sjeODEb4TSc/AVBlqyLVJbQHAg7DhO0N2co70pdT7MJZd033xw
LF3gEGXi+osPSUFu8FMnyJpSJ36uI//IaixO0Ad3HcCdo2l8H8cquisJK50zg2+FeTTjDAcwxB47
Nu7uSVMvrVlM68czaKXiJRNnBpUMPQfwdeiQdJkCv3ruzoH4YxCtDWMGG1Ztqng66Hd0/SIDqKBi
dIo3l07OMlssnpQGaNxEdkz2fMk1PdVDEkdzkpBLw9uwhVEQKe8wLjYA+4nf2JIQs/6BJ+m7ihS5
wzJwrPSc4TmRhulT9P2NqBj/5x7unfsZ3U5zbk/k0lUR5GBmYwbNy2kCTIjU8gm3tLOHdRK3unpr
+jGJal+tMg3Qv8xCZBT3tVzQwh0z4GrFjuDTX5BbIh7i7pprwqWvMSwQ+VGORfSG4NShZzPeQtd3
fPbLgo+E1R40ghNHjkq4f5rT+ASKm+Ql/Tq11MELdgFWDkDXLvY9KvN11fGRKce5FVV2u/VobwwZ
iCYESHY7gYin5MvjPyX/bcY3WdiMHCIVxd7RhLsjPVkRGTGwYPwkYFyEYTpMj0tBIIO2oZM9cjZ/
DMeXK3ZketxFVsKxIPfHMy9l2q/FEbAd9KFLsa0F2IhEhiflGSFPlEQZprXHwvB0oPyBLXVidYbs
9dGulWDHEdJrLDsU7MFf3rYlIB/ZRUU3AtGnavtZ4m7/QX08DImTlOEzWRLlujfKzXkYTrJi3ycZ
TfOc6o9tNz+lM3586oKgWj11fHjCEzfElAgsAq2xzXrivNncqyuqFSrL6p9F4bIrIkgsbpNIAtgy
rfQHknH7UL91ZBXtiFyZ77GlCS4FxxQAkNCrcxTblFEHxkDn2Uc6rlGAU5B7GNbPsz1/XWwLaMWV
McAPLmpSBMnqZRiOtuKcjnHekurGyGuudYil2JRsYnZeeCQCWdR0FY2FSyLxi5oimPjM3OeXyjn5
lsv4uFI0WSwE31KhLWmhYJuPNhKLjcJJBv6z0Wtwr3U4DYQ6zpg+Rttc9sy118l3SgAPaATcpoEI
3eizpbcv7T4vr0QUVGLr/8lMUmKsCeOWUIkp6jgfd4mamvvctGbkZFwuW9/sa9xWh7QIaeq41NVJ
Sg0SmOOIZwuRcIohED0N8YCwTJszI4CD2NfoABsoT3956xl+s34HL9xMoYA1kVhyBtgGcKfBRmpJ
a+AgYsGMbEYWs9bExPq8gelYGm0kHZZ6ijOwtMkJ1P0qUVkF5nFaqbYcLVFr6NJaexxx4494FXSa
/SxGB42gvJiWn1Z5a1kEPOQtGkgDWqBTWzL8otYAUX6NwO+6Bbx4RrJWD56+8ZFaHJP8PUgUkgiG
ESWKuewGpTqbKjgUD1gGUYuNBFc5n1IfcrkDbt3Ctq8b7cr/owsTIkRf8hMAVq06OnuI6MX6ghvO
ZdVXhvXzXeXYaaJ6DhH8mDrHQUfjuG3XuP647+npNtSbV72VaFcFmLHcs0ctBduMkdgOOv9TvYHz
GG27jL2pJQ+2vuXZdDEygxU7FolOHuSO5J6UP71xvKz2kScyfdmv5LuDIYcULZzmKD2BLH93lHHC
wPVs1wFzeFjtL7/duaJPiOVJbqCqKlb8EBLpSOGR420X7TU4nFcepeBaqIwS6vMraqZE0xYiegav
WMs6CeNjALlr9s4agOXeaTvTTEaGcBoEqddP1MNfy/WtfzpKjBrsx5+iXYa/ay3wWRvhMHUOPkIo
Y3AeDcLsRjaedkA1sf80wXcgFyGMYchWGQbVQ8T30BxTQPCYuhZ/VrP65h3MHTsGFcYKsWhp0M46
v9DIR1GjTn/fi+9msvu1klXYfBMHji5SLC4b4x4Goc/u4fVIo4ePFg5FiTOoB1Lrff68rE1pMGU7
8ZKub0NB+fOFD/zotcl07133nPdFUquCYzZw0xSVDva2+dEJRjq43B200kIhseY673vzHZ8KfVSn
jSJC0LRUEvs5ZuMGtlIrcrfU7V5daz4vuNXY8XNS8Xo+Z3INAI7I6gRDn9t1bPJtLWLxndYDqY0W
LmoY6Y8a8AcFgoM1gBZD+XWKoqBc6gBavOEa7zncpa+NsaV6O91OeAjRyGuisNoljq8EaBSa2PK7
TTH0BsqyHsHn5oZCALVZE4yLi6YWBBLpTOElr6Y5j1eA5ug5jO+2W3dsgMGCN0jyPjcPomSY1s/q
oQWOjt5YhLwo0ZhVI+kNkXdldj6LVPnoSrJlrZoD5nNRt/gUdfFTK41pQ/Z6cEBFkwaiGX+X9OSC
3UtMx5/0/r8XX5mLCIEA4ZSbVauEePcvaEk0TfdWgFIOctrzwp5wVRbP0VR9nZIXoilqDHuf10XT
ynzCmyWKFLCJPmkC74/KhW5ueYvJiJscSURPI719k/5R0y2ztqh0gKutuynKzFotEdaKXImXjRO5
rtXXcXev3P7iJWyAXqhIo8ZP6d9h+kJfD8tlEl8VKAFwI0YeYlZXYI9HmfIrjJVqd+ohccd4TlAx
X+eNQQ6m8gGRMvraJFDG+E7tt9hP0ynRUhRBqtGtGXzjaa+KtCEQL5qLkA6KmEuRN3ljP8k6LsDO
/VrQ8YaPDDKcjl4jaCZFfAIPs/JZn3KWv47IHp8M/6JyAS0ZaLBYf8Qin/xarIR0Z2Ua5U6Qoyc7
hbNMtmX5CJ2q1vG6mZENfl2sICUHLkb0tv7xhT/9Kd9AjPrllHYtBSOLABWVZcWZG6Mqs5umxIaE
KXfhTZlbTFZaFS4wYBPS5FhTncOVlWIUFK+ybMjVSSqs9iqToAbP1qcjUWTyvOrlsTp706YkVnLm
74ya1AauoDZ4LmSQOMcgpNmTyIgQ87y3rsrRSxSWVLLpAEzrP3Ypc5iKAdkVboNh0r0+4Q6B0TTD
e3foVaU/yFcfRDT0T1966UTjJlFYo1V5piUnYvGJLFNmaSUO+Rcs3WZEcsVc2i+o/EtcRMJLLRFW
N8cnStrSke3yltWNx1bHkqqCZp0/73nJocXvoqh2tcvl5xh3hZkbns6DLxURAKAb1MN5GvwHrUef
4znAWvdGiHPLtOoNl2RxX4xqdsY/wQU6/tdQADG379R1nRO+5Kn8jsxNEKq9kZn3oOadAK0ePRoX
K3EHXmcPvBa4PaugYuIPJ7ZIS+uDrr1fxqOXIFK37gCuxOV3WvgMwaVoeoDmG8jTbDfCOPZ7Un1j
NLkD+mgp4y1KeYqemNJ2f9DY3TyFh8oUipzjLJWst4mo5hK2LRrx5541pU7kBFxnIOJBRgv/nCMu
flB6Bu8/s9ClD7chLm3hs4f47Lwcr/7/FWAI8psStyeDhxyVbimeOkDj6VG0BG9RKRQL5dBhfkRn
H0Yeab51z2e5dF5L+8dpR3rZaj3IWbGgG3rSrY5Ru65bEjoAFoZljX2Wyt+v5mLk9kaJBhClSooI
lPh085V37H+uDcG1aqB5dcC/2ohZlD6ES6N/As2QwJV5Ln/gtfjqSnqtHBXH8/tmo+czhlr5aw4f
ClF8l2u/rr44fonLxuHZ+n3Huagi+Zky5GRum7fXFXbJw4lre6e6UrfR1e3nUgyZs2zwfHjr0SnP
U1lY+Ae1otHurjomqmWw8iDt5jSlfRbn59WrNU33eR1rVwFS0cIAf/Nu7ZHeymC/18Fy0hQQPNrx
uOWb0UljS0w78UhSjrnqIBKyjUanyZBdH8MG/yAoz5h+plNYJSFGQg1yDtEwfzK/fP4Uix06Z2He
6nWmzeVk88mgqJOsmsbfRzCkXj5WfaXleJHo/RaOyiYpvX/a9ufDF1l12UTTY+EGUZGfcZiP1t+3
rbwZ+PiOQPIbXzDT+Gz0eX+ECDJTP5ebefJZ2pjaLYP4MmTLxa9ywA5a705yOntDIqsUEVVZ0FoP
UHfS/WyntWt1j/E16rA8QdNAAZUZAmSDVvdJgzr7RB+DooH2ITbxxaK/kh12JNkqMH8Vi+7thM1F
a53ik9cNKMWAOyE59F9FHMhlQddMfMJm1Z8Lu7KPB5arhXL23a1gZAgF+FiceC7Iz0MKWpnGOv9e
YM6YmRa6r0tJO4MdBcBX2qo2FNFpmImfJRSkCnc5T27bZz6+jVqAjx9xAC12Gjk/ikPKEVT/exAg
KxJ7+siI7kwCL9TYBrXVw6gqsXwlYbSdR/PDqXYPq165SMfSAGW0BrbgwnoTVXUivE4gEN6Ian2o
fBmgGzh9rO2Bfy8y6WkU2jVgFLIhvyNnQ43pgnrdgC2kfqNmrETcj3g59xylTZBT2A6/M92KCJvP
O4OJobu+1iXohiU8y2Xg6NgMbi5HtcwTbQ7E05YRiJm0t5wUwNbcJ4TqNdWx38g0HqsmvhbMoQ8w
Djy5wkaRnOP4OJ4I11OemuCgHP0VND6j6jLGewGziKAzbIt5TgW6MjYbCwEHwzK7wCMm3WWbFc/k
PlT0e/VIUVnh0WqOOD9oLrOrtmf0zZ/Or4BFBekB/rObWYM2Vu8WwGqRIuQIVS06mgiXXk/To87j
ugPPjvcYPXYPPlTCjocPwxNEpRZjxeYgTIVHB2PYM2bRl6E1IiLjiBavdHdk6FhUA1tw5cibpV1v
VFPtBHFbJYseGU2MgBNUyavpgNjbZjDz8x3NnPbhZCWjuV3UgbpcDwAz/7qwkniEYleDHpcwKxUd
BeJXDReCOe1JIgbIcwUzX7ijQcH8MtCC8Gpzo6p6KzghHwfKySk4jmi/LkwFvjvVhW+5co1jLR7Q
IqL0QTrSBNFkgm+yFU1NRff8SXiJLBDofVWQ1tVfUNJ82nAOyZtQz7byhPUR0MdCn/5V2/4ghFNs
pv/9QzDYBjCmVBwgXrTLzjDFqquBWSA7nSQj0bRs99A1azufF8PNMmStsSAN/dlShyqAzTrVbKwU
D0MB+dwIn+JHloHCTntdRDX88XbC7nfw8OqG4X00OeZ67HAxqL/X71b8hJ0WCSweSMciK6hF2+wm
s3zp8XN4Z28GYEgv0vQmlKRFmIaVF5LqPZLC7XqICslWLXXP9Ogm1nmeVnWk/ko7g/LgaStDXwXm
9QEyTCDzADlZBAt+ww5ZjQLHxa//SPWdhGNkZzqzDv0roRb3rFBQx7sYz6DxVWMWdVP1cI1otKJU
XDqTa6W8Pn4mAK6IMY6JmOJERqznfKgigPRmzrrFN2MgngqlWCFXKJnCkMPQiYLR5kHI8C/9DWVG
ZOkjf+kmLNxgfViRxLdag+krfyPJcOROXXIgM8tF7ygTjFhq5fB7jneKnOvaBSJGjuBAhcTl8NDT
D9AOecmXjb3TcBbMteMNw3/tqwTUJlYu7M5/SA91hGrfj13RJoo/ua0HpomWMmKzbG551vhHMk0t
dpQJdLBBZkUkAN9XzvDoNS4564Y4rJV2LO+XCi3tRjWt/2RgeMEtf2yXtnN497Mjgbv4IvYKaASv
0o1L3zi5Qyzfstr2k9BlDZfWXx+J/sG8oK7gc0YChHJsen8xfiaogmnGHIMU8A0yBZbnF7CDQt9l
cR6Yi8csRoipaNimHznukGBpsEOwL5x7ot+ME+mnf30vja+htnVBMoSJexRI5A4IzE39VSqLB7w/
HSJJ+7bNIpIyv7lR0pVzpQ7CWlzYMG3dP/YKYDSmaLlQpOa9bjjbxMmi5bmRSdxeC7f2wgsI013B
OsTOKl2w2lKzuIeqXP7OVA/yEhfr4iuGwkho3RL+DeLobQNak7WL7VlZjfdAXp5gHSRZIVqF/wk0
Vqs0pgrIFZ6gMDo6BLmLx0F2ikn5mPMJi4bphAwKaS4073bXw23Apl9E0fqkM8DUoOr3S9rL+C1v
BKD3rhKCB3FFSL9ogMY/pQwwVpPq5dvc7iKw33OJ55VLkUNoEmx8YxS2m2Y+opF2bw1SF7/3JA3I
vxIQkaqKpEEZ1GBtfXeVbQXfIG2aeN5bLHqzrKU9D5j3BZ/aKdCnhQwmCfIkhhWe3UKqLaHsgKj0
OzahH2ZnhdAU5uH/e4dT825VULevfsfE+NB/o7aUWb7DXRAes9VBLQBeOTWVHSMN62+frV5et5h5
Ut8qY+Lrr5lylK0C/4NowvinbhgCJFaUNFvJ4pa8+NUJI7JkGT5UF7uXdP5cL4Qhm8hU/apBVXvx
KIx7QnVBaevDR0OJX1L9fhkHXHOK6ZQajuzw/CmpFAcpe2Bg5yP42cDTyi3aJeDgZ6cGaOa645uD
jbFahUwUmcA/CZZi7GpoFP2mkLo+m8c5Alabo3CQf8JeOaoHSe3DK50re/8t+WLFGCuP3s9xpFvm
IOYJeF/3XKPp/J509bqQlm7Z81Z1euyN1IN7mffLA7Lp/dCySyI9qdHEmNEDKxzu9NaoVSgXgN8R
ICQTKPJrQE2bIgRYLg1/Pduxcncf6myD9pZdt5UvHkjYzpZyBmtzXqtgw3OjEaqNSQ28+P107wOq
KoeNrBXqe3xNXL+oilaA4ZhWL5Yl8THh41BNwCIGFwx06JJC/QRHWcsrqpbG2dyw78JdhxZym1BB
K/DUIOZKkugdU5k1S7nlt+KJZyXhvfc5aAhPpiSQ09D3i+s8k27Q9RKz8PBqoqzrMRq7e2N1VSqm
Afg7Zt9iWDOM7grHTWfrWkgEbLkiEEq109R/3EOAG2MTAu7agVhjP1D2ZtxdIueNAulx1vRTz2pk
ceWr/YMreYBWS//KPvIC4WAD99jxdb/UVnrUlZKzsR6XoaiOGhdFiaEEyXgELhM9seWq1UTaS6Uz
4moURfowgAWvJE8LqhlmEHLsXr1mfoQEmphbQ9EKTD3OMmI8+DR2bQtq1zvc2+gAdgEiNOUp1nb7
2vVOB+Lyh2IqKHU0CLlM6iym+JVwLeElxqNDmqo82ax+0JlUQDzQv81kpacGvRQDIYphjFBhFeUA
YyDuJlmYGCcPbkOcAZ21SEJgpdyS4hdiSDsD1HnaG/0CnadLzDCGjj6hbEjxL2VRNEWdWHMl+AoK
RPhKnU4Gq3zLU/qsKCjLm2NdMpBiZHk8XWqrfslqnN34/WLauOkf4Nf9twWEJBc9VSclBy6sMekV
ri81gflh1vijZfKVfwqMnys8Vy9MJZmCETniTDhDhGOx47ozcPiYiGxhrh77mPFuchI9YaL3dIMy
UDi2lpj3Om5wH1k0QqQoViqfojzeTxB2N8JhQzMLf07vN/6pG+2ion+HyvT9FuKfQPd9bUF0/1g0
TBkx5gfUuvwxEHdAtbINanewuWkmyU64CuiGqIrqm9rpKXRVbHkRiIwC8m0huEpqGjDvIYIV70cd
JFN3TAGn2k4uzMt5tJ3XMwTYTjce3cgkwRgsmV4j+PWhpcy1DTS/EAU6ErWKqxigvzuBewmwjFeR
FZCn7FBC3y8gMx8oI5xK5qhdjX9x3M+rqNr4fTYFIeyvwYP7VqCfDRqyyICoaPCWMvo0cIUXtmHm
sK2BwsNo4GuwaRKNtl5StDZhK/FwpD1ODVTHER5faHSO5MMCxFFY8tivvr5dIFzTzuKdF9SSY6vo
qINL86xd96SzSgdfny5qMumW255Sjwxtgh4tFs0F3LJA0tp06uA6A+8/NSF/6HQOsoi4UHdTdm2u
bVP0jnO4o3YdDi0+IYwWYPi26OeuQdR+0P+feaYWlqshhwrhwpnYfqrKS7+gnCieVRrPXtI6QeSV
nbY/JusyUDuMT9q4ct77CQngUmKVef2XMHiPe1PCsIg1+9XgH8gMl5BWGWDkBwhjx/T5wfClPnRy
SWiZ2JiH3uDB2fI25XsCKqNvQF3cba3TTdx04kDxtNGbv03/r+iMw63uVWA5sSP5tpDEgkCe6hHJ
HVpXY/rlJwk1s5lL5bzjslIMEFG00ZvCNOVklBWMc1J6J+tEfxLMan91NmRleUyaNGNcm4sokxu8
yKqQcSAsyGg1zNzaCVieKL4cqaVkxuZZdQW9q8QUiZ7GitWR1I1e8DTBh4yOIfpRUfU1l7dixP2J
t0UZ+g0O+e5nERgSjHVSF8+ON9fxYVA64fJtQiV3oDZqUNvp0Z1cibUHxXAHmTQmeEpW2FJtfLuq
B6RVdjGpLWXdLFxrBe+lIHX6ZpEJjkr1Sd7P+48tv7MS8dDr0GgmDYSrc4gh+iFuADePEBGddz2u
bxyLDm5uEussTq3Y8J1q99hM85/WbJZLpBt3i22Z2puncEMDZ0+wW8RY6RW6p4iJcqY+NBo+VKeK
uxWs12GPEroDyCrR8M2ylK0NZ4h5Sk89B42iY7gZxtQm5VacZK/HrbD/MZAx6QHJxJE7XRp6aqfU
AM3D0F3He0HMdxpX1RTSra/VPsLUgL89eWf4QKOMinpXIEkuh9xL9nkpoDF0YNBju1mNgnssFhXS
e1QrNvSQyBijYzVaZzA1u0Mmo81SclXlUwh8IGC2DC6asmb+AKU828IcIzf59JFWGGYZuchMttSI
m9CgBRlVynI9mnNLnaFYSjpeYyouFb3wOHHb9RESK6XW60BgFTXxe4Png00UTYiD960eYDJKVPLW
f4t9HdlBBd0lbYJu+32bMEVb2VW2E+Q6xkV8IoWSCQkoaoR7d3OH0aNnwR+jFSgBeC+cR5YpZ6KX
2JFC2cgQHKkvGyi4rxffrOGB/7TN712dkJ9jpRtCw6LSF3X5NgRvBRAV6gY0x30gkr/a7vndeuxB
tEmJX5qsbr8ZD0413oMiIY/ql7qqh8ESNwH1kwPZezf50kMVBkFWxB61QP9dT7RCL/As6uz7TcFU
N8/v8fHrf8PNBkxql36LtnS+GwoRIhlxVWK8n9pMACSHnnx52QRlC2mT4VLNmGCMFI++nvBbcsjX
zW2vnHIDlicebR4ilW5236d8Wuu/qLCA3TPdVpCPUbUvZ2jox/AcGpHnuLjUCAQYfrJA9XYfQlHp
mTd9NADusmesV+hG2PFrHySbOO3m60dP127j4dsu4pAXCHwOd9x8XYM39nv9o1jgxV+NogMnOTJu
WaZtT8jHA5ZP6bKngFWcHm02aKNKqcPVwr2l1Hp82TfHsYwWnx8p+gQNVtxCJVWYtdkoFm8Rrx6W
4H4BEarsX1Wbrcqe72qw9DMRsLkQmwT9Nm8lAq8xpKWB6O5j7l/yl6Y3/Gi6pLHEO2KPAER/tX/8
iv4/zWfOYBM/nlMzfunPTS94RItT1tRGarZJZRSZtewtD26QWrxW6AbXjqgVn94Y2O0Z7rviPg6N
pFpfjjTcc2g6oxjbr7lvauuIZPwlJqlmxjeIMhi5GRSzG+ru7/K25UVvo+pE13nQUpI74DMXFl2i
ldSt8p7JiVV8QpgatbY0j0/leLdZOoG8N5GSo5+dtP1GHTnMVyfYpSMnU5robwmZAFo7kPLER4qZ
gPHRxVcQ6/ofkM0LLVm9t/8ZOA76CKEdq9G5pOaSpcFtZ0OYenhB7REAu7Bm59Iprda982SL9HX0
rCwWv/Vk3Hn8OjCT8FzNha57R1vkE7M6PDFGtnhQ/980YyeWZIKNccgZU6MMRjOrcv3Qm9+X719g
qD9ZSq+avlBMM8TDLtPMKn02TQzMHAAjEJgMfb2cvbngH5eteeTx6PX9NMjWTVhvjNzyBiQ+fIpx
yrLs7RHU3Xsys/X+88sA3B9l6GIk3RCEdTAKScOVGfUp8W9hR9XKSlsVGPtMP9Ndw38Wii05mo8d
vENsEMydB7nLG6D4Zk03Az5lIHYouzTiLskN4c2UcsfPJMZv1RwD9Nmg9SiHJs7SkpHr8w2xIaUB
AvWMkFzVNnLm9yyaF0c4JnhYrxteM07O6uAoHUNXe3WS8zcJAve3iv1Og5KwM60XGTpOee+AT01r
ofFsTiEHedPr7m2Dw9uLcRfpLA56hLHpCZVowmTJTe10Q0CRv+/sStn0zjdUzfu6pWwjC9PgaXXG
ZPMRDVNG7ENz0UFksWf4rCRNpzVBxL9iMRu40BvMx6p495iE4h7UbrXrO8FyrMHybWJuWFusI3uB
GW6qU61fTMx1n+S7PQw9bTVeUdblizvGEhUFDsQ6nH6WeykD9NY7eufTJrIMers+4xeJysvluflB
9irWlHovxbEB/hmh6KryJ8GrmY45fsRHaNC6LUsnWkWRKV/loZpfBE5We+yNVpZXKA2dXueQUwmg
CWaMPWQTJHqiGnuWzRsnkWfahZJgx2E4yjlej22L52GSL2jFFBj+On1L9R7p388s2IZs+OtDPHF3
TmoNwdDnvoWIWDn7ygRumovqhQE/H40hms0RzOvopRVIQ5ZbOMaK8tq2RIVDCaIPalhETv1eiarq
pqOy6BO2agotfNs5/JhxfiZqT/72fwMKZyzmSv9gseaRmVVurjudu0cc8qiDz+PZ5lpdSlDHonVF
Tu/WyJ9omB8UbHX4xAltDyf4Yge5vkbL/Lc8U8vZT0HFJIPZXeABgyDmcV14Wftkr0JgW7CJatlO
M75u6Ptjgx03p1A/0wcI9VnmnGCTSa9jNlrIgkqWBbuc7l2c/CVkhuJqapNiU8QGuR5mtkeZYYHL
nGINRnzzrCD/kgWOvEMXEPJQEx2O1tAJGWRXE+EsPvj8DzejsAymA9MiR4vvTcYuiIlNsnmNV+Pf
5wDm1gSA6yC5+PgYBGN7Rj2Av1PLLZt8BiDI3CQIgnMafIyFPdQfb5ADHLcr76frS/4uYTnQfQwZ
1VPn60AAiWmivDUhXiVxGPu4liGHb/2IUIN4iLZReS/YZiO0/FSByT88SY0LgzEjDLm+ZBznUvoL
lpzBffGqlCHO9Q4th+LJXd1Qx0j9Ct5eJtgBnEJ85CceOHi0BSH+PJ3UwVZF8ulGxzJtApKcYi85
gJHQ9ztFed3PrkwOVl8DehCMwlzOU3u42HW+Qs9Vze/gHiJLAcAIq1UgSZjKTbUaMXrcnHX1r36m
DTOXMNmZ9fjM/PJVBEdsYZrNZ9jYCxg1ZOFwa+Z8lciHNYneALY9rgZs4RuaBZgKoYImkqr71NX1
IUpp/WS0gmaAqOfdrYztH5dHBuTTwCgDWz/eVquVC2Uvd6CFpJ453c8Hgi0vfMATQ3DxLy/sdhrH
DAcYJUbRMhtamfWTdCIHrdr6i4R9yDmRogBmQYiHPAdeCVx4iSVG1HoFMbOc7w9FqhNzS0QiaIL6
4qhFC1ShOQnZFL1PpMTK8e2XH9e+M075DA7McePkcrnIU5vsAlMChMzojTe68aSHJeMv+lrKEu+L
mOUDOKpxzsNTX9pRUtunlvQY6/0ZQARml7RdogIIa9UfCDxnN+Jj7RcNY8TeN+/tJpB++yCmv/3q
5ovgO0esdAc2/T/HQfBxD8+wQNSZzC9T3EPDxzZl/yXMC6f93DvGpSTJb0GK9I2dxfZgNSceCCAG
aFZvRaQi3KFF129H1LgjYdaPtlr+f8TGhi5stjFq2Bfet9arOOzVTfEy161syiW97KJOFWrhA3FK
3ituD/5rYggH8ROkGJoboyOL3VXIEPtisMpt1I3wcucjyZ5SPUGbbRrF0FILAMxu4tJufM0QCChm
HBMwmU6K0rI35KB4aapiNMzP3RTSMfPQrbIiBzt+M/jLg6/xg5ELx88aT59dmf9w/wTZ7ry2PtNV
xu0R/Hk8o4N1j92Tk5ZAhtlSCqMx1nL8oqMg015XfwRrsAGXDXRxsErRoXZcmEzKNp1c2FVQZT8x
JVvdF5WhJS5VhuIRWb811sEDZfuuIrZGWOewEn0WmuOXYOCqOFT7eimFkv3nn++dBpNINgDjHYYi
P7nJaQaAqkM5UM8XRYl1VYaZw9AuuAHec5pX9kckU682Dy2SleKXqGVimIqiM+8puEfkPY+zYImI
IN5TrotGMWJK00PQmk6/EyFL7VlTe1yo9S7ldDl4+pFi/ZkKr+nT0N+KfWZ0Sj8BfVYhUNwg76zb
4ueDfWWBdF3Ci2xhUSOcOw5XG32UwTO1gNqmsEdK/lEcg3NhECAyfSkeVao1SFwMVOSHpfvCwxBx
3NSlpQtdMa9i/rqNp7Y3FqpNOrXUPguMEr2/qhAnhXP0uv1Us2Qfgthp/hmVVaVvsh6KFKzh/A3H
Z7aB7+typEh12D89vjQLlFZXZNdj8EbDjS951vA8KZMO31s9u7Gc6iZuOMyRANZN5xvnN+oy/frO
z7KNCX8+N3xCZX9yo6yH80LpQjHwdLZYdXUr0vioupUBUQEasFhD9FfqBEw6i5AAziHkHLDj099V
yLswVYnkXuKCiE1JNWFzYibYhh5GOcs57u4W1iqc7ik0ZvL6w7c9kyqJVHzB/tOEeauOc2bONStD
Ne9GG3DO1rVHUJM/GCuJs1nSQ5Y74wPbIas69kcZCbTE0F5f9nsSFH/JyYdNEYmhmEG1UkyAKzbe
KFqdbtgoSEPhMrdxE0FZ91yqOBOMKJtxIrcQM6z77PVhyxhmj+bFtOGaEw2+WfCmwBU4iCKiUZJZ
nNgkP5pG4jh6jaIhDRYdZq7Vk9Nc7KkUVFH4j1mrQjoKbfufargKpgN1gFnt7TjwOQLYyHTwOIAT
r4m1O2D1j9JgNzhBAYMBe/N3kQxAM2xeN11nm3wn9Cwt4946n6p1Pq275R2vMSf2+ZxeOuygvV9l
1cxUrQKGBuXj8CJRQ7OLlkKlY4Vx/boGsjQ96WqyBaRYkoY+9MkTHTJhrnYNuroIW6ZAm5TWls3b
zj7gNJ1rfHzmOEC7BSNhU68bROownS7vfS8r/dszKvYcCvZ0QpKMXQpWyVmG7FDAKiDvYiFV6FA2
LvWwApx1HOwHdxoceMimgtog5K44KOqZ+ecut1EmbT63dDxmtanYi8qyCpGpkhd/lEdBGqz7Ysq7
6GcdTUIsvq2iyfml8ta9UOItW97pyqbO005Ws/Uzkfx3hIi31m2YiB5iC4SH0w2kSQVjXTGkF02n
yIaEoht/KxI2MlRHEfG+wKMFlxBrCS0emYsMqlon8vwUvYXGGGzRza8yIRzxN8dil4orctDlMOP7
tw1B80UPe5bYTUypSyxXXE1ZwqBgbOCg46E4rG017im8qcgbFvYce/WXHWzjHFFV+yMT3aAisn1C
KrpJrXO5kF1D3zVnJmgzKG6hTFK7vTAh70cpJR5r2YFEsNMp/y8m3PiqW8ABhufK0GBN2zzY9RsU
jndiYvaxCZeN/naNrX7lLRRqnh9tRBudGCR1lHaB+4MlECcnRcF3ai1dTZgRYcqBn6wc3v3lRXhx
VYAp0UvzaCVeyTOOfHVMDmzvsLJw/RPxLef+45otIHqR0EGC0OTiO4/iK1naFXcDSGwENDw8eQ8I
CNsEQyAeqQesXmNPKcPWDmwe+sw/kYhSt12uPArxuB2s5Tv8e3v+MMHu+ES6KpjgjparB1xsGv5g
lgDN42grdxyGc96EEUVeQyvoE/fKg5gpSSzjkEgR4+DVn/rIqnOour20/DXn2EltLGGh0gxuXiRV
vxm1IpSxe5OHz6mQgnfpH5X2z8+ppuwhRoCkUgxk5puwjECIHisXyiQAiHniMNV9o7ZTs6DJT62w
mSuXWn+y+c/H3mc3j5R/Yg7Vb72Jpz5/UnCcbssEN44cKztsVySC6sm2Bi/pWjFkSiHN1lpq+RRI
nD4nANukKz7/a8l8ZMjrVpfv6L992Woix6lGj5gA4vIa9pwHPlulIxprtIRdX46RULFmPG4d5x2m
la6yDp7zY2oJ5tp0eCQx+mlOkfiaQIsUUebgJTcXhdanbp3W1ygQILLeOENOcQ9F2sT4dXyda/jf
c423RjUS1U95h0Y8oxzuR0vEdXfgZQA4q/W5lr9OnnwHeAM6swXBzIJc3bfCw6BZwOwop/zvG/2/
fZFo+AqcbQw5YU1Yydw+YKEaGBGYV29UmvZryOiMRi+nGXfb5EzXPe+54eP0No3d+oTdFdnnfyjF
HW4Vc7HJq8/vR+oOruUIm29SgIarOYnAQOiacmFBrTZnqFoVomiKV8Vm23pkzfF2FC//TXQSuJA4
Y+/ibcHXVPa8n3no78sj0FiSBDkNJU/QWwK4kCRfW/Jy46XMMZHRgWIH/Mau6qTghRvC2800cviY
P+5RpH95/RQJitiEnQwcq1MglR7ImMIDWNZbmIiv967lnKnkFKZTvn5u/xHgkJF42zRb2crHhiYH
kLSlMJ33XiYOPiCQyqvpDg30Z9b+9YIoIWA9xXRk/nWX6BdwEgz9Z79+FASxxp6MLfG1k/S/h6Qf
Tj18NMYaI/S+qoCtBKsXkDVhnp3J7zoSYh5njnQ4gtV5a1UkfERegrqKvLwhAatZuipCtSVIMtTC
KQ0pBC4Bg455iLJlW/Xl/vXWsIR41qGL+Z1HcD9gDm8FxC30xT7tHrNYA9AnrKcGoFzK+sM2F2gY
EBHSvf3awaLXHmX/4wDqKL0gcTfxaJn2T38xWi+cEwdZ/+dsFU/uCDaTkmt9KuoX4yY2NAtvTrP9
nupX9tmgcaRmmajNJrQTeM7r8275EfykuffAP1avt1AnFOeMbXgVYfbDOnKePVYsRIIZGA5N1Jj+
C8yJ8Ue9vLkuSqZgSFiYVfnbtvpFhkSXCodXC9kXZy02dhtPjNIGIN32nD6Dn7nomU/bD98U5pRf
ur3rVShi5606rkZ1kKwYCXN5geGbNzZWn3JMgkR9hDq6cXr6QTFzAYqQEEj1+KriVC75FPfa+jiE
ozXTGsYUQDgS4Zgtn628wW0iFYVlBRakesrEAkfiU0eavvyBJLTvHq7W6xWFFXrI0y+wRSlaxOAO
g0XKz/UH+b4bvdMr13dhVYzAPDGYxn3eu03RmLERLiKLD+GfpZxKjKzcI+5bOOpnkL+e8gFFwWXZ
dw+Jg68MIwXCrjsUUeJbemSX5M+vHq85JSLps3A6424qd/oAJW7QxbwNTXOZ4yruBHRfY19zyUQk
7zu57AgoZVEchs9l/AcE+MB01XEjxKtiABu8BwAleiB48amKJQRvr6Sx8zJdnwmNpQTRdCkyZd1N
PVUqrJbp1/s89HeKuHfP09rU5aaCm4V+H5Wziv9Jv3PZt5dBP9lKAmOmtp8VtVKPPocz5/2It7q3
4/veT6IBV2CNdg2s6BEb/HtFSbAo55hijTiE8Y6ampJc0C0xw+yMM+R/pUaHZx9kTSwWCNwqHMPX
qmNeOuOfkKtmNNxBTlFLvV19d78Q1YYEnUiOd4hLQqGrd0qEAPFIlakSq5OmE+sCoUN9d+xFDqux
S0740/eCe679U+As2lPUmRe84q9M8YxFzdxMjO6h6fqgYgOR7tdkC0ktnEHALQNaf3bpeXW8+G/h
2+CSlQicZPsBpcv+aSAPOhIJTt6V+ZA6vctZAlg22dBcezq/VqzUGaHzFJ2cOvBRaXo1z68PPOt9
vr6eA1lFR8GGQNXGWM8uv72hX3yySOkKoRHtwgHC74e8uivcxpjWDfswkHfRWpHYyhblc9zZhIfQ
RIQR8XVSSuXzU69CfIEv7+eXFwSBQsboDNy0yQnkXPZ4rrxDWHhiTPjE0D/8QpHrUySDBFDSAw/5
WG8YhHtJeS4ILK+Cns556EKXp90fndhQf4V9+zzBxGppy/39SS6pNm1oVJoAfbqyV0cgGEqa8TUt
32brSVEDxPHQEXfxm7w6zXDMqqyGKrbExnsHFD81SJoxKgbplLnwz5lumdYiDKTK29u4L7S5Q+X6
xfQOPPLkqDYiuGcZ0axpnds4Fnu0Ee7CfJZOKgJJnG9tTSjq2Lt7ZbIM4/xycJGaadwiLDBTF6bO
RmpH5aqNkGbj/EhLKaAAcDoFEIGq0FvgZOLZjvFetqCd5MxYU7GU77QV5fu7XFwgviwtciNfSwhy
UglC10xFtMYQ+nVsz19oa5Sw8QBSM/VPC8S0N+MBEuXeliOOfwy7NmazeYmPoohSB44I2svaRqoa
CpB4gl6z14vALADEuSA5gSgtFWKwfpbV/isl9vWmckXvpAfoL58AofAWWsxpsd42g2B2cgUCLgs1
/Maxs0p6chl8KI5vO638eh59W4P7rXLmR6KdZtAxgxH4S9EZ9BuFRzY6nwm9lBF+eAA544EelgzV
kzcocSqYBtvX4tzJrD8RAZNsUgzSjz3obJHuSwRI+TmgftoyXmFY/HPtdfK7Xk7gJ7Ca1htir2Sq
bn2UxZZwLEo/UeyNn1J1yZMJVfPui/DoNXhOiKBPNrjOvuCLF9lsujHLPN/2sDwQiWTe+YkH8xY+
yXOjvE+z+LGPWtxH0BKJO9CnhTNFhIBcXrmovXJ1BvKX/fVGtUY6/ehyWAhpBQx3TsORq3AJPgXt
FJa0Z6dAP6E4HukfuGXvymFceZErrwKRe2r05AdXy27vsIow1TEsWjtOTW0mCh1fBCy4AnmawGx5
aMPWkG9GCXrFiyB4VnA/Zi0OGqoIaMsLOr71bFPjSEsqZ6tMwg//E2Lh2oAnEUrh5LriCploRwNY
jxl0qhcQ71y99Yz5veVCWCPi8NzQIzqCcnRTIOaFOO/Lo/tQCDd/YVhpaffQ7c9CP2f82ZfK0Bk4
qpaM36csZxD5PrimOp805xC8HqwzPpys0qySQZX6LOPx0h93F+EIRfttKnSObvavf8FJJMD8IBrg
Y4OGEsD6dhE/yqkclaO53QNGfcc86D//moHAq+KXtNJ7C1PrvDIWdP2lZyIS2Azcs7FR0CnjrdT3
aLjjGYygHM2krFvCHSCnJzbO1s3C3NWdCC9tc1/KHvV0UYA1+Fkzs+Pb29VKd6Qh/Yd6vpC6cDPM
vMlIPL9Qw+U233hb9rK1Qq8NzCb2zSJbFrLe9KdIw++gKkemn+fDdly+s9zhz/JedITZNcEPGTJo
j8q3np7jyy1Mxe5DUF5f7pInYa1X5nSfokFQc4VpDKKZbRkJdxlVwsKSvygmZKIUhTTEN5miOwRd
pySQX3BnW7UhhHi7aAg+aLjCULY4QJJJj3QaSzxQM6d2y2IXgclAzM6ix8mV5QxInqq9TiBiBWmF
gFMS9Fh8jPwbBi1ebQgwLoNU4H+eXeH9fXg8hgpeodunDJBwY++B+UTJIJUkJ9ZWY/DKl2c1GWkv
P7XFtKgyCPy4o+ojGq7QplJOqDuDmYQiSukXmNOn1Kw106KaE9erjAfxRDdvyS1YI3//OZpklm25
YxH69u6wLoq8Ifre8hdD6L2vVxfxm47A75Q99Sz4xvG8oI55KQCMK7dSHRgVvw/SmIVvtZN+eO+3
jZgLjC1+QLBp2CmunEX8wwPMTl0yIzixzHmVbDDUnHGpRUvulkkqfh24AwVhKyY/DwvM3tof4pyr
OOb/TpY0e2/aqf6VHOg6rIOXvPOr+1/9abn3fUz48yNhdRgPqyhTWt0dCC07ng+Wy1ztqvPZCPji
M3cgbwZy7CwxZcNau82qwul9/FsNsKBexDjI/9hXpAVGALfRlp+0wG8f6Mn3FEs43t95FLsLvQao
NsRFtqWubEjRERNYhZoMnEn+JBNIwzO4qyzqr4o02VTfuoFhyYN2GNMzPEU4+CrVg212ugY8K41M
U7QrurlbsDsZ+R2pq7bnNNASrm+ZcJ94jaVBmy6RAQo4iaU4+VIk1a0PEcUR88o8BDMA0boaGFRa
WyCOEniSQZMarrO2PIcQFmHxhp2jg9WsXewjC4CYaUczMm/aAOP1YfecuHIdCf6mzHPVDh3LcHdY
XYNP9jdtUJLD+EgZORFJH2sIn4wXqEuHtQ1daGXvnrfbfsII9VnVrh0ejT8b97lk+S0gXXeNeMmJ
rajGS9QAd5uprKYZwabjUigAMmBzT9FrGkt7mCM2WVUaNSdt2tjF9ZvAASHkioipcddBcb0yUNyc
fHgf1bdJOG9gJgghz0UkKOgD9HpBy7ps7hAukHXVmkpXGK1juxOMxUM9FrNCqoxQuyjdKiLz53ZM
Ccy0AoDYRzEmVaKDEvw2q2oGEERPXp8PbGXStPdbfidAMaaOzZ1AvE70e/wa67dDXnOkN3pll4rg
P4wls6JKVQyhdfRx37tVQDWzWgA8vj1i24p/IrT4x4pQ0ZQ8UGqUpusQG2FFTWTqEQLpo/EAqQc8
CkH/aMU73wflwf7lCOiLV1NoUul01uQ/LipGdjW0+ZFH9pOYCTMsa096sOBUYxRME0zLQJK2VTl5
8SahkJpunLkZESfNUNx/WcFYhFwrFTQ21uLMrmTyjkZZEyv5l59lYPM3ZDjpb8j6rldjkF1EGssO
TN+E53fC0iDVD2WMjokaWkxpoBnYh7UtnjTYUZfIBihSMndrQ2liwauvYJJsfFSj9m810oiO9RR4
aoUKU0pN7R9jUkL1n29oHlYt6HYoXgpbKdUkzv6m+975OoE6E3w5ymgsy+SGcJJwUiF+/1H6UlIq
RaX86yRpfXcKN/P4ph7so6evzob8KFRjo3lpKPEOZGcB07RpgH481tlDSvrEfNpbduYQjfc1/oxh
8GVbhwTV7y65s+NcYbsNIYXfZy1U+bVdR+HXE73xgLCN0gDl9oFaWkCmrEGgFc4/uoP1wNhd/0h9
4ismkpagWvK853ok+VgiElCGeCGtm6H4pkc6VUTGy+YVVUQmRH0mBPcF0rpmhCJHhuzaqZKtatBo
fve1mQUVjxh1Vkp0DIfA2GNK4qPv+mNo6Rq4SfTMX3soBSNTMGAd82h6z6+b5ptNYhf3URKiWB9Q
zL09DPjrJWnOPzyvcCjwm3+1fj0taudSQZFiQ5kW2o9tHkQWGt7l6dpPXsdmmp9wDDKA09ic4LN9
Gg0QTalP+P1pXKiSpMbiGLBah5X6hyuUFCrA5/7Knm1odmsQrESLwWRAxWwXH6mTXeJA8GDG2yGI
Gn90bZ4+9Udb1PdBR86YkTjsis/95zpJtAikFbZZjPXpO11lEFuV2Sw4IdFC3Ah8GKGF+G6qCh0V
kgU8r39O+DyFgwo0CDc+nzjyddxlCUJvH65mPWj7R0OhOEniL0KIe4M5j/rWY8Ce6zGCY7mF8YGL
isQ3G/SaeH+5tHKlLjc+6aCr2gWpJ3vqSnvCceqS1OAVYPBW96QuBsV5X15wfwMqGKgQMAMYeRK7
PQ/yRBwd8MXP0xnT+oKOWkzUKUNQRkxHhEVezcoQy+DEgq7ZeD3I79KgZrnxIEbs/vqeBJXRpAIV
k/aYkzMmZYz4P+c+3fiZAyeInL7Z5ZLa+ecKdSx3/skrR/7EIgWl5sdOL3sNRGfQ+40tqmgbaodd
yeGKHeq0zVA/f5d87AaPGJpDv8ft76rgR8XxmpOfPYDyvZ6ZP4R68ZneNxyZT7WRyTe8LYIPmwH0
0Uxe+X6sV45Od37HSrQYkFlmkaL95IQVzBumm0YjyERyWejR1d0gzATNbWuJb5IMwZSMcBj69FO0
FzEpnstAVBBekPBqEALMaGpWv8lhfvlZJq6RLZnmgktjktHHDkhfSLo1qZo3lukqpDh1dlE0BgWd
ovnBbsP/apSYD5UXD9mcko7ue2gDc6MPxgS5cmYZoPjMiEA2pn3v5Zgnm7T0RHMWuhOXx1w1t7Vp
R/Rwa6fn9v8xMtcyVCcjCI/18bAlM6IEiOHc0REk3D2IKegUbg5ZMPV3evOhMz/NUctDWat/fmc6
OZEEMewkMfoy380jY9Z7TjKLuqjlz6z82480alnUCmyU6meNBqrLqKP15Galdlt5QNTzL4fz+yft
Z1eXEt6bGogWfOnZrDYD6Ena2tnK2GSeQLc5P+Q2MqKVCEde0UMMuRiZWw5xaHtisOCOv2D4ylqv
n4gqfG9ycJfPrGIKPys49Wx2whPY8KAIklc6bvHWJO9TImDtlO69VQXHWnrYRM+VSeeNYnAndsxb
LRBkrJkz3VITgmJF6kg1Vw6PJ6xm+yKfVkXGNUdPkIzYg1vqBpYrp4W6u7QR6boA0lXnS08MigMn
+ZQI3UQK3sKRoloCjFgMwF2xFL5f1qdIoHlqP3mNcLM1x6+beUznsBMIbpCNF3GboCcm+sHX2Blp
GsFCifEPkCgbQWMU79gRnVVWnvI0aSwz3tVzU5H8302YpAjjI1akDkcw0Z0hsBKxUJjDWqDGjss8
sUjVIyFsMijStq02GHNbP9+DPBK2OpurWM9/lj1yRG0a1Va6yOv2t1YJa448L0MitwXPcP7E901y
gWOylMNUcW1YoIsXP+FxLBS6LBOhJL56tVTqbWmdk19lJLUXmvIwah/ukNuRJatEHTCF4FMbTaVZ
h8R/byiZcABtz220DoN2W4i/CsPWhspSCDFiVXiEp0BF8qMGtbZLX9lYYT0vEXa+DskywjI4M4Jo
Q5zHT97n+C/3r/lTVNaxX+7LYucQy5N9i+/5lvCL64Kkd5au721jxLAuxqPLypyvnMGscEemsZWg
0wtJ2q6LCrNPPhkHeYMKVSrrffsSmTbWs0pYbnaRT9hXZ3Q99f19frfXNFXmttPYGDblgiEDStVK
+Z6zx+LlP5dSiHJsUclWUoDBjJ4R4fD7zeg4ECWxWd5TcIWwWL9UAlLg7VFfuwBKIIwH3f7sFwVl
vEj3Qyc8mdo9YRSx2+oRs0IGwhQRJ9yTFTEfJa0pcymF/tUAVDVVf3sL4k5r6tkiF9z3pIXE02SR
xFHt+5DtFJM7ZDZNltL2TGd6mTE8DVjlgIuOwwWLdRdBR0F2EaMYIlfvqwgrSYvnDpapEXvqGDiX
hsq5xoNIDHjRZ8BXdrsK2Q2PfMl8yx4m8wvrL5PFUZjNRxd58RyNZ1XmX4zZ/4pbxDU+MTXv6dP0
uEfU2dledKW2tYlrlIxd98NZysFT4u9jFxf3SAUCQZY4fp9EiFqWV91KsVIQvk/qY6Cg25RTchO4
fED7WhjqJaX62LZzJMRiMOEAjl/YP56u4L4U8BMJ6fgootysE0MzKhBebz6cuBetSEKmMpegsdxH
SGRsJjC89ItF6hGgtnoMJbKyJhZZSjeV6rWkimR99gh5W+OE8YjW60i5cyiA0VCwuNbbn9mQlkjr
0Vheod2Gbnet6tKAqWmxYDfdlAX+mJy/RqVxRnWTLNgE0SrOUQYn5Vc7ZR5hoD2EKqr6XVko6Tqm
vDTkDssQcUwoHbgd24o96YINyZ1G/sNA9NoqE7MAMkb7jkb3x9tk+qGzH/Q0w2jr2XK8DRYOih90
Fi1F/Xt5gVxrcD/JtJ9oID4MImqDyBiSPq8KrHXMgQrUBeTC28u0WpO3FpaHyXGEfcTrJMQ9aA0E
/14X6eOWKTqqSXS1M9v0Ga+xfkSx2JRMPa4KT/OjuVd9oPcK1N6mCZNWrfvkk/k109Ee+OmCk/u9
zhLHVjOSnlHL+MgPuCkTkBMYDUuMfeXG7s81SdZ6b1DLQJievSKYY5yIbubmhtztBUJk2wdVBShH
3fHA5szNM13fTBixnMFj6pzX8msc/d9fxDsfEHeAFffZcaxFii4C8e9DXub0SnVSX1SeN5ky34QP
fzRQnVBHBc2kcipr6talMkYytrjcmomlViyKeBukl18t9oP6YkoAiQFveyc3K5Hj/uX/hGkeNMeY
wBMlb9q5cU9fDuclHNwmsLTiwJX0L/hEcVKlMRdTq/CK4CLfzW6H/BlCcfxdM1HUdfJzddBP6KAy
fCger4hxh/XvvR5UtlCy65ZguRSFvhIVbBobU122rXTGnOTJtUm/p2oK6MqUpZx4TG/wesfled9U
vZmeEcGkk28BvNOhTDCITROJLVi4c/XUQsMYYL/nlhNG2h58TF6r/qmKIUBULmslhazOJpC70QS/
Tv20hc/NcIaFmSPZ/+Aqt/sjFfuME+o34j+mNwrWqlNbiC/S5rYBgB8dlUfe4cByNMKdOeEgen1A
lExgHfzaKkfiTZUn8VF+WZW/odGdSl0yFr2k77S1eATrKb7uAAlVkgfbbEUW0RIQOvH1AX2FvD/i
0RmYYLAsaz+z9MAf9DgsMEkPEU0K/NklcOxlWlkE5QSyqKAmzeCV6C9gQq2R+beaqvJT7h6q7oSN
oCththwrmdkBCN/RpeE97QXaJ6Qs0hNfkci0TEnZTGZQCgVtiHYbK5gQOTzfk5a6kg9y9kBxRqJ3
p9bZinpHI2/i0Wx9UVsKV/Bu5wACYl7rTvo168mV4me/Gy48K2gqSyHdt1AtxUbi/kV7QvCV5zN2
z5mLAbhQQM2JxRmSH7xT5bLqXXqm0Teu473/kgAmz9lNLRupnCZGW8Tis2fpENsa1OUB+IrHh1BN
pkk9CcYGWeubaMb+NlbEhEnIhHO/26r1BqHXUgWv4PGpEI/7VL1MV2LeyFvjIeNxMFVi4QCRCPu7
Hd8t2wYXHZpiJr1ETvHIwj2I6qABQ5qpIMHdvFdmMrqeQX/4vwbawS+lWvpGuGMFvQiw9xySwIse
SX9ro2c9x5rRP1NSsbzlD889X7WAN6Ru9xXLWwNPmfLfR64ALJwLbv9vayYPUt1orCIF4GawlCcd
UfkwTkzDBaraXd7Cz3ASGFG48MqngxWRIrwSWKaIhz6/AO9emSWUYyq/a+qgZlDB65SWYffIosAb
RSFpyeHPMIB6msdD2s2GEdnzV1SmbHf+6p6Mia2hxy2oxBD59eWU1P0X3tFgzx663G2sRm5UnZtt
QsfdGFo0odEqlYyHbqurDZ+kRC0nn5bMwHf5gbVgvuXj3F18dJzIlMo3Ade0V5tj2YwAP1eUvRcQ
GNHfCQVsAgnEaMAZJyrGstm/KO4DumLcY+qVrMcBwlWP5OlCf7+4jYlz6/S/DtYgaVZyiBop8O0m
7z/KIpMN7EVEtT44iOLxKVSzl1STXNGVjx5HYU1MbqI1T0+FPDrnBIGtw3N6rVzfklW7HQavaoJc
oOSN01OxuCrKLXkplCqvDCK9zHht726eoeEv6BS0YAulJoseyZKbNzdz59MGEi/silU9ZNVAM/n5
4nfKAdpAnj3rp67+uSRAvetlt3qjgZs3rXynStWX6/+rM3RZxLgs+ABNi8xZ6H1MM24v3ALUdZcw
1GFLv3puHcXXG7FMckBGiN+BC02maNAbCxynT8SvsnIb7l5Hsria+gnkjj81xhPGpKbErl01SPNN
yYxZE6cjJK/kFFZhG2NKGdj91SbchWxQGjb/OaT/cKvCyyjUFxEhy7Ajc4UdFTdgD4q1FhBDKDyi
Df/SLcWWdU9WkFJdYJ47mI84NIMGO5PrAaQIfvIe7HGWKAWqKTzb5+qmPXT5B0Qr3048gyoXj8ez
4TNqDp1ITUgugKpruNuE9klgIL8jyzvqD/ZSXoXGrdWC0jnvE/2pTmkX5OEZ4V2LXBoIkH1vY4MM
N2Es64t7ErAndYFWXIcElSxudUS/NglEp5VfIbv3zC/pDvM2k3jhOHqd4D0Yi7lmu4/9fb2Qpiob
RPyh2k4rqMQc6F5juO/va7xlciGQUGYSh2R3WXIJrsQ75ECFeunpW7voBhHUlnSkQStDqvtCAOGz
xpwchzgRTV8Amhpbd5ZR8vEaTUD7zWYc42AGBdNaoPzRJQWTJ06F0brsrxVsdiOKa8TeYtzp5Rzs
ZlCKHnx84haDZAmx7RXAfJrwCKeutLd7U1VX7XXVaP1yw01mjBiYDodngceeZ64G/cZOBkcE3guB
/GKir4TMYUiFBGTE5TwZT0yYGTL7+srqaLCUcd8DiiskO/A6iDr7r/r8r8noE6PblchTiTgcaUUd
CUe6lcFlXXD5HvgIAbOpDWpM51nmR9JJVThJGDcfrANJZTUpFRjuSxFKUcmRysaW8CrISQKKsfkd
4bcu50ZgxezoOX5YDfDkybFzZJcQ0mqhr4MDkdlnp3rGeZ7i8Jqb/hLNR8yQiBpsrsK2FoXlcYPe
8/NG+sWzagXCITYvH+eslJfKPk1gkMDmEnGSFTdFPNpGFgZ9Vy9h5AzjmddIHII6cVwUiCUeRrkh
1Utubcn/Kjc6S6ukXXobZ9mM8vkELK2m4Vhe2RG9nY//G1p9PkcINxexkyPCHUfmi+qjYu+ZOO9s
PpPxex/2wyxL4X8IQXiv4Kgc87VUo8CJvAZVW3Y2cpfEB5is0M/Z9vnwtmfwJlXrje/qCa+9xB5t
f2kunGHOUPpmpPygWj35oR0Q95fhEIx9fSsJkcDkvfgF+PgWAwnZ4aSWE9VF/XO+qC7MfJC6Bkxh
oV0n62ED6WO2y8F449syNfyg8wwFev1MG3kOVFGJC0o4A2KZn0CFy+s92mjtoqMc6nrI94TYg+Eb
iz3n6bAgoSmTLSP8mRApgEEihtBnlzOqhWAWn/OT2rhcYHtfeERoYBS/7RFCsYrcysCyXhkAh8nS
DEyZSWnANP4y/pTHAFnqOAiGz0psKfs2q7CwHk4o5P9UCjfX3zKYGk0LG966PjnrULbIcUnwxcN7
1nKJJJKdhokSHA7EPkEthxNsmeqOgHobn4PBv7iMPtb0YOv9od/Wmf0LY0gu1yWSQX1yVFHrWGdz
lU1yE5IMTuJ9ZAu0i7dG6RIQ2nQYIkjqn4bIQLow8mSoXrrVIMTo4WxmPnF5WZ8kSIiRltKs/uIp
IQcKIVAJm81bNY8hYznDZz1xgBrVkgbcZdIUvxl55uI/nneZb9QGZ31hQ/u/UffQIDL5q2bV0EAK
dj+QuLI7yIrgzKEhDm5Il4OPNEgUyDQ6TsH37GmbQj/ifarblRc22KyaR4jGdOGKB9hksYaQskF2
qp5PKg/SmGnNfNY6LRzM3740RhQaMb+xemuGxdoqpOpCuHIdcXt7cg4XZ3ifl4aeweGV/9Mw5WKv
X9fINUn0d2y6+JYKIm4PwVm9XhnyAAVnlBlQ5eg6nRNoRLlkGt/NTo14teymHLf9mCfmB2E608fT
teU9NEE4NLU5l3NvQGzCIVwpwuUDmDQVGzfpfwRN7aeoXeIhbHku+eHlZuhClYAV0CzoOIjBK7C8
m1YzKgYwBWragxqxvI0IkSkSGcvFaCqK3d3EImcdA2zQ6yhDzj14BKp+jT/Byhv+UWr6lEnDaWQA
0BhpvDqh9TRUIMamEmcYcRvB6SJ1kHctb3fqVu8THYicKVOPgwlTh5hbsgOGsWDa3m8FZVMJmHIu
SJvikrI1mIICCNixoA45I/hDkCV7ngXM7rNF3f648SpCgh8XTF1hOxxZgck2VhTjmfSew2iPFJHm
vFbzIKwexswn/l6HenYZRgado8LQOntq/1mqD3QEreZEAEDMxIvY3qJb/wLjUoWEHZiyR//knVGh
whX50La9cjWBgSV1XJCKjb4P+AUwnYEDcRkmB74AMwpk0SXqmyOa9X6LnjdN/bsOWNGrpggb5cOj
92vFxmv/r/10xuic3HzJxaeqSlBPv9KgIzV/G/B7/y0h4Fcoot5hRqMtAk5RbpCZYM/VlDMl4nuq
uTJX+f2SWOCsKdBv7y6I3yZhefvMvOdDCXr8qz1ib1USKUEXXAtLhohbyLEfh3ybb5xtz1uTzMRk
AsMsa/P0AcuWq+sLRAtfx0vh4doLjgRib/Ilen+l11+/SqMjFPKvhb89ZZUaYZi4psOBShudtNGt
TycKFmHDFR6aCToWANWMY6e9sVXT1pTBg9WdxRy81f8Y+20ZRXwSgL/Cmr0glbqiLl1Q/U9Ko1Xw
l5XgfJAt1h5DUW9OB8a2HCB9esZJcWufiDuomdpxRmKRXppbFLleA5uTAy8Fiw77bPEKTH+GY5Xo
d4sEVIOuaRvMEDkQ9Reh8RkK2DmqI4UTaf8jKizJb+IT/E14fJFdQ1fvfrw7PDQxgbBoZG45k/fa
SEqZ1hL39djvrG1YwivVvrnJO6ivWxHrrmR2RjwL1MOH9CfgtlW+xkIISPEGmmJMiSfnrbZZiGJK
vMuZigRrLGWm+zxUudRIOJrU+rOvbAKWr/boZzYjDq60iKcQXi1xyLlSbufDhuCVCM7oq9lV/RXd
Oz1KwJrAqrn0zDRIGWRQOm8tcmSEpwA+Bb+jw4mquVH/F9QL0sF+9cP2Hy2v6ruKI+iJWf9rkg3K
dgEEnTGtAfK42BIBZ3GMd/fUcCQCp4upOVu//R2RCoPAkxSJ+q26xC00PecKEWKwBvucp3YQI6My
vtMIMos66voPjnF0RQXTGirBJ/4pDAj/F7LevahXT5tzCNOgYpe0PYwGI1A5q/DzqS2yFC/GQ/xB
ZtT6OyejnMFxSPIlDv33z45j+L7wXLcvrrwAaASfHkajE+WPL2qEfaC7+WdOyMay7BRBdkpBnxEG
U4zwAQ4C1EtGA9sdwwk24hCFzFjfA0oUym5fseZb01Q3H8k8IZLrLTt3WfNbg/Nx+JTcUWo6uWzV
5FsWaatmj5Vf6cGESMjDj6A9JTYxYC8E4dzUOkSXH4i2xSY3QOVd0KJBhaZUrF9Y7p30wiMtpwh9
dxf+vJMkPUZBoFvaP1AxtPDUIk+2oB4zi5OqN0lrcN2qF2ma26Vvh2tg4BTSOtw6HlsgBy22T7LW
P6omYpNKmaLunfLtiA6avDEtnrUIEl8bm7sDeUwLNkYCVydGN+I4CtRH129Fg6bHFS0whontpiUL
F8AmjwLzW7p0vO4I2Xybn/66NKarvDl7krYhYkoJtTnMUtHMBaR7tvZXBx3/P7btmtalGrXyl0bN
GuXDxTem4yFNcS3cr9400UzZAfZoyJmRCk1psLlCFa+MyyOU8uMoJmW29nY8xR1AtS+oUWe2QqnU
uSe6YwWHkMsfaytrqvR7HldaLAGfsn2gGBExt5rGwtkttKT8nxzI2QgsTbA611dg1p5uM/mdxDOd
7WkOGQcMjkYF8PEWWrcqxCZS0MSaXiMIFORvVNuMrluUWaGj3AwStnwHJm0C7KoGrvQ+xsHcXycE
eC7rTjOa4aWLefJaAaOOFz8mQu1Vf1wrUbX3F7sP8wWCgb5Cq8LjrljTYGl2GBUfmcJWEfhfoufQ
xK2u8kAboxr7/NZysrFtqT6pLNXPazFdVFNhp48+ICF11Mk+cADjeXkDq0L/NyFDMGoPVpZnVyH6
ZIkE9fALeJI4b2D5Nqt9SmzfUtF80QRuLrsQ/ahWqXW/sPAJWjBRbJeWuEsdHvxNbRdO7wgH9Rwc
ryVS0wK55AldKVqLDXWNdYA+TGQp7AatlsRV9/ZobQ6hYeuOVSuPHDKcGavJfnWHUczqRJEgF3qT
2uUeFhpTlRmDMUa+9y3z8G3pN6fQjZAN2J+7WIMdrOYUB+DwDy+R8wF9orE4SpFcVNw+//DxniJa
I13hDNMKpehw2GTwCzfwcVega8ZK+wzUgR/j/ThCXJY7RV5YUw6dNEVEWm9gS6IduSkQ9lPToP+/
nO5/a+NrOnlW7w9Tw74FgS/roRZD9avBpPAVhforp76e9mtMvP9P6FaIrA/DSWMbiJcyVDI0UDo6
FZ8pPy8k20otxZp+wJWRf5O3p4yqvR4p2AthsQqdrojftym1b9YPQ1CAzZPKGEBBxrU+KCEutgHn
nqAIn0v2y/RZWYvfOfLBNn91nwzZsp+trt+c3ltXs3sc70IHoOvgkWY6wf1OJXgfbZqwOkTdimsQ
wxvvxruVenqUTcro7UEi+PkSA+9/9z8phNEaYOFfz4+29p748v19TJhnoQLm4g9SZktNx+b42mQo
skgTvoluaLmk9P78ObT9wlIUNHh6I9YVrrUlOSDPk8bbDjwEPVr0Wm6TVMBF6kaFHegBaDS5SZOK
Qp+CfkX9Ew7zmwnjFSR/57aVgs+7zgjiYSuT7qm8nMjlPx4oFISBkzR0IfIMn90X1DsvypGEPaCK
y+dOXDXiYuYErrbhB05zeD7fSIPsAgCe3NqNh6pRqGfvLZfqrSf6yc+KizwNjzHymjRvAZzt23io
TuSoW+Gf++xDl/+novMqDr5ft6Hzd1DXSVfyk2+bcTkn8K9lFumPr2BkShLunIbwfZWNOlGYpM2X
s+skWxwqqR2oZOKYKZskrhxsfPaBXdD1oTh4SODbrYlnyv4cyLyOKMLOM27f4UfampixTFpOcTkM
wg5TfoUJAdM/JqCIwMbWZrixxanctRuINjVFekghEMP6S7I46jRq/24cdusbldO3Ut3OxkBQD0LE
F7ylLKQB/rSrm2WacWeJcQtROwrF3RF2D5em7K+GwApBGPmC8QVguAhGjbu75V9g0xOIdEzgzmxB
Bbhd9hDqXiEWtf6W7ngC1Aq9WSd2YoGNioovCRyI5r/cixknwccJmxTZI3FNZG8h7ioCag5QOndm
TNZ2Bxu9j1roBJKcWOy4P8mco0pnZUou/sxf139uGnCvbPiJAgyn5Vd4r3k12HUCv0DRJ3cgkGNv
X2nWAZj8fU8FAsiaR5Xosf929JSMFtq6HcF8wcwEmBonllekx//QQ1PWBoYd6SFRLjk6zDwLvYsH
4f9soZ+rxofyVv4Sq9xAMQOaUgzycE4K2txA2l/dkH2JrkD1wOqlN2mJNp4g+9Y9FatMk/CHyl0n
6xSyk5Aa8R1+99Av++D2Y5VlbjWVrU1PaQO6OvU7IhNsAHSmA93owPyb7hAlveGgO8ycMq0EiR1/
HM2yY4vcwG4qS7cxh+oOfFmt0Mjyx8U07BZXHATbkTgmY5nEqFy+ASomBvs78bUYvOL/cFMlBeaQ
JPqpyvZ2AaRkR7BYxtrTf+98LzrdmfQc4pUeqqg5XzHA461NVMmXNXYhhFuWFbPu3LPJJf7L8j/i
AukFSwpMuYURNnoRaWan3C+reiC8hnDXOUPFShW1WC/XjHGKpiojjkzeUkYHuv6gMLqfeGAEisTJ
Xa+Hlpyu17D8Wpo7/rRX7RscPG6yLrcRUjSZZzge/Jk9IwONP76JfJXAM0qJljZGaUWQKt+kSgZI
2PgKWVT8kjfhZaqkQXq9pnD+dn1ilwwCQ1gwSc6NrQHCDvTmA6uRDsaWl7t01pSHFmv94AdGTxB6
DUm+9+qj0abwt6rxZ964iEizs4KmjuanmI2NInylTyL7lv7UpPptOWqWuSoU9oZ3hjrIzGudvfre
VgqNXAHy9booUechpQLeL6+YH7TNtMeKhRMMQMhshPH6CCFtJfJa8DajG5MG6J4iwxQCxDIkiRs4
QJqB1SH8LShu7FqcNi01aJLZ4u2MUr6KQ26HjsJTptMc1GkN0dDNegAgkUMp6gt2w3mKQ3ED5ppC
TDBYU0yEdVgqJwbEeHX7FTi1C3RTq9WRRXbfcve3gRla3uqlykSo4ZQzNu28D5t/zaKivm/5Lmrh
aSfwabKBgEq/F8E60NNzbbBse0zmh+TzOoGbr6U+3D9cnLmoXY+tHT7IbPODfcb/1IlRiSHbDv0U
FeBDeRnIGzBC3lfnB0Rg8ix/0olEfo7MFd35VYD2+6KCDJlVP0gAWanVTOjvPYMR0h0AqwyGMfrN
4Us5zB/DTILGcvYlGDMxJX086TT+QFctTkBk6L0USdiiTD/LVGkVcyXyrVXuPbB5huVEJ9ohYrVC
nYQ4wi6jk25xnnahGsKxUOqZN5NiP2AOKKWKbp/0cIrpKgJ+dxrUuufBhWHHlhU7Ohfzz/IEerfN
/UlftL6rMeJOFXxzSa9N4FT6AX8NCEXC7PY3i1damJQK049HXpZbWFK6B+Xc6briMvjSov46cO4s
rF9Fo6w615gCJO/2NruLZtRnj4rB51F5eWuF0zQPtwY75ab/Q78PyGpIzRTzJBtx9A5mZJxHApRv
f3HUR7zIwe0ZZu8BY+dUTj8dplYslVmNsT+kCxz86GowV9IrIkr38s0U4v0EbcN8x2MN9cbV0fqd
fdiuP4YeuBotk4QVCdaPW6tZsfDnKdN6fKy+hO7t93/fzm28PR8swM+txnpUOx50jsQqvNBEtGeb
csyowizLyzTMOWjVU1FRYffTzDxBQRvKj/C6ZIEdl1SPRzzZD/XnZzwHebjNOZIik7zJV4E/N2+D
yE+xaB+m3p5xfPIFuvTRSIdbFQXsqgpCJ9Tw1rg3eJePAFNiCt+SXMOtD7dLPvloe21N8Ow6TUyI
hTVqmfYkE+qa5Bu7Z4MC3I0tkqfUtCK8irzWh+kKZF0MhStPohOrkQMA/e//pMLeIYchGgnddAAC
AwoU6P9kofasHvnyL2LiNuXDbwyF6swKdG0vcCGNS4MLvP5Y62MmtEus7pjCwIMlA7DNkrNdWMP7
tyNWGaKgZjuY33nsMa2yv0yjJmdMYQFuR3KkVb/7NkMYQWFE6D+P6VTW7KJ5hDhkgXRO8gzUjFp5
4X+3iPrtWtQXta7AtwrA62MLY09QAMFu/qe89jJc1gLyrbaLprNt6tNIcm0hypWKAXVO+rl48xmp
JZKkMUcbP0sFBecq83lGCGECkcFYXW0U94QOVE0R3F/rI4cWoAw/TKcb9K98aO2G8AJ2tkVGRzJY
UOfnkPPe/hI8g2JoYIZrF4Bdsi1kkf4xjkWkSw3HJOTQdY2ucIyWaCn1D/fkl7TkqeGig1fuPOkM
KmfyBXwP/JFkIWoHLHXAUnqXYlcYtFijsVnyQuVM8rX1uydEPq87RBtFiPGn5KsGXVjih6gfiwhP
ueKcsYYo0cZyGtwPeEYn6UHCqufD4zmdmHpyN90WRExyk1JnnrwODPTlDi6eFdDbows8y6nISgPE
Jaihqek9aepAEnpapVitZcJSNT8b4p7o/P1I750nZc3qRo4jrchM6LfQ912B7vvhgdCDRkQgj/c9
Vv8I9su+RTmzUDBDKeYIkCoH0zakOvxpjgGkJACpr+zAk+0m6VchqCnBMOTlXUnS89lmgjKL2JwM
OGvdnZwPlWfvpaRWydj4bTEuUyJewakc/e0TfwNX5Gvowg2A+4uQQJD0oe3qYJS6d/RmD3/mnG7A
AUMkehlXVgE/A7ymvTnS6g9KhrqSW3J8WV5Vrlmc+DebZFURbOAXpolAIPkw4vsDsGGRgK1IT1u+
tLxlFtcgoXHQ6r3ueARuIm9GXlY6K/qAQWZM13NHVKa+G003flfPKaO1GHQd/P4TeNyauqYtNO6I
Ng/kMmygLrB5ukK+nPLE+f8MXMSUjmFKAI6u5xj5FsrJ+LFax1nDPuj/HSnbjYoevJ9NdGjh3Tyf
94zD3j5gKhNIC4gNmz7MiMdRJGee0qAc8NLkTRtz3Re/ccYwQeygQElqr5kRwNZY7aNFSqj7yMKG
H0zW1zoWmW9ZKjTrLJEcgOqoNnUBPuvlZcv742efemMjPqIfyiew0hEMnjq+X2hW0DfSv5ic0dZd
iESrcp2/heyC3LcSJMsVUmwbEbykwdqMQZq8IBTqHhtcfFIzSOaMYl68s0gzViRHrEjDTRUZYK5s
/lDUanLjJBvg6Gse6rL8RTbNeHJzyZFBoyC/6iBoDmqRuwN365fSvFyLiDMH0t/paCQlZnLGjvpG
ymSWv3s/WPTxuvvkJwQNyHkeHjNlQIZq4yojblls7zIir69m2oWuYed/eENITXPB77NsJMTveD2g
P16ukx8hcyguAYDVw2HXmnFIV1TSt30sagn6mDWv2hIg83YxLdSl9kIQiCNid881avMkQNnky/yb
33yiTB65MJ+7zyJ/OHiJlTVUsmyxzBzrr53ihSDTvni+jmYnXkfUk+aOcgHUElKE1Hd9/MHChYNS
hdKausOsUOoMJgr44Qur/2xIaXL4rJ6hBPRtR1VJ5hFcMRPVFUyA4Xw+hHh5vGZzkYK48QRtcprr
5QPYWiC7OsteLI63grcmiwCdXy9kSnrXpIz6E8Q9QWxA4TgmrXcoZgeMcgF5xX1/dO6Jqv2xRMot
Pxjg0SdTmV813kJRO5JHZf0Q3sYo+wtbthzfOUC8QYWSoAiOFvX9xPJBrmzPmXaz2TznLb99qKeG
HERyu0z1ZnHuj64ZhJXFejOgLzuGfWz8Ri9wIZmSMM0zW7UGoeVsv8PRi/JNw3G+npSWYU025NJm
Fi+ZkS94ySE+8kkhm/vP0lPJ/6hkDQ6hHrWZzUdxZeYx/rGHoL8ib5iSafVWIOE6QZMNzMJPIW+C
To8bvZeNRy39/mlGR8tHcs7wQcjvXxF0YgfBbzXTXHfYKm1chLYaRU/qyIwmdoV3E5hYOuPYRBbA
NwRbGeGL7NmAvAAzeolSUrkiZB6v/bKs1zj/wQp/0RH8wrnj2yDdYphmUgjNBN2iAkNHi+Bk9Z2d
YneZ5K9rGrbQRHo0az7MDjK9CmywJagTITnr9PKbY+wIkBFtfJKYloPmYtBrp4cjseomprtyp9Zi
ij9A+JR0ACV1lrCkLLHi9wsbFyKZFUBmfJKP/U5kl9T89A8/JeC/8aZQ07j/cTy7dW22aH0vPxj9
Je1VCmkxSr+iNfwE/kYncD0Bx/2lD28q3hrTU4MbHmR8tHVLQ9yqB7A/CEPLG9gcRHs0GAICCXyE
cR7f2YV2urtIJI4G0qTs/rLHDVvU+WAnbaugJWlwh7psWpyU/bvxrV75hG157oTTmENsbKvMau6A
wWxhwNsVMY53pg/hw3nJo51JugSLh6DYUjb0EEq2vBx20Cf/q5Yn7MaAkmwWnnknMYPlfgNmru+V
6mipjeGs66Bas39EsOWvv7HkCxsNNO92skrtIQFf4ulE3i+HD2NIpGBr8lEvEg910s61mthQhXn5
eHxwGXy22k4zLJhW8edSenUrSXxbErZ3kRyaPEcWT4hVa7afv7FK8czIQfKgDPIM3aadhqdYyL05
hH8fb+lRpq/iUNm2w3gnvINMLl/d9UReslBj8vdmh5b16un2DYk0IKqvnbj+GXUCk5XlHaf/syZg
KvK1WQs96AJIsfeOg78ed/WYEXDAZadPYV6zfKMpChpoagP6hHbNSNYJC9FO1jOkdOEziY6lil8C
pvdH7Pafb+Dv8TtaFKiuIEFSwGGJjoade8zN54GkPL1s49GoRhzitGDKb4o+DV0zIKk+8zWfTeFT
vMMgJwcTANTpl0vIOkb+3g6g423lfp+OGgGJw8VdzXQeWw3AsgYCzhAI6KvZohzfHkHnHzcLpQI2
tZ7EKL7uRQAK1OOiUPehd64blWSBQ/34909bt2xqnEZvSEX63z/d3LGCnZ2SI8t+IzTqJRAnUynF
0bi0ZpF42/XebDyFGT+ZN3eUN/dFnk6o0i/KymKPI6q0WS1N0E+WA2XLGxVX5BtFhh0Slm7FYyJh
NRQ09xvRoplJlHaoLKjVIx94APziOWhjqmPKGOMFgsrDD5M5O5kl0UiwcQYTjiaf7MWZmWHhGbhc
D8x3d++4DS03jqiwiGXBGw2TXk0m+2e/TmhZcwhaD+CsEpTqVi20JRr0+6O6KBcF8O0jzNAOMQXl
Gxj6Uc1JmU4G7Z4Hx+8U+8woYMyzheagR0uHOKqzE0cMQ8Sq4a9hBOUhThtDda9H71uwQGQYEZhK
IPw3BF4kKSU9sRoDGC0x7ZFzYtOyc62RbKSDLOEoMgL1YxPJ7LFZwmqLGHn8KpPNhCLEGK96e+H5
QLDHEpNItWKMCEWqwV/20iVp01eJaxnZHnNcRZTqKr+AWQhlxBPidM1DhJGe3FR02Jtrf7bZffHg
G7WJuC6lbii4LW8qON0emhx/67OhRaprMolj9nvtX+USev9K/bwm6oZE08gAQSYW6hZCwJRu4sbk
dp6uAeR19nF63xUsknfhlzNmZpv2UfDEx9vQ4VprE4bpGWUxfuGAOubG43ju+l4PNIrG1xgTP4g/
x09bNDZ60MPz3M0fJCq9vRdwf1OAWoaJQiukKw40grcXmMO6ts2BCvILwX7GvMKAf9Hrm/Kre6O5
KJyn+iM6Wuh+teeHBUX5NYC3A4OIk8ybOyoO0FbrFaXaYE7PYIDgOmd0d9VGK+u7ufHESmhkDKRt
6r3tGX1fUEa7Z+GkZadxVDkiTo2EAGVkjFKYi+B3qTxTXZas4BEZSiEGgIdFzB34sX0o89EDFj5p
JdIrV+dDWtev0yVTyYcoDw46AFbwgCdMn2kvyMlvq76A0hQVRAjToqqAc/0H6N4d/nihxfK48q6a
AmsAGZBvAF+mRM0ZnF6E5irznn8jT2KjPhTv71pgZDMjwhv8U9FHZciII5nUJINhlSMyWMywbSZz
38l7vgL7oz5rnzzp5Zhg1G6MwUqSvegb3nTWVbr1fB7qjKpiRa49n7rpRr/zI9r7pn/K7L4+0AK0
KFkoEWaL9wxk0u3B+NOfaEoLKJjGBYKrpuBfSpZwElp3KmEM7EiUkYRIJku2LPeApFeVyqhdvWGR
Jaud2Xn0oWyUi5ta1SHz7MbgEoaEceh2g7AkZqI2eTIdtNxv5VgqrV/sQDsbKzXIRiMp6inwOQjQ
K165/HvhoRZXjr17dRt/jz74+Yk1Uy7zuIHgQQJLiExzjDVmPS766892rh6YNNBNTlCKq6i9GuBu
EjGYm6U8v+pQpGaJtL7IFPoJpj7Orhd7avul5K4rl4Z9Vd4Jok7k2cL60pVnHOB9p4Ut5OSHT9xg
xQ5Ylroq3Ddngl7nkNMjDhX/udqp8+97h69BUCkBJDYVpY6IXqjq1PeMYpApSRZeVhIMHyEvd6xI
ezB1hYUGrHyf9OXw2IUmTIiUr32lQU6pu7VDb4VBWi8DTnWqGWUdEI9ZlWeDswA+AmAsubsZzBGg
Tx8dJ38nvKTkQgGlTnZ/IOjA+Qpy2xK8Xi60DmEzagqkw1FmvX2tHOwSI4eRDuMW9AOHNMkIdrNC
O+YolbOGVq+G+H87w+wa5kyjBwKcXGBXHdaupTq9hF+ooxJ9Io9Wdlq/ASKtZXv+ZFxJ3RecmGIr
2K6j4c1kHfIz4FlS8M+Ok5SCaUWjdKs6aEEYtE+hmlmEowb4zYywNUhdnPuiBYofTaXpg8aHHg4M
vOQ2Sd9uSpgBG3hSmBeGVMsC6rEL8HNtZIRA9BmP8wnWwgzh6XSaTCpE9iVQRSb5NVLOaGPwIEAg
X/wzQbTRs8cLsLfLIHnEBQ42HzdceN+c0DDPn6qsZwtoFGBRB3wHD4GJz51IDx21cRRL4bew71t5
tkIXPqjCOh0dxIshtNqgnyX1ZzRi42KGCagPfcUlz8YznjbLWuH+GnHoMT+Wu4MhVUqAfUXELyUm
n/16MaI8XpgXvAIfFrsW8+GVO4ml4UYEDYUKfBjMas+cWu8flVBlDTZH0VTxg34anWTGDpVZhBWI
rp7B32RJRaIEo1qk6wYs6IqnFRNBGbc5puwy174vqcxt/O20ikYcjiHI2UeDhWwlhe9XE/L3uyXD
C7c8Wuqrkmt8hzbbm7WjddnWjRCU8oQb6axzYtQLqW8GyjKEyRxmrMyaKxE2S8zasuXyD49Elycf
6q4+hChn6ah3IyNIgtkM25ORM2UhZ4/NBAgSitMfl/Sliuu9jdUs2hXkNNf2J5YDMM5Y1Uvfjkrg
H3gRe6Ufu20DMVN3uDxhADE/i6UJoNd54d5xEhEzYwbz0UBWWptPuFwd4uWDgHWt+77q3fgaEBr8
KldnhYfkvXyAh3yTjlcaopun+QdnckbdD7JQw2DLnP5x+lmnXMhapmAKs2dYpd0UYI3tTZ+czxN/
Q6kcITFOnuKK1TGkaNMUz9iX/wywirb8dcIUckCgkjzAZEgQoZTp5Z2XuMn+E/GuyQh6OSWMw+T/
vcNBcrwTyAqbBxl8gBFTQq6esxyDnftTMgRigQ+72cF6eirNNGHC/c9CPCQFTtnNuhPDl0UpU+ug
iIkHu+ofWrZuQepgJDrGfQ4AmiN0vDx6NVF9SGet0yw+UjIpSh3FXc8ZH/wpJ5UoIk+5CacdDPVp
EVWbVmsnb943lDHqaJLLL/gBvVT2SID9ZfnvR6+HWUxDh+eE+xTswkcUYgSWKClK5fpZn9Iztsb9
I4+NvxS+eZWSNkIZCmtUpcR4EfJCeXQHUi0eKbINhBMWfqMF8DiYSmSQ4BpfoGNBAMAdTO2ibyHW
9dttnR6gxd8h0gi3NBvfv3rlsfr4D8CwhsjeAP/JaNkXMgRmXb+rHKq3uY9JtPWaog6rxUoDR4XF
xdV+d77MO4LtFIIMEn0ZWFHV78vkzmhzYLH4K8t7HbB7jbRRyaa+mhAya41d1M7pXR1QaPljBveB
4lVOJpNQb3Vghk0PSqyXm67O+/eYTI5dmdAXLrCJYA8DaKKnpcSUUQe386ysFjh9REbpCUJybLDw
+ZMEwMLUC/XsUxcOMumxun6auKl6E1jTj8fInmNu62C2MCsvZjH9ETYvbigtfVWGZ79+OzPLlPC/
6l5k78CxAgh2RkeDJL5DEcUCxqJaDZ4ONGOrsqVFeJNW/hZOHwg8Yl/jSfD/kkuyYMybV7ktUdAh
u19GxAQeZFhFGLu8QXDx6OQIu+Efn5diThNhsmMb3MVRRCpj8mUYD4dFVoazr1NEmSyDRMVuGYdW
s3PnFwZ+S8Xl4qhP7j0E80BMZagZ0KTdjZgvEuneBCkMsq7HpGo8ZOHai7ZL4du3E8E37JMOgtM7
oZ3HLWPj8DL061RuvLRKqBhvs70vdIAyV2JWf5q3wlVCCVXTuc5+VBexWVC2Yku7xlq4CLoS3pJu
kE5nDruNh0Unl5HiJj+jro+wg4CUiim5wXeMNKsoCv09AZPyYcZabMRBi2URuNz81kUGlgHAKiOX
UsZ1a0wVGJM+BCN6io3PpuipAEz/A/w4ySVVVb4DiUqim+r35Xo6ZGUZ3cZrPjIDQFktGZOMGMpU
Gw2WhyPOjFq2C1KlHLNCXkST2U3e1p0vCOcBlmW0sqdUH8g/gxBsdGiFE+qjObiWp1Z1rHPF67fp
oJsT7gR5hDwV4WsawZ+qvbNe42UAcG/qiYAPE7ypmH1KzLNJXw+r8A1gWOdUAbxR6gHEqNBQxJLd
tKQmvNRg+wHmKFy1hZf+tiISQdvJjFakZrT6tcUoMGgLPCfTqEgVNzfHHKm31B/eaO/LSYc5vRuJ
9rZkzi5g4Low0pWMbkYkUUR4czd98l/UfvLGBGitPIqKVnpJWF70eqb+xJ+/X2DTBAVHSVA4tUX8
wy4dV7fU168x8GykDQQmMsBc9UWuyRSvpkJUjz9f7AAFcFXx7EUmDn0NpJSxfSXERqOtmQpI/aWA
haWRsQkBxTkoHV3gld1DtAZY+t2WfmQbH8TmpU5Z1ftSfhfSZaoT1fRrxfkLRHO0K7gCFQ/bYz06
g5oiHzH1Bh4vjaBjPule1Q+xYf1tbWWiaGlTNT4z57fOvWT1GnAlPTJX7o+UHWagk+e3S/O6X682
V2ma4HKag/TcsWLPCdEQo946GZA69wl4ao6uKufZog68b0KuSgeuo31BcTn3MtXFmA7M+vyeaIl4
jhjlAEITT3pZdQReyb7drCWjvDPgMM7pCorC7H0IFK3uk30jHjBhJvWTSfCohanlwLxJZMYHeIRg
3Vi+7XkBtUfizSN3c/NePTxPQBS+p7xc+cRBPlIPEGOWCWBRb5UK7X10xlk9kaCpyfnfc6SCwpmj
kHL8ZpKa7xSbVoiTFSi6sJNJUN4QklOZjT9qa7jwYVZkZ6tEPHRgzp6lRx2TYRH6Oz83+lwmlBf5
quctpZcTsrbgPQ1TxarYyOdvqSLnnyOEWFHNW4wwFrx37SoX0zRslAxtWXPVssPi5kSI6VRqBLU0
HbtQghwerWG73NXYmsSLwJfeTpVf+SRdv0u2UxJ3XD5CfibZtdUqto5KX2zxKqMcdfuqHhI0IIPC
Xmu4W8oq7/8cL0c3135SaqD9Q49oDx3PXTL34QigqILcmqjqn1v3tIFH/oP0dakaPC/0q9wj2Abs
ZK2R6pBw6uTSae5KTdIJeSxKHVfpccoLsRnp4JFTb7WTvM7muTH8e5r2l0KXoxew6ZWSeZO95wHJ
7gJbTm8IrcluUGkJYb9SnZCvbr6pegk79+P8SqdO3sni9gxSUpjEgUXfhhVmbZXH9jbggcVBM624
1g8Mbeewi6VC9EBmhA0zDGm8XxdFnMSzwfPVuSddouoYPOh++Lx22XbaCMvSPirsir2hjjanbYXn
k6uw270IuFcnw/Tx0dZiCCkshJLI0nAaKAAqkSJMYmCb2NCEQEEMVNNhpgChEnfEkuuM1wLR6kKT
rMMr9Lyifn4blbz7hzZBmUv8T+QPfwlF/2BSWjxuiuECFV138vz7sIv7EMKewpK9g6KJYF5tLd4A
S71M6Rvj/CC9zqQbi/4txx6MyLq+NAIicoHzrRcZSyRE+bgVGAzHlMp8vdW7GbO7I10Cr1P/IXo/
BMOOnAozc4IJox1QfRTQpAjTkEk00pjz9iBAmLcdpo6HVSdSxs4XQK+ep/WpXS2A3bq2khySOKeP
BHgZPhXpI7DiCyn7ErecOHzg+je2c6yUSqOG/axufrYgxfjSTx6Kd7XYLDubljKWggW707oSyhPg
a5MDDMB5ChWxKNOjbqp1hWq+NPgYQTgFBYHVUQgrVBR67j9x9R8C4cqbfeQhy0jB1NzajVTz94Z8
iemr8ZgQLWWOZdvgeCeRzlDwewg4Kzgbq/1AUDofRdet9O2p5Wn6vuRsvVdPRrRXZL1XngWejCHA
H6KnZhuyla+ByiHzX41hUIKEFQvyOhZv0ZmV85i9x/nqbWh3aJauoh0r8G5RhYwUgqH0fBLtPYR8
CphlUHRchIqQ2V7U9TrQsmoSAnvAW7D89YoSUZLkIBYtSw+aFF/+UngdwIS5QhJokHMGn4/usaTb
9ZYBlLx25REhFXdkmT7kcR9me1krK3MyYVsdSLqQd/DkSc/tVKTvDX5rB7etpWzrVfhl7euVv7lR
iNvyayTAWQQTEWN7kqEmjwpodX7SwLjxocOPDF43+2hhkJlsmNnxkrNQAFfGBJzB4knAKZMW7vMH
LAaM2ngL2AQlQwgcaLXVjQmRvn/NOzHox4/M+zHWO5UjZfg1KsfqrK9TqeDbdIdXhYJVcbw/rYKl
sp2k1v9zCuiBfK4nZSySepSnFgGD3KtLrq/6coRIHWn9P/1R17TsQC4F3Xf2dtW5rTZUd3KPX1XN
jsFIFlR1rF0YiCfmmPyh7zktLkc689yWMyEiB3HosXu+tj3UomUiW7Qj/qeJ62cPBefAwWulp93C
2+gee7+Q9Defxmb5lp2G0/kzIVId92ozYTrj4wEj55gjtUfPvUU+5EFzo83n1gZF6eCk3n5+umeH
5Oj6QeFiZDdYti+qpTOM1IGEFM+1i9AdhpfedHFWqsMhB7mbPEMwuMln9WqVfnIq9gs4ygCVVd9r
NBwueqT/QH7KeNz6SVPnG45bTN8GBAuXIEOhN7OEL1Fi5T8+bYGyLz9QaB6pKcPEgA8E8jkXYbeS
QtRU3rVplst/4RAl+4zYsUt42CqNDNZ7NL0hYUjjaWVtqHlGno4Ckcgn1Notp9W9Ihe3nnMJ8eGp
jYr0rR3toiSwng7eRbRH9xFAzgasFt+fW/llpkBoLPPOdETsLHRuBnHvnJaQMrKyfZbghWlJLKr4
MoeufzFSqQAMyjV0Z1jkB4fStvs8MwkajcLC2gyhN+50pttmzazmjxOQqZoDxl4t1iJnPfOonXNO
QA6+13iXZ/6twe2IZWEbp2hb/Al3WelmNQ8kyrt6B7UtbRsNdIwJYJ9jJ2O4889qZXWm/FRmCYtP
bKgRdQqKI06mVsbXrO9Q5QrZYuXw6cNsB6uSPF/qyaAevjxJ2IHSZV9UlTTB6nZOxGZgQ2Bb2WP4
sD8rtm3K8jxv60iqVLSCr+P4w/jI/djxUKmIuqq3lumuEbjjgZqsstaE0Jkjp0hXkc2wasSI5F59
MXin2I9CEiNKS8TTv8hKtyZMcw0hq5xmYBYln4G+qVRk7Vam3BMqr6CdVcKZxDs6OYek46s41cLi
dZ6ncKF6yy2B5mLWU8phNXe3eNTJwbbnE8FSukM22HrwRSQmx8t8siaoV4I2c7XwO9yG7sjUNeVu
XghbJ+MphHgdWsyhnHqKJRJMLrQ459+8XLYrJo9d8g25Ls8cpKHo2qfbXQE+ROGvo1Adwysh3Phx
7U+4ba7gonIzG4W+lK2TxW9CnCXEn2TfqcLgIiaIPp5W1sYWriOG+eO2weQ3UgwtN+VnkIzFJYAM
Q/MLpsm21fII2kuY0GHf8eW5oqhJdBYfMeSv4gYUBKXwETg/SyZGwc2d0pPT1qk+vYgR2UNYJsJo
LNBzqkQXPDfJxberyuoyGTVyF1OIFTQZqjaNK5/15WvpKsdBUC81rlf3rHuya18qNx/kzuSQAkl7
w22PeJoPjrwG6C15sdSxIcBbTYRa1W+xG9460B69F0Zk6SJdzevqUdKTtGApoaWLPodOOOWTZmwG
NwmGibOO2iBmt0RPGPXvQ5TFnjXtr7kC9FxU6/EcfkZmn8rLPMM+MjdUIWOF8/X052Jvsu+gqa3V
EmQ8FRYpCAbHMn3uJZrLSyrgKEb0uZqbbuleZhO7ju2mgvEwFDXJfluD3hohPTbEnxEPdkY7X4Wc
6PL++Qe5KmX1mwgXJV9lbh+I+MbkOV3NgSmDUM+ZjQNjtRM3bdGqXuGR+xMMmd/vjImjdT09ktUv
hRoUHpMFV0wQp6j/YbndAWMV7iTRk3Lfmveeg4RbincSN4CP/UGPGGeh4+0oTdHZ4OGz9T7ceYV0
XQ9lVNClUs5Q/x71rP2t9Mb3gvvAhg5ZN4KYupcJQeLUNYyAMgtq1pOu3zF/QOFlvmwFOhtJMbev
47tHNuZNW8j74IwF+WNBiuM9sUS0AEz2EV7RAgGQwR/CdQdQGk7t/7il/of6oaxnR7hjK3HflhM/
DmDrK/KBIcyRaYQ6YiGKJMggS9hn1r8+tFZexZoH+6xxVYqblmb/Ufny8Y3ywnHNLlVJbElYNx2k
+xdfRyH98I/Baky02KW8tYiij0gezQ2WUqd+LqXYtXe3j/+qIaIAQ1nIj8k2a0M3t0WRI/DAOVab
ziE2NMlsIqwrRqCMmRIqqh98UyTsKEViQMfUUZw3iRZZNa0TNpxZIlyxPcG45AO5w6d99JrbIw6m
YdOUGZMxQgKKoRIblg9PY2eb/bU1vnAGTt3ssiOfrGCvVc4lbJXpKah2gj/Hd/cSoA7JT/Mxyrst
AVBNUWC7HNn5XqSAQERCvVsiZsXb3fKUfWWEvjBBWAdS5QKDyTV3vQOlqyRZF6Op/q2KkyPuUjG4
0PzsMXcA+WSo7RJvkTwHWQ5CBvj2b9adCHtQPqYdFBIjSR33KAZ3EAqtio2oGAgmtc3IgUfZyOQI
7MTZ1HRs6BsAcgTmfL+kbQ11PO7drgcovevBhfroeXXv/C60HX0rnmPolzg8l3G1psp/IuMfmEzM
w6pYlFN/gWU0kc2dO2T45flvYcvqo2xOwz9++FDHLDQcZFFskrskSZzzLySJWnaC1SFsgoNr4jw5
Mqa55kXXOnS/dyQVioRZS7GGRR7x2jqaCwNzNoJnF7z90wipoH52yUmcb3HHdIsvH9RcTSCs0Dqe
7No6O0kiedbMncXI4tD6Dy5p/i3PyL6fAEj+gKZDFOoD998c598+krnzqM8OJ+OFm38eyN+zbXMo
YwAQ4vR5UDz89t75qQp8JsX58DkAWlQohOfyouREVW5P/w25nzezHD4RYZo+ybvN7FHA/u85GU2Y
xotAQ8eXq8k+4YtNNko0i6YmYRFcv0MkDdk4IU25KmBko4iREmeoVTT609rpsvVk8MaphKdwNv1q
6I+NeXMI+wGgp6o6MV/PfqNn3su3QKmGcFEO1BK8BcipL7kQhB1gRUZlqK6jfSJVLaHsMO7c/vQe
LC6akjfG8LjVT+1YywBOuU+oU6rcn7QbwT+p+xYCACLfmU17yK7/HVh1/BIjNWIggHfDRztcHwYy
O0SZsuc17Pjj69kQIdl5hfU7a6ipJMgR1HKcGVMpvifv3RsTXDmEYrFmZHnhOgnwloYXeWI7TDX4
CsGnAvX6izv97coEX6PyLVkCQ8P6uXn9PUzxPXvoPzkbkbHP3GIkxTNd/BDAGYzzCn6gXu3A8u4C
j/V3q2BXk9tZCsZOmPeW2+5+G0zTHlgwsq78JOss4aiK7CoOFKqtDOI05cdQiOk6WgvOjFYoT18U
VaVjEJ7B1aSe5l2eNXLcRhmRT7KIcTrOMtfkEJ7KpHfKSc1ogrPL6KM0V5oewu24l6M666g+NyDR
MtBwLY7vhmyE6bqQqTt8DGHhb6j26Tu8Hru+CUg4B1L+xcaPBvPyMTNtNVD+DeCpG8XGAfCRFC7y
Fwh0EBqHCmppP31kTITOchuTRSapLOE2Xt/x/P7hzoKW/Xd4ouEyEM1VBIzMzpgxvFirGE3dFbPr
5A11fV6LTqDoRwmRvQRg7DiLNvH2r/cnoa00q9p+CL15T9ROu5qys4tzPp7fiKPwK+T6hoSULmPk
yEJZZaRlxcGSyTDmww3YIdd8a1Ply2T3C+W6FPTr/xIPzHF79Ff0cn8YONs+RNnjKuWP4TJs9ZB+
3KrEMDcHfbFAkNsDsPosfO0wtCyPPXs6NzXSXVW8AhjkcpJpQREOxlqYwS3TnjtLGE6SiPYKeWLG
ZzwjfxVmUeflwjpyqdEfC/M40b8YKOD7WdHfZFcA8C/IrFdicNDUhhvw1AvW+y/YUMNyPslFJrGZ
TqOQtdPgiSth3n8QLd3EbQHHnIfP5FzepaYtT2IMxJ2uwcyQd3IogZVzHIYPvJya9GST1y3kSGng
vBT+uSL8AGMkjE+iX2leOhjNXdD9D4v8yXSFRk+cJLVOi6QxBYtfESWfR3vtNONG42c7/HwZUfY+
PqLzCuMfLf9/POlnJRteaEsTlMVRVyQELUSm5R1rMttJRzsiujjvrSr9SiO7fErHImzrZ6IhYXYT
aanc/y3XTFz8++tBx+n7/fa4CxhaVW4oXaVjoPTbeWgbGSGOMfaySxo+h2bUS2Tk/CXJ2YXoqcO/
q5mnkIablwc6NY918BT3L1RgKrm/Yj8sWRmIYiHKoNjjBUzpROoA9HSrB/3xQo6eTe/kqGSib+Lg
OCV7IrG3wne500oppT9HLQJIAeSf6AZYorDclgZrNp0xhMkteiTBQ9Uz8OEukMcwsA2eN9QHwL6l
hnw/mV3/Tr/6dpIlIJMKKoleByLiWc89QTiVaz4od/aZw1Pxlb/qn0hKoASHglZq0jV2RX40ZgN7
qvWhta4OD4ciKM/NTWB57YdMuLK9UKgzUKXUscHhfJo2ZEaWH5gUbkku3345iaRT/Wt/qh10M07N
V6i9Tj3UC5iPg5vxXDA1/3QkjnXe1bESW85NMbSGKqhKeEkCNZNeBsLUbOhS339rj4ibCqCcGogj
73U2qUKMB2trsDbv5oAkBtkcI3nixpMHzBZQ4ug2x8d9uE15R0ACD8GO4W5WaztvVJwGWCJEAuL8
bOZKugxxDrFQknhw5XwVQH9bFQMTIV6v34XK+If51xCf8geJQil1ngEOys+wGKXcmhzoF+jrtQqU
nFGZXHVFFNajAC/M0lLZnIKPZwGTOiuBX2q5txO0uanPtQz/ArKZVFmkqTv+xeZBLsJsE1tX3gZN
BfJTshvByo3+aojAErgFzz4vueMWhRUa7nC/XysbsWt78cljCuOtHLZOVyB/CALDLgScrR1eYfyv
11htynt/LrucZw3DW8skXnNY9v7DXvH7HVgZQ9Md4hDtpF4OZ69qNSPPei+XyB+XYzB/DABnbTlF
VYo19GoLYjJvlVLfw7dvMvjq5yjOvbLBHm/kLqYZ9upD8c5zMDG5FCS4MYhs9WNl3OGiG7SV4uoi
inuyufcNCoNvePdgsZXCjplVN/4S3iAkc89Jrt7g1zroP0xGwf6c7caK2ajetmE1Yrl1d+8iEQwl
fi4D03dAPfqB0TbDIcdQa9d9MvW7cl9pHGrN8OqdAnv3g1RLefwAVz4PluhSFc6CcVmSjXpjDm05
HxNlz2kuN8D9IG3xRPRfWlnbLKoVUghqCphoNwfljvZY3gKNWBQDL+z32+gAnoHiPgFr13cCCtjz
gXrN0q0J2hEXTMnynbEwKtruFwgbOZWtZQND9u31LhfWF6XXnTwUtLc/N0OvClpfb7oA8PH5x9s2
oca5FblGsaEqV2bnAArYdfDs1fu2QZQksYxDhD2om43IkGRuUji/RRqQhbDYThHajELqFsQbJWVX
wteNgPpFN26zauI1KctYaD4sHuEBcQ88YCHvXjjIgtiR4/pHymG6+Pa6xA2ShqRAuB6VcEowE8L7
7phaAI+/bs6/tJfr/3eFczH2xcZa+Jggb0CuhCzSGzGegGHQqK2foD/BDQlpn42d2qoMeXOovX8I
q6O9OhKh0pouwhYQsGikQI0RrIKYcDeYBdO9NZuGasSSjWhxLOfURkYVJpIVgA+h9Dm+obNjSR8h
uj1fZjGiszSfyKKmbqq6KjG2gRvxY2pHYpyNGJwFy29sVyygfTldzprycJbFbgW91qEQk21Gw0/g
OBthl8GjO4p6pkFd2w+eJ12ENvdYUHAADaDef3CUPEQOX4vDl6bqWyK2ujxc4iWZ1Xzn4g+9WxHo
ctIrk+VO6sC/4Ew9DEQp63hvfY31eqlZ7wP1qEKBLar8LmGKo7RsXapoQ0zazhDIBp93VjQWjsu0
a+q6VfktUvSz2+aebB4rpYDqUBHMKn/T+O59zuAkT9fJbQRCON4owmPjAnuWtZAw0arjfTJJf7fz
rCX7PhBaFLuNl5vE9dagOjEWe+qo7qptUT9xwpdXlKoJLaKnErUtdFMwfiFPLR5vVOPQINmj/mTx
3fRxDXNRfzWww9Z/tbkl0ZJkz3xcGQ32XfFvQby/NhkmIOblAuC82g1s0tfStWjnVd3xQPf4d+gh
RMw4FCoyhRfQenKTZOhHmbT5vAObCOeNsTd769xUUcbpZm1sPAs6aC/iqmiEZPCsURBW6z1LcyYz
+fwSvyaj+mNDV1B3aCyC2OO8zKBKsSf/giBM8MlUxLW462Vwk+17wX/3Ln9Z/ZuLIJ7lOWzsRSuJ
AEAj+/DyRNwTa+gOCCoutWfHAJ1lsMBL1BkXGVr0Q9ff6iCFXvD07FbRd/biA7tnFYbXt62oGQV+
xBJ1nNpYiDHwfbvHxWHUms0HQ3Chj/u17u0flOSMC+HizI2ardRHzCwYmnghGadnhBeWtrBhxrLQ
eUW47XWibzNCL1W/epEEFeKiOQi1A9F9R8uw+2tEymIgbxunGhj8hjN9SFmjkPw3U2Egdck7E0Iy
QoddvPhIijUfIkl7cWRlb1jvKI+cQ6X1Wsh4MIOeqPbHoGclJ0A6a7F55X+eHNNs5MJ94R/Xw0or
/uu3a1YOCutdBafv8hR2SeJBnxGoq//Cagp+vkgaPjArW4txYR/o0fVB5DtfivzqyQqJ5bhtWjL4
vIfp90oZZeOb0bp/BJwr2d/fUZrXLSk7/ttkHl9RBKlj2qmkdD23TngVeMYziTqFTRkmWXTx3CGA
JTWPMQGBXAyxkPmuj8EfwVHKxWMij/nBtUQXsA47m2iAGbS9+hNaDxPEBiFW6BhaR006V3b8WmpF
Nf7r7709hIud4w/k7YDb5j1s3x8e03Y/o8p/p9PKW/ZwMIwLkwHAAfuug5Peb9ZpQWLlw7PTooRC
ER+ceru+JSpRWtRUnMtZoUmZKEZq2vlJmvIg247F71Y3tSGhg8vgTuD/uSlDLEU6QaFxxa9619SJ
zEPUGT+Du0d+VipaxWYOvVIGHXA9f6FsFC8UvyYGkMn8j4N3I5PX17zVFmuSSgrxPkYI7Kz6Kp9m
OK1Go7aW6cwHPFQTWfpF+4M/F6FlIVavv2Ok8Bb7JdEQVjAEKUMk/pvWePNIajTKRKljrOa7dQEu
Nqnq+5h9eQKVPxjWjyLwaCoMtMZYImYt8v/JVsV2QGa396fKvEZ62DxMtH6pK1rqvwF5lOUxFGYs
mPgc3BFqlY+fPfi4VetcxcCRY5pfP7hsBwPmypB6SHjgKqkH2HipAwICU/GwZMCeKSeddt+wFvbC
L3f2hxd59JKyT8Ep4qEauzGAwuwsHef0JISkSj1ZcOr6uRyV0wEoL9ULkuu1kThZQR8aGtEcDO0a
uHohTIEpLMg3XzPH6FbH9CKFY4i1UqbVI/Yr60KW9uLxYwabYxL0bUkKprut5Q1qyd8SLvOc12tL
2HCCv3KhnA27UINxdubFOtLorPiwokofD+Y2XrNlRGpoNwdCnlb+PrX/WA+IKcCTWaEf8jI2VeoU
Yod2uREknW0N9AYBUcYpi2yslphyTh3oZawAgBwVPvN0Bu9NHT37UPKd9uHtYBScvCOgsVF1cbIu
OVwLUiiV6KSqCQlkwyX1f7bifH60x7ORVnb4sdYa2qFjMXcDPgJiFEDdm+uqa7elW9PmWzTiUneE
cdXzUaAd2mha1bnjfwVkd8/lra3JD3CHB+2Kf5vVvU4NXciyLxQ1a9jtgcYwyGOuHe75B017/6ha
dohhRXzJ/RwhcwJIcsB/bTbvRUXxy6mnRgc6B6hHfYvjpIBgJmhiG/0G/mxfheBe2cA065Uysq5i
rw04Zkfe9VlpONJDw2ymBXoM904BNoX1wD1luq6dc42M/luJCcBtqBu4c+XvbRvJ3d05oZLDwVSL
3Nf21fBWeJfM4jjlteQR1SVz+80BNFfUiyTapLmKAwKK11AQi6S9yqAJWmNxoeQTNQlB4X9RquSo
CcFJaLQeXIHzA1vaPgcelA3b5HfoR+qU3yHAcy/lijR2cbyH43qnZfV5mIHw0OgvDIHHRIL+Af2U
XnH84PPoGOtZ00PAldmDzoojC1HFlst/h6pgK/cW+tO38bKN385hiXJtHQypuvtMh2JSOXAllF1O
dCsVFAK5WydgoQsNVPgBdaUxVaiWJ/x8wLwO78RiaeO/eRRX5l/w9U4CoIOjRrz9poKooyUd3320
bNbhFZHJt91Sg6FIxS9LEHs2AqJENkgrXFfO9TdWZrQV4JkJ1fDYT38AsplX2AdRdYyoUBOMrGZ6
Hym9WFi4Rq1+mdkskNDQjXdIqSJIkSU6xny6QkXRC2U/iUhOtZRMt+OluIJUV5lYdWVw5NGVVjXw
goXP5LeREczV2WGHidydlJ7+Dt+IP7Ekgr0nnFZ7x6ZCTv02CWEzNNBdqiewZdVQ87cZjiR3WU0H
4D3E9O5MGF3mKcRmV6/Exhxja/3tHJV948LcSWT/0IvYGBNTKRgNpjAvZbe7eSJZxFH42deiXOjw
/VnVRB5q1xZS8fY9V1xb57VCQ15bD1p/tn6K2wYFORhzMkGr1JKYIrvIwoc5HmFIwrHMLirpZ014
NyHRUuccXXCS3mH9XfjRdI8XgMi0tL3HSyg+p32A6JszQpizMaG1koskWlNHb5UW9Rh8O7LFyqSb
ey6+nqDeFkqtXZ/rUa0a2REfuG78I8t0s1cbr0wjUFZfRCk8jFufXC/uZNG/lGW+5jfeHCFh+fQ1
hiDFSLlzEmhQYWcgyPkn/WWXTh22dqmOWQiMyEznin9QLbxKnBdFELnVsMkiAcRg+IbRXZOEbX3B
BEDwPB7Fw7PaXhUfunrx+Uu1kStDm0ggfIM/EAjkf5Ji0tdP1B3c7RzWW/T/KzABxhrDMFfu3axz
/xdr1wQvFPYZe77Z0y5c+zWGlaavHFmTrpoIH+8BzEv1juafVEUePzP2u6JLAtgqDQJMsuIKk1d3
ZQ93FJc2O6zafAA+5VxIvqsk7MPwN7arbqmHEFl7RMKP68Wlm1UvrqfgdNozgo0X/gBSxzvEaTF9
S8PJ6eoUT5mAFpcLpWdBzEM6tsDrn0IMcmwe8w2TxQ6Gbk7WwLGTJJJ84h7MiTOCUT+sTbcGPH+l
IkgCL0S1Kb4T0/CP5lEBd7xjnYvM0gveP19wjhuRXO9xbEDSUMJDmDH/WPGhsbVkDbUBufo6/iZ3
KY3qYR9yEp1Y8a9u65eW9nbjl0KLKw9fYIKRl9eHs7v9PcB06mZMBAni3gaPqdS1RsiCpVwwTn1w
rsPzfJh0/BEIdfOMnQ9bjN0tkrHLEJB09+RTxyYzeQeG+X1c083RUcq6jd6uHKUewtdh3NySRmTy
C3MM6vyW/BUdHNr1eKXwMVBQE4hqSmqznWMo5LsFgQw3+c0EfzKpuslhk1s213py6XZCaOtrDid7
yP0XbCNZjn2Id9sRivW1+veGhVJbl3gWVDNQYwgh5ZOlykajGjexL8gOET+rJr6NAt05h9kyejjR
qGb1UtpHjrlrepFGFWNCZSax8QUy8kvOOWODd5fIB5Tm8t0E6Sp0rHHOjc9/iwnX3w9wo9OgtRDp
Sap9WaF33/VQ9Cigo0rO0H9oKKBl13A3gbO8QSbzTz5B2W8Xv1Yp8DoPMIQHAr73bWqkvEnB1Cb1
3w2cQvsmRcJEgOYO9yK1eSL6gHWNf6criduNboffVGIMr0bl4Lj1vh12Zj+gzSQhMpDfvrPmUdlH
y8X8YZ5rJaKcIlYJlGF+4xs34EfJ3whvFtlKfmd7M0Ml1KNtxsMTKYCapdR7uPBNg7vtahdClZOX
blLSVb1lSOx8FsKbgUgYEdbsFSRCwbUO/sK1Y7nu2yrSJQikulg7almSAmdojWXxSg91YP9HHXHU
OvR+9N3MVpzM2EwzWBK2rgeLIoau+OSSRUe0gxVJSRgvZ940ZqLZISgzd8nhnZYIDkVNejK/Sdiu
L4IXqNu0ieHAOTM/V8YFXxiY5c/Rq7vbAhcAVgStjEZYkl1oIXbdUjhxISjdxoAOalzdq1IIgnE7
Pgvk7exdcy+9QF8uv7Fi4A6iD4+Czp4vrjPGybvV4fKAv8ubF70cESqEO33jp8HloX4n0/xSpqYV
MQqIBH25kIIf4CB+o/9GujaNnD5VaK2QDlyTXrR120ku+ot4uoJf5tFGTLSIPo9rcsHt5I2u2bSu
O6SMXhbfvkz27W0mRzVq2BBDyec5s2CfQbZxchHgcm5mdTpzCew9/jnAfLNf5Q6BwDwC4PWelNKs
7rd8GK3BJ8+wSplpupSXHntusLyVFWSFXnVPKTtMA24fwFtFPwPDr/PraLI2ILJUKThY5kcWpCcf
0HWa1xWHqM+FID0RFmkIgFrnfz90GzfeYcZY13j1sBL5pQpc7AxEWB/VuAKTpo+L1uhad+f+Z6gg
Isy1PiXzLEDCqbOhBFDqXAmFhK7uNVtaeV0BgY6JtKahbQdKR+1SOtABE8Cu/+YjdvDfsWgfBqVy
yqmtL/1sVTUm4SbTRg0ZgoYqN4KdikZfxU7fvS0oZ4yhPZulvnRLNbcG9KNl7RdHMwSWInhhVQev
MbvdHZ5gwULUlXcgaHwSp+9MfF0u6EAoYPxn3vCWAZCUOmyY7DlPnfl9b9JLm8yQ4FkRLusJaLkn
WR+QNsip2QCMzEvJj5IoHgzZHub71Be2Ptiq02OneVldmESmqPYN5VDPYuXZju5vODO4uKSkWJM6
Xfof90ERa1K0cQLH0r5ORiPrmZSkVmUl+GCc2HpAPs7SPNLPihmKhZNfk58oZgrEFjzzd1+YF/wT
hs3iSvEQbqO1xDniq7CZ4MAdqO0mmJCsZ7F0klG+O/pSbcGBnU/00KGGj62VpTt5aELSjq3f79M7
0xfjpSpgY5t1rbO0hs++Aa46vdjT4QzAoucc5w2U5Q5KJasteBJC5QAiXmKNqA/UNsP/2HunSl2N
7AdhUKtXPy79khF/a4kX1OPQ8YHk4McM2WqfZ72xqJEnI35gQjqskE1YbGxS06DflB7+IkitNAy+
G18OihHuQCVIsMRpe04J/jlSDGvOWNdWMvz9YDUnc4IXatDrNLTbmJd2wAVxapqsuxMIqZfRXKfi
r8N2z64xAkJFXGJNnT9mQtPC/Mz83dwq1ZAnXldFWSgs0rh93Wq2FBZ/eaHKD0wmSHgPHQ/uMG4u
80WMBc2gEC3CVIFP8G4FmoQ/02ynbBX+g6EXXNi0csQDvIswaq0IWWc5Xjlv6hYu7jAlES17WdaR
zDXBHCdE4kxCNntTiL42eK/6Ezd0vUVTC5kNz6+EQLfjzJFljgzEOh2HLoOU+xUh7d/EuHcaZD3I
OG7aiLI2aa+jsqzgrkAjby2TrUyaeircNNxOvelSu0N9Gn0z8ELcPuurkHHa5eTYptb0nAcnja+5
Nf6IVdMu3WZUccJ6Jjh7O/phcjCjJE0LEN7Wsug7/Cjn+bl9Ij/pjDUjN/lqdEaTLWVoqxjKtSfm
2MURdvWQz0hzUzWQWXhZy54mzFVrk5PGLpx84yB+oUnO7LFq2u20AM8hYPbHGOP8gRPwH6fY/jB1
+XrGUlN4+NvaPPP5VvrmiFaJe9gxFLs6J9qFQa2OxdvGl00woT0Mb8xVBXm7m6nkcLsVBcYk7DGa
lAn3FdnvNK8ofHui+M8XHnm+n27Q0I25NbVAaQ3faIT/MOxBGOKdrWZIGO7DI6ReiwW8+VH3KTz1
0NVQTMMBTaeZqvh9NwY8oCMai4HOJwEDnSVOdzQFXY/Za2kGHXNUASuCJsLHOKiACfsZSLWskKOT
rWD5Db9dBOz2L1lclsb4mTWfTsaWNXtFCwwE5M+KgDICPVq2FROJxeCMZARKtnS0I1B1iYra51Pg
WjymX7RA2hBuQuy55Dlb9n2yY31BU32kDARK0uVHYfAxJTPELxU9hlEn7+7e6mEEfMqOmz6pA06I
BOHySXe4wfBj5DNXjvI93cvMhB1sIngw0nSpzPof6XKPyIPuE/qhcPgF99+4b2U+6ocCHY7hvc7c
kBORE8iElYCeKLWnWfN5O0Ox7G4nwWbWwcWe75He7LaDWoM+Fu96l9X6fZ4MAwWWQr+x52oSgOp9
z5oG+dcGrWm560Rw70ePOALayjjvvfyb245rmb+81swWvjD4Q4y3OKtJY05WDZUZxbmgrIL1VaId
Yfo4ICSeeqWwNT6sL6xM0QSkSu0BD8sD/7X6TPSSfIe+L5jBgFHuBL0bGSLzCQdMUe5fBJc6/Au5
dg2xvgPSi5EHRH/x7A7YF44mT4pgZtnOO3SV2V+DFKNT2wbH+tfnbYGVhJ5qY8USIN61JktWrddh
DMAWd0LE/IfuwC4lfbT8uFwHne+fnGDC94UvvyAWPmq5J260lCPXi5CrvyoJz4EnRCr47pQGanfW
4i4tVhJOHWJSljaz3YiDLslTgprXx7RncVOczAeQprGjtss+3w6Auld6QsVqLmz6W9ZMpVJhzKpR
qBf9eBqB2DBYmCNvAqaehn7ZDRu4Od9hn/Mxy2VEfMS/ZzLZT5LyvOe8W9z0VOYl1X6s8OcffUMD
rRlrx3MNpHMT3fOnLRhHnAQvCy7lbyQ+uWnhBfQ6pjp6jbpCLhgQccJgSB5iHbmlqNE22fY3BmTz
4ft3xOV9Aoakg/Xywci1Di3XwSCp0fOobQ/rAAeHaH0doCiDyOqtUZCnPcOZCIsfaf0FVPcJaYzt
R+br9LItw8yOFz48Zph2+cu4RzN8JntAvfEBQIB04G/93recX4chkNxHav7v5FT1A7Y9DGZyZv2C
qTAYdJ+LP+dleVjEMowzHnnIZfXa6YUAgz6t3cBT1R/dMnxLXCF7jn/uHlzdzOzQ02MBaURMtYgK
KexfGtfaTahSWMGqXYSGwnZlcui32ZVVE8mxcCHb0Etw83jyEPrlaFK1Y5yYa6z2kvewrQJecNRF
XHIEqGXtrM6rBd7jJt+2zAKBI1ike6Ea8410ju2lJE7eDgoJn2gfvkyuJVRXUmXcbqaBeXzwnclQ
L1X0n5p6FadTsfPPl9JjGU4C/Y21gCnsp7fcTTlOaAP4LDL/ZhHD4Lld63zvdur9ZKf0pVaufayW
teb2yGwczLmX8I3NesKSumRJk7x+ftb7/SLL4IsGI8LJLPR2A7rulnRzLjKJsXEEqAAVBmP6L0Sn
8env4U1NljEy0DZ6yni0bb+zp8bRWqIiY7lakaUZJ/X4ppNHuHYt8CgXIaNlDXssUOWWI0K8DXsV
oytfXAh3w1p6Kf45COFdCPR47M8oi17Cc1yMaMkoKFfuuBPAehluzfmtku8R5037doyAnmiT3GMp
XZhmyGG7R7lyGooLP1VUguqu0b7pIFoot8AzN2tSDnmkZw+iBsixuNrARBCmQI4DxC5HCi5ou2ep
82Zna9ELLMJ43WbwtbrutmgnOIRIBVYFWC8oat2WfGFwutOM6rJpdMTEhlm3/sism735m+nBpISH
HXp5q8vAASym1p/ixwi6K9J7T28q7x7xTT8mEpukjhYEhL4aA1w6dt05U1Hi9YPpgKr3E9Mz5nI8
URN4r6KMd/66752dOqkgB+HgEojs+v/h4TVV29aE2tsK8xql2AEr3M/UYl9Ek6K3YK4V0bEc/zp9
lFoskALQcdphAtvShMBx1Cs9C+hfzhVD8fP6/4vPAdAtE84nG8xUEivQDuuDwPUMJRlpUchDDPMo
BvND+K5rmUK0W5Iy5ZnclVaaqX+SnFLWpX7+mJYHev90NcNzlrpqn6BbbmKxV30aaa+pbbbPELE8
z4nrAaAPBbejkL8P55ToHWSrkbHFhlPZUDp+1ljjnYrOn3eP0G/hI+KASvXXIFbn+FboNzwswq4e
wU4TZb0INrUJ/7FfRIkozdBHRNlXvnv4sIFg+jA0tGYrOaw9fLzCqnXHqSkZG9KDBHY7ysjO0F0R
WqE6jce/nzzSlVGzVXfcaCZtlK5JK39f2R4GwczVbVAyZk3/nzg26JCOWYqncvsWDnQsO3liWnPj
KyVOYlH4PYTM1yj1zsyqdonMiAAzawrD1bpVtQBq7CRaKL3RpsJ428qEdJkJ8sP6QFf95bngO7c7
byWgrflzHK7k+98utQ6zGBjJJAREr+Q4oUekUr3fkA11Uojcn37mbATLWjilrHNe/W5svQ3rSCFd
QIkT38tyOTyrxrMsdODeJqZc7Q4zkHLqQM510tItZmvXWfayk761DiGJZjL8BOI2CYjyHT8VIVMY
8KEtNTR51Sfu9UFJRBcOfCVjGhQRoMtAmNvNvrUa6QNGY5bKabyA0U0fnZNPYNgerGTM23oWPi7j
gr+hMjo6613KqACqfgocDtyQW+C2Ife2cKkIl3Of3u5VHexYvFNWoUrosNQUKzBA5qlxMVd3+ScK
6IEfYrIWPyxJRL/G4fkqeBiJrK6IVvfBmkmYTqJ1qP1R+BRIlKrfCCxvlYaRy/Rtb8pGnI5TCyxF
1sc9QGf6Q3XjZTpnHvK4/QUwRCbQJq8fvAJJzoLtb6wOOzWyqkiZiW8URBiIsotmSdColiY8sTYx
CyU6YrvClLo8M0HBb9YX66wq8K3gVVKoB4aGY+ec6UNi8ykHMaGLXeOyZe/djyY56n+qDDXjqEkk
SwL+DnW87OezQ6mBh/yVlPHNdLpVYzk4/3nFC6wHGyGqC627jIoPSN7jcfYuuBw3HIrItaYLW9lS
f4i8/bFF++t0V6AMwbn+FWYgE/dNtHQo0VXtB3XBqXXLcGSMIpLSyskufrITknJRLhkrk1JMnhDS
hIRbQpIIGwFYErhpASTBPQUlq/UlZh9tUYZIqbYIBA+UKx5vNwMSnb3jl1/bLk7ZJKtacVIhqRdW
4YG2lIxMb5r26iMyHzr6sMwMqAbAs0QtfCxbBITatlft5vWXbGOmVnUoN61NP3UFtYWkX3b+kWvk
aazdesqRYMLL1MrTiOBUqGdoQMosyj6ZFjWh0mdNfbIQS3Fog7GDBvP0JrGgzX0es0+kItyYsEMh
y/lEznJSVA1pCbC+mbegIHRtTC4EaikspXCIND5C6NFdU6Nnu9+k4URUrJu77X5Ckyyv9lvtLfWp
QXfntp+Eq16h4gGtp0NnMm49eKiRhOKwmYFFljH5PKDTJstIz6V91nnqqMcFinqd9KiCx/udL/Or
lxF6xqTHg+uAd8qTAFkvLQyMI/9PadIR1TOqFxFX1rXYx3WaQ4k5xfbdRjroRmcpFieb1UlQcN+4
IxLDVRUbZ4xjkPNQj4MiMMZThGbm33+HjFbaf4ELWCyCE6vURZ/svRlHgaPGA+RU+lp+uNI2rYGs
aESAGdaHtCihLus4/W6wl7DmKjuwoZD42m96kuJVu+Za9V3fuB5c7wu0+5xri9fwBNkk4ZKD0tv8
7nbnB800fHYu+KMlFbJ+uYLAQ6OuahmFz4ajS4gArzBjjRM2iDvM2vyzX+09R78qXjJeCnNvo0uq
LwOxd/UzG2F3j1EX1ZGN7LMOoypStxIg/Tx6mncXZLdQ0u7b6qeuu+ZnE/sCyepeBX6Qamvr92p3
4TjdMhsEBMjA2+eL+pfYnat0u20BbgTuoMs3OMaHpffmjG/PWqR73P2vLE2MMt0IT2n6kMEVTfeU
Mdb/Bd6KahrOxoXfxeNfLRgdHZ6kfb4fiNiuJBETKbRfN8a/ohb63OttLr2cB/Tx+iQVh89llzVS
oUH6GsAF1MeY57oTEA6Q+l1CmFugFyyS65R40N+HKxCl31J1oU2JYwxbHCUnZ6f0N2HrD9I5Oozx
oLXdN09mEyqotONEkbST3FHVTtXq0wRSxwkLPJrG29UiovYIu4/Qcx4SFjAiNV8AMmhO71+AtYSY
kBI0Qv+qE1ztn3hAqYNRADmUzXLVXARh1BsURzE6SXmm8UsJlrMuDBrTBQxJs3uiuqOecAj2po3Q
chBKzgqmEZjIHXYvu79+XKOeiv4h0+WcnENcnqjw+REK3iorHITYYT1EEhwDEBiWvZpCxpHa8WT6
TTXZAl1HwCJhWG6a146KKQUN/Ebm0c3bHRpvOrYTPWGugai2PBG/jLUYPeB57R/QeLFzfOHnQvcU
/tV9pLaTNiCEy/TXaGjreRa97LNANXdq1rNhOIgJS1Vjf1D1MRqAzJj39OfvVFvU4Q7RTFEi/fDy
dS4o6wuWLs7ruY6o+1KWFCWVJm5bV8YhZ/QDmzhLLgtKqzV0DIKHc6+tw1cJLrgWOIv5kA9DBS6P
9CCN7pRhaj2+APWGBN+vuTx0rEvrbE+fGxHdZUZElX8Jp1R6WCHpWyF49VNAxz0Rlkf2FNKQ9cs7
G8HoG5hitxVe5o5Mq374IMcW+VJ8KfqI/P+5mEtpKVYTGUV3WkOu0QMB2NkGTE7h+bMO6LoRRwT9
xrM1FTSh4l/H1P9ddmKMCJZxk15EJGdo2eLNxs2lReEF8TqODHBzA/KUKVl8rVPW0x0XdvwRP8tS
1/+mgL4DGPDHZ4FgF2/jb/zEwry8gxtjOOAQkhVffWKK0KuVDN+Gm9xXtaB9jxkdAK9ZfCaQCdGw
U+UtSeGol0LuMCb7gGEGIYoeWldyLZ0fJGd7tSJn1Fn2hRwHCaGJetlecR276n9hNm0TV8hAXNQw
rghLridugJrT3VP8eFcaIEye4Ev/7q2QZqFvydgJKkhpqOe7CCiTHtf58wzFnLob+eyxvxUYcPJj
at2W4oDoKfQGz/tSa6bkYh+JHtS0vskM/4hKE24LLhF/ONRtyzZ+1CkBA9qRSe0bcP7DQVdNe3St
qso7ILMYCUvyHCq1L4Z4unq7MJAzQt7DaKhtd50Y6UDTejnil7BcqoH23uBaH5C2ohHRWjFLeRMy
OfiqJKYZQ5LyxkYogwgAQQQMzr3UX92muzbFSV4OuoyQZ6GE/sM7DCmGSyXXo0R3X+Jfr0D4W2vr
3xHapdG7w3AIfOTwWUW+EeJlPfcrUpXZK+jRhInkLTY2Yf8gRI5QerdHtNsZWDHxijE2Nc/jUf9M
Zt0NLaQau1UPdpxS3cvhAsmM42NQ23o8UlLF0EGad1QMaXIG/VuXLD6qY7Voi5AjODRSADXZLG/D
MajOm91lYb0RQypUlhtj/vb6r3pZRayG3mGfAfBdH80n3pqDa+5If8/BbBc6Rz7LvZwjPwsKKgkl
dPRgjPqMffqTckin9nni0VS/Ch279IBUtO8lRxQUsEV7GXW59vKto6iwmz0pd9Yr5mHWDSJyPwGj
puSOUWKJJBQDUXaSGL7uK6neA+yB8DX6sFG3psSjemBEd/vB/6hx5B7mMwSlpRShOvQdlTcZ8pUe
ut0Kq2TQafwvDnhU7vFG9RwztSdMKHXA8m4vgTWXWXiL4Q/W2MO75Hpvuslk2NAWZaCBpIQV5qyf
H5qlmL3F7NyYqAkgdbmVsJ8PZJsy00Zp7r17C38KrEAq4PDPSc4cx0ymP3oLMFHD7hLM51VacCju
xz3qi5+RpEZXUctrEVeifluh/NMfw0+mHpl/52n8be/Q/F5TiMtaQcwFPUoO92KusbcMLZCwbI4k
PIR+AtxOQCfg47y+Jfim+T48HjZs0r21eJMGUy/JIU8CS7WCaACafW7kQiryjt4ctfqPm/rx5FoD
6HcWWK0ufabPN3mar6Z0if+Kw0f/D1TPQtLlMfnSmuLNNhh7AuT2hdItBES/JB1risQfeCoIcWxg
cJDWhPkh4aqabwcVKvLUTuo7qV+/aOVD4grn6vI76alOFvumuZDSF6+5HPiK4ZfGZ5puPTEN4lup
c8Mb2AQ8PWaLWd3GSaWR/8s6E1Kn9pHx58LguwCiEGzYBaZvTLyKjagTvQMFJkOZUIXgeYKvi4+v
vF2pEoKFT70gvYG/XNNPUlyJsR0eaMsmsSdnPRR7G1B38jqjBd/s/7IG03WRAnTctSI18QvDg18L
Vy4O2cRLNiU5KATegfV3tHRgu743S4WrHDb5i2mLCiH6BpnuzdhwxOlAfE0g1fTi1VL9vMDJajYV
u/1WcJwqaRa9l95bD1QZW6ifhdlGyLKEj7H1aSKNWNeKpjiTeaVdVyb5TYYKbv0zB6KyltgARsch
NA1SyySAbNgLzaggeqJyCMUKAwdvjHwLKwMCllx1hRQYdQMLwJHYm/6sOc2qoTjkY4ZZiAN3VP3W
lnKB07hiAe9qVFb2EAKuvUkSg1CGw2yec6N71XlL3perunhhOpJGvxRxDhjjyj28QEOQD4ayvZWJ
DuOb20UXaPlQiO1Y5rVe167xfWIDE+bDSNLtFHyHz/1iCrrZtqCT3ztgUSPE6QWZ29A8HDMP6a/U
OP9RS2c+V/dtsTh58NCLLLHoSccCOtKaDbu6axjXv9clqqxcySI+R9h8YhaaJEayVfwE7u72mNwI
I4HfYgQB8RPiVPEWMsBmyRQwd2Hy+Qh05CREWKo9y+tfBgWCXVw9z7rX0ZFMuf7/9skdeRBiADWR
cP2Wq/A1iuiV2hze9s08oLgk73Ig6InKJ1yaQW4MR/SFeHYGhZUCnYxAaskErOx/BtlUbq0NMLxq
jzEXfhSa1m+tR3ye0nnYwGSc74GIDIwaQXeqEfksaby8AMxj+/A2QSW0FQAYUrug+2dOzJ0tl1Wz
z3Nd9KbFBDWT/tD5Ucf+fUkv/MDXJGa9sCXai31H/15AStlfVBtFgRqjw9jMXLRtLwxD4SchiSwJ
qTN7Il9Fy+iG4pT5NKYdBvNQGnKqoMFxC3zyxEduRYunHa0f8frGzcQxtXJ2Y2OlLiL6foUeFAo9
m4/6fU2fUGziBjZ8cBcnvmDNKNNGdERpTCUd8mFXw3m0lL0OhqP1iEMQfIswNCFxhineJamIIbK8
5hlp0I0SOFMbFTXl/JvmpHoyM5BjQOAHKf/55OssCiZBaZuj1py45+10hH7zzl+jXuvYZgHkKOvX
F3DZj4Vxm/dFmfYt93+VsFw9RBPz+hj+E9VyuDQt0MW/k/PFdDsTYWwu419PUpFeR0kejbI6ySRD
Kize4wROtw9hxMwyHwiuV234+TnhivdX/eTjD2ibqpqIs1JZalAkQDSx2uhtWIGZne1e+jXMKOjo
CZU6TShyhHQTdMcQECC+AUrsKfRMqNn/qCZeUQ3nDhVSF9A1Vgt1q08zUQKtYIhGgmjsLnjKKz4g
/PNuV57gVoss7fBIOilbHtTE6SigoOhbAKhwk1p2NA1z8Rt00qHVjHaRHldBAIrsWB02JikGVpCX
/804Zni7/9gKmnWTW8abC2repEpWKOCMjj+BpVjvtcSQg2QmNx+UODvcSg+6Hwz9AtJxEBhhs7mi
s+D5vcXKAyNrJYrjHQZH79CRJEPuHpa1uP5hQ+GFlP5HNVn9d8BQDreh9creb18c2zTitWGzr11g
crUsCtKBGaOAnGMVfYD2kII/E53PbkTW/l6jDcx+6kkTFV7aqjR2MR0VFgVjyC5VVegwm04IElLU
ByAM/54uxZhrpeZHIQyEmNADjurBLNIsY5SXgqSumilOAYslbZlAW4BLQbqDS17HY0kn696LnEFS
Koy1W+NUeGTK6CI1x2jfHYF6URJeRqww0M9DY6eNid1ks9vvj8qJqqlleaRsfhyvGhppnor02YN9
QC+lMqJ2s4fd94FW1RUYfTnRRjaiMflvx+uF3Rswj1/DbvbAaezjrYAM0YJTQvZqWsxOjFM9Ou6K
WC/4yVe1owDOvk8PLX4hbeDhL6jkJkv87UlE1k+i+F+XhO5LieFtMqDzcTgriGwIqtX+qVFC8wUg
W7k3z0d+2OIQAY7+wMnGQTiOIKJ3KWh5Axve4JBsQdGejEY8XAxyXRokQ0R/X9n0pY2zSw7Nqk1r
8A08Oy4KkOyA/HJSUVoIsU/zxYRIMeL91eHa32BmQUMNmNBCsLr8PxQh6Y9jdC+AXZXFlJ1aCpEV
BiSMAhSx7hMA+g6pmDFQgvkE/cpG0n8sjyJfnz8NuaQCUIIO1y61jNRsZbxkhoBZU1Uu4TBy+WGw
Pyldp5cLEeXvY3kMNQYcQJDFCXJapW7p8FnCWRSKkOHi4FeLNCeViTGTL/eSmqPOKD2B7S8O3q9I
CUPnvJ4oHeYjj3H9Zr6FROun55/OBxZRyubGgqZGKs7HoB4bNjW9EkUsNsTZJcpXIouEEg5WFsDp
i8l79MBFMLfZRvoy712kCXCsOqvUXUUce53Ub0pf02C/J73JCyrRLnyGDdttRDSPgVJ/JlKZUcKv
NLmO+bBPk6qZucH3BnINb6xK7slPiDe0yZDdTyQAs5nKK4bAtie+axzdCksEsFGI6E+kRvF9P4qs
+rSYgfnFUOI2kajQ134qONBxDIOtXVUL9rW+toxk5jQg0zFrDe+KhRIJzlCdB44W9jZfZnXz9cP/
pCdxy/U4zc9sdE5jJ/U1rDA1AzMz5LkCTzJrs2d39uZ+0vUC9qs/OrvAvmc+JLm+jYYK0pIS4puS
H/X9snaouteetG8WXKgsGV5ZxECWdwntxkEUgTAwGyYd91V/3sOpqbVF1NoAGtUDaWRrXtIeB33g
PRcMLHhJ2EyxLjsPLI6d4YhX9QK/J5ZRHQ7SzmscIdnTNkVus5ybXvzhpYUckiNSYKfvaNGOIwX4
ATw7pN+nFPbkYTCom3tXEtB4BeqMp3A9X3Hbmz9YiR9NAqi/f8WBq7nQZpInMV8FXK9CdEDx1qG0
66H3zsc+pCeMHcVg/oODJGL5/xX/93s4PU+lWzM8kNZP0dvD8D/vLGvxXqSKFdcVDSErwuWgvlnv
l/HcjPNDhjAsKaT+FvKCIZPvST+0xl6G0VKpDj99iOfEJmhPV2PT1n7xUf8PWAfOsYegSfztwFPd
PWXVs6sU3aXjv5nXRVPXnZ8kx/r4XRKtTfno+1TmmALXImXK6ty0lpMTUNZC6uBg1pI63n+Br10D
QJu0bwUF237OwdbGEA5hUSwSynw1dDlp+t7oc82KESlWp8js+s8JX67j8QIxRVkm9cdeJ+KZfMHf
6QmJXCaIDbiIELzKpdYZsSMEJDy2GMOoxvdmBX/mF1hKkyUNg0vhH9KGjNy6yEV4VBE4KKtAd08F
3jfDek2EtTvYTWxrjGpAjNN44WSSawD3+l5/tqTEdxI0nrE7UTUeQU5/qsHgHep2uOmj7ZcLuFM2
SmJRgqibmKX0018SxvWYjcmuyyX7g/PrlS7JHthPMX+dUIQDBAAkLnJzMWq3isqIgRn3wSR3MIFS
ZA+zyCSjeplq4SVUCDUqnD7fXPmB2j6Lpxb56hqlIAPlRbonJ0lif1baCIzs+alUj47tj9YLx4iZ
GNi+7df4dGNwqLWy6duzs5UBHSpXRrZarDjvoLLooF4+xVLgFmCBuctNeGIpedebsp+Tq1fhzoi+
QycL112dBG+Ne6csE1cAUtQxMKEeqZWELK1Je+qQm3+Q0Oun+QX21+8qhbliYOBp5NBznnW8sKuP
3RcrpSqAlhWcv6ufQ7fftcg57lxld6XzNgWnvE/cA26HtuLCiJjeqyxlJA3SeJKMKD/71Abtwsxn
Fx3SzbxTp7xYT446rqumdE6BKr73OkBCEgd1v5nCqbQhtuSwhD7WP+Ulb53WoVMmecFAfj5rYBrm
pGhBSXWg/FU5dkK1HCQLo//lSmUDAIjhPDMsu+IoUPikg2WkaUhOia9RGCx91Zpxtt+LDDhMfjKN
ErViC0nIdqd/+ze6q01NIZCu9rRQmJhvizoxG8glXNSBaArTzwG+sZb8O9Evg+HuRftK0MHbmDeO
NR9NgSTosP8N+qhh8vawHva6259fVGsC4T0/qp+dEAqsJCLaYKZo5jfyywJQUBb1Idx6+OUtqv1r
/fHNwpQsxWw011wBRHUcPf4VGrCoDyQWQnorygqtue2Aj/FPpQfY4v7D8yhRxLHHaETztrUWVsVO
QEGur1DV3Q2BSIdLwo6S2g6OWtKqUpmOhVPZxOpzi9XkumbEHkfAkeIhELKP8wmo51P6xtr8nHzf
e4rPIG8BFMdPMKPuKCVa2IwsqdfdzfR0ecSlGM7krzHcpH/aY12SQCiPOiAZvjDiGLH7SdGG/Wwg
ROK9+E36X/USuQfEWBeRWhyFPO3CNQWQEFi/PkGgair3wWj9lLiECnIr2l+vLJjQXW4AbzLCYL5v
cHgfPBDRbpa2gdGQuqsgq/YLEsVfnkkbuOFdJFzWODOXsS0Y9iztYz/mOcOApAAJLzqh1gN4AT6G
uUfthjkT9XjO7fjSS3EIlXbFY46YSj0eg9xE4zHc8kzcKeob2225Q+Xhv3QjqShGsWDGhnxSyhE9
dBYV1Yk/+QxedpF9cERULAqERFWHIRGmZ5m9M0aF2vWbHhKfC90MTs/UquuqNxC9Zj3uCZh07bqu
Zw4maza83cKDACfg1sWoQHfc7THZMKRzxDKAJWzK6Rk30knBd2rpExPAkkfk+DEPwLk9aDgrrtZ2
DkErzREz3iG4BXXm1qAAYPYIg/pzzqZz9X84Xb2Wzi6nk+xzeQC+rnhEMUKJX4AiDmAF10Lj3Zq8
ITmhpV2cS8Nmin9A5UaI9h9eZILRqLpIz3c5BTbR3ak3+CEB1IA0vj7vxCULzwVXaKGqOXC5iNG3
IIB4eIi/yL7dyz2+/nRX+oZHn6QN9N7OtyTB5f946aLxVKH/e+wgV/3QBNcL9D8BgbGz5tjqK9ku
q6pyprnLgM7fhlArrasX+BNJtCbxNueiiw3QN2KPtEkp/lDD4vROBFKUq3/43bsJmJ8tu12itwJ2
NzQBM5ZKYun2rYIwQYp6BvgpiwfSvZi3xywT+Ug64qiCZfVkcmGPOPu4dvNYIHf/mK6Cyutfd2Wj
bTG3Yq9ZDFyXw2jGMtwczr0Kl7HZHcTx9h6umVuF7I1r1AzKf72pmhqKD1t08PIv3ISBP40J+736
DJ2u7z+a0wqDbfoHwreHEO33UFbv8Q1kwnOZlYsuDIxw5uuMVUTItHsnuZfNAZZLkegsCP4ouPzq
uruw/vyCaS6Bay3Q72kzlrYJWBKFcvMGnkXwklimv8jg7QnWzJcpYNBsOPktTV+9DPYb32OMYXTp
I1pXzqYdo6iSvf6mDTKbJsPYYnbSlpoUOQ6bvSZmtpOnYzpmgYdYGPYfwDoEQjLVKZopV5Cgq6Uv
hs8cXkqc/MD9sKHsK83p2Utt0A/FP4HIpO67U9vvmWr5TGUeE72JPrOUtM+Kex8UjO6pay3nQYOU
jWGyyLl7RxSauEN7Qr35Mq/qUUGLr3mDRVBHjuSy7dQCNGinsxu8qN5Wld3bM5vKuwykPrwIBB8Z
cvTfZa9DJvobI2FSKtCZjh6E2IZ1VhhBnL+WZbxLgeSM8tWhhXaTHruNaSxrwvljH6iSJ9RsSGp+
OYHBqsTYROjpn2t0KMlij75f1gT2zQMODxd1BMmS9LZLVZ1xWFY6z9Tar5GEUuszdX2swxCMfsSQ
lwBozPrRIS1yNJRYAmPOYaTdlISMNqP5MCAQTtysidv4lBiIyONJoTbqlzzz5HiNQqXzqpS8jjBe
kM78Lk0KMtzqstGe7mOeD+Cqj4kG62xJz+jK3hxUYQhobYrKjjUSexwUDaEfQStkeM6VNvWq2r2i
Q3AeyF1lxaxx1+Cb5zEmE8EvxPvEP+1JaXXbp+I4HUB1tIP6FNBGcw99h/yhqWj8ubfvD3nxX7Mk
KgOEAoZCTS5/Mm4cQ2jsuCvpaWQfaFYzq4tw/GgOS1iGaoQpxRl5lsklU6+bPEwbMH4FW8a5eJjq
zNHy1tvbiB6I+QwFVcdQE7WN+HkCvSTNscPnO9h5PNmGXQ4H5D9GNBa0eoFCdSzMxPSViK/uCY57
IvZmQC0WV254XfhcJjYl+cPbjQ5cBWPtbuEREDEMU45V6Xl6DJyXeWqkzn4N0G6QlkuQlsOTEinq
yl/VhKGJunsZxNlubj8NWxlTDgpxDP8E+zOFs9OrEamHlw1sMLjcef46c9TXJ98I8IQlNvtRP3tw
70+i9gB1CzaA4PHIJEAkaZtqdEvwV0WYOOozhQj8r9IkYZOQlAeTjtgdzsKs5BbPG9U62HK0BaJz
q32tN2TU9AqAFbR0ynQEcHWlsJTnly8dz9ceadMASV7z1RyzCzSvhHl8aXdOMYjiYT4N9FPeqjEJ
xLzFYbiVcZ9HtTcjTY6htEp0XQS1h/RxS0/5VdUhEsxeqlllk36EknwaYsVB2eqKmh9ZB0ntk7BD
hTfswbIS6y3OGHl9glOqBkxHNZMh2T6dfSYxfIQVtHZ+mbgCkpXh+NKPsfzW+548akSpHp5Yhlaf
NhdVYCaIaJ4uy5wjhnRGQdNAMPFAju+UnCWx89jO7XdL2NbGzlyWPTCthUwlja2OwpCOWk9xKq7G
7umJeNcZwypcAN+PChZCD6hrQN+WYuB9dXyIeJEcSfYk/n6zj7gnf9YvN1nBW5xTwoDpKPzUSpeu
kndL6tUkFRX148DIEHytpARr78+hpeF9gUbR89F4Qt/Gvi9aYvJCQJ2Ul7BssIf/5abxIWERybGB
oxY73DNqirjTicsWYXqJdnW2Z/sknVl+V4c0vc8ouSvIG647H4y5hjbjr5aLpASRQGqO1KVMTB+x
s4CVBeJFlcPfaRZjmJg2ftuRahEFDvIQ2oo8awk4eDSPwqnM08iEmbvGXhmljQdMklPP8SyDBwb2
5q3CCAvARBoYZOtHrbt8CgQH9zxVI1hgmhrlgoVUheRkyPFC8XxnwXs5cblSWwgTBavQX9gi4vfB
tEJBSVWGxVuw1wHGNZe1X9htD9rtrGLwZN0s4NgXTTV4Pacp62Q4UBOkBTZEDVpYTHxSPEeO5UNx
JPdkxue3Yn8nhiu4fstGYI3fOKVUvwoNsPbq7NaZ7I1eng7YS3UNr5s4hztmj62NyxzQw9ct7oq+
OhZA0WRRG1RVJo23YO6z4xIfe6I7LNSdHxPF4ppqoTG2epdnSpgXlEXUlPy5pqYUKIXuoeiGb5Eb
/QSagQtNyeAOvmEtGGbuEDV3Wm26Zl3byFf12HRz9S7tXyQMtpFswVQrx4GDo7x0I+VgJpHxy3Uf
MhXvw4SHM7E0KSWnp6tsghfq+yIv4apXrNXdOukOBzB6+G7KE4+UpiXr6wBTFnvdDxn5VQSwNjoo
hFXA/BmEy+vjSO4tn6pgsf2rWAcNnpyfGBMnqS23d0vjK7ige4zWLcWFH025+2scaABhqj2twOe/
vr1ZAcfN0gKHvWDGyBMDwvyjB9V9MDECMfpc+/JAdBydJ87MPeU41aKj5wEtp5QPtiH9wK44Ydpm
DDhfhTUSbnMVFQ3V8j42ybSIGo9j0dXU8RrDbvyO293BG4lxjTXf+lw3/ig2vsVscV22o9TC5esV
0+Ka9moNHaznwDaNMA0SFOHDLu+uaeSt/VWICpO/owlBr6FWn9ZfojGU750tBOspVD3b0dzMnkCe
HD+v4s27BPsA4CgWMSP0CL87ppZAVmgrU+JYO2RI+prI2v3PzLz+FbeJsDQY2E4PYkTsiWY1WQps
0PT+x4b17Mc9OGyePj3UY0lM6HVkaqQl1Bry5vNLCPiLk8G4vQl2XUSo2+IyKg86A/IjazwNBCSW
6CB82c3CGLMr/XHHV0i+R2F/sfqr9LrlqY6jKJR8EEIJ+ErfyjdV4CrQENSQsD9sljqmIwFNfCH7
75l2Ju4yu0fQ0aR6XX9xXQHLJqTWmg14azMHIQG+/axCy6zoE4G3OFw2ZoWnvFemQdJHXBURb9n5
Rx4488CnwNQXHPt0ZdV5ViA2fLm8EAUBnQyv95+RY7qmCNGNNG1Gf5qzjcicEaenXGgn/6RtlFsO
/voIfY8Uv8sZe9z1w+UsYir4CwTo7OB0GcX8rwOMXbXUA7kDvw3lcRQzqUCwqB9142nrCeJFv55v
vYBTw107FOt99JoYFrPB3CeG9HL7CoAnbJNrGJo2uu98xSsioIpJPte8HtAqaBs8yPeRZrGlKTVo
ZcfwLik+uB7a20SwUPOAq/5wJ0ht0GR+M2cs3Rl1Q+6PWd9OMwDaq4HTUE1we0h5lfMdNAH3mGR4
sRIFUPqskDw4EY0s9lweyvZkwto7mod5MH2e53tF3lHi0nXAjgnpwcCmn/kajyO3hIZZ02vl2D2a
xC/c3nSonQQaX7hJ5tboymh5LB3P1ezSM6cN8JRi8woMP7w3xjzYsvUy2EFttC6DKH4cqAu0DPXV
o3FHq0VxPIlWUfLmArfjiKYjsvL5Xjt90eSZhwPYlR40xPtBDd1dYo6Y1TGPV5ga8LhXYF05m7ht
ZOf5jDXhhorGepfvAAmCpQCwCNS9ATMld+3DXR+jJ9+ee5oO/qUEuSdgPHgKrL7uWdOkIshhHCoD
8BRisGBshOKTMFRzHlUSD9gCe/cIojB/ZMKUgjnoM+jAp9wLiLaCVczcSlQi9NGGZfOE7BxZnvwN
hPzM1WU9cY8G5qTpdCM0IT7vMTZHr0LeMn2RA/YdygyiHsHUhlBGuhvCdPgfyMzzcKDZm9JxETU2
83Z2vLugyYs87cJ6viieIVgq16AF4wVzGGiNNcpqf41nqaFkhAQ9+XVCQhmLlOA17KvfsA6J290T
XgtJ+ardTYd7GiYYn2SVhVkyAIwJfUl+pupMEmCpC9VYL6LwjlQ7FJw3k6B/Qne4ccws28KRiOWR
atGPqI1edCJe/tz7qNXT7AIIPiuKeLg45k8VQlpfAycUQQtOUVtYRMwOrwnXTickCdodyUkLKpxV
WNjeKuihYPLS+4MVLhsUAh0Yr1Pjf94qJ2Qc7BR54c5kxXvh8VZa39yi00Jy7RNetXvC6bthH8sN
ikyU/KnUS4szOIm81IFYK6HeUJHQJKVWxEEdhn6YyFwOT26/N9HHWc48COdzpuZYgHAgcdej+31u
VVA+P2rMutjlifp8CIXcCKjx3CmeKtpqw0PYeThq1VVefuYRsLfqeXyoiKdUEFOOySCdfZb6I8s2
XDp19Vvzuznb2tnV1KoP46ab0QJ9usgoXZ0cZaqeJtjDffeOUc1I8diNdD2mHnm4wvpyogRJZRIt
FVAu9/jQi6Jlr/u3wCjGt4DW8vvwKMYm2xBNvRMWD/O+e/1QqmanksBO5uumVPa3nbwMsVkjFdak
UtgLyjQMgsSDVOlPTu3fwop41Gda8HLUzMR+/I1lzGwVhrFq1i3G1cF2d3KXg7qypcXxCBe1Wkr1
hupIb+q5K1Ht0zDos6Ihry/w5mpwpB7crb3wiFJUHVguiLX797dyWoPYeQ8S8fEcuUH9mWNg7kRV
Bb7GY0OtzPVO0seYXaO6UIJl9IVXLiHACYFoZqxmLdW+Aur1mIJp+MxDzqDoHnmRaEfW/h58jsEc
8oYO5Dnt1po7ZX0DwGkcF4I+hl2+Zr4eEdOuQhFehsjVb/6EC1QnaI4qqXtoUU1GIix6puc8SaCD
ZzF43t8vaVOejekIwwaoMeXGhajlSEGgm/KpJ6ob1gF61TzcMXh32qGaOqhiklZweI3ZPzd597SN
lnvoKpAGAUdpFXQt2DIPc2J6A7j9s1tyNRiyxR6i9e7MV/KnQZTPxtolUXgBEOK8nLTDkO8VXVHX
2rJWOKnGAYDcCtJ087A5+6VPxk4DnqG7Rhh3RELfAvSCW0KlTSepYIB2vv7Ba0gkOric5cEj/KqB
9Fxo2kwBTENTgUFX35GicP9t7pMYVjSBafAc4erT/GIIPdU7u5QqBTqezeCnBbBiAr8tVEfHIST9
VZ93cqS5i4EyQWTTEL2zpTbiCbfRnqYqVCCtMhJW/xiITIeYc8PwFZgztLdqNvGw7LqIlgQ1conq
2qr9WZgQmNci85eMFQ6ENyS4C6qnZ5k3ZQapcQJB9C8pyxsP4gqJI0HKaTzvRGLxpLynDxXaA0gw
h0rkkELPw5veZAje9RhtjqDrua5DrYRZ35EhQxTZwa8GTWbmlmKVPz9Usd2vsP9EdAhwuQaNgcni
jW1aoVOnpVNSTBLtmXsqJoh3ioTZoTHpTForhNR5Es83w4b2HBpmB/ljk9xBjUKbB1iZ040QTuwc
r67Fo+9rOqrM05iIJbC+L59ODPtsc4l0lA8X9D5Yx3idf6JUa9dUBGHd3eDzMuxV+4p4dZ/mn4qb
hTplnpylpvkNO8bl+LGndqRRI7YRTU1QjgabAleSPfcPPbI4LmzhKC0lv9MScy2AxUf/UhM5UOXp
jAvWy+qLCU749+i7wV65HAH1mnnCykaIRXORy3fppzJumUnNgS1Y0htJwVFdRKEQkmdVqw5s4vyJ
Khj3LC5GKKBNsoTvnkjqQ7nifT5xB4qaHYgVSGKm/VQ0IWswW1/5erk+IHwB43N8ZNqm9NwtJDmi
q+409I/wO4/hdZNesAw9VMqUiOXIOTfDiFWEUSl2tW0nZTC+PMrvFW+90OtjBgGRP73YtPS+hdz9
K57cwvdD63mXxkOd12uc3y4myH9vtkSTX5iadxoFUO57CJLOeT1K9hK5aaIhQBOfTLpxWEROtwSk
zbrtl4RtcLdN2IsrNvQQp0vVdyDc+qnJxH6JitjBU6Yn4n4C9tZclltufUC3BwT9CR6Aliw2g+po
P0YdMbEJAaj6ZgVvL0T8IjCghTq6xxRjTdvYslX26lfqq+wvsqbcM7p8njfN+Emahkda0hBh7Be6
9aIFOZazm2ro9mjwCmRzhVY5dCIN97KJXu/uGxP1CLp6b4kjjyZvj1O87sIdgypz47cC0IBwc0nL
VSwTQILdinqh1wb7fxtG/bwf+d8bvZT5bykhl7qAWOGaQXJ8AVPBo9mdkO6EsoiQlYh/HLsaPiv7
N/cfCprUNEguA2Buqyi5m4hFsS4mIEgqyPD0/S7/aGV4uphXIq/ajjSIVzNAjVTxK8wk7e7nT60m
XeS/f6g2rrY1sPs67bEt7VZBiNDbtG1b3nDAEczAigaKn+tNMDv8b/Uuhvhwy8NWBZxYnvBBccDC
6WbsR+xIYJwKmVHC9u8U+wojbX1/BrB5ddXXJpNrnx8EGrvDRDEh+SbPyswMcERp4mC1xB1MIsDt
bapb3i6J2lN65JTvGTehadWV/5zZnf336nLO7n5e7t9d2K6+s+82cPPzBq4AbJegJF7BOgzchTQz
1lr6SPW6GNafrJikCvoeV7L/A2iSbkVs/00vD5QKHj4EmkAPNvNM/YkuvLipoPqr1SE0f9+ShfS1
ZA/fKFOBJVMoHDywGsef/ZdHDLLDrZV2lCP9MXgpFNTPwnZmRoGPwMFnWdDtIvbXo1xddiFoFJ0g
eokM5woqEOZPuxLicgGlMaC3BECUJm0/vCxMraFc0qUdUsvShhvBJlxMg7vNx/vLb1Dz+l0BkV8B
X/s6LbWZpOR2oJETdFo/lSVup30oQJcFNSeN70Fml5NGD3mTGf5/xc/tiovL+o+6WtL3r5QM5lZu
a/zKTKeTsWZqLc5aDkoTtHAqVf1KwWE23admU/wxVgutBGZtPrJ8eJHrxr2FQongVxrge7sQcVpb
ixt1NEi8d6GUg7K3zj/PumRpQjBrFUAEFSzd5AFPU/zxMbqlUCfA9X0HSA0rMSTEPhC6vz6LiHaS
RgnsvTFgK9mbSwPW6NjYHwwLO8zZ3cJ5HBJarwidlZxyKvRn+iQR2FMPw7+KAXvAEnmu6A5yHVJN
gPxCCnvunWY4T6vBtwGKGDCu3y/Xs1Qv0EZTHLkUncz0Q4JbzgUoYE2RbWU873uhnbG+egOHkUfU
ANEQRzaaaVH4ZD3/ZGIJ34/0JtOn2ENnFgcSagmWdPG2/QfdCEZRpZyz/UFSO7cS3dP4cy862ZWK
TYXHu1c85op6Z1trz14S4NUYsXW6qM64DMWFov6fvcUZLKdQfu+aNtgU8EynOQMzevl1TvI2GGhh
Jjhqn6IsexF+O08RwTHVQR0rsit/mE9/USDZciJdqyF8GI5otp4+PaB0J8CMxhttj3wmHGqEb7DT
WhHznCJJPSHF5rE+IzWDnz77bt6Tu4v5UbZu0GWzoOjiFB/ZP0UgM1b/AhzGClBLP03i6OmqFpeT
NUd/023H7eBfSZETogDf8Kxf+9s1fx+n51Oyak+NGohS7r1dTXtMhQ+hUkMGGrRmCgYYtDdwLEvE
BkbR4Kg0mmuAhwobNjjJnJW6RbEt/rHA6RbSG4kS9qD+0w8X249NSN1odsPNGWPmImvbHUeyniDB
bjvIQfEw+SCyHIsLORKNbtrz/V5W2Ms1NWfT4s9NyxhFYyau30pAxZXFsHd/kWBNm3TzzpaFDQ6n
mlwMd5TJReqnzqxu64bZ/pTbQcVsfrYFxuU9Z+cjed3CyFcXz1IjH28XySmVd8gzGQSNSFc9Ss0X
ZdbfzMsZrGlbtchsvPAKWNPwAoAlJKbEO9KH+USjaERvdmuzEhypXFfB/L0G5x5QG491ciMP8z2+
sVw0/LD7SHoqMA+7j8RKCr7UKOC411Rj/4203f2zJZyxSM6WrLUvOQ66HSNMsxyBF11VWd6q8pVW
Ly3Rrc3mlg0s3mM/EMpPlN60ekX4AajgdeOSVgehIm05OPj/6gnLWnr6snidk8wMfhjZ6J3e7gFA
i67G9mnUFlkMJFFSgSP0D9SjdSWWD2puTxIWCbYpcEXBlMeDM2uYCpL6VybMIKL8XMzTj35bGLkW
rnIGwnn26HvLVnBYPTZHVaItKmC4FM2Op0TLxdsakC9T4ekM5RlmrTiwTJN5nT1M06M73jnHnWIp
B0VksNX5ZKNrfmQyA6Y0c43Mys2gGbCsc15pCJG2CKCLB+ksH66xxtvI8zZVSEHW8Eyh4ZbBcg/O
epbgJ4uyPKSuh5Z28LlXBh7wq7eboSvZn17tmth1PLM8daBMPE/nZ/p+mLWFBr+F1do166rpRHxJ
Q0uA2e5g3BBM7FpCEuMmN28RvV+Xcee00jRs6v2vkYFFXw/Rz/CuiFmiLeOXcgrKYJE0uQUVxeQU
7xXCguL2SoKrDt/9+rFOGAd2mA6lsNw2Ib+DXrloDYkX43Bpiayd6WYM4YHgyBO/u0Y0Ks8XxLQ0
RlVs7tH52yfHynwNLvFslQKwippIHor41X+c86o11OaOeuPXxN4VCfP5D+isKRWSxC5WW92wQtKE
co669p46DBMvslqrp2sz2vQTWXjN/AZOuZendoUCTx5ljkQeBuXiKyVHpmdXh4keDvSiJTR2mZyw
oicXi/gyz7D0U7B3p219PjUp31nxg6Y1eSTVaqpTYQ8l9gkj8lZXcEFtrbCpIIeyUSK9za5jB7rI
vGv44faRJsjIBcqZT2LKU6d1IZYnKlAZV2EHsd38/icWSyupqSHScTJJb0mrrRWJGLmKvr6IDnvQ
+qGAerr2qkrU8QNB3D6ZhBAr1P32+aMnHhO7r+zk59jiOv9qkr1aNlkg4vBDaUB0MtxQtBxFBO6D
BcKc8vOR8/q/vXzN0V7PtlCCl+dNhDAwlVmNIJs+dfABluuTg8bqQDSLW1b/9PRSJoxanBLs4MFa
P7ffc+CiSCBway39gtKCfFsg9oXsF11JFeo/KxpUgMySOagkTOIzVTnbkK1aWk6MgMASdVPPk5iJ
M+QEbr77aJmYseL6aiKYBDn/0+B7wPndv/Y7sfJNT2NLVe39c2nriisNesfcPIP+zefj8GnUIigh
OOuHu3KCc/mA0JCgYCyC1vkdr5MPltucr/fBlKUutKgWNV8VF0EKs+PqtUHXtZuUaDyYlV6iN56x
5MbgYiSKxjsiJydm0mJiJX811w3GcFbyWUL8W2A5tmTjw9WpYcqGjahYtUbyATQC1Fykx9dE+9kF
qSQfKeaXx0yJ847pdM5kL8vcDwu56h4KhQdzhTOpzt8BP18/kTQqpx7DyQIJc1Cpai2auGJE/Qc0
jfDFXiniH+6C9/nOuL4bsS5nhxuOmP9CwvMnUbE2+5nibMGfZNOPJXIsinkV13Y4B7NMos7pZdv8
NgoEKhtgCM2cN2eRR2nNI2Bqs/gCbYOYS0nO3yzGTRSlohI5fQeNnYzPUAme5rjcRChquG+wdCls
y3T0UBWs+QwKFna6kPvJpf0TzCHgRnQh0rP76GSZA8i6M2qsht9ji82CRAfD3Yfy52hy3I+ZcJyc
Kv/nLyD8Fu/G0WWG5zg1VSPEjZuMQPo2jeRflORqpkK7WGQTaW5STsCWiJSJYEQWdvvgW5TBi9xR
n/xCMn+ej6MUtQ4qJeeU6kd6sUUWbfloVFMu4oqndVLmOMAfPeX6NtcSb30O3THQOF3rN+9fkGnQ
J3w8Dj0d+7guUMUuLtVGkoBrV4N6dzG+8mMrOscYoLnPsEHW0lkEO1XUZQgXKZUbXvD5sIyM6Rt3
dDziP+MU+JYT4E5BQrbi7jlnYAltKbJUwEgwcoVyM6kmwJSvEWgjL88z61sh4Htc+O2DPeu8e67d
yxTvi2GVfKg5mKWmopLax+3ZWITto7RrKWCxC0OiH93nyF+8gRmXdNU59RFPgPs8qEp30S0afhoa
3DrAPZRhxYZkbbZ3jdEeUoU/Ym4ltBdj3pb7yU0VPMI3n+09/0fpjrj69gnx00XG2/aVvCN0O1F2
aY06jUu22Po7iPglQYwTkDWzYBH5KOao+wSIhlLS4monmv75bJQJUU2NptqBl1s681Jq46VJZ/x6
a9JAMDjq+ZmUlwzz2bg6ufudqYM1ElDiZvIjJc7Gi4V4xd8rlSK6XWmBYb9AU+DBXhlfbxrL1ANI
KTB6G6hMnuyVRBWHDUKfQidI8IXiVMJ4WxMeY8D2tf5yqzlHYCQYj9HOLo1NBcgIVs0heJQwLro4
Af/2Ff3b3+8SH7npG0BpRIm5PsTWLjiXEVkXhtXEa0PGT/3rRhK0p5QWOMbdWbsMYYS4U7EVxBOS
URUiCeocZgF2Z+YqZ193aNxxkKJo1ne3UyvXwJngliQYphPQ03lw8c/GP4+yVA2VUTZnewGhgB4c
eQ0FoGyvotYgwcx3tN8RnKsNPFFzEAMUdRe/hVrJhS4NHWLqwsqn9SgqF4v1XbrXyZt9XA3k9bqM
nGZ0M6gVu1jDm/lX6ahG94XgH1oqkfMwYAlZI8l6qNNa5TQXAZU1562TsoiGIAbdsgVExES05Rja
Vc+7YqMWFWYR8Y0MtO74edJQpJufsux2MzUYZcR6OxCWqudnfre+AecLUX5u2iinKmrM3/fG1HxD
FqT2+Kb+tMOz1zyoXfLhVyEPXXYusY/PJJzJfujwWMJaQmEvf/e2CGg1q/1DzrciGRGdTeM3+6ln
C0nKBCY4oCOM3F+VFJUkYtLuEp4K/3NxEAjua437fkWoZNgxqAXmWBW+ILi24IXh14pBd4ms01l/
d2jb6LSJ+1ZvDCcFKWQtUuLMfCA1tQA1vGetXRFbcg2pfmb3p5XJtR+uf3DN9PD0ivSD8a77m0MU
/nCgbnVZn4TZwkHT88nl/PsbRmN2pKfkFhSkFQZ2owTtTnGacyteeA4h40xVdNmMSdlP0QWjvvsa
qFahsy3MZ6kXIM+M/H5DGajYmGcYTiO93DgJ6A8dmcfP2BBg8EUaF/bdnI2jeYRJf5oFHbnIgiGb
lPyi5UR7vgansTvZbiaPJvROg+P4g4YlfNADw9845y3kB80Y30aryNG4ZIIse0bMtweRedLKZ8qj
6xmhG0U+MSQGqRsi7uZ4EXFQafCq9FtNhuj7UngSub7NPSgnP2aC7OPJWtxhzoUhryMuFByAU6Wu
jWCullpKVOe6dCxLIGkXwiqCp3idegW5KawPbntI/5V2XB53Hmx3nO1sTJHwjfz3xiKplJcwLWMQ
iHHI+wrtNg2uJb3DLQ1DJN2eIuw5HHtOXpgMpAus1pb+uCNRR1wdAmEK0eMCbvV5mJVwM1wXsuHI
5wwDMmAEjDZztoEOBUfuTaFq4N+MH4IHwQfVDCsdnugEuXHOxwwbdXPtXlTOVA8W5gzdjQG+qphv
wk0EJUQh8U9Y2qDq1vKx4Vq6Ruogg5IgFbZFNtvoLIcLzwsXaGKP5P1sJouBMDt674rMFxApC6vS
RtpxSjyfFee+IvmSsZRtOZjbCYfb28qj5i7g2l0KqFg3D+foKT3zD1XmYiQ8xK3vtxsjl2nk5GXe
p2LgnruLeG5nTqU9qc7Bc7oZ/INftcY6tmQf4q5FflNg1ucBi7cnyzc3ojaRau9l0GqxbVANOfMO
h8yRMKlKkb62H7eQzOttrC9bf+diYzTX70U7XUA/Af+3VpC5wPcuYP8QvwRe4aRhXkn14QfvWUUQ
zMGxFuoQeGJdgedhxL1XzNH6sutYz1Qa3dhozKfMRTxrgJThNZPhKnaxJWqHg4xnZkEIrv/Xm23Y
8ftptnRjM3JKv+QBw/LOUOx6ah3lDtQytr3drp6VH7iFoGVqBdvUbf8wkJ1jfshZWMz3dIWKVFDR
g7oYSrE8Rbba5T+X2grkWHbwQkw1q5emEs/w8Kb+oQE2oBP6yvumdP4da7FNa8P47SAF3lUuFmt5
uBv6kPyg84m4gQZg5CqXFxZQ9rJl2o2MJRa7WigljIs+FUMOfEtLQzaBzV9HPqWTiKxnUVm3U4tU
AiJYWTdEgqPYwiMG8xOKnx6/0DbLsmwVSTbFck5RZp37VQ6PBQVqekJ0Z1zcvUU+tx8PUI/s8wIx
W9sMYdwH7co8QIBvF408agzWcSX94u8Z7qTpA8gN/LevG/oGaBzI0D4rxHNjiHiEMxELdr5x2pxg
v0CMDlc4kuktQRNG8zQ3hLKTjUMrNmyrYpK4OWjYC6h3UPIUx5MAmCOv/pdpnvg9P3VXBNieimJI
S/ZMXUDepY7nuW9Bj3+BHUZN0LSuWtX3jtbGHMFZ7hz0pZ1CSkVZ/tQyvVNUGy65BIEnJC9HoHHn
lvut2WpKvChGIJmA+ha6csAdbVMxYbKNg//rVsXIRgUQKit7QXFdU5oRVMMoBAR1DWt975ymhTXf
wyEEpt7MVGZ+IyPWf0xoye25iMJ4ibdPhpL+3ayqGhXIh5bfHSBodtfmYd0L6xThW6FBxCkntYn2
Cxx5ZIEK6bXKNCDVsTYGWLhM8SpRf8Yw3zEF+2nSuO5Y1GOyhSHHyRXsCkjrJbcAemLPAaT7mil4
4ZN1AKoZ9RCl8lQL9KcUV9Jk9bDSquMPJDCybeDPs1L+LwkbB2bqgjhNgJy+YBF1eFkZrmcmqiwe
0FoOS2UK0T08SEDUWH4ojpnbRbs9iiQ0TYZGyUb2V6k+SnPAse5Oq9otO9lGBwwjnYS6X9iMQ+KF
AI0VOy+E1faI6O5M1dZVSNgvCZVKW0RJoZoc3x0fZMUIekbPgM3QZYTHMIyQQJ+O7zvXuRqXntzu
vcEkztVEwlW4pezvq2vZaP+4zTJnRr3aTs+H3bSOcWcz0dNXk1vXV4Hs8eAyyttwWNJhNSPFyYRd
fKcGSX85Ml0XGyMQdDG3yvmx72heSWqNFXt39tMW0t+Aa64XIeyRv0jWeUPtHVMBPXpl37bu20ZY
wx1cleoq6umpgg1jArV25iiTyxxMPCYsbsYT5IE4H2wBS4qvS2Sem2OstYmx/TD35NTon77fdKSg
oTSJLZqLfOLrNJwNNSZzJaPLmY7KyzH208uPD7+TsnW/573DLOBujTV4ESo0WtCqvxN0DF2inoPN
Y5OhEcEGP0FYk2JNk6NYjq4iErN+LX4Enu4lVrC13NiI8TtGueGLsu6g1I9HpEB2xybamAUliGeP
DeOBSVOFNmsllC8UVmRFbDdUd5zlbQocMKOXwDi+aGA8+rZJTrBxiRajFu9FJ+S5hkPhkQVFpqRq
fnnpFdCrLtrMZZfpwCw0p67wBswMiE9vr5j5weWyzbwRSM+uPy/i7qMiY+zWq2wxeR+TiyddPhV5
Bq0oTNNaoVmGZ6r6bHTnHFQcMRvJuyRvPfflryv9+V5yzzQcb0mwoo0oNZQR6TjxVUHFWKtjj3np
fv2USGuHwu8S16W9gMZUIh4Y3Gvg61dm+Al5VrgRb5Ep+5XcLFJwXxwVofjiK4un4iZAffi8BRH3
ZgyGLxvIvdXlqxYIA5DCxNrCXkCbYFDqpXx71xBEW/vhNatdGotVNUwOiq2qtrrLogN3r2ch1dtq
A5r3rnjKkXCSAIVwEVBKOALQGQ9fkEVmEqdofB97ETWFgXR9iv6HqnSC/gS3ap+13KcqkBvZF8O3
+P2qNAxBbygmTdVzJfLpOHGut3azO3exqAzVsQJ+aPwjm+f0SOj2efCXU49oaMTW+mgVECgicmaP
InsR5cJ8CsVF4VQTmFZYEeheoL2M1e7Y4qV4fhYItJU/4bFmcKcJRvDIdAqKqivZMe3aKs2BSw8p
mNRVIlCQ9lvJQQR8tyjwsH2Gwdb4owgJEOYbTwfarNsfz5JV0kVgDgSMoH+NVYLXvlivO5XqQH1t
bRqo1O/3WkEf1tA4FQc5aRnNzDUU/ZgfH9CMss2Kd+FpNyEwSn0amkGPnh+NZ+/LjTDY1qaGs1fs
VX06SyZPn15BTF7cOdAx61vspKF/JKHkDovU+UmCfFD7fF2oLqTu0HLXj0gaLLORpayGS75axdsA
0tcdYT4lquOsB2pUlZvvqmO16qdOiFevUDBptFQFGj4eDsvTI2+RkGshQbki+sW8A/zC8SIxv6wJ
OqpFsRLIsSBtQ/5m0WK+HWJQnLzsr8v6f8Z7To5Gg+R8IMuqJG019blu/rZd5vDrNpWiFOYvfK3m
UDPucGgh9anfrZV77S0vQtTCVTJ/W1+Zl2p8/wedZKlRoRgwS/ZfW2oQEh6OY85cpjm+mAnu1Okb
YOJuPLxTcodHvuGDAlfo5bx1uOQF2rKHuFr2OywER554rbpkbZPf3LvxIV4s2c9cUicmEP2xMId9
ixDwg0lmOQnHrbRs03mmMkYOeCiTvCXvFz224OdF5pVv/1tbGQiqXv/kd7qitR/4Iv+cNsKjxGdu
M02Pa+X7hyhHCKL9kuoQCH8mFj/EPyoQENZB9pS8tRgTtHh4dc04mIwg7oiMjArtvGHHdMTXBy9m
ThdCYfIm65bpedr6ISZZG3nzEhK2P3H1uPzklyl1ySckkg+4K39UAX5VEeZwJmDeXmAu1iOCPFBS
+YZisTTWUwWO7YhZoRFj/oEwXOY2bTEPBEx1+Xg1blwDnreUHJ9RhYBTZIrmW6l1ologwF4nwpM8
BkfOyEcCt1I3d/0EPSLLmmcJAkeCIj/smbr3Iks4/y42nir8gw/UPSD0d+pVVOx2SaSVwOLGghZF
NUtWOispsFSgBYuoJ5EheQN5jB2HzKbZ81WdNZpIqavPZOntzD9ptdtBZGJZ104ox4lXGZnseLSw
DBzso+gQYPEarPlxZ/0x2aGoPgO2TcHmM6UBL38DPwOk7fsCg8uaDcYwrmsMVhXhEHT9OZBjOW7P
zdynLqjb5/ppO6VA1aYymBitWna5dHgB+3Icp1aCgOq648cpmRDHs8zdmYXDnOyMDEzILs9huw9x
/HdFLAOWUw0UwYJI4xzbLWNcP/NWkQeTGJIcQv1BJExZqtdLJq635RLw4GNpxP8yzh1a06NuBOBT
1UtGwubVH4DgDgHal1oBLSArPub3TxMx5XMuQBECBcxdvWQAQKqzI32LI0qfzGsztHZmpPmNkbcW
U8jis7C0GpjLEDuO8fkoClQkVWWxTh4MsgCVdPBUUYUoP26EJMthjysnTuztO2VFdUSd5y+RJtAN
OEsX3xEjVpJIurVMQXfFagr9GGRh852tNF55n5D5GeoeslWU5W//fI/aYsM7pXVbjvWQHgMmCIT1
P6kvMe+LN2wbKfuPrwIMqZdjSAsM1Rs09wlXlm5GD+FseLwAvHOE5xBhTQjV0/dfplpAFamish5J
Py5wxLe1sueXZlYJVsYGA19C8nl9NNDnF7X2bBiSlKAqfPqf6f0d2z7Tll1Q1iSs/gmadEH2MAva
vsJt0N2lFNww32H2UJ+fHjCnzbvHn7zKsxQUksJBfIY1j12LO1CG4g7ZnIKVvSBXDpjO/4AtcLVa
QyJkru0zd/FTkdxEbi90VDMRTPEVGeB4nXAYkLxn2SjQTSiiX1C1ariCCs0iZXTdqDNciUHfwU7H
dwBV1bJ0c1WJurxBSq0I09bW/K3eva0N5AOugc8RJt4WGlN5Tg+FNhoisCnJ1MJvmYKf5U7sQ7rh
OLcwEcTsbjGVsSQ7DTKouZVsaPWQ1Fb8kx8Ct0K+GN/ClGAtS3et5NL4AhvFkL8cP8TUEmL9bJX7
CZrAJclTmjuCwfcANSUi6xybTvyGIftX2dsRb59KYNonlwF9P0D+xpdf/8VIwfDDYnQl5t+9mqBL
+FON+5C26fesLoUALhDyLN1QGcMhAqj6tXBOehpyKgGdfE1tgFKmtzKRV2ZH4UjZ+Q6HsYio7+ww
+14kE2TX0wG17O+3DUbUdaxMlPkD0qlJaEzW0hxCaAsExrNEBR4Dvo+Q3zjozZHFcCs8leArLLAx
w5p9Mr5YeM2fyYUcXitNKAUzP5G8unsq2SmwpERfNjEN8uo02/1ggQ3DxocBZEUU6sKPUvddaEB2
Mby5u/EeTDWJ1kbtj/nEFXdAtu5WwzYh8Nef4fxiNSA3pOzysCH4ssSjIyZl2DACLKBy6BOaZQa6
XL6Ks1Y7juAv5XXgnOLkD/7B6Ksu1fDW13JY6mFpZjrJiBRUrfxiEl7iExAUrihbAnQrqNLdUyJa
YkhCCeuG75mQTIkmkPgmQ3Ub0Y7ecJeSj9zN4hht1212Pwt9ZuLTiVGNNRuavjCTV+g2ncq2USYn
XofBa3L1E0deDzMlW4d67kYWAE9jZ/x1OOO9Sw0kdrPoOhiErvO7WQC/EsSm4qGDNy/b7dS8Qpof
XP3gFIIeMeEsnaOqspDeK526EiokNSc9fQ0Qdz2247N+OVROEGq+gdGeAUFVOrkexbug4Wl4aCpQ
BmBxOzwN9CA1XshcfxIY3byVHOjlHn7h71SJOFtEapbEDHtTxwmThnvCaWh0EjzU1dQAJue3Za6w
8AN6ih1AwXM/b3FQ6fTYZF5p3REUT2NaoJi/zwbNrzqCVpiDrPdBQa8bxRZyZXZkfFSLNqRCRBZD
xGDUW/bjapPDHeRRfvjZsyc9RwPUg2xo9K8LHRJfjy0uJJ2geD5CTaQAT9yIABYzlXlqWAVLCoE1
1EDGRvd4R6GcZNBG2129/8ok3GR+TUcljzguko2wsq8SwGtU1rRww4kzRma708Nc8ci/dWsYrPPJ
k/AZdxb04J2Ka9uBasyW4rgb4xUXqkYf+CiiAn9INwj7jb82fSzfGDsdPnt6hX9iCiqjMjykggVN
6NPa+gc58ej3T4k/KXhyLhN3ldu4PTzFOD5OfsEAhw58e1Y/CrtYX625z/GoHJOWbyizz9GwcSO5
GkNV4sjRrAgj1CMRk0tzVnuaaj/IkRCm7EmVHTNlYOlCmRINJUbdaJlMyN8Vb1yjxBjDsTpr9OWV
RHMpJ6iNzfZaHh/VNyCIUggPMgE/BiTtdXi+zCiAkW5UZgqAkstuc9ZrV0olmANivjTtWyP4V/iF
Qzlv6BJDwT5HbQXuKvt+eIJk5OAyAYvYlnJ+0NuyyQ4n9ISzy7ZxDL8UgqWLtL/fycWXeOF7sLF/
xFRSy9xRmLZekzuFJq7EfNLY+iOzKAYGlx9ei5lGsx/kJ7BDibn3YRhtmL8Hsyuo1n9Cf/mSg5/p
/9py/Xm4XoW/7yP4NwVqC6djqZNJZ6jvL6VSHZuWMLDYgQx1Df8pYCE/pB2JJzE9TdfmWyX5J/W/
G05lc5PoOmIEVSvULjZECYh85i7wS1AFhpBPId+BHJV2+BomY+yZs51Qe3ImLe51ZQ5GKNGYpJxg
uKFj7PvrK/qAkVhJjHt/g0aVcvP5PCafsXBJs5YvPOCIzcscejwW/MRt+GVJDHIChUiVsNGpwe5S
c7JEPgGztHlOjNBr3irgsKUtxZtV5mt7HXOHgZv1JaXaMQe8dKDIUxVYW1ORpqTJSa4NoAI667Yd
lEXVBMsrhtt8C1Sil1UvwYq+AeV5b91Wql3jLpTcZD80S+5VV0eAlM+nD39Wqs6YAl/6aQ010f/F
dhFPOe79lZqkwLIg6rOevfkP1NA3EYU+sw835MbU8m/PiT601F6/foshZTYOy4iXzZJfjwv/Z/ly
rM0yhedps79xYqSk0mYYN7NOkmEyRVeybdWbM8PtSO0zYWPNSh10X/x7B5+d/VS70w09s28dM73T
D+7FyMvPPQGkpkQ9d8Gp7ppoSHnewUXz1pBWmLEjbW0jHr1lsdcJqwknBbZnOrTportktSWuPTBq
nYO0NzaL0hInu31fDj98mLeaxrWNtnfXQHuDnFyujEaLj1XAmkmqlex/T43oYQ2YqmCnDkPHYU+7
j1g514RcxR/dMk3leguEz7Z36KYKugUl8+E8NGRbhEGnUcWdmsFzIhtSzPebB8bqhNGUCKmB0HMF
hSASiONlm2/GyhCR7vRP8CgnnyyJIYyG55QYMZdUxxg8oh9i3xC0CWdm/Dh20HiW1ev+GsAYMoK6
aS1YPJy6XKUyXAXBCO6VL3vgr08g6+u+GMjdj0cRHHvURgvKtYYlI29iNMQT56Kie6LPIzH2kvLf
bPm/y2PRM+k9nxl5J61nUIvpsg2n2x4oM1FJWA0S5RH8N5yKs5VFrGyYKwfKaW5BLA2gQoYRu57A
LihiRuKDqU+cQHAujrTqhkEb0Hm4kKl7MtP+wNPqYc0nv+ufD4BRdaD6KjQX2r94U2Amj+gUIaSV
9aa3X48jkLrEjt0rQdS7RqgaGjwsUD9CWOf9o8wSOZsiO/qSyHEvQiqHgMCzK3UepUOYfENt0KtP
8ElvpzSaXcS9Jr2wLJ0SqkD6G7FwZupzZAoHwpmSl3uuSXxIEFHRCAx9DPt3A2+wPpDm/X5Ov3sF
7BdfQ5l5Pt3AM74+Qwe9F92rmE1XATei9yXtDhXt0Ibmhtqx9LnfjjOLMENnqkPf3jTbK1YOGsLs
5wv/GTeMvbAaxpCAO7wKhJCFH7EfphA/37SMg/+idwcNs12vVduElw7kYE4Hxl+YWLSj/NgFtIlo
KCRqrJ15FPbn07Hav6ccZ9js5uVzyVpi9RAQaEml4ARSnWnYJQCQRakNppsWOihlmVOXkGJmmlwM
IIo9dLTPJzvyIxciPd8Q3JecL6/jFgp+leCbqcxKO1gtlnUkhCMs9GTkdkNUH1ZZDkYd/FCaZopq
Z8xRSMsJ3JEXKQ+gPFYfmxmrpQnNzLVPQGhpMJ0MHSBNwUFTTM0qhx9HI+GnewwSuVvBJWyt7GAV
nnyyiC487MtKlewd39IUwBoBRt8NM0DMCm703e/t8+MXE/8ectKhKBQgntrY/e4ZwrZD1uVussrx
wdq5HhqM8VGgHfejPVf99YvPG8295IC5D9iBRXQPhMFbg3LPnAJUjDYRFe+tK7A0Dpllg1AAZ1JI
FwdeqfVjawHQ3oQ6RUCOpnf5Wref504XWfexEPXHM7r6Hb/WVautc6aAhwLvcL2Rb4SgRT262u2z
fMqbhUxyBY5cDLTKu1MFuoLz9O3g1lB0X2ihYKgvhCE5Pq/wcOIO/E9nLAcLHzpfpkzkccr/SOjL
C/RxM99XDXrf5pRWANUX14G4yvR0zLtEzVpUQ9u/kFkX6l0JNKDpSOIm83VGIasrkNHnQemrBst4
hoC5peMDSlVmRzVnPD9sZJnPUsCiNxnXITYM8hpt8PoaQJhdIqDmBDxhcnF0uBmOKCZROz1Vpti5
pFvkqMXWV1tnMFtzCmPXPVTO+0jDXofTIj+n5tQ2lagd2vVKXsM91epUfOTHnoj3DC207wzzq8VH
A918TmDAYyR8CpNXwnaGogq2qftTfunpp/k+bDzEjKUWIWFzeh2hvTMF/dBy76Owi8DoAPzQeBYr
YzT7+iVoWmQpv/9o7ce94fb4zWs1oZ1AfofMcLdkDQGdt5IgrJ5DE8ZH/CnV4vhHYiA/z9Peocea
uHd1soZy/yQPxaJeTvc7CORBTAGLC8LYxlmYZTU8ccxI45p24WEmgT1I2aQG44KiRS1SUggx4l73
+9RGR661mT+nQpd/lJbu/hhg3yY8IJY73spJVS/N43hslYCDHEWUsXyx0SN9QDn28i0s/9a7MXt8
o60f6S/HmDU4cJqumHWya0Us5TOAuKiLuwmW02UUgSJXSULWb/o1J3/0xoQofeAnHZnlnKd2VqcG
J32md3wZu2vgdkeZAFheQGYGDJGpvc059WqQbOEATDTb4YxuaMW1fVOfv2ywrUS0TSrgD/blRqCW
+SLybqCSxRWI6WJpGTWt80ZWz+ymYrJMd3EWlgG8S0iMAXEaehyyoMizaDqxOamBlWSnZ+OXG8rO
wm/Q6D+dFbTmdgreyL0An74vzmEEBmTyil5LAgWSDc40iMFdl3+gNlrOINUu9RUMJDikElW5F9CK
fcKPEByq0IBareYRYP+4jASGNhb2mCZQcfuAhIOYoeLfyUaaSd9nFRXOJzDsbS7YcyLWQbWkQ37l
jkcaO9bkfj5P2JbVMUIGKICWFONmvupCUSWTweOrDvxOUswRuvm09tAriQ0mjrJ/oukQ1/IEzrr+
tDihhHdYTsr7c3Gi3UBrWMHTPO31HiltKNHTu0nIBVE6jguPsghJjnjONb2AF+7zrPG3dBkUb3YQ
nxgdRvwvVJHNjDgGF3dFI7WDhuy0oS93fWOG1vuVvmCzZkxpt+5UNy60eM2CNSMQvbvXN1sblMfZ
rWxh+LS7fm+BrehV8wKJxbFXHlKi/1OOadNbf79H5OIr7Bl/HG4D/6ksav+9AB6aIJTzr5trtWVw
is4BS5ClSyuUazGa244YisS5e2Odh4PZOZdMAGvUJVT2axUIHBo4ksWqeJp7WXNv5Iz11fAcIawP
ghCE2wCXPZfTh1Ezno3EkW4bV2o2NYtFQ/XDCqEAKGEup/gzS9tcApp8zanecWTrG9tRLZuG5+VQ
CisRXwy49rCe6oR/pBFevRJPMKYOviVlVSLcY6XRGh7OnEtzmD3M0YHRhrFZ4JS4DOGTXiPEsZO0
O62m+tfh/AougAShVlag2s/yTRERSSboBNuVJb0Ojj9+Q/FaKkzVX2iMk44qEaBgizR31RjBzZ16
xfywZ0RrGf/zzOfpiulb4E2TS0lLUorVd7e852zvyvA0p+fiutlf5/Ct2cnIfwevgVfaLzqqF8kG
76nAKHJlzUhBKC3NmXnQ6J4Nsyd00UZGlfXeK7h2AL2QbEqTdTwdH11SSfWAJnQwqE7PcDYBvg2M
xAEjVpV2JeMsabs3DhZY6IHEtyR7CFQqHaEwGGlJXj4lCxtY6h/2H9GFb05Wpy5RrKVpnXISIDhq
+Mn78CB2x1AlE4DRzT+4ouQcJpZtUIcf7tM8TPZMaiR72wkWxBScxXJoFFpy5LjBs5P+iKdSMubJ
2Nr7X7kZO1rFXVq+6hvZiyo53856BWpDcO/hhU0FGDj2kIp+/jsky05lgTWVWul8tjxfzK8ovSks
93QDVIeBXzWKGD7z6qHAj13l3iJI2EpIls2mvCS+B4WG9yELPxy8E9Z4WZ0tSodLBJhPe4rQ6ZrD
EYxXXa7/GDZ+SXgyNZcgigW8spbixhNaVdF9mhD2TBGGwtLLj+l9aCu3R5SGlHUsjIah80Tztmzy
J+bv41uJQam3WbpOB6oB0y51zCWeqhG8kLwurtN2i+QFG4EG1xV/hJOWn91e/k2zzEH1QSqW8Uji
/l6Dfh+/8615CL5m+R2Fn3mdA86lM4VNyVWFN8bdr5iGH9NZnxRYxOCCU4kTzN+ymSArghwE3GxC
03lPtxHtdBbJHGXtV/KiRScaXweVZi1l45LYxzAa2gZ52af/mME1cDYzin2poldXOq8SDgf/QOiV
hUz3ByRYIbZCdfr8z/IV209OX7AX5Rztacg29+l8FF6H9S7YYQnSa9ee6wUhj+8v7A4MdzCW/57S
MCkbEFX2u4JF0DWewjCmbSy2oCxzGtyDbZH2fNjsJj/SaMcgcZ1b5PWEkGDXNl1zsCJRlJspG1+q
NoGPP8uj+L9l3/2ch3ZDfWB0NaMKMsek0n5+dt3TKsHe+44aI3OxqqQQAeEmgn1aYMbolm3VxrDv
n0p0YHkbYIsaaiQfm5tfIFQkmnnFDL76ht0qomEWNczjtWwNrC9PwjZu6q/nVfz6t4qXusYEV0VF
AQAGUkCyH6nKhpU3xxc5zhIXwnK9FJgn1WPzAe75fA9Dp0d8L4PJ/6BcK6UySVi+x+s1Rm2EUihd
I3dKup/SwTCabESI5OlxF1vfDi4G1N5gpQizyik10WEpA5KZXTDvF9probSNrDih04i7Z//BOoO6
8ShTzTHxRBw9v1Q6xCKwqNyXlKcPQm19FZ/ALNMMU0952QvBMvTpDYgscuf/KjjIHQN7+mMs7bjM
mlHMmw/X7hvNnsP4/2rHkL+ykvko23Pk5QFIG88xw856Q2GWM+QICR6ArrPbNWCkZhGT9Ow+MrMC
ItDWpHb178NjpgojicxzWF2I+gVdDHRaKrWZgbqZJEfjayR9p58+u6aEIEV/jhINwyja1QZTZK8C
CKKKcZE7tY95DrMhTWH0oXG/8qiLUBTF4O/w9zQoq4tl1CQT+QWmC5YCK383S9tGHxKvBoJm/3gf
9AxJbXAgaYUHKMnnNexjtMqU7TP1D8k3t0aCUvypO52FwIeNQU9aZ56DHPiWbF2+DsYv2KM5c/NQ
KyeHcIEe/tNSUGqmg8NSszBGE+v88uFLPzEyBDj/bqSb5xJ5hTZ15KbTzNCJqez9g7yJRVlsk81p
IRWczAuYIapjnj407PKP8DmwePCwgYYYzDaOWz0LxWuS3vC1X9BdJaShZZ4hkSSkfmY6Jn8Fqqny
kUIheYgeDVjOsTNmSp5Vqjhu1OcsbYVztaxWutpv4n+ZXojWN0aiVAsnj+RgaEIxGaH+E8qOU+sK
Rho6rNpaq99sGwsyP4XrPGWRYwA+0TDjTveRI1zepTC0yXd0Qx33hgmWp5IIdgAryiZ8Y1Ax9QIP
dUzIw/7nbl57Ek3MquWYRSuCV5lOkBVUXXpjovYdL+29hUAwT7+rMzsO7sUMZU1Y4oWzJz1a13GN
VzzGu/D6lZxJ6uIg9scHCG7Ue7a0E4YgTU1hHZtbSKEbLrZ7FQjiFwk5ED+PrRTBND2RKt/8hnc6
Du1P5yw7tlCzAK6Z39BkSYKNLGRlTfuX5GIO5MRJWWpb5DStPQaD7A+H/pxwAHDzKFShQD4oBrGc
pgemgQhqz2Ge1hGuCYK5qXU2ohf9wUFC3xmGjqQzJYf/tLmY4lM4BBviCK1cgp89750fY5ig5DUa
9F2xpnWsb5Qk8mbbrY8UUAvW1/SxVC4oz3KvmDs4Eo5cXiGlF1SAvHMqdSgU8a70VP+p+BadjlwG
fQsEvfztb854ND7nKr1vqHfLjYwV8ip5qTRDZrPP8ulp0Q0npBPmnZHT3oTVZDETRiN6rce4Te+X
pySSx08j5yzv6lQHn95iCn9pZUiqZh0POAwU2Ki6ZhYk05qE22R0iSXpz33M6o4gULUAOXX+7dH3
sHkQEgmtoZLDiR9Nc9m+khxCfPospNe6LIOKtoQt78ZJOhm6/zSOjNlujyaLkn7xwcG2GPS/L3A4
JQAzKkgo9sXniEpZ8HYV4erbTNJd7BNtA0zdgpQ2GVoYNmKR3unoI+BU8zMECcOO+bqEVeHmy1EQ
eu4XRImaF9AOkn3hS781ggd+Nl1AkLXgj4/0XxqT0yUkwRVm/ShKyKkj2KiOK7K4VC4aEPgOmBqw
RsWhnOJgZhyTi1KuRaGvFmIALIhov+QBlgpJLLgC5QYdQH75c6omV85PRoK2a+yWndZQUCWnDQnf
gSR72aG8Ei02xNIrXS18nP5JxHC+8Zy+bE0VsvlYB1PfAW3YrDDG8i8bEqOMOks7NM9aC3RYO80O
ZsORffMeIxTmRiCi8snMX3f9oP4qFJTZiuJ4IXwnOaZUsBkYK8foaju3EMVI3l9vcGN7S19G6y8p
aabZwYw4D8RDFROifVf8DDzhYuhM5OuC/XSBiks/e3AVraThVzgtfoVlnmQ313PJ0DExCTHdw1X9
uF825HP1KYjm9b5uZuPCfJyBT4BG25MVrSOdfRmj32hw+VH8bk0Ay1Gum9vpDpcE0Kibn/WDhNgY
FqfYaavneN9Qa5NIaaFmAYrOUge25vcXQuASmejfDtFm7Z879VK5oIfDL+HSCfAo7GJY+BeSMqDb
FcGl0gYTLMJIYpN12pfQeZCwNujjP5O4cqB+zTxfX2x5tch3rJ8ZdB2tQsLVNU4pgpmhBTCgWcQa
hyAuKrjfpa2lOjGxy5Kyzcpqdsm75jDRM7qvR99/jc0DTd+JK4uSfR8KXm9fY5d3MP712w2AiVet
BoPRRDoa6FbjE4XK23mm/Lmt9QVGQwMangJaff6Ti6d1lEuKqfQSOsDcPEnhnj1rIAIta9dEMjto
rpPXduW4zaoYIR0sZYBzpuMkMmQKlo+hrH8kL1bTEDuzO9gs1YIQxVjufrgKqEaoLbQfJlKKRIPP
jimJoKghMdspD3zin5BSTxYEVNJP69MsM8LOTZIqEKcNhaxRnaI6XRwwx8i/IZdl4k+fF1x6oy3O
ltg4Ngl2mUigdV1UngOkJVcc9cgVYAfJKiCbLaLrW3vZEAJo40l9JXEgEmLe/b1q9xk+gbGPSqat
QSVc03SO70C6PhbDwvG5KIyscuBSxNAKCzqDCd6jeMSK42w4Ifd/nwK9bpde9ayAyv1OIyNKaj+Z
HlymUTSd+ZFmwXSHoH55LFBVPQ/kGBWczQh0krebEpMQ3Hn+yjEjaj5YWgfG9GTWjboLSYgbkI18
yU7ETppXsda33Jv4dVbSmvy+PBC2uuYE+MffNc7aEZiwZwOFrIzRxwzoOoTvKrPHxnUchCNtzCbs
0Ia6MTtaUj/mxVPfT9XkKd5WeHlzIXh0ZOmNg3zEILz+oQXBHH/D/anbbA4l/NtvEc4vCZu995GW
LgIwDLXerXzLtiy51yZ7ztZ6n15i5XJiYvFpoShmdfWlCVGTiF3qfxd8uOkSr/i6iVHc5gs77Tsv
klNfAIWJoCPWB7j73dw1yidtD1xO+VE4xg2SEQRQ/pJ51QbRB7DBca3Gek6nDiAIIAFay4lqVjnx
FHsoSmd9yUA/ZfZAA8UlXj3SgKFdOg8D5WJHUi3978g8WiGy30Suc+YTo0Oau+uRDSEu+/uJfc/4
jSeVdSpTZ6D6K3oDEVQHF4mg4vPgW7WcbjF8QzVaEyf0f416oV4r6rNejvM7MrvuvxsJk29IeiU/
IYjth0c5RKYFt0+gIDhwBbUMEmpRJAhorLtjbbqIMMWBf+LkfJvlBiFdrX92iKBQQNgD0fynoe+V
tBBOBIXgS8GVXYfUedy4bO7quCF2uwalGP/B5MrMbBTYiMFjUCdmHokYwvoQKjtt5FkCFYZegapO
oKf3meKS05+hhhkSxGVC+aQjzfy/rIQIBMbDMqHF85i94Dh5W1864UxeepCvOK4jLOSJeIYfLo3p
kz/eh++NRsQUdhokyFqdg9O5x8Pwym1eVYWK+Qeszqa1WxRVDzGPPQJ5+930B/FK2lJzxbSkTfqY
JrdzMVAYK/8VsiTfsRBBQ7ZY76e458JF4Dh5TXIJZtcl3RwQwCVqqGanMJ5nKihs0HK38CCwPqp6
hkTHrI/Mc6Jj3eHMZmU88dIWfqJJgia5VsUmIXq5TslMh2zWVr1VtwrbpuFiW+ErxFlsrogAIfwS
PJkHnpmgTzjxQ+KwXRGXKy9HiZk2zT+hdHtPh4oFDky5OvbH3yu+D2u3kV/Mpm1h2K1PJK+3KvPv
/fIYoRpXvU969bfBE69fXgE6ItBGy4T1af6PiWVZM0e+mCYsxEEjcEQx3fepKSruZZHNEml6FrIm
iJ7i1kp8C1PilnWVHwPGl75cxWy9Bq/c6fDSDZimq2kvGMKnPaecZwVmdtfhFaGKBlguuSGTjTNn
dzduT9yjca9/rJnBGkdmkslzhxO5/9BThsd1ZL4qxZ4P+YVVBwvOcA7A4kTaLr7DjYBFgT52slBw
RpSt1DAlN8LlOE+BYV9oChxAEu/D9u7sc2j9THlFgqySXuLhgoa8+rWPjXrhQgMsHMmrjejBWPfu
KUbeXDZWO8Ohz1GFdAvj7JBmXKIePeAOtvVALUSJhYz5sRqpfluLWTCdThQzQyHdK8x4BH4UvWob
xt3OAngJtJEY91zh+6Br2AjQh0LuQHrzz1ipMHG7t1ceqx+jZ/Z6P+1r70DuKmOmiJ7NgDfdo4q8
gD6u/8XN+5n5I5eN6y1YuIGngsEDOW12snOKGnoTTE63fS0GbnQbRWkohfbX8tIR79uGiDD9kRLF
hi+cF6YjRhHcnohT6K73tF8BPfa70QC4l4ABilb90vTQjl5CtuazTZULA8/NcF62SC0IxYgvngan
gB6njVK4VNIOHpTukd7b0iCpj/RQ5X7OThSY3lqraOvbTFFqEHF/lPjRqZgddWsnIHxzq4T4JGTY
7U1F2K+zUXdMlSoHNT15hgJyc+p6dt9BT3vHudqNsY5CCQ8o44QsB+W5FA/pIXZdFmKGxapbfvqh
mP/us+yYW/lNApRy62Cm5z1Y1qgKjXB8Zr5CJyDCb7VnDAD91eBTWmMyUpyHQlnUVLqEFn9wQRxV
u4Mw2fREHjuY2Kue/NHRWrTEYbVc4Hkleit6mcsP1ApXQcRpN3Q9qtGaiS3HBeYKFp2BUC5007yv
ULWAveQ7sjjdnF8yDiNvBm+7b/bMnUsd4wTBzyz3y8LyXJ9lq8ORq6oiMFbMJ/kqR/WlKyrmgK8j
nanrLpSjgLklmF8I62kU9axHtLz6kzzxPOdZ5tJezjKRhb3dXgN5q5NuP9JdiZPEusSuB2WPICz2
4kGTgSOdbmmuNiI/cvRuNxkH5C7QA52AeRjenRem/8HDaax7x46QrMuPFAA8dRye8UkXtxRf61Va
b4yBZI8rDvhPYau8VtijBl4Q6I1hj5TUdJBxc0DG2xByBtOUZ5FMsbNJ5OetrBMoIG3EBR2TOnUY
7OMaeJFdeIyZrkzlYKlSbPi5xodfZffCI1g0rQOxdeANu2+o1nLF8b1KqYI4j2BuOXmHlVwnDSqG
XYhuTJiDTsKAwsgEGmbE2RIgMj402pc6VrQPCv5TQ8t1DT+cEhIX+VDGtRjpTmp8dqtmyD9pGqoT
l7Qcx15FeS/I+ImEMiaTSoaASHIC0JxznXmBq4yeEMhRDDnzWuK6rf6SDd5ZHRgx0QiMwTY6JOhG
I9dx56CPz0Z20O0R0UfTcfNZIm+YcjKsTVYvFyfd9TNI+yPP3UJGUR09UocgrC3gPFw7Y/qOv5d5
3uqb3FV/6Sj3Nv9GVb0Lh4pnuMrLGj3x0tqpd3WytpmD8iy4sDSR4vXXfvZYOfVP5hBROrTAx7AK
2EGJo11NKvANgql905klOE0Q4O4K8nTFcEZDzqhXld7i2u4fgy/Wrjqw6gq9PWTSaTn1gRjBdgYV
gXeF1H7RAiNkeTAYPNVcOqUBz1kQp4O12d9MO2a/pViwH8M/P/V6xccBIC+js5ipC7/me2BNe/o/
uTh1oThj1n+4v7Zt/iRQWJJCYiT1+Rkfb+PeHTNCmV1OjYPjZ27sLacTdNmb+L2BYK8v8meKbVsg
GXwnJerR4gkuT1/KMMRK+sZ7px9I8SZ/0viMJuRPe4gHC9olVYwmEY12NAEg/0ItOSxVAZczRQkw
i21lA08QnOCZPgRVEzwn4csBCVISgP8l7npxfVqZ9inwx9NRm4/ElE0TbAfr9lyuae1F5U5fOsK4
pn7wdwJFwfq9cqGaSgqdzbY4pKOwxhI2UYCP94oeFoDdsPnZwM/qs1EZvaQ6eyWW5a9yD3KiiMp9
Ox5yClHyxEjlREOjEZLlS5kl14tM/O+FwAN/6vK5i9d7eJ8ZOraUVNojGNimwPjfbjqDjbTfzqhd
ynbZNJKvhQh7WnEvNJCRBx2x0UNQUZOFcA4QMkjbwvAVPZ09ihq803C3yWkgjVDYqpe4xg5YDCmA
TbK92EPN7pCHvZu+Cd3wKi0c32VxdT6kpKmUeC5vh0g+scwwAdiN42znh5kGd6XSsteSRNHYDmmZ
XHaa6KVPCEx2VYfyZ/7GZkyxocvc7vbQwOnJsk+WQcQIQgrEIylOe1PiPicGeuE+RK5NEn/KLibg
0V4W3qDU5euj1QaA+Xj61As3HeWSs2WcBKC1MIbHq4AmCpTCFcVknSrnkXvUImIfCUGKOD7CzEOw
iPS9Q6Wnt9xnEzEEY9znlOdL71FACRCCjQ+gms775esndK8r4HrKzKzHxnfye0BcGOn0JSMrKabt
za/RzDLawxbCDDTnnCRi1UnoEDcwTelhaGo5kRbSxoGzxPTVBPnsbNqkveEkqAFC2phQxhTChHCx
nwro8cQeeKGwT5ExGcr/ePHQNgLn/55KiCgOoethccGZgykSRzzMGxZjBGTg4LWH63XF61bu7smI
DFEdefNqbmeHqcWdkeJmaY+AVN1RZ8L/TFauAI7fOl2GgpFDOiw+Ra3C/CtWu9eVUauYUhzJBTho
ceY0ma+gZ3SE8V2eFZbiKSVc0wMXOMAvrh0qROeANk+0fCKYopH1s6qL6H8uH/TGkaHwkfAKtJXf
kgdGc98paTdMNKAu8ceKMjGn+xE0mHo22BMyiQIOYDE/5j4JwygF18EHfKWpe1x9YEiYumUo345E
f843p5ZSKC7YySytKjuH/ZAbViqMgQ1ijP0URFgoxvrOTVgT2C3aOuUILRiMuD41wmiSxa8gbOy2
p0PTUmzxOQEpWGd3F+O18FrZ2IZCRGHOTl5T4CzGGTRCv1j1e7ZcqxkgM182s9Rkvnv4Y1X60EB5
/HUwNLsvMMSHMY77IA7H+PXPOT/YFjao4r8ACBIaUnd0Efnyl1pDrTDjL9f0NRjX7rTp3I/wM88g
ZP3E1T3Uh3Tqqn/7Z2O3gXjJxFS5g1SRmRcm4jJbcac1lluLO3P6osUFIZ2LLcWtcSfywev6UTsh
bigr8HWibY58Ju8QQ9HaLovjwR7ldU/BLsc1ULLY7TlYTKLDZxCJ14+tlGGNK75WWKGhgPSmcLOe
s3zliDFUa8FRd8yg4utJIzyaikRs4FQICxSfhxVaQbWSSkmTi2foK08w9VCzaylI8ppoHIqJcMUX
Wfge2qB9evpREwTvI0iZY/64VTH64kIDe4QTl40KUlyhga0JKM81xaSTwaXRWLa5200WXxZ2N8PI
yKk5Z7nB80RCdytqtjZHxYWVomGAz7ig4VPz08iwGHrTUZLDerSjWPkzSB2Z8T4kOXRR8wvUGJdX
6JucKoqW0zIHg4CIRoOhBIwJH3t+5Ff2vLYRMILfWOPQJyFhTy6D8v0EOqEyvK7p08407cetTbCZ
A8Bl+ItUn5H9wpNTY+4PZaJrkzJSKA5gAVBaZXcITYwtNFmMNgO8N6rAKMKVc9jjIKTsMt7izi/P
+PLVqELuZXN/9N0l0AEYtexMubJyNIa+m6VD0SOTwBcgsgh7yaRzcBUWIFnIH8RVbWFn+Zej1jqg
whRx5RrfEf2+jU7uff0uYNMXOCRSr59bugwl4PPcI9I4VinREOpv/31tOmWkSCdTRBe5sA+x4LsR
vbJym5FtBixHiZVQbwKZAy0C1vt2TsdIoVSKoNPCHFKkFm7n2KYaQ0wtKoFKyirVXoC1kR6y3Ywa
JEZF1CxNl/9dSi1MnlWLxslLFGdh7YwilpXzCbB8TCbtcW8sl8+K9Cf8a+PRnzqkhWtvRnlC2m5N
r7bXDXD8FfBtTBHMI5qqrP2uDktPaU3yTM8HKIjRkLb916z906t3PQf/yJa247CzOnOGfGBpCb3Z
r29zffe2lxeS2g+DQY8F7l/kfN6V7Kd9WDI5azR8FIf6KsuOwehTz6S53/r98HNKwTKRDRU6AIW3
fw0RHgBic97Pj23979DqjpCqa+w+2JyRiShxGKh6TmMmxusy/3+ulfIBDe+UA14gIk8wlNjZUQUj
DpoR/Ziwj2Y3lKGMtcv7u/E/9LNtQ8/aeK70enSOx+J9GQhQ3ZwlSap775KAH7fFYgn03uHMPcaO
VyyK9tHAi3t9jo9Wnk4kGKgmDg373QwjDdIqRqum+8j7vYeCB0x4eHm3QFiJB3IDyT7HUBjFvt1M
+EBvpeN6MZ004FfPcoEPOnUp7o7eSJ7Yrsv0juj12zyVnxEqLv+Vkfy0ijEi5lpvPyOyTZ3kIF3i
RQtwoBLQAUznGCzINGd+wAdRiCia4OP+mKm7Nvxd2bGuWSQTU8njO0CJIMN/3okbPwhspanlfoac
E46sFeAhUriXZb8ahPEGlRujzBSiiHUoYwBhomVl0WgJ0ZavxQ9zqctbu4xNT3b2dnQG9N7BrY6R
x+k72qApL9+hDucqasMzsA4jDKpviRN4gifMNAF76SVdtDtuwdnyGOGBz6OtuVCgLwIxamUZG2xm
KSe5Obz4EBVkBn9tC4x1yJ2S0fbnaruy1rB2TjhjUSJ5JhRZPmMFKuPAcBuxyLB9e3XaYManY5Rr
ioxh3t9aFbuJzmogUHxVjM5OHeNqAYQC//y01xxUVK48ClztI6JSJfUhNpJZJtrs7UgQdyzk/xrN
/3GQmrqs/YcqMgb1FtfOQXR8KGbX4RBYfRUxfYrEmXKUoM16Ab0JbGsmRVOU//hRuFI4Gvr/3pGb
2/vOsTNJGAhJ4e1H8JItOLUzJdXMGOn/wdvXSEo03k7VCSFfFgoK25BxeIPi+6HED4LiBb66dwyB
McgHjH2U6X+8k6Ts7TqSi/8EJznGpUYcl0Qhk09COE/CCqNTJAbavEdijXuFaXSa0iiAMQe/kiVu
IrcjpIHCDQK9gtXIotqCvJicQ/2aB8lVUDcRqqsCrozdPUNk7uykGVm185etoX78turUJ/E3Invn
Z1rN1qnO7KapK8NSj3mtfRLi/IcHqFtdXwOgFocODHnMPvfYTkaQ01xBZvFbr6aHUz39QBUVoaFk
+twH1h6q/kbatmrLUUdKWnJCSDx8I6rt+/1PNPDuQ5giJQ3LrSphvtxjvWJe2yx1PW9Ddnj0CJOp
XoyA3pLmTQO8FEbYVOKP6YKVUemgMDHYdgf2WZkjecxl3rYf4C7eoIy3ouXn/Y2Vfbs2RtxlV5LX
SKoXRGrCpXDcgrmRnWuGxAidVM81ZPJ7SvklU03Dyk07Moh1uBRpk1EImPv9AOViW0A1AgzITDOT
2XQBAS0NbrFW4BlchL2lotRsEzVo7tygZcD47+zZvorZAzyuEReK4jVykAsjXnqQNX+yFhMfV3X1
OI2gQ8ttgt60OTD7aPccT2JnDFC43OA+3S2JLSZ8E4GvFKQtO3l8kZFaEcJD2qhAL6/wBVJW1jnP
jouIVw0Luj0tjtdn8IOjkQE0Zn5ljlaH0eWbVajMIcTufdeFV0lOvFwa8V6nu3VsJq4sn+LuPFiJ
YUHj/YHtBehuSh1/Nh5ZmJw1ic6el9RcQx9J5ew8g12M2PrcTrR6YMFlmaOAE6P1xtjoNFpb7vu2
XOl39K/n8MYq8It25VaS+Jk2HdCt2TH4SPD2l1AteGrZblagaNpx/pLGXroOZcM31rLmbx3Bwi7Y
V5ZJFVtOSbB0h4RwkrAegepQe5fggMlwLFOyBuNRrhCpa1NQl2aPz1nJKuN0sN8IG/lPLAU4q+ua
X5BLBkQCNXocblOceWLb4eXipea7guMbeBnSLdP2n+IhO3wMc7HeChXnod+mfVjoxkWQHOppNECT
tuGs8WyUen26CeAlKsoJVzrFf9Vu2kW7f9gY7vj+dhapSdGVp2adfUb47RGj7TnC0jswiKQw64In
8SjmUTdy+uOtNOkXkrlyLg3T00lGek6+Q6uR2+mjwSaD14M9RXa3CXMlnQtkVOtgCYo9YTdt46/b
SI+9xJKMzE4EL5k/tyNO0PzIU+sgkoeWwjfPD7CCdky/V0ogcd3LPe7vPpMwJe6P7vq3W0dpTsdP
JKI+kqvYg6N2HqgmVbHLuTyl0BMznbd4PgnLiTuBWGxkKd/I2kpiucFNX5QYnKhqWIF9u83tjvQS
Ne6pQ75gzmFH64qGBODUm8Lpi8Ubvr0SzN6NfPBOfiSfCUknKqYOcfkrJosbNF6TJ9u1SDyurS76
bbcSA+9PJCF1LU24Lscys14a7ta3saKV9nTprpQT1BuMdUgCnv1ParV4duBc59r3zEwx4sruXyyo
iae5QduaJzy2rbWe4FgYIwgnR2z34YN8y4xuhTrLwrIvbs9m+s6j97JuKEI65mhu4jKlr4CNId4s
Zd1IKWHYiDG/z/yc5IFLahLhW7h2m/Q0gPVWiJj7qKYcT0/sQZD8V6bcQ9oBVqfjk0HUWtyPyNth
QiwxbJz2pVmdx3y2wo6fip5ug9Xjhl+XF/WLJuqDYF+58mFGuu0cxNGqZ/0uVsBjXIE9+KSrLAkq
DrqOrd8L1xwnWnvPXi38q6+quEQgDkll0Z/VPyv7uDoccUfLNBI0kjUmclDc4nco97cwcgCjPP5S
BJmBmogu358ugjg04R41cOAcWg+BSmHZSwKBFxflnnHY0wyJZ5drbP+ET/frlM8EX2InDGNvbYmq
kiXFvjchFtrXlRPLTQI9qOB/iwvvSvIzYMTu/Pivd9RJKtsn6v+LS6DZJRfxpnt2S1ZeT8TBsm4A
tyfQ7Ulxe/hH9bwQxTbgc25o/QS8B7jfGGFKd6oQczIoV/dCmqpwwQ1dBqr/+mwUcuNmR2YtwJji
MZXk1RFnBORMqhxvzV0nBvbNMmDewyw5OJ/E8NJtUH5I1UafOwXvab0Ap8GWWYk91O3IeX0+RsSJ
VFy6SgjDGF/dspLK2OakmxsRZSj1U8eNjhrledHNUOEQ0Ol7lfca3ZYqpJXjK6Sl4wyDNVLpf1H/
kwHhdhIUBVeQnchBHsR5SyhYYmWbPRwTAH3hUVUOcva8KG0OqhSImOzm0nKNFU5I2tyM1OXNjJFF
NxOVfkCQU09jMVRScgHVZZ3g7bFEy3KjM6FzhjMAln1EpLsfSYfuCbJPyJqDOgwxLAD9mNUe23vU
/dgf3p/dz7pOQuGjujFYHEgDD1xq93oU0bcBQnQwWId2PHHTMl1kEiBb9ARVduZg6HytHkuDswlz
MDZkscK47Qqeix2c9DkBtCQtXd1pSMNJ+DA9zb8gL4j0+U6cSSOLGDXEsqlTKMWFk+sbYpECV9zj
su72FJ5WmrfzTNix9Oii3O6QA3AZPyTmhhKrxtE3DdXgfQxbk69YKzFrlrIXg9BpUycx+Ib0QmK9
eZI2INgpncS5J9dcPMYLGgqK4RBJSy/LiOn1+WW+adK1w0z1X2Lqj9BrqE6B0Dhj1yp7MKXslFKM
NEPTBfbLJCfa3yUCgmpmT4R0tHbQy4TomiivZcyTJmXDyr09qfbKa8x6AQO/H+yo3EoeZlU3y603
k91+Xf8ZAgO0eZvNtVXg5rxHiS+1xP2nqtkEWCMblkMqMn/mlrSgEyepTkinGqcVTf3oL0H1jWDP
s3pUaI1BpOzqm0pUEEk39c3Qe1//88HBgsZCRka+JjY/WLndLls/1VVuu46ADFHr/rJVr8e9Hkb1
MmUe6gJOWszTYmVvfpRwTVUEY6uGPh02r7FDkXnyl9dZ9YIV8nJv1T6vjFO8ayMJJHSfgl+xl4nz
ApV5u6+6ZjHlYUcSrvfnyOexr2LhYJ9k++oCIPfRZo6kev4rI/emWAmu4EfSwDJgN0khhYTcK4yh
gma8GN9qoYUrukwn/i+buuUkBC7GDP9hhbN2Xho151Glv0iVmJYcwxlLg4F2O4SNAKS/rcPO103I
LDTdthLmA9DyBYz45DPPcTExIRriMpQsFNu0S6M7qXjHQ4k0w0WupJ+2Bki+rtMoKUxyL24mEG9h
kXiDdEHawQZPtjttgYHtUABakWGmrbJUc+5InYrofBmoPsR7q6mAbSJkbQh3da3gXdWLZA/NtXxO
nkeMwbQPivvDkBD9gChSkLGFRfNJlRO/T43026ZlnGj1yL135WvIx/ad52z7i0v1fz1BYpLpGcDy
XxfvGP5YJ4kqkQ64AcqVYobuFLeWS4bSQC1Os8aC48U5kqjmb5WmGF2b+pQViE5OZVf+DstUYkSS
F5DLRbTnFTpupU6VxpMLiDeHXnxv9mL5MwCC07kTUCTaYqKr/Bd7Ggck2fNCHYlymxjSu9jJc6tH
fWPLqVjiwOfhI5Z5yQMv4EJABGaSUhpcmH7leVbfhcTdItKz8w8OmZqRNfhuIfqUolb65sKdprW/
6pyUMIqXmAdcw+I1ai7xHoOd+wMLdVD/f4n6ZbdYV8vIk6owpOtgvTi2DMKoBBGG6JEVUUgyG/cG
mTGWgQVx+O4oVHfNwfgI99v30X09qpAt1Sj/KIaX98HgZQSnXwyCAio14kjx0q2P/kmytwdarCrt
50SDavC8M6aUlepN8/A2XFeb+dhNyqTyDarlbIQ22iH0ZD8C9Irzi6RBhOTs8aj+QrTVwf/xBWrb
3q71VGCCQeOCeb0te+2MAZv2Qb3ahVjqtpf3dJ2QqcEBehRulCAxQHN5Nxmb3N+ntlUOm7DjSNS4
0YlasWwRn6ashLZ9gscaX/0opfL9gNClnEOtOH8aUOx4H52YqSbFoLO7bUlnjdkZuRpPI7g85+bX
H7INbxbBwRQ/eRCST6AiWWOWjOt0+kJJXl0OXTtjmdVxgT1pn9UpW60E/5iuRBlsTIZA2cyrA8X7
uHSYLlUbDMab1xfWNriz2Bgw97yHwiTBB2Y3oRDLZYIGJDcx/L7kFuF/9UIclbW6p9hwiSyCCdNO
5bC4R8ScXudbUHrNl7tCTeZYDfwLLNg7BsAxvrbrbinOqAaX8rPCscpAoKKm9fjX4pq0MMtvEewM
mYRRQo/i++96pufKBJUpCFcRFd5GuP4F4HA3oCC9QuO7xaW1NDmYq5xFy5b0mKPtmETFN2qkM0Pv
19AiqhFKnnZrx6rTz47rViSmrmGThrTD1dVeBDdDMlFX3TgqvY2kHB5DSVFtvTerWiVEPcZaAknx
bLk17aJammE14dZLRKo+9Lqe1wWu6ftfXnJbFeLEoCr0rWO2t7KYeUn+Mm+J6DcwHM9VGtjljzeh
oCVnT9TU6YYmuvi/kn2pO8NXyi/pDHVCk3g80+9JRss8hiC2zOmRhzFYP7ZFZwRR56MQWKl32/Pv
dkffD/BPXvooMG6BXMuSxBfyj7NuTvImy25VvuR3RvH3221nc100oyD4wQPsYSo5OGXB/w4rgl60
PA2Ras+9ymFtKZr5V7FbB6I1yK+5XDHBP1Cm0x8BPUSmSsx/3t/JY9ScGrkM4TpGzF8gHIsRFTor
KZqF8yHJ+BtyCFXnGvmDdwMW/GDbjil+qxjq7nibUeEA3/EBNSQs6C/WKPBqSVkhB+5i/XTu322g
ifwyg7wCtv6fDMR0O/cU0fia3SX7CNZiQreyZm7OCU9fed63nfeySCoFXEU6t3XXWh4alXWGZjQK
7lzD47fHk+75UVE74+aduwxQ6RmObYa3E+iyYJu1HmgQq2gdVI1gs2icYePlTE4sFQ7sdFKm+54f
vNKIkF+t86VBaEI3l3H+E24/J8J2hy1KJq9hBeKHcFYwy9ptyEJEDW9R0YwDTMMGBinzk75jR4J6
bxV4C15nYY2EErj2FwOQ/RqmPPl/m6Ak4EHoU+Feg89/IJWn50IQuUlRneZmDqRxmaUJ1mqkNhQC
rrNwSzDPNRmlqtccTuF38jqaU+5misU9GoXQe1KHXO5T1IfJEPTpdw+EHzr5Cq6FSuqs5FIaii3a
n3YI6fNQpnOhjEoGIKpBIc6SeU+TBNhoCim4jsTEDh4bHx5kyHIJ2d77JbbmbEq4Hq3aM2qLh6nN
ey4D/NsjAFIMPO8+gwOGsCq799onXKKhOT2b6jVDoA/CPCdov7/edpT/cpjBDQFg/3An5l8et0aB
VYqkmTLuUwcOLmHxlMqZ8osIlfpNg+Y8TQUkW66TTEjMSFkR8HVuMsgNq9/whsw9M+Y1p8LpHH45
DA6Z/H0J/7VEkAjeGpfu8btOMC5vfTHCz55mniwCeGr/y2tj0fWlZ08yx+w1D/XmHM5Yx/2Zu/Dc
tnCbNETpvDboh2XCA7gPLqLR8gn2+JBhFpdyHMKE6hfpsP9ojO1hXLZ/b6QM/rDtVr4AqVa4CY/+
eHHaNa5za0eclQqUg2rvIywyvTdLqb8cTHX+1TUZsIwJcMzeXM+9SPw7npEzkC+awSga86Zd2GCm
4/5maMXWV7Z69dqMnIgffNBRfni2g2XNNZuruN5pefGDUZoIqqu3o1DOiCT0XL2YmfAy995VMnBX
VDI2K++gbfVO7MSCr/3i0cyeW93u8YZeTKtSG5uQ/p1M+/MWL5G8k6yj8EcUA2J4h69sWjf6S+k3
ecnr9dQzeLREMHOWazvt3Co+vA7mE5l/ypdgfEjMOnCcSyx09c3hMRpq2+02FqmXmNEGUBte4C2L
87b6jWQLKkwg8owCl6lKP99K8HeVcVwsVkqt6d6HwjBQN2jvWG9HTTSAOtYAB8OAV1WNWSRpNdbS
G8XQzx99pO0w72LcAfGd5/Klvps3O3hdnSWXGI0dMk6ZdQdXv31jgNiRmYWXJP0D5REaiKWyP5QY
tp4IPXjdPLguFSwSDSDD/F4LcLYM2V+Q9Q1x2FAJl5YVDJQxQXR7jHdTCnp9n31WYZmRRzoX1ZXB
NFRjGNiqOLwQeGfqS1pQ7/2Php7HpsSCryakW7YffpihzSXsz6051PJWwn9g46USLOVlVjYICysR
p0FeEbjv4t6HbKLv+iv+YXUfJCwUae1YurRMbYOFYC5KbBjvhiVWpVcx2zH/3+32YM6slvH2Ddkg
OTa/UmvSltsn88fCIYjGXQhQK0Uju4LCQkYte3fExuJzmbp0pKa7LW1oT6qk0SdAAMfjCmDt0qQz
dc2QVMPubNSUP6pzTbnEqhE/hgXN5EHUHul+h+UBqg3tKR3h7x+WwQFKYFKDxbjPYDA6BBcAaSgd
LFU6DzpQudn+hL/ZhLlk8xzG2bOYvPl295xkbP2TN5XNK62DOomhMOMyqnREmvVwRKlE43PaNVB4
qlVXtWWZkpA+AamF7QFMlibfIM9quRsV+pSh6neLwT5DQ384ma7Cgt/vod/dp+dlSKO4ySWLwI3+
NTZko05YwlNcCV1B0STe48C5sLe5GkRxkwZyf+9e7q0FawHB2ZdWLTUCDPlk95o1ld+XF4nBHG9f
bk5pmsc7acrByRkv4+60R2RUl5+NXiwXjmIN7C983LC64zqxzmcQ8Hc3z86iZ+KUbr4YGK9zt/md
QX976keqpVx/nkNuR7h+eV0fq3lVFDcM/auW26jsvF6fh/b9KywcfOJeonn4l2cQ+i7+6MEnvyD9
Z5cebMOTdc+lO96BaWTM1uenYPV5QYOI0I4lyHnfKnDRlVXDdDbB4qdGXArscPehRLHTriSkoQXm
DM1VVUNTMnp2t/cLtIjaOkE8MVRgL6Aylae3ic2iTS7Wqu3gByUg/rBHcFYukTGTginuTVPyYG/M
zOOH64xhXEsWAhvwLwIjXzRa7wVNsXEA75Odk4cfaXuP6bAkU2P1zlnB/1GEB3kM4KALUYhdEHqN
z8c2WxApFGVuPG5B3QvfwaA4KSj3lIbhTRGAN00E36GpRAGZ17gmCtsWnPfco7zCA3aH3os1Hrro
AIsi9dUvz1WYhmqbGEm7EMm6Ay8KAj44st4SYxBWxI5bPznyy2V3/i218dMF85KQ4KREvtvsUVcG
S67gCOa9Xv9S8bHdAtOzfgaM1YsRsGpS/iwc1bi76WsiDJQFfhVRxvQCqeHsYe+8DG00zXvXOS1F
CInr+DeT2IhJynrtrjfdC/2M9uevzNy+cG0nhD1jzoxDKaXhDSNVvJ9OSjeHDZBIHdRLopcObtnt
wQDBscS7lrJK84xAolcd53Alc8Q6VxmODlvCHM2CA7adfy8zAeiqsaAz5dJ1+lwf2fXHJCRbG74V
3PrsmCOJIXsef7wbLZb6OZp4XgOI6rDQt37QIuYxTQd0EeNMxebRYbyCnNwH5j1azu+u//IRHQfn
yN/96rMa5+qM03La8C46Z5CaNH7IZrzP4rZOuE8DSgr3uqB7hRv97cubFzqJeW0f934jkJJKyJYu
74WPa01avhImNOhouMbrNs+YBGKcnKElix4OX6sswWsEcZZ0Xe54EQZbPMWvSiZKloykKLegvh1V
GcaEzJfWRgWSlFQI9Ksb6taeA0wWj7sdIubrPbFixiF8gY9+Qya+NJ5TfU0bDJhH21OAsTbCGQxW
v7PsOZ9n0FcUfCG6qTxwVMVeTE4RMLd+f5+ThdtLVjx2Gsy3r6rpMONB6JrIG0QHIbc7dUaBjxex
5tHjY63FHpAqJg7NiokTc1TaLW2Lc1b1pF2rRH7wTCtozxV3LRJFLxFvVDe4Tsg2OfVCevq4Kz6+
iKEQx1Dgga7l3wIen8/EDsg8plqPhzbFnJjxvKc3TOz8b5VyqNIKLDtVM0ANR6rYBbdCAUJLEjIK
sA6UygK+fpfWIiUXtAZ/XzCD5znyKXZUyiFG9C4nMWRQi9flY1JBERHOYusy8NIP82V6RCCW+wMv
yU7H33vsddyxk7h1fN9DrfrI3TnVYp3bobx9VyfnmGOPwBnrpB7/YUhq/0BvqVCfuY2eA4qyIEtf
BFpByl9JIvOINrbAYxQkhkWYrj4LN68qCb2ktV84N0H7m1P4G71MEPg6PNdnq35t9uZH4PWGHTyB
IhvDTR+X1bwBCsKUfPnjodGYXdDN6LBUId+UjYXjpLFBOYqmPIyLpXUPTuV0ipdfxc4jA2trm3o2
ErFHLy83MOBxux2jVkddtAqbKOmxAXE6aO6sOBd0C1zC2QqCc+YuSqqu7rMiIAVjU7a6GSF//Wkq
TZdIuwUOf7Cm9r+RuRgsNWCXsLtfHVSsBrWo93VjabKBkjLS+LqKgMI2b/dc00qhqC0Cx5IbV1QY
fBm6uG93HU3IK9GKaCfSNfE2COSj07DmofgAfZ6xEPZmfno0w+YrVRPAyySn2V1/mcqUbDzBsrds
bDwr/iRmaBTeGhD19exIO2vZVd8Zxk32BpZDCNoeH0uEuLcnkUEdJ6QnMC+BRh/HaNqtYGQiDFLT
bd5s4fjd9rQN/Q/HMFluWJB8730jVx2d+PapC+3EcIF1R0IuPSrgzdglMUsj5Akc9EYJVHGVyMVa
e/9kZFxIyqSNTzBIaLf6WG0cAKbYumhED/bwGHuHl5J8guxZlatYRoT5HeTFeURQmdDGmDDzvoW/
rJokPOYiE0gflu5f9jeaCEJY6OIwLys5lzNwuAgFv8BuKoTVHSGVtM1yln/HOSi7QYc5AIDjWp+d
MYyYSp5AlO3PqpbC5ClYk9kxxv3EYqzMoey745leWLTDJPYIAn/yLrJyX9xI5mGEcaXmxkMC9myW
dlX+fXqvL3mvaoY0Jh3WXOvjGySWtnZ1rZI4RIeKFiZVI5QOfVeCVXUCdV8BXOTzEZlLRZROQX2z
jHXR+hbvOjprpDo19QHP/Gj6B08h2mfCNcSBPaBBhycXg8P0A0ohcPxNjoTRQz56mUvbWyame6wC
WyR0IQ+yi0Md9/rxAYYwDwxz+iO3DNsDgV3dKE7GnSFfP9qnyRiQCqQQVgUFeM1jqTXr7cCh6tuz
sLSdV4f71w8Fj4BAc8ie1t36CJjBgIa/u5iP8wn7Kl4cg9oTmQIBqcOqpaoRbGNTPUDcCAKnxiFu
N7XqvnWCuQHzrzDDbbZwRHytFlD8PiEGsMBBMu2vtgYZpmwIL9P92RL0ALRk+XYg69Bw0EXJSMxy
jrrEMjCvi4pDSL8QXIWZJcnyVqJAT2pSrzvLPVbakFMKjea9wGmSeixeTQcsrzrJwFLlowgRPhEP
zXymQqJPRwH5mTK1lXc4KXjM8JmP/nrw0jAfDcLTOwawwhrm+8mzcgIrwcTjQesBzNE8UtKMeRNa
eXGACChZkBCi2rC4xx5p2jSYvD5UwPk89y5FgCsMJ7W6j9h4yRRje7AqAcF9ZDrAOCXTnPHA4fSy
iPgbcQl7AP35dvzuHKOMH6AZ+NJFt7i8wZ09AoehIy4EzvSF+DsZyureoARESV31kmGBOCb/IA3Q
auH3yOF26qnxX+bvEM3u3JM+dOthAXBMb05oTHiji5GVR0tMFLiI0h3zIaA8fRybXBPgYJ2Yrd2W
pNAS9HxB6ZcUI0Yr/3d06k+WTJYXHxhh4FBC6v3RHwTEcAv6OEiu76Q7naxIoEVJNfp0dtwo5+dK
mZzqyGTM534cxg/5TOiT0Zvq8SZvgFCGPfW9DYy5JskgWjoQDAZ4hI8DMNNd3dr6ohOIj0KcwHfW
kKB890oS2DFkbInbl64qQWquQoUwAxkT/n9m+qp/CslyZtQFRd1RlgmF9wVAItwbpKoEWXegTtB9
W0T346E2Vap4BFanbtgP+H44uMkPEdxyeG3jevJsBp2m0yRoZmuqatqWh4EmT977DUfZvhURtcmc
4zqBnEZsb0m/+I9WLAqhdS8O0ApfiBiWB0vYQQmAp0Kej1mCUSYAziVnPiS7auK8zdnevLagpwZZ
NEUxxVtMUEYhj1c+AxQ7T+OaE7ZBITwMjR719qHYAHAGmaEjyfE0HmVYTSb5YM+LNJc4zMFlt1HY
sb4ewHPj/f01A1DJJD42OyW1lbz41RWQPYkFsxyomMBdlgU870ZVPKJ8ufDUF8QYaQEdnGvJRa9w
Dr+9tB8JYjCiCrTdiY7OazZqkIAvWtD1nmztzFH0jdLvIXSo8/zOBInaKQSroTOMMrcqYPoA5OQt
v4blvlXw9Qx1RO0Qe82iZW8wVK/RZAhEsmkLzShobr5927CWCh0y8zrUvWvHB0vQKyEBLBabcRfi
ekKzCArYQaoY1PKoqfOnft4IScDrTf3KVuxWAhNRVcMvxMcbzojFV/aPPBH4D2o02OnY13cN3XT7
On+CswENruOI8ha3n0bH9dhI2jcrHFdsBu/G7krpTRn5gM3TIHdh1avSdTIYubc1dtaJAbKDQKzI
vb3SMullUCU2PmINpMQKPW7jlEj2cBAgIW7RSCeWto90Gaxb/SZuDVzN35zkLhqFvZ1k4q/q+sxy
WvmFECFyZtMMfz6G1RZ0ToG5ls85kJl8hL+G67Ho6YiDRh6jo6X7R44bDOFLID0WR1YR4mp0zFMB
PPvtnthmu0TqxlphFkkNMvFANCHqOo0ANjzDa9VdmxOUfIm0CLyBXx91KFlsMHRSHiTkrMlS7peB
+kl0T9SnrTDaLdfGRfEIecCpSSqPaexIadbBmZB3WRM6DZKLjJmg1zEmhvsTTeoeEwhzJw2t5F71
TM8+Xe9v95kfKtNqFOfdzOxJ8kknu9rSlpy86Ek9PTevvZ/tkfJRu8NHQSeblXuZnA2DnvtSxZwa
+HhWSSsAmwWt/15pLG/j8Emek0xVXd7CQrFrmYcj0EUmWj8Tmmr5Of9WlTFLfQtrLWB17QAZKXhQ
xBqB/t6fZ7JdbcjO/3zCjzH2D0RktdEr1wyRVQcxFUzRtyWjW5zCcrq4XeJ6vo3J3/cJ2w2vssHS
G9HOqiIBy3Lx7H3/zne4+zDFgMgS+It8HTg0YKvbr9ydozuuT6QFIaEjwLXplZpx/1NOAl+N+cBY
tsaSawwMoscJvtTwS137eKXqB47E2j0zIdVpEohq/3m1ApMO7ZhNjkhXvHUn6tMxc8kZGBLfPX11
Udh1NAoReT/IJPdCE57BfSQ/ypIWYgh1XcCnwPq+EG9lp9ZYmRzzz93+avr0O3B9o57dBTd8YJyT
17U+zETUPoZfO+v8Sf7CZt2SeXMlFjm1lDU52QAQjFXj02UWJEFvpkL2C1rucXfghM8v6bSVytV1
HcuLXmfn2sYX/+L5BOzUTOV23TmwCxvZ1kItsrJBGGOSdcp5BAhpGopkkPCTCR/FpYsWijeuoSsa
NdE9GwkZqPtpfCueIhN735v7i3ZIqhI/LgT+rq1gPZn3A0BiAu4aLXekr27QrnDFJmQL8FJ8wZHQ
gmqR6BV4S3EJ45B0CPM+MP/czrA3/ZffbEdtUxNX+VdTpWPE0Vy6Pdq+zTPDh2ayc4ABrUNkkTez
tqBWXwZ/cwjlSe95WahqStZU8U6MzcU/+6M15jra0gQzE7TJhRzWJRukiONomvhoEQrP7RiTDoka
HTGjjr9KxAuK4kEOxhEMxdsWg/lATw/lCdJVlu+PZeaSXqR4ymBIyutYpYamacmOYfvKH2XDBKhC
hNilGI93GU9XLaWHqGw1Z3UaBL8aFwS4MJaKDKxwB5NTadhw133uDsSaP4PHAOGXlQVKAgt3UCWR
pJmH3nSp8hgqkdA4ZOLtQRxyRhHwMTg0KXFyO13w9ZVNauSTbHrzG8/paIu1IC2HzoxVpC7qo/+h
7P1amgMlBvIkscUZ3pvJ+x3YhCs7ETyLXamPZue2OFzfUNHyhvn66A82AuYMLjQnB+nesPTeM/Ym
41S/3VJ0cuFRUNIc/Lok9SqeP4jYPfYlm22XqbtqC1RXTQcJghMzERF/OZ1zFuMeGblyhqfleHKl
9ZvMykZuKS3s6HYnj7FJrG371FTurLsXhYzA1eyMLiCxu60q5SkOcc6ETO3ohyoYGTTovaB+CoHR
hfUrC7UiiGLNF0lEIpmOwHDECfRPCwGANDt5e5bPTpNSvgj476xh7lRf1YPSANlN9lw33EdowMNh
zneuRXX7qhx4JLuUqn2mLbldFMTl+dAmDRLyOErBqQGvpCsWIO/lgUGjs/kTaGKPr4205Eh0X7OE
cd4Iko1qI838tROu2qq8T89U+RmwuBcTezArR8ThuJii0LgHu+WuqQYyWZguNCwiJN9yUeQVZBsL
qZlLeJgX9lPETzK6O5Gg4rHw4UYbXwxKukXgxUfmoawcxrKyWJrq6O5I0Nqk1/4pMHUy2AOz0C4h
if3LETCRDUjU/o1F066s5C63z7TUS9q96cTq27MzmDfePUOebUZS4xfMC8L+Gfyu+ZtqXwIKCpdM
OolDwPngtleQrkGnRCU95MmQWwBJzPLwUWlvAt09jvUNJRrz3HY+fDi1ZFM7Q7BtKKO67Je6vWZE
9v+3lnQiIvb0ELFYSMm1BJ5s0o5NseqwRtgIw8UYVm5fQsmS6/BVKFSFZxwp53vNs46LSXCTu3Ca
OyTLrATAP8iqe0JtxAUx33fTpbzhro/QuZcZEPOea3hhmZ8emgyZCyXWvxqtVDGghVfhJ+Mx2LTz
p/dnZbnLcYt1SRtVfKmZV0RAyd/rx+Cd7l/azZ+flpTqSMDehzpSEDpil82Mq7W9ktbNNxVllhSm
CeXEgAPJUabY0QMcmHQXtwzw5Wx8oCa7GKja3a5gSYkPuLEi4O6+xHgNpe3O53zbWoWWuGN1XmMk
bumSMsM94EXZgEPIaV7CP+r6W58g67hmgaVX1PLTzC+Tign6hQq+8kg3hBPRJPnL0z2KMXsgDwId
jcU0ABtUc2eF05G+08WVJhOXH+X3Z+7DXnvWAGqonyGQVnJYMhjnSLS9Vtck8qUd/LGNnY6Auu8t
mUUuVSDWrMOr8G+p8RNnNQDYsArqjMMQcIldQZa52bABlkEhff3Sd9RM9BIlhxPpYQCbHnlIxGPA
b/fCy3Ocwtp+/zotO8Rt+5hgGZofq8C73rGi74vYRxo1DqJVoPWc3ZGMJhlpVC6CgvxVJ+97H4Wm
f50S52RD75sUDsDHhBJ03M6vpqlqLVI+NY1jtYjCDZCkcwGr/8Td2qezChjX/Fp1kQyt/FMfppxO
v0jc6XVH64sY2jDkvR4rZbrdXrVwAA2LLj1DvvZPq2r6SuHE+5syPmxu6RCa5HoQtxwBCYVBXa/X
oVjICNGNjWaa6Btwh38kbSP+4TRSgOCChGEJO1GfVdEPLZBL6/KA+GMhW86vQnoFUfIVzAI6EpVC
ww9S0sicZNzbW0d9EoYwdfI349A0FXad/HJOudaUWpwtto+FMiuOWKFsXRA0KEjOe8dTAjWMfTJB
layTKjPypJLzfArUXOnxM0nJDj3Aa8cgSUFEt38yMUJTREnXeOwjdManGPAohzRjxNSsE2qswyqF
0gYRcYQ6mvZzKTCzGbdqDjaVzQXPOi1AI8R0GLPsUqSeot+aGilqJOPWL4+M0ynmbaNXZgB2Su34
/Z6QSM2SEucDcWZjGyo80jiqGdy0F18ZOAqnPUYc6voHJTnUnq7E1Lc19LcxnAC8+k7lqd3sg6g7
76+/2PYea90o+ZWeqVvzxdevdYLGyT9Rgjgl843nFAT8TitldQitMaUIZmXDoWambhF2yXAdLQl7
zK+rEG3bzzztoeBf3qslwJJssiKw2Kajqkj262y0v3bTVR+G6W7nRMc0IKE15N1A2THcwJHFNMyV
o3vSDZLTkUTJPdS9ZdP+ddM0kYcIjZCezCUkjDWzDMCNbnivnQPo5WlM3DlDCUZW8g0I7P5DY6vu
0GoqNOOsuJcrCXB4BcchH1/vcugZwCIHLrcOE8nLO6VqG1Lzpt26vw3iISE/pfT3aYjJUew68njV
t9o4ekZaIONua1vZ/Pz/OJtPqSWfGhXb0t3ti8L0MoMiCzMu8Zaje53+Zq/bGoWgeOp4jSJckvUR
C4byI0vM11ndPa/xRsm4jxhJrpxjBWhGe21C8zgcmenB0DDB6tRmZUtBhqnk1g/Fk7R6hZLkTZG8
Ea0CvRbS5yqbrZkXROvjF68EE3jAo6Zx62aUmOT1eEYDr9DrpDaqWoXaQp7ojbLKpq46s5jhpfDc
hbo+CiyXBe82bVOobt5XEz2hPUxg2Kb/Wa8I1SINoihn7LtXEfO9pj4MITtldnxawzeGJc9WwGXH
7eqqNawpdsxmlbNobL1XuiioHuO0bMW5hT4hVAw7hmoCpcYJeohnlJh89p4UQ6UWkwGZnXGAvJ2k
4bWxG8qSt258vAQ8XNywwLxwig2llP7NkmRdqxQ1gx7yiFy2NnKvRVn6ddonABXCpYZiHwpJ4BzD
55X3pPpU4vAp9OiptAixnthkFdciHW1v+cICSy97mLpjL0WOunELiKncpjb0E5f8VteZZ+KOyyCi
bI8F0B3lFvXo4dvJMywpwnq/TYxw8/3SMhXvmbA1PY9MXZIrP1Pjr1OEtOgkexHN8Zsbu5KzG4++
oy+4jOiY4mVmWX3KOOSPMHykGthdGju1q+ZS4Rui3E6jahDSAxsl1BhNXNzL+AKBOKkUvJCVYb05
99OJ4waZYIFhvY/OX5Dl0REaKtu8kksx7jtdan+VsQxN6iPydR9f1IwL9XOJo2D3K9dl8GbRKdxx
/h1tB5Hxi74XQ86hoxhyWttGjZdK3jMv2briKbS91x+aFOT0yiWQ1ZVd37/C4pKikBziRinho3jC
xzEv5UCscDFYKDglcSBHz9HAw1ptRdQN18CQ9Z8Q8DSztvfP/SU5RCbarym7w0R2VGbIxPLUioCZ
MZr20GYtWFb06siAN6S0UUuk2Oi7tfCQpZt6kY4IXtDnmvofdH4wvu5e2RtMRQnsN6FzcmQmnHLK
AMCOnxyAWiicRcHgWzGhekhWc+Bqnrgg+SL/81n+gIUreC1Q8YDrH1+sOajfPoFnoYrYoCJERDCr
MPFDFC5rfSZPvDkvB+uAn8gdp2P9v+McrypNiXVsf7ypAmw63HgetHeAMvfii0AHyuYDJ2b81aaE
GdsQ7aC4VpUIuZBNJcTjfAdH1zP1JuQpLVjC1vygfu4fOysRe1fuG+Xw7+S3W63N/+DjAx4FhHRF
Y2BNSO7wXOYHKQzPOZwfPDl2WAnakrL8l47qlP3gpB32/pdnXKxM/QfkUZT5/2ZGbCeDSmKXjgrm
1WhAX0OJj8U+hYCF6v+1bS6MQPoOTHQ9o8ED1TNc02htAzMjGWSfdftcCABNOxyrlSz0vUb8aoqV
WiOOhmzx89p/6O8T6D3FUB6uW7VA+hMm/ghAf7scJZJTgpHYaepkeBYC0uxK2xH7JZ8K7eZuZCD4
MCX7IxWMYDPTY+1VX/0ULj8lcaAk1862RzsrdiaRJHaoXjORHYqQ+1X8EwGsxFNWryhKxWau7QXC
B8X1dvPF9C33XQIIZwRRwLJmPIlN7vqc7hF3AwVy85OE/EDyKtpF89aCzxIb+5fEEBdaiD5V00r/
NLZiR4eKuVRUCVaASGIj8l7OquecL9eCTaULzrF+OevlJfPAstmgMYDP4S5Fd/I/fM2jYupfdKBv
hETEGxYZfvX1YQxC8HJeITr0D+Gahzp48z1p+1MON98ZVFwCYP1C/uVtQTrzACqzfOwdBptsgQhZ
NECTZ1dcI8+izoGr697WCwDvesY2ujOfG+Wz1822RQoZOMQlQkbYvrKeLPtctPyOlvBHeUUhw5kR
jSvN4s1kigboDxPN7M2syZfgq+b6eD21pGiabf5EcVy4oEpxss9gCokDs22dgkXFmlwukwoQK81G
ZdA1FVgUXluZIQlnwUBnbwjSnsBIvOgDYu5hO8oGHRz/ttY//+pYPYLpcFH/v2bv+Ajz8dFhCyiz
QmYeAQeNfswAwevmx/kZxfJBhFpAdrkRVF14yZvqpBrKyp653U9fRZ2yxmnRK+LJCh6KGSsIcBPq
SNP3s6yWzplDTqY3mZ1AzHbRPW8spqhLqS7r6MaFINN22ixaIKGGgL/6mTySPP+gUu1xVYqHc6bC
5bB7HGHbYkjNaPg5gOSLVJTmcGSADwg9Tvan23eF+w5MBNzTCYQxy76mQegR+Xbp94BCPNzPi42U
vD8pCPOO/P+bt7UI2r20A5as00svPa18qQEpikD88Qs2xLScrhpZS9RbLelypqGq2/+XZhz5yjOp
z+64rBXiQEnJF8Hp2ePwIeLEZHIGm6x+jwxvTs9OTHumlmTcO/vrrGERVwp4ZTV4zAALPCFf3RHJ
ekfnAloazAR7GNj0Hi/I1YxhRmFZkJqNSdPpDO1gNSs0DrI5Uag+zhsLoQWj47aLtScsqfTlMdfM
LapU1vcWsQWlSGNbp7oxTtDNpumrpwlr/aJ5IoSu7w2Kh0tXTwvg3GEbbauMKDagpA3MRnZvnxKx
uQi9EWmfNZxcSLak5WgAhkkJCLCPobpQYBSB01Drs2PztbMC6EYRIzTQeTXXAxLWTKSRWHwAlmta
jcXXaUwwqEby9HTGMMhMQtsLULYOIdOKg0UBU8o4KC0hOu5StHUg8QDUR+ZgrjDyQ3jjHKNDPTS7
osbrOnmMjUFSu6yVIj/oGufJfSAtakcSc4TN0CMt8fZ/49sjs8687G3gU0OrxrxTPc9YN7EnBgiK
hqSQYdbZ2zGqldjbLfm7O88Upvo1uDj7b71fJ5vGdhBjQeEqX10Vz75VWJ5Lkk8OYr894iidPqVb
w+bG5oXGYdipi6BjyDQdwHnYe2FLYzF31Wx6vbRkZsgnIyWoT0ZTfF9mNlmBRnOK9orj/QFA5tnj
vpdyJLvxvn6l3qV/oyIiVfL7OFo7+bYRT5D5tZvZGTYIoMCpOiHJO1sn0J8drYqzv5BbIVfSBbU0
Jj2iGhfZcBUjL27bDxryGGXwCxlAuVFi4Btz0TM44M88FCNySvpJr9CD558JdPY7XTav0DP3GzaB
/iHw3RKlBCvlozA8a20jnjysuW3jL70IJBIxADmT1wAQbioVgTBk1NO8YZYEmaOGjGbcClD+yBFh
h3HzJ/dvnl8oAM/09xjEvZuYBp7rfpZFKdrAAqTsqml9c842tGw0KRvV3vRN1Xuj+9Pls6+sNsiO
eskzaaRQhQxo2SOx6qWR1L7voQHnApx8uZpMWYtZOsV/y/hQN7geJzpX4D03oCz2TK1UL7gPBz1l
pEq/3tiZeXUv17ZvHzAdD/UfSxFhwtl5jhQYbFu2+p2aUlgPVG8vOluuLtil79X4D2lo9fBeK9Ny
1epPfJzdcreV6aYFdsgNCKBZ99b21gg9vMX2O1CtmBiDDPBKOtFewgR8/CEHeXWJU7qiVuoKnuIG
twLRuJrl/SIW+9johff4u09e33aZ0NvaQZUO5VU5aTHLbNlzAfHEtDNmQEXV69raUuH7LpWuTUww
lbzXh+Py2N75KtlfviykwqXNwQDzS3ht8+JR2kH37iZ9xReH0c9NpcjyK5AZYSARpnz4AhBK1byv
fJiuW4+fGfYGDM44l7jKE4KyOtOTJP/zNCSywHvFgn9HyUdWVrNxBHpiCDnqV1ImjAm8pvrA+Sws
mxNn4cR55ivgSfKZ4+k5guGg+G8L1AWV/vrpABo9t9fEpKB7DwwRMuCgSA/oxHO2LaJLjvyoCiXN
LoSbotur90eRMMLMik0gutZyDe+CKtxPiROr4lr2qtih+CttP6Ud1vgMAzTXrPPiUNSZQRYRMw0C
9MKRBxNlWw7F6OtOiyC2ZUAOfXWbouklOca8hESmPEcQ0B+Czut4F9ybfWgBQAju7ckJgJrymjLD
Suby2S3bOG1nKWsj7r3Y1x/tqe9JCB2I8TAuPoPT6aea0PdnOqpiH3jl6vnfbNCb3Cr0c/DFPLif
A4GutEJ+hXFaj2vECa4bOfrK10139OO5pKvxmKTLurifKWLjxwITVXIhspe66fHcLkMZQWfk3Hjw
0FnUhD9y86mLzlWAZa3of364mA5fxeM5kMTNP9ogZpyyk6GjUHepJFshzrNLcdeuFr7CXqioOE8U
w3noGLzUUXNrchETGSHNKnHZsxY4nBg92+D9Pb6Z79FfHtArfA5A5uMzwhunCjrXuTRQC22FDt+x
1fbGuOQKyYulj6SdE8EqgcSk/gPL4vFc35RMZeYmiKSsGAHZCbORAEDoGKoe3FAPGnxDfcU8xRLn
vSeRXdYjNrMM4yt+myNhs+onsWlNngUmoJ1XRJsPkrkNuhwZLyxNy6yivNfU6FbIgO4zuUMk/zSE
xDzGYvfsqRJQK581YnhlvGWN5Gi1ohWUnNFQ8OhInwesRQtiyRHSeEEub1EJ/g0T1awbUTmK1rPD
bhL2XAbkn+YUsJV0MDjqtGMbSeMJwW3EisIhGDWICQQ1sux65vrNP9YGmJ+xmPNpEwzhQXXM0XiO
Vs/Mk5WPdK+3hYaeugkRBVIMalfa8gIprLvFYKPOHY73TzT3alPTZD10QFso+tH3h3PCBjHv/Q9z
rb1E354SRypZE+kDvzxXstDZ9hZM9pijl5XwBxeSgpYhoKlMrectVQYWR7iJhMjBTB0EfqxBbbX1
5U2xvGbqth57ZJ5ncPZ8A4xPQsf9za8XBOVS/YFOILow1tsKIX9nHCfmAqvUjEb6oXXGwhHUsBFC
COYJHXFxDax/WHVC/S1CKqc+gicecFWz4NYpwIFrrvj12NuD06/iVIjBABAPpxPtUUr6EPJeTJTl
a7XLCyyFz/U0zaOKINpxUbr4qeUPapsHmeNnWmmqcSWQ9+S24ApeEvXauWomhVydSdW/+owLwlp3
GsCIkW5GzTgNGmGr7+tuMhHytZCz/vKtNBSJ+Q4YRP1izgtp3G+rFIJa8x2Y/Wf+5lw+3DpJV95y
1W3pjZbCvLJRwrQtjcerGJazrfd9n9FGvB3oONO0synBvoA7F9bNrPE9Syqi8Ynjnz3yWiV/hFYA
ho6FqpaL+wCJNf8lVLmVIWoWDejKkcPOAunAWQ4eX2YDr9Aq+5wOtMWNGg/UzqGyTjhMTQIkHKAX
kEa2jaZTadWhr5q4S3i4dA/JkLZm6jk1vucl6tbFdfdckXFGR64h/vlDzMY59HaqBEZoyFhUDbK1
uFJpM+JpjwpGewAfeLdKFGwjJ15G9vl5BgSOjDNoMBngBDNnoQZ/mdxgiX7PPaaIz+xZRw+zqXa+
sZ9Dxp3zFXt7FEBAblJ48gUKqjKbC/RpVyWQHlsOgJmzh1EV2+c/IVKxB+WT7JeGnJ35WlG7VG5O
GF5B2saLvjXo91zWEv4kiT5VfvT+cPavaYp4Yy2d2N5YJbkQd9lUN7u2r0CBpohE/OnOIYDkpZo3
mCHn+6P0gY0t5pEN1ddrO8/4zWjg5F8sh2HREsOYQQVDA2qBSYCtbt+wJvT0omZKUiyTIV9Sibcw
48fmJ01IHyZY5g1mnbyS0+4MF5rrRnkKZCjh9D4/o9qrAkXLSEb0Fo00sVpXvEXnIdCLDLE9PBoO
tGBw/+8a2k476ZNjkpFFz8w8EAT9mjmASBbojTZNrSmXMjq/B8+uYV5MD5bcPMiKRaY11my0FNfV
APv44ZS2+gn5qcBpqOaPL9Opm7e9bM+XLXkg4yzw4Q7980k2I2aDK+MTfUGbCqAzn6zvr+kNgh0I
fn+T9lgpiZn/K6QP0FKb/5vRt/mkqbntj/2Mlq57/sBTZqR509ykfrCBEmBqMNSlzBXdiBLDPb2S
/q/5J1uiBH2hbk/FXsC0bKD0Hf2PEIA3U06diJzP51/kvx/8KBqa1GaCp+TwM9QvWHWVDZS+X9s6
ARu982WKO+c0gPZJ/ObrwQzi4wXHchYsEAsOmn64s/rSCdY/livnLWg9JgJ2CjZJJ9TCDrS9PWm6
NFMizDvwRBJh3fQD/B7Ifn21lOgYEDl6Rz6mQiE9RnJVqk4mLoJdFHgjVgDIjtW5zVVZJqOkbXqd
a+lkeoLLv9nDD6nCh/dijqGbDK3QftI5LTjPnmjItlP5tBMrMgJ15k6sRkhgz2gY67qtUicrMY+1
SZnfimgAFXbNyUlJk8TgnEK0pOTOlQP6BEvNvllPe/nbHbnAEjk+BH6sj9coetbNuNd/8ZXyoCD6
pEHR/XzliquldItadLnPtvrtW+nmsX+nXcuq8yb8YjxohU/AoCATGSFzf04nWzzX+fUhPsgyqbcg
ZN0TPb9xGna6dRdzlIP/QQ4fME6Z2n6uRzhrA1UQ6575zGdey1E1MnwMAcvbulZ6qltLasWbJ6B/
MVlwMv6dkF2ozF/3+ywhQw3Cw3GGBqJz+7OCNGoiK1BP8M37Bh5LQB6ZoCcPnZs0YxHeIky942KM
WyqQqcOfzxCBRqL4p2c2ZGT3MFWRYjGvY0fRua+7gT8sqYDNdfLEEaAJBZM7/fYcBHQfCPilnULR
IaHUQkYrBJX1mR7N1wYRgnIDwfXmPaLbSRfFkFfe6HC9iSIVge/BvneK96btn706UdQXaRBw6I6O
THjNFKxpWpGgXViUGihKmGB2OrhZYCHv9L4VZAjCM8D93dF8kZ86m5H0CkyeOJAhtmbPHbz62SIX
YeQqZ0MzS6bbeQyjdPm5Yad3DtpVVudQQdXtzuBnHpUW35Il8l4ipPmhQ627Nuf6qwpHvDZdXmWY
BspIqepx3D7LFfskDD1psT7DUC+aI0eXeF50XPQu4CPVUxsE2QI+P64gwKctCkrxk9N8wkJKWkr/
Y4IMCA6xVvmx38FI08Dae9GeuhUFMgyqjqwK8liYZc/cPllhnzXRmbH8e/LF2mVhsG7CcyP6FILd
DvhvK7PkQbGKdg7XggC6wVF8qHu3fXWOjsArkxnJC7u/kPXPfU2/R60U1icDs2zCmrf+YPhIlpvz
Imdpokm+Z9cBNcyZULWs3Vqq25bOpWtq7it0FrabnMBbXIcf+WHCJ2TozbvojXW/PN0LewAFx3We
uDz0Ul2tT3XSVLGwzBTFF37P/mbJ1tkUVR1LjK348Oron12viJntIDw7PkH21vO3tSIAurt26zrd
7j1gsX0z4pTm801lDD2nkuvwRuaT/K0Yd+Kzua0JA0nQzorQZZ90dKI349ca1TulqrO9/csVDy9X
aptE+93xA7JgQPiAwnB7GbFWKGoLu6tgSJA4EU+4cTv+n+uRZ4zYPQ4qtfPUacfXWFy9avNlFD57
oSRJx7wjss3Bio+HxbNxM18FsyP9TImtSiVPHvGSQycSZlssL+I/22DW7ooWmOHdcbwmqrye07Dq
DKZsKlZ8aMQyJLzZW5rFc5xUHYz+7uK79YQzae/qE/Vmy5dgN36RsiQhvVpSLsVB3l5/cU8IXBC3
anBPUvBI+hvo9LQZVS7hzusIyYtlSa+LfdVk1UTGF+l9EKjz/ZYga8X+9MaNhnhiJ2SfxIV5hb75
GZw5fsQIetrSpRgga6F/SKvI1H1S4MVouYEilDPNkQLZnxGboxKQ5oFcAaVRR8FOGHYh0eCrPE4G
AVgAAEaqnjERgEOTBAloexyDyvHMdFBb73y3iF6WpqYog2VNONyKaHEW2vejBsYZ359y8o1eWabT
31zFhRXuNkN9YOTBVtEjPGgdWhGmGzNlEvap0Y3zuPhZK2z6rupsynOoYyZhUcYlseRvfmLOnPUe
6jzywU2CGLqUGZSHw7MhFBCP/aqU23fXBaXZKyjJNqb0iz99CwydzVAPb2D8VAkaVtOB5629v1th
pkRH5+OzmKsIiQb1UeEdxFCQZRtjrkN6bl1RMxnqnro5xXgxik40xia1MxX5IIXomtZ6SEbcCOuO
j/hzHPEZwj919Vq8ZjG2otLpCwbIUcA1XjS9mBYC8ORFKKigXd75U2eMS0uvtEHryVuZEcdrxrSz
sQgqeFHi+aW+RxLIvDW6wyYUMuFUzJ7jSzNMviTeUc+3sq2d9oV6bTlUreFdQiXaNomU44CyTBP6
lBFELKPduvg6leWLEYUr5SWE4MFjH4z5+bO3n0FmIfC8fuz0hPyqLPf9IBFs49tLP58OXInUpsET
NaE3zdQRX2BVFPMfsgWCJv35V4IbWnK6NWskbAXM118p3xt6YVtGhoj0Y5OHWxocVbXzGWNcrlTJ
JeN7p02n9q+UNjUA6Rr8kh5+aSkr3A7ehTWkfr3lwd5Jfs6dxxskaG5GZgsaaS8sVmI5hS7YWlAR
dEiSAxjPM4sYRuG+XATX1a3PTbMQ69pqWq8H2Q2X1ZKZTEX1HuXF6l7NLw61W90yn8lJWCWt9x+o
romcMayLVIzvGLcqMpXcMKHasH2xHuhx8Qxo1DUhIzcb0L+adNuznJCtuuIdIwyTJN+0LfnQz6Q+
4klkBNGwci9ljI8swzu62tF/zQlyM/9lKTHndRQ+04C4gltJkIYfORhfZ4HaTM05e/wrP0sGjAa3
fiqt1nOXHqdFWfbfmz64pkmgVnih/PEW7lBHRg2oDhro7g6PDDUyBQplnSiF5m56Vh4NWuvwZIwR
QZeLdaRHvE+yWA2vYBIT3go6dU108lDtsYGn+pdiAh7bLYrGVC0XmPhLy+AoY6b/LvzybD/w+Ucf
HlOjRHV0+GtPIyushDcif9SDlBU/oXKf9PqUlkjMe39NcggQ44Oa/GVdYA/IVtRjVuVy81yUv0i6
xujhqrfDS2OKqyY+Z/r1CjuZCaqvIxFGcE6VU8hSdf9YtBQtdfd1WNG58CueGa8YNpmjSIpgJJ4K
aRGvQM1BBJYaN7ZU0OAChm1+TeFfBhaKqRt7VjmpRnosdOn9uTb0cJcvmsiN3TqpdiAODKkhn8SI
32fI8CWgTZlSTCeRNV59aYBImRXB37oH/YKA3lPdSz2IP7FKXs5njfv4+QoVPqR1vKA7TQR1qud8
nYHVqb6204psKnjJLP/NN6YUsuNhLN1PhoAA/VCLMal6rC80N47Ebj7OXrNUHmFzmIeD2RM1Dyys
e807nQO4EZEbKy08r9KvbP+/4ebAHmL730nh5IHEBnNl5XPOm6R7BGtbttL86ZjheuBHnobc75N5
Gr5QuVH7MoY0vXvj8kRP3xKHvQ3eAGrDz9nzs5LYLfAombw6/EmVnIiBG8MaqxtJoDYff7qpgYXj
i6JgAhVi9hHlT8sbHAV8l84MYs10rn6fr/jxPbqH2XOSSmm0K0H4bS60y+1kv6SjuizQa9gBNaMJ
9d4zBS8Zj5QXM5JNoT7z/n+9deM1veGLFzZKviyuunoUUWNt+yxrfT+Q840bMioqHRnrmzzicDfY
1FRo41diUQWMl60jAvPMDQn+ZCU9kYQkzvdnhRG923iCPuys0FaB8HcSpiwHb+CaHdlpG8Mg5ljy
XUOkr8tkd3pPugyB/QyhexSxc6VPLpc1M9ycVvyZ1zPtvr5AdqaKm0MAEKKhC2VE/iMYJDfCzosZ
XAVvYdITkX1GsuP9lTj3O8ZDnAvpaXtm2WeZ/LlbhPhuf1ZNzGcfc1/46mJvo1b2s6PHpTlvSnJB
otpSPezuk4YYdnQAL+BJD++MJIzxrJtiyNPh1FJO2ftI5ELmK0zFplgRv7osZ/sAUj3IIWEzmrgs
8BITGvOj6jRpTUUKVKSO6PyC1MbXphyfRyOV1j9iSdorfDYGIM+TW2XnVDJ2xtIzdfwmV43rZ5X/
xegysZPusZNiaMkDj+8l1HII8TT1if0O4ziO33x2sjo/jY/XW2Xfw0X1xneeJgTQQHa4iOurSQIp
0MBwNbryUP/+t6xEhVZilclHyhZkE/8pOjeWxu8KteCGPnQaanXFfs0dVR7g6KVt8ioebaujImWG
WrrhQlanYgHOgZnyap5nHo+jbNekUWmLhLgBoyEwXtzhxN/MgM+PNjTIBAxhjT9fe+IVd4svKAPR
Gur0ASywScOjZVtIc9ESzQoRtNiqFucU3vfhHjbLlMYEg2wgZH2FkpfqCvN/KXLAWMOy1nIzGUkX
/TEozPaYpVX0LoO+jOhODqscT7JBEuMIMnnwxSMvOU3atgiG0Gpj1+1RCv0bwAlWqhkuhkA1GUe0
6gks5yDCpPwx7fsIXwq+FbgV24ni+QQnVweO0nIVrQzNVyYcPjxgTrDv4G4kl1LEXsHLJ60Y2IIV
tXtMzB4sVeYgQoLSkbPriNc18xQqdZh3ZnrakPnu9LedltBPp3icPVGA8nE3r7G9ePIg1/sHKTFQ
xPouasy4IIyLWndBUp1VyHqvdG132YZ0MnagvxVH1BKl513XTeJOs41HSLTFUp9dgW/Ez7xSbn1y
zSZ/UXQlBgkACjakXSaL4hv+spm0ZJiUjF2wZlORUDPR2Hngq9WjOijbizT0ACO3IFb935eFl/x5
VCpERn+6FC+oPsW2M1WvYQUD1fCeOWieRkvpf7GBQs02YaXo8RsxoXN1nx7itUut+0PR8LwyhccP
0+fbFwTtddSBBad8pw2LNEVRZWwYvLFGCX1yJDouvznps3jHovtsD73S/01eD46Q8qI0xn/kc+5u
LBAqc5FeZkjlOK5jt4bHLzQE3vDAqCXJ8G1h+kWRvq4c9pSaXWH8YuAgJtIknDYyKLKycVvUeUvp
HYhsnXFyKrpXjWIQAVsGn5FvffFJxmax2J0IY4wQOF+NH3rBp2Lg//GL9EvTwI7daaRMXGRdp7E+
xo7uFk/Nc48vBedll56MAm6Bb3S2dPkj8bfeucgTLLsnn1wR5gQYWDv7veTXd2FK1F2p4hp29hZp
rOGdfJlIik1sbj4WD5eyKMs7u0U3EWGennjsW3u+U1VsjQdQVTdZRVR7xNtv73a/DZVi+GDbPuqz
BPJC0XcVYg7qK/gzxJ6+rY6MRTQGtJ1+6yqBpi79uvSkQY8l0dLCdmRuY8uXZtleWFAj//yWvHnM
RcAzqbyBs2f3uCKagg5OwpAp/1xf01T2PgAMv8YoHwRQEnm3YvCdSvT0GP+0wTJm+9Nc0GGc/XFU
rpxGMnNaG9lKb1QqxgayOIqbpFsZHtmhjiPur7zSriEHs0MkYBWDD9C00dmnR6RPiA+l56vRrXZb
lOrwZjkB1jFCwdXWVhjC4/t7H0Jogs90z9iHE94BlxzW+lL4ApL7ZXPwhlYvDcFOz2t0LEUSYt+z
37S/IfgiOVSKRgjYZjbUGky/dgoTvySqVkr1xqKkVM8dZhTeW4u8uBLDJ4lXAi9BekvZcmO5NQ1R
0CK85UVn/n+iYqUHQBitv2khRbpTi5ygZ8iLXgc4qAQzdmYMsKEJQI21PVASxRteAvt0UnhKWZuk
x+GOSCS4L/eLVrJd855QrA9rgh1CKnOzOLXUuQniGM8YQrJeCqICr4kA2DPk3h2XRaBZsylIYIUN
ktOKtQAfh4i4QRM/yqUNWtzuHMz/JF3MFnYr1N2owTMY1JrKL6ZvGA2gx5H7QHNryzBdb3KAAT4n
+WkwlKFVB1xznUfzKtEEg4nF86vY9li3WJMOXp9cnAhcdoBlynb1q7jzand9hE5ISGT5Wa2YysyK
TpUMsrkaGjBVQHP09iSwMwAbBlGQouid5Y8vw02mmO3EYPb8ShxVm+txNzDPfMH+AIv+CmWIX4GG
SC0xTv0dwNrM6YFY3kDyfLAMpcAwqxEbs3UVix0D9Cx/HicIcaG+OrSiw+j6p76uMc2ywGKx/i9y
jf2zlyH9ZVj9T9hyuEp1ZrR4fJF9IhBGMGDtNtVV7wOTuEUaTjePw3xgyMBW4Ens9MnxpgRxDzAX
RAC9P5n51b019fkqRZaZxZwqmH1cLg4J3GG8I+LqykBSb6ABlTmnvdYipfxadREslYeuur2KQaJE
ZnfiBn70NZtnGjxmE5f7WRC08nl5pBl2VXewRA5CvdrQVtAKEfy3BZ2zRzk9dgaVCByloBykyphK
BnAfl/b0kvAc3twdZidcDGQDfuvMnyzvKXoEc4uj5p474IfEAZkls5F3D0gW3E1MpTbhzBmHX3D1
glyB6gmDQ88hRg4xmDkDZ9iasOtLYqo9HCk19pBmRRQ8EF4enYsw5039Uf9jI7AnlWUYYIetFiAs
2ua+7eyiQCl0gCwBE5scEkneFUSnWWfVS1EzCMbKyKGJHcthFaMD8Ac1vysQkH44KrmLTGy/WQhv
iwclZB2zTM86f59dlLnKqNPpGF8HKPfstf3rR32H7tBjmdXSgEFhv9fzVw0rNBSheEPho3MW2+dT
JkKwt73w7hIG0Kgc/uu4NYnN+wtyCzL2oK/ti2VyakqUPiWY7JiLwGVC0IzFaxlmfL/eZHo1NjSz
adAss6xQgWOGlGpP1FyDvXJDDGUW42sXdrrP/zOolnP4G7FQ9uVTxhNtwsJhFz4g2KDnywetV0/H
GF6yIKl8Zpn3c44FxFcpokhzN7dwisWIWT35M3gkaMzJr4CxnKDVNrj6+94P2NjM14TDllyX+3z2
oIvqEPuRofgtcxNS/izOt1ReAp5i3SX6ofylzHGWoXB2+bsjbBvjSTnr/vUg4qD/4ScWxoGvDAej
QUmqef4oqp0bJwO9O44MKz7iuXuR6Y4RakFaL6TQexl9/20PTEIp0n7AzOVIDvH9B3Y5R+4KIoso
2VKms0Pm7zYzvtIilZ9DRBXdCltyrtCd8kccXpt2m4ZHDgwoNz5PgVM8DwqQ1PPm9BkVpH5Qvviu
hJPLGlPIqMAhmTx3kJ52gNjW7LiE3ZTMTKvojKlfbRVeNF+RwGubzxYXeJ+081TzEp8Dbg66r+50
pUcpC5NnFuT2+qyTlUEMr4g1pN/LjOmIixP7U6zXWQV2hJsZPL+pot1WdRtYFTKpq7NolwwPuTiT
DI0i5dt6w/xhhePzpJg5UwSv4ggD8lYfMPJl4o91pJ05rl7gc+QGovZ41BrayycZdYDkFU9UlpI2
bdKrlcTS/bemQCJIFknBh5ysXsr/BtIEssFEzuco/6FH/mexAR28xjuocJpVQi3ewlTXjC6nWVxq
tEpLe5ckgHTDxmNtyqTVjFI1+aRMHjrUgTb2SWwNYdDutQ8Cs5CEdw5bOnr2bgX+BM/qJNCCEb47
yHty5DcFmZ8Q6/XNnqdKB26wii/fyVlzaxKW8EyhbIqlTVwsI/gvahUkkJudabxCtp3xYmBTiG6r
2Kwkn14AQ08QBy6SjQon97d9+wkLpAQ39Rr5YUZhd5H0FCrkVyhpxbQvh5d6qp18jpArbYdEk0Ck
Q9PgKSoOnKanK0v3Ba302aUYM8YyPc3EKRhp9cxFgZlETg0+M3e1kTmKGn+uWKbW46lGIr6BPTMx
WhHN9VzQeWdOIuimqYkEVSFoNahCe37LbMyUYsMXlvnCT5+rlE7YJdnoIeDeh+vs68/HvXCaIhBD
VhR32lpIcSGmdrAaactnAjBOGYwb4/tEx9cnT9ZPdyJcGLrXR4qqv+/JMGUC17bPxno+XRm7Ag8+
IM6Pjh5QXUfg3w08zTogJTTJzQuBPe+P4HlzT97HZ0YJMe443m7N2RRBOqFegqSOOQoL+bFjZSyy
yANqTT7d8Y5e3CwaDUGB1oDS9q4rRvu5w+mzUPQ70tnj7/1KD6G9M6/82++r+EdU1V+3gIlR9/0e
eTUubUEjBrh3GwfsL8QwMAXYb6zap1taZ647ie5BYlzeDp3Y7RXsQaUwBfDrV1tQGGF4KNTg5O8J
ERm7gc+FpyzEPwBVvvEKTGqo4r1DopZPiSvtNAhVvAKplLaKYABlqcLpppFVGsGg5RWI+jIT96HM
dRyqzzBx6iJluNMemTtMDSvScgfnvLvhyd+ozN9DX1qvy8Kw4xkP0+uQmU/3hakDoFPkJvka6xUh
CyCb+S4f3ULM2vPd7g5pD5S8hZfFGWnMjwVTPipJ4lvztfhFDdrXq2mfKFgDWzD0Vqhs74pyJeE9
kaGxFde1w0l15+lT+lEQDRYDrq6Jza2b/LATeM58P1/IOdQCb0+rS1EO6mN47dZhIXmbmoyIXsem
MEMlwqwQJuPBmj1YfedRrgYPzGwYt/SElfIqW8GUtTDXWHRpgLZbAPVFD1vyYOYNsvWOkiC8va2M
/GTpSV7Jmj3q633zC/ggxv3CgUSaBI+RUTMv/mioCEV93xxt+YGtqExbqPfuM7j6DZrw4u69MFYc
BpSQhge9hqp0PzeLYk2BBisuq47Mv8ZozRa+Q85MFvfBQ2DgQK/NbyBH9OP/DLkw5nGB0QR7v67i
ACLMJwBiwDDiSUr//rgEtn4hFrjG1Wzac3Goi1Z7b/pMBuuXLzoOU+PqpL8USwPZ0xbZwKzVxfXD
nuEe1t3EC7HSwehfZ7dKme2D+vcVP4s9H3hTdQI43Clw13xsDlRZIO3433fuCcAzvsAAzYjH2IDr
heSu0lXRUkf43PidOLGcVVilTYjnMLDAgqn39G/9d0Bmr9hQ11CiBjDysv/5pD2cfzhnosWK7M2e
k3syKHbl7IpaW9d/ocApf7Wliw4PQZdiDhBmGLNVQ4P7+1vt20rgtA2LddfqDoWWkrmhanxlzYGu
S6T7T4xS/eqRIqH4ldSNhEa/O+L8MazlsFwITB3RCydgcscbvTSIvCI23OA7ZfW/FBr9DO8Qi6wq
Kshdw7pWHXx0CyuIEXtHCn3ONqaOrMO9UUSRI3ksjYtXvyTnVhyJw/QCVf/2sMOF3Ql97EwAwqjM
nXW33w+DPXjfXAPtRMP0lW7doscVDQVBtCLGk80cX6SoKOiU/tS/sE3ERFDQ8lCu+Yk2/0iP0QtU
NdJpauhv3aujE2XxAXMIGtflJ/5DrkspjPU/hudCYHogteyeFdKEITURXow4VvOGROUtqBpn2Zdf
5iaPlz87BL/gElkcCD4/oV0+YpeFTgJt7eZ98NEib1ArbQygFcA7Ofu47bYWOTLzcyd7N2yJgwVR
KzlQmXhmGK74w3N/d2UcFdp9jwNUqrkte3q0+r62YCv/ecR2iksFdoAugRVw0RUXr3amcRQIT00H
Z/zBR0NwO6Z2xOkE4ONFPQNA3tfwZvYc9pHR7IUOOedFdHRrWO80N5Hl0kerw7OM/LRWkaVSaOB+
ib+LJV3W1C2oKip1KpQgMUhCMwSaLb1BSx/HxXFKOPJa6if3LEOAMz1UJ0RCtjTUM6LpmfVFeCZd
KIMvAfUj/Ot2Dd2F8rpOkE5IKOpPYxCLa/Eqqd3mTwUmCKQ9DvbsLVHv4H/H63qGRaDMnftxOyF5
ghDRScecVZW5BEGNUG/+/Wqe4bZMPCebgrEaIa39kUrxgq5+V0xqzxmoh0A3hZCtr5VXO1h0xU0t
MOEyzvuuntRJYU5OXih8x2vGRoM9+GNOwO0BfHveutSmCNM8+N8c4Y/ys3b64lrSNsB/3/XFGvXt
rYlCQTGMFuHYNdzLC6H0Ric2nr1lntwchb5SpePpcGAPIRYtqkFAza3OL8rIl/M4s3FjAsE3OEIg
4NAlcF17+iqcn4jVJuJx22Ttilopqpt/25owKdobmasomLz5ANaF3UV09fyyFgyGU6giRF7iFCAg
nlNTxOW7ScE0wSDwI5E1SwtkgQuymu/wPdvzW/O3lruidCwEfevr3g8f4r4/KtitX76k4p8lU8yK
FzH5jEECOnVJSose/alVuWATgBYCJReu+VffkNE8qhziCwlEXx5u5052/tsDNqRTQD09kJaO7PeI
FgMCugti29zY9f1kC36oj3LszLHo9tFT0zCLBOqrL6GD/tR7ZU73123AZySOIJ8ljrWlXy9InSFh
QxeeO50aFTSM6TQJqDCX7uhvPPJcVNDlh7yUSh/7ALazXzF7gH7Ez1SiIWzKYfm7p4q2WdK0UjP1
BCrnnowRwxgWbc0DHN9C9gE3s+IGST8eWKDPumSGj/OlOInK01LTmuLKaO13ePbHL49VA5/WMlAv
NNvDyUouUsfFqYjDqpT2NbK6SyioL1XAMep421W8Jzfi2tsKaygK+yChRFcq6RrJgeXqVbeu9N/O
AmKGEfU9L2rUCsrhBQtIjjd3GaysxuC8T08w8doCRcOmh0QnqYlkx3cwUaorrS3oZXbQpiQKQMe3
rAVuccQ6+vfjuPp1G3Pr6cUja5l5BJejrl8mnY772zv18nMztTdyeJhNdfnbFi8AYALnhvXDseNb
CuEbzG0Yc3I9JaaeI1J3eSUgv9CDbBd9xfpjQcpM1hfhjUgtGO82REaJyre8Fxodmcx6INZNNs34
sw5JgW3mjfr/9PXiuiE7aEPoqDdVaXBVOKTl0g/d7geCqlPh2llOjHw+hU1KBVhGViO2gCNl4lAF
/l9avm8jCrJg2boILM8YbnUHU3s/OjGB7c7QZRYDby+b1lYw7HQ/KAylBRrLuU+3Z+AOYRaXURgL
yYCZDIGgCfYzELpIVrIudnoRAmBNb3zuaDc4r6E1h1i1mSAebVLFqrfpao8hYADdmx1WVucGbmJh
WvpD3qzkMpxoppthD7AbnzQy22VyrLrpKPTBllNUCUZlXwQphA/tFOZq0hpMi6qwj5OjHGnVw5Rn
O9TN1QI9yBvU9o4kOj81FZPRtB+WbogVhpDJjoGIc0QLWHNm78G2cw5yOgAXoblpYzWnqT1aYb9O
e1z/wnr8i70PpWmV2+F1oMcIZFWoMOuHJZRFILFItox163qbVkOGLKB/QfrvsV3T3979nJJicKiG
TodXxFRixZf6VK+f4eEEpvUoQp7Epuse+2kc5QZ/zqdYr5T7mMmhB/JDMXoGxYt90r3w62Va8Y1L
fVNiKitpLmX/jVsKHKQcx2t436zp8oEr68ev54kOHRFmRYBE5tCh2+grtOY8tuh1L/f1W2c0ad3x
6jeNKn3dh51jLkeF0JwJtX7dQJBEYetMj4RAXtphZm+0QA5Xfnrcy3L+G+3tMiVsNbgNkYDOKMhl
c7l9o0/KbL4ZglUSXP/cJ5r9CG+RHvwEommghMzgvE8XtWWcmfWVyZZqva7nNt6BWl9IalBaThmp
RuBtygzgU0kpbOdGvNxLPPYiG5DUToVCnVzKHry3QYbFfNbPngTKD35oQTSXYzTNTkwJmjoN+CYn
Mx/5+ImZb/MWiwO5KZUHy0pXwMjm02wPhlWJ1hphdsou1z/zwkrCHXrQRKKMtutH9QrXMVFdjtLJ
7d7ukuFW9lf7eFMVZnPDA3dSzPuqenEWBBj6Re1tQytPwBB1AKxLfVZLKGrDSp2EESiumhisRdNP
uaML2Wg8PkclSHo0xxN961e5XUa5fugvLuCqbJp+mywLxrZLpZdmKTZnkpa10EomP1PXPCHCnxaw
EXMcVoxrtdsIQ961GDHdxbm5fFtT7r1iVuZYYywnL+Y9UuZIY12o4fGPXcsMVxeYxyMw1frG1BTx
ufxllpmR3zzUGDpQu38pSXjJQysaxEkTtrJK30wWpJwTk5HaA8GdXPLjhvY7M7CeWI1QIhqtq2r7
cmmaDpbEXgc7AYi8OYap07aAbKvIBrqCsBg84GDntbnO/79RAi8v/TE4v4+z0qMTfnUdyhEQcX7o
1STl0pBmzB1JQeIX3CBQAaZ9O72A8XWH2jmKk0lBKC1gm5z8E9OFS9fpcVm4xjzsuUsFtpqGQpNi
UAmPPFt5f6Q1SxwrhnSpho4luGJMf/9BNVrp3/VFQjpXC3rl9S8nslklk2D59mtrdP7C5N8SeSIq
7bS20W7tQ1TPUQNc3DadYX9vQDJ6uEaJZJrU7bC0qSwCNW53MWOJOl4UyifR7kqa28jZQXf/55xw
a8GnUwgQ6o8UmO8Hpa6qjJXv/tkoWkHSyrK2pzH+MEGpVTIclwN5MwlFpuL8cXqOktBgzps25pJB
wWMipbG9RqfRFHqc+sT0HNmBNn9ityzwTDV/fGo3MdSvukpVNZ37V3GCakrkY6mg3dnrbUK3uCdd
kjMnJbpsFrpnjw9NntDIPlu9tunAwfvRponvgi1+Ej2gZQxVwpz6/e0hbGGaUsns/nNDvnzNfY2a
0eeOUu40209XqJcDxC23Trb32HSWYK4EFzER9pa6zznHzYYyqIz7bGajwWMwY/B7zI5voMrj2WR+
Go6hg2jGro/L9otYgO+UU9j1u6GprB9l4TYT8Wd4kfRzY0opt/0cJl5HEMr4Cuc6MzV9uimbelRu
JGR7p0cWFhKTTaWv6Qst7ZfLT3kMY5gNg+dqneUwY1SR6BqZJxUADYtqtVZwjQPHc27SvSMfrxwl
g43LUmdI6zhvQb0gZe48rixUvPGnldVTdVkBq7b/XGfZOuze2jkogWCjr/QFYSDBYGwwxIf1yvnr
+LSCzRH+HIs4CsCO0gei8GA6+u/iXKwQJs41v0707PoiaQFq8+9nUlhldwTiGLgA6lWOiWjm88M+
QLbXF6w/Mn0bJGOzCDSndn00yICUHCwOF0Lz4esrSXEsuB2zYfMkQDtb6Swy37H69xAGeHLdIQUX
bB1GAInSuspu+4lNNcCKR/oWCbEXV+FWzzYT8xdmSMQeCyDHbCwu5PClovrVp7eNWsHoOlu5Cxty
QxBNu9UNfJkKocitsWl5e8VfILwQDxx8u2HVQ5zwNDVWvrffhJW/Xa6h8FCisVr6hF6z2LQjXtRh
3cdDIg8nhhGM7P4lNlcgrZQ9BcLbwQn7S6SoyNCFLFbwMkahiBwT2WcvA+hx6q6fB/IzocpX1b6T
tt+fJ/18gLHy/WpBlYLI5S4VMRZWpB0vvbuWi0kg+UNg9PpxYfcvHGdNTNFWZPiFgfX1I5XpaARp
5ODDK4XTPOEBm8ruOJywVgjHakq4gaOQwZBYsJfaINuKxN4+EwKroXKAsDIcQdSN2F3bTad58CTh
3ajYl2Mp1/bRrI8K6ImP4+DLJP04zkhHcDWtQYL4Lxrjw49kfu85JWxBQMfeLxxBuZujGjad4i0a
H26yc8GM7WjAuYokQXYUO93uODFkSsdqZxzOiL2t93Jy7LrZcDz2IXFwt+7Lbs6NWr76U2xfn00G
iZ1vD9l9moZGMfo9tbI+eQzUh/W15EMrsTyLExieP/WDWsi7ZFKhq/R80vFftnn8BNYDQ0mK2Mm/
VTZ1nH/cWMf9yispIST0am00x1c8OrjZVck4L8P4ffmuPjtm9jYk1HHEzUvP1AalssSi7gbqfbud
7xQuzr7TSF4eyYoV9xjRuhuotBZtXqIgdPODQFAi6olzCjzmdG9bItq1dwGP14bPD5v8THxNAmD/
s4JLTp9Ggbp3v4Okn8/yJi8YyD2pJcCAX4WuYYxojchbvxNsXBIZnwhIFpvTSJlsZLBtEHPJvwBY
hW9r4giTq1hvoZ3KRGZr5mVLfVmmrsT+99sr85R/idfyMq/Y+5C5s4UKFXgzO8P+qVpMDfcLmDef
X0f3ZP5HfI6gWIoWI+fslPP95Jqr+M9Fgi5V0pasvhMxffBaed4/oLpSqkFSoZ0uI/pCDb6Bdgvf
Hy1SuZB0yim6UHYFcc+n8F2Z07cqFwvgTbafi4LIUGwxBQmwdqIcdkyJrl08DlLlXfKuTtVpwBiP
Y/1KyBbFrKNrGmMvQtTAlAXI698S6lW25O/+vM12IzBqthQqYUbHwSMdsodWzzuB1JcpAEqz4l4d
cCUgtpA6AbK0Y0VfeSnJ8Nr/Q3I9KnS3qJiEAijrVpN9dhkgYUQ3oea9yKPveWoWGu1PukjBYrgn
nMK2tI8T6s+Lhm6rXwEMKVVLVXXnQFp0UEfcP7u+6kOBvQRocxV+R5zacnJ0LEzbXwPnJxZehk3u
yh4S351q3q4IuiIsMIU9FBDTwTtoFj32sH8zbnszk3oVJfb04QJGAcG5kAHwQUygsEHO1N61K026
WVOzOK8H0vOuublgp5/bEUelJN2zx3ahieG9CszK69/i5CPl0mQsPNFflHGn7AfhLJCtuCCvTCCQ
QDz4HYJ8lHmS+tGHww8abtynGF1KLxgPVGdS2qk1mAkHu22tbGZHRsGNIfDb0vS9IRcqT73kQoAt
fNBQkX1LyXX3yPD1ED2cPVfBaYutlH7FXO7SROKInqiGy1FdWQ0AfGAE5ftuk5qJ2SGWxDeA3qAw
DewAwlCrNx8S0g9S1262vQv2ZBaZlMlpvr4cl19DKpnmdqJ3EIC72P8vRoMaRAY3hWZ7dz5kk9t3
kGxNXIK2LtekNsmBEJXRRJDEVudXSO9EOmsuZKHEbZ4V1YqrqD9huKgHKtwPEt7ncks4ZyaRAWLY
P4YWG8TA3qH2hiwYJlcPYth6nYdUS7ErHfh9Rt7ETvgdCKi6iHTq6mcjHBSwzxR/dNpwClf8xks1
cF7NuGi6ZGI8oNkFuHeNUFx6q8ZcGUbEyJtOXQFkiI/598MN+grPJiO3bW8HZrzhAZDxOPMTHr3P
C3MLtE1yhQx2dLSSBQj0hjSmnU2pGOWQksbt8MspyDdpLIbbJfGaXL7shs86U1gUzOiqnqylr+6Y
QxPCOGvqF+3pG9DIB9mlduWcOsJNS+c/qdbd49XWfdI/QOcSn1lDY0wD7+oiIxMZw1TbA19pHUIA
Orwu8MBkDy8FtSwTzWQwooePQVupKUd8WfBebgxMYZbjBONx7y3xXUnv/mANEVociZ3OIIiWS5l4
kGAtGYCmm8Szpc3SYFL3jidb0J0znulSuXGdvKo1xII70Q2prmAvh8Apn2POcI7aC2RRzzrlQ1wj
oGMBClVYvANGkeaYY/dPdmYnGPRQs3eWT1hKAejXvd3VqvBDXWCZz1yAOTc1+b5ccJfinC887p9j
ZmgpmfmlKCWVUO53JrEjRvIUPTL7KgaH+9fwWtcmENUf4Bp34Ph9TQf0moXO0hMVKA39FW+OmDyu
I4ffDJdlc4s7jWuxzjNUJig6wnLN7dAAN+ZPC1mCnjqOgYL0F3im1/k33nO0maU3xFHsfkHtFZ+o
xXf40YYRF3T63vWoSPIDLbFc39LU0gwLFT867Wkzz2haVmbNJTuyrkNK5OxIc0wuwFSi6ghA6XBX
op2+7l295/C2nsMEKGV/gAMZnjQNvV1aORSyNoUyqiDowvoNs/eaoa99pqAKVyrFMI/6euyUy3B6
bZzd3TCMmxpBFlUnuJzcj3fA3R8VZrPZxgQbSNGEFelRrHMYLUaRVryZkAQVftccYo3FsxzBCr/I
BMALuZ47xdpsP7M8lvPsrzvFyh3VxxDbK3Tl64UJZvRnxg13PIYi6QeOjQr0dKVMleVDkAzv4A1s
7hwzWn5TEEy0QjteNnAmQPBgjf7KBY+M2Rcr0j9jfrpyLweeg1ZoAyGuF2hUq/toaOKDLekRMe7w
oD1KdGVMWO7fKj+7yRFCuR2PEfGP9Ahdf5P1UL38xdBOxGzKoSWpNHYzR48bj9NKRy584OuTh8bG
kpEM5ZLzFB2txBh1vfYE6AcZiYLPVgAMF0zehUB1BOFot5EeO/WZGBtqH3C/sd3fXC7+RHyXxiTR
cgGSK+UXXZ8QyW91ErUOKY7jeRq0d81rTS8fAWhU/YS+MR+3zpWVOVhm2SkocIs0sPjFH5Yg48sq
IyQDm9cE2Qnjiy3qX/E6pbx/uh8o3G6mNTqUgRshylyHGCSO+MNTAwM1STxDjWjYJjWcf75xL9mn
X3e33A/EtdJY8exC3RdTlWeNlqOab71ivq8NKzPMqWemq63F0qRllpJljS/ipl/CZ077my2o1+58
nneeoAu/U0lhLZxDGVLKvPGNg57haCnSgqSZKa9oLFya7pgKCwkWwRZaP5xVcfquFazafE0Pxk5f
b3i9a8IZkMcMfb7fhjMs/Hxv14m97XQHdwikgSeGEucbupqT+e4ulUvRpX+KXvozqKz4isdH7WuY
BZzHq7vF40WN39azzs9/D3tJdSmvNQbrXDm0prmnTuS3Rz9IpPp/mCHkX4/Ix+8slkmC/0zX/tFM
5WRqS3biT/0JBjvNPJ1qnD1kXH6qRw5FwgsESX2iEsUXnoLXuA/WmQdZko89pa/et2Rvoo8yEz1k
2akuYsRsOhAVLI35/b1+g/STNKV9DMgGHSp6l/YiXwLUgBuLYc7/EGuhuDlHRdTuQw4E6IcioxHC
IGH4Zl7J23/Fzs5Qx+A1XYWVhysNxb5fn5pIuQfmC2OGPu13zVywP5ESS5+DEFg9sfcg/xyfAOSP
Rs/tIB4+xhLLtXzHbz4WkuJld6N8jpo6Pp43XX8niauY4QnGpDE9aKUDgxcq+iEC1NJ0v8iWZJpf
WSaj+FJSRP6fJoWFZOQX643yVElhW3Dmu65SLDXvzkZ7dEezRHDwiv43v9wmIpPqIIqtzbXDMusy
1iEZK3PIfRTaGr+0a0MLwCYiomDOw/uVF77vEJDLJiHkggeh7sq5Pe3/8flmXgdrT1tucRmiwoig
8SjXcMCmBpdfizUFmOFu2PFf+eBQcl5JVvv24490Hgz8mSk/jZI3gNtXUXMO1xXxa7xpN80E068C
oR9HqMmHobLmfO4Gc7wATBjYD8NTOqxN2FXYcbofuvIvEgD3sHxU2OJC+dZrRMvGRzBQK2Ul7tpy
yTZrYohZuDssH+GuWT3s68/Zfyi7jngb6DlbH78BruunHl7GUfRBVjN1aUKUDvVpZE2nr58oFogQ
mtTUNDsXEpD/Aq7RNND/3BaBPKveqi6w52MYh8lC3ohDDm4X028VNyvDB7l8lgZaNzim/WOpluYH
IGivY/XluoV5vdbX3wlH7BnOI9wrKsbGRkv9QwhX/0pIeUGDXuXtZwIV1F9VSNbcsAysGqLYz01R
0p/5VvOejX204aruDf8D4XHyqzZ0hdUS1Ng1MWnrU2rVjgJOJoj45c1+/1qUlCvxeOeJ9e3+N9AY
2J/EN/2O+FC7Vbi5BWnTb/obnUw6lzDZ/1kxRcCQyvBpjzAQ7U0yhIe3xQhxtZSQfGwipfCLyhUz
sI3MlcxRmwVU8f118tSOSz9i8a/0eFoHO4lE95wtYvNu2Xp0aSx9ZcKadx1pPmZ/BIjQMhJijfTL
VT+joStkSNFlkZuUIyQ7Q8h3LJxWLy0nsZWHLKJhcgiIT2WKLB7C7KsE2GMApkDKArWYr35sPwBi
Mz4GyOAoVWtSUfRbWzPF7rSRdGiRowNnVEmtlB9vfqT0Mr/QqvweWeDetUgUcEvywhAyurUbqTal
oTLEKHdyBigGnqysJs7kLGZOWXz4R7ri8dvendsEiVzv68S1DNbAqrDRostRRfW3opCESKxiNFB3
DZ4lkPdeGakdsJlg9W5wenKklEpdlQhpdOHtDlRoiraO1lizWSiiYJ8MPEvfJTneHTXNWeJDzXwd
CwtM6uSu6wSS7ZMq16fkLCkbUzzCXHu+hl0kQThfONf1mq/Fj+huaoMbQFnDUfn9OHMcZTth36pT
Ls8/dtr12P7jrCd7rxJqjTSLcJmSxq9TVKqM+gvxaMWbiysq2e0ZRwBNwcgOLh2JUNdjngLkOX1x
tzX8MeoBW3g0OfU7hQLky/ggLRx3Iyb9hGGGXASwJq2FsWzN3/nEoxjj21syz33fZ8d5akFFCxm1
87J5YPnQpnecdDfk1Bu2qc3mE5wdsdWrD1jtaqlGbaBoZ7mxeLI1QEEcnnIIHfGgs1dH7LbLX2lu
0xmfBIQkR7YsDHMiKtZfTNFgdmt9pG4JsarztzIh5eIUYm3t1EEymDaRanzwbPCvLqZivR+ZCuzP
hmeSVdlGVo54AzhaqMauui33xB4yhIRZvrY4nIzOYKcuKSdVf+Jjt6+iGuoHyCPLQuLAsbkLTWkc
X7l62/R5/zRcs+9g1pyWeuegZR8YJr0K0MZO2hV9iqHlK9DL3IylU6JtsTg4PuBtUgUVLAeTJaz+
i3F1OTzwGa0svy2LvcI+T1+mUcb2erfSVAuw/bIDzBkOOs8KvvU2dZBNGNSD6Xfwe76ae1JLLuxx
hZSUBq3QNivI4BXb/pGig+87ryqdJhoItXVtpxh0HbYP0bfLVY8dJOoipZJdZfOm+4C0/oTO/l9z
fTkfZ8PpGNwrNDr8IgngsB2RdDoSXPrOueKwmEgU9EExSTxNSnz6cVRxd+okHp7vcp56DAMq4ss7
2kr06C+C7I8uEm2m15B4rr3TtpOVVzxwy1cPE3viUs0ggs3iUNWARMnfLgzWyhkAoxKYx29NECmp
yORHfkO7m1/JyQU57KW/bcoG57mIKx9qH6hILtjaDoiTGqZYLs3bY76qSSlYlfq9jylxdIvWsQSx
U+4jYvnVrqRL4L8dwaEqCjDLgZbYySF5cl03SIg/RWptbaUS8cRzolNTyLvKqbm92eyLBpWveyZH
4As39SxYOet6UH1NIz8Lo9FrMasZf71Cv7MhhUNCVJhTyAermLhYu0uczHinQFkA5yrABpZStZxO
lH5xqHdI0y9RyBw4dPOp1GPDTCirl3pZdXfhE95Wg4MpxSzwy+TROuM7E243kXhMzTKrKbl77IHK
HsMZgv/Gw781jv3cHW1tSaAfH5X/qxOBD2dfgnDbQAYNONSLP/nb+UKgU+fwQAN8MjyCttPIXxb3
n4A+jqjVP7vFxOOB9EneGzsWXoePOKlsXmiXaG4sPL0M2riUrTFFuNEy6z8VTOPtRlzEPVmYKg6v
q5NUcITHj8ipPIp8gfV2+Ta0uDM5IxRLBMFQE0MYhhcj0VFKqFCqws/jS/JZNIO74/DBnVewFEkr
KHYyWBWrhTIiug+StV+cwaf5kuviA6ZdsRp0A5UIUpy/sA4La/OxPCs8igT4l/xjWtdAz7opgeMs
yh07JsYYPvzCqjAYZ5LBsgK6ViQKCTYy0rj2+tHIPLfGAlWZ2sXqtJISfROHYpMnLLV7shkTWtwR
GxRvPqOjlKmLb8Wpt466O8MHgr4fWkMLi/X1pTHM0PZotiadRijR6T8iHkuqUyRwOTVN4+6V1pFg
S2qAbwD1G6T+yqXmOkklU2llqIIDcspEJuaBqmiayU03ujWArev4wjKkM1nEQBXCP+huOwC3hnZO
PmGOgYuDs/CmLN1UNRLYz/ob7nDSJ380ncaQWmnPnB6HYlHcTXWAx6jIYRoY3/W//xy+pLiqRgfx
VoKnanpWPeg4SkQzhImI5qEUAZ2Q+iHkpd/RAA/APBu4Q0b6nSXStiO6hXmBOB0ABXofc/Fv+uUY
zBBwoo8+IbFTZIN9Ts6nSIxYpfaLJJZHWI2v69p3Qq9Y8aavLT1vZeRyt41AZpkiVyYEfK4E3ffN
FoZe9Fv/EDB2MkgYjyoNI7Z+2IPV6BTMfY3P5vmUaWgivi+GV7dXYGzU0uOfn7h9zrXJv6VaICZ6
jkC1U4XqO5u3uJ2ecAuYGVpq8g7EzHOJUn2pp1W13ZTD/4EqKCArIyD+TNIjAYuMfrwyVTY/LtNv
5BBhmjflREUfMM8N75ILKneXL7wvMRYJrRgnLJnX4YzLPowDR/v1K+s7qgC1Z3rBZWNW0aQ1dSsL
l6M5+MWYqTSKCNVz3GSt4//AaSxLEvgTkn4GavT/LHfFF5H8FtP/IkCCsVaBquatwmgbThW1lCRl
q6W71x0F5CoXoDCrWMbmeVrDjhcasuwREwbduH4oYbiSe8ArMOtA3qAFNyA6sHhIlPQSMmK2LHqS
KUJM4e9a+wN1TL3Ir+faA0EgRHtPPP74IBT4eRhM6bmF6oGQbR2wieU1KMn+Gt7EmNNyTWS7A8Tt
eWNvabzKR/cHw4QRXXQuvWQ5azBNXY+yrS68mwgMKegPJ56SFIpzfZh5tngm+0T0dE1DHnhyK7fE
UbpxfRQEdCNoDowtyMZq4D0d6auVytIg9ltzgj2D8z4EYZ7+EdtvByAe/+yvBxF0B4/kN/D7IUcy
UWymRGqKoWqm5XtMQiZdBgyebZka/KBsVfQi/hLGaULCDQ5zjN7QYl8QW0bsSrUDNOZZ6Exuz2Fw
mqGSYP6g2tctcejigJeSK+Ol+YYoSsyLfjRvL1rQ+DR4dvKuVy/s7G4BuRLXPdbZJ+DhSZzglTqy
riroofd5Scpvb+QuqnqAXX9JHTqb9+HcZBqaDj8xDm9SRGRBNXv9XCzj8+6YFMxV6OElxLOqvWZz
YfIeP3fbCfJX+HEF+uZ9dteMqA2ELG9uy2Kie8UKUJSbMo888YWGIYYgoLoGozFh/8+FTFJ6XlRP
hBW5hzt9ncGsKSIl844IAqrsxVg9kRad7Uv4/qK3Th2NOfHAY0bK1pz6NkaSnbt86u4cEcnqXuRU
+OIuDCD2OyVHQIwT7kX68VzuV8H+zWtp5bjiub/SStm4hRrJB/AY3K3kLZJBcd1B433G03NNNnIe
027B/XWTbTM5bGwhNgCdbTTaM+/PSJfHGyY18T48mkYGjdt+CWe2sBaU19k60TJxWAJskS8jNrPU
c/oKBpwwQIxiGeG6O6N8XOfihug4X4s1aE9//jINlQkJ4H75D04FZsmdIk7mPF1fpHJT3Q8najrd
/0yCC2dFtrsfG1YmTR1kRWhiWBuTwpaQ0jr+7WexsQSLAcCjHLnXSBUDnAlGpf2iC4m3c1MKireR
s8uGneI+3vfdsyw+Gbjl4fP8/POE8N8hY4UnYbAYugU9YgzRMupefFhhPECmf2RWPs8J0zzuCf2j
DKYo72De54U+EGh9yJJe5kJ1m6mFZM/bDs+nVziUp7x1yVX7exStYQK/nQrkKrrB4pY8Dw/xg53j
x2me8WM9n2UtfkX8pvvdmjpkBDzk1lbtD7yB7xF/IVmU5xrUW6USuosnFjiwAdbioDvz3w7+xo2m
WafA0U5xqgzhAoX68b82QS7Hyn1ZRnTo4YCisgTsk0MqNT16eGJPfKqj836cFuPsvmA4yYReUUJ3
3LdWvS+AmnZeQQ5Q0DPF8zvn/824BBXTYhTex7CBRhRPlQ93Y+tt4hHpCM/YB9KWNUB0bQFSXS4I
u9cXFcVXJ6MWH8ToNXaNwUjjqzvu7t1oO1375qBPtwY3GaNcOQANb0aoxerBZUYN/jXrvoLliAkz
hDgSQHbnPUZflBcZ0Jnl+0fMuI/ZnO3h9f+4QO0kes3s0VopkByYCNXXCXdQ9CWUOI7SB2r3Npgs
R5FaGVfsOjn6Srj9h0zi9zFtM4JVPnyHofky5QP2kOtYvfoDZvoTcnvlmM/MmIdhMcRN+Vnp2370
YBn+az1bngIW2fhlU/OdHgYoHF2vSYZ+02uU2OPPJnxRIfXjbPDO0gqa8f/cw/7Z4R9Bdx+V4ovV
6us/EKqWEPFAimSi4wSXjnUK0DQUf1ScrXt8Y5qb40RtCGRyr/DUOAhCxCM6SqZ0dWjUVq58TRTW
A3a9dXP1r9iLxfhdAZURWb1ZbrcsWv9CsFeRsJ1aNQBjCfP/1e9bAFluqHD2t1tWFP0IdfewcGqY
4f6wAP80bTDTpR9OyQW3vpWnH1MwrQQ+Zw8fU8kARX6vJr1H2Nn9wiikoDBWhQI8KRBv0NohT3Ud
3WRLxfbPGwu42tgg2bjrkma9n12UCOg8KpDQmt9Na6RvHGKdX3smSm5sZXRjwciGBpIlPGM2kTGB
nXMkz9NeQkQ94nVo8KLnYd3wM1bmak5QoVhBE/b3RfVvvns65AKPgFt+Qa0w8to196DNiUkAei2K
hEkxvUU7i3MlvEq1Igy2T/BjNWMtOQludFMrRzenhK4uV75r5/RlP5SvZk6JhW7bDYIflPNqdf/s
g+cYn+4sN4IJ6eTeAIQPKR33T2euyzXDF/kksMyvixBaBNP8/10wfRkwqVIlht4wQ736uY446dfa
EqqpKYnepMNEEh0eUe8qdqXAoBmM9Rid7cTwj8Zl/LWtmsjM4lfceanaaMLz7E8xC0WhLH+K7eqr
kB7bUZZ7X4OQ6D9nHjcZ/3w1GzGNvPX76M5SpH4ParoQ+P/2aHBHK+E7/emmEZuPaPtWZdoMiYwH
3Ax+wp9SR+gzbRGOPz9E5RW6VOY2XzppAD2/Qevh0C+5+LnTUkeSgbnJcRY3hG88U2VmhdhZcfYb
VMec6wq1iasUoFyDXA4/GEKA/NJ5lXKbQQGnUej0v4mishXIikLiRjyAzwjeqbCTwP7bjeJDs0Sj
ueqlGu8eJTEDl8nHM7ajfxPqyZmEwUfsfDbBHwuMMKSFwrHrMllEN3rlgIvGuxmvV3+acAtR4Y3L
ONpqFbzbIDwoJq2gcDQI5HcP5EG+u2jkSLxBOJpqwYyO+G/qU5+dy1H4+23uWu/JJSO6tQOoltpU
SXoA5pBsQWHuSn3nUUte9SnZ5Gp0bwemjCNUJFsJIiv817PU5zEn94PLvfLVeKkSq0uVMF2Lkuti
k3DHQSLqFupM8pQjXbsvJeplAL9qOgriNBmGFe0vHWkMu1nPfcKr7joF7pui2cnWLMbZ5WvuDnxk
COUmK/BQ1zAx1iTRi3vuis87ceUN9LnU+dXkuhXS0Z8QarMBMXev/nKxVa6CgavgfdYUH2dbgTsa
cxDSFgxt0epipIxXLTxYqUimiCW74F1qSYDIQopQEYW9nj7Rxps0XT9YqFtVJpJdknd7MhKGkBBU
92VXSgl3w9r6UngPkWosdYGf6DENyJlvGKzvPhQG81CjKPjEJu6/+ltkWb1ImaekardeQN1IANZU
bYNfGzMgpSIoI2ugJZEP+KLlzZ9KQvD3ty0P59vGmra0ys7RTSoGk8bGfRc58LhNdCUIjHyN2K/C
vYp3g+tyGbx76DX99P60ydgItJvurZXnIdrtusVe/TO6e+AkoqPqkJUAEPTwZqrs0QkDFXjiP+dx
5PntwH//O3wj49b56vbejzvim1U25xh/0idgTRWquJAqwjQUAN4Z3H/zvsZPsTyr/ETIeV/UDmck
AiqB1blzOt2hGVlgNJND+3exiX4VXUFEySzhIjtI5yXzaIRjBZWPqZnAhNMhW/1jlsJA+4oImriM
UFV/TgYynDGgXuWGRuQv9G490VRClC4PtSh3Q1ZQ6J1XwHiRM9CqHUUglClhmbzQvA54/hlW84AA
OozLjSO3TzNl6ct679cvK1UZiqZsqncw2cfXHdSvfSADLyOsR6jHlit0cNjzhZBNRgfotAW3sdTJ
YOV3mdmvyGROEmNzTylxylbrbtQO0AlhRFeTLrJsDKPMe4RK74CVuznIFF71mYiCb4X91Q/eIHxp
qzOKkLpgwgiyCRofW/QKHWb+vKqziSyF0huyst4Y4i/b2XD0SE97Pa7Zv+qf4Fwd3IaQDUE59JV+
68xj9RoX2JXNzxn8uUH0eTkWRrpq6SCr8U6z/1Pqj8XoaIY0noV0OPE4Xi3kQJ74dfG1HgmeUxQh
8uLH3UsPwHXXtZzi1QzZkSEGoHxrivLckAXJ4v/Y1hVGiwOI1JSZxjfcvyRBGH1TbWwRfNLm2kgL
vrOCDVekmzd2kRkARzS7O2uN7djEPYaGKqu5fqGzBSxDoF+XIpNJ853yrdB9ZwOCWdbIQYd/cyPz
KWIiBI58eX8YtXy/k4J7J5gK1tBtjjM3LvgmaWOTDX4OkA9AWcPuIK2ox2jslYPYZYedGkhDdw+Y
zJmAxhIRYFclHl2wZBMu5Kr0k3f3bueSslfciVhRKyPckWyiRWaeKDO21z5Cv6XJO5bOg9kOnfBz
Lx0YLazbzslBhD+1RbmQwr99xu9KJTONkUpsK+wj+iDzN+y2zuvrZQ2x5deCXu7jZmhX810Hcge3
6n+OxoqYwPvV2imGlXPC034DAD5VEIaOoCzE3wZTVQ3ZXUINIxKTzGWcywLkknP0/WP5SBfWzkL0
dPrscvLMYRgmQ+L/jQFSdFxsj3A7leocmG9tiajINLc7SG1HSfrKdLDr4vhPx2Qm8sMR/cUF296E
JKujaEFly5nNhFrJOXHAbQp2bKl6eF3jqrAZVr5DkBnJqiCwk2g9cUaPUy3fDp6DO4Be4mJstgOG
LUE/FLgJ5PyFwwyOG+sGk/+aQafwOHRC0/431VI5yIcBXB9YDfOhxZEpQXO4imldTQjuo6DuqcCr
9aX/y/+FwZg2eppSg8xpbUGDWePc6H1WeqMeSsF2RuUouiATNamWnIN4u7xxcQhwj/1ycqmd2ZsY
QVuE0Va8KrMoDTnLxjjARjDtW4nJVmF4Rm8eNuzvlqHDAOe3qUX4kmCSgifLEpB4RWZgB4QvLTaA
FAec2XFO47g3uZyObzVij/ZM2HYJ5rBtqfgD5JUWjGJbUzf3oviIkC4x7+51maVNvC+cK5s6GM6q
m5L677REOoDZcoZFM40x/8pnNC6nCNaxQ/aZhu3D2lq2scLPSod1X+QPT1MEyfR4ik7JuZ6yMbxL
XittSxw/XVZyWI5QAXHSD3AERbLi8rnV9lAYu4G5naPdtoIZeio/6FcwyTNvH1WvcVWOoPSknHaY
8B1em2dXeN7Wkbp9+JVdI95kGTfj6I0CYLMzbkrK7vf1NC+8UD8c8Ah9RJFXmjBZSndJC9SpruRY
zKxxe+qNVBAN+ja6sg1/rU1O3XYc2T/R/xkqjKzh6xUeTUZwuuf/7dyu7FMwptTrym4Af1vhxVC9
6g8rY5z3GaDunbdt2OW8kNBKt4F8iynhByJXk1kOjBwIKekr/8iMv0ynD3CaDw1pdPiXBmo9fQ0G
t4HnTM1WzjAXUDRwway+qk/evo/XfwIGY+97Yd+vT9/FN14OdY2X3PEW6iisQKLdFD/5ficKLvQ/
gnCXF/BRrCo5D42a/thm1OY+THsFftek6zcC8u5mFf8Io6l2aWZ+1n0Wf5sjEFZpNvREyECkfCnK
z6Zu7yo1YhqwenOAQWEWVvchRG4aJXJv9bC085TZlx77UTyNO3tYyy5H06vpPRbN3qdJLpS5bt5e
RRAN+JEebKB0aghAJflhT/U77N0o8IA0oSk05H2m0/1ZORIhFB4wxBTkYVhrvQ9X61Hw9AGDgq6g
rWcKzB4uS6MLaZuQHtpdKYQj4JQaifXBdJd3l55f+XV0sJx9FYz6iAcErhGE4aHx+r0AXxn8vlqE
ZxJiy/6m6VAem2uLepE1k8wsDTyMcfr3DFm3+ZshcR3VALKAXABmzN7tENMh1WEDuRwWb8f9nPGL
xArMXvCoIi1pyfGAyiKj2JgoCYotMgJLvJpLYgv31M2FIsc+nzThOfSUUCloNGOW9AAxnhbZZdgm
rhv2m8ZiDBQGcNOZsDJpxAHMT7uesxPI20M7mvxqzqLnBYFC6GtimXU09fdKh0ohkbWZwK6ToC4R
s+31U/UN1Uf2pr5Ahr7RnemvC5rvjdpzpBw+3BewMs3FlbnWrU2eqXfcPRP0deh3OOgz896VJTo2
JGysiQcG1pF9ianGb/OreL9e1tqZu2cJEODDVX9Z4Tp9BgBz7114RoEaI8gVc6Gj+NvRqxu8Rpv3
8mbN0/ZAB/s+4+LTxViDkZM74CuaLujqcjqQ6j2pVK5PyeZ89OW6f0GdT3kFJnGkV5jbCXQtCZ4A
I4S5YW/Y6sc+PDbTr9uLALWODvs4uGbZlQwPHjXa6D1JfX8b0x+R1OQhwtDLB+MV5j65DUcaSy/u
VbYq9cGz3w4EasF6kmllnb/lB9lv+HMFBU19M4GZWNShUfqTtFpX4jTB61/bm9VuCU9EjjDfJ4S4
UrSy0E1PRfD/eqF0oMKeTIr2v7G3XEGPEDheJS4SPoT/sgtWj8vulKt7MMMbC5LdB2CHuIVSxQlQ
sf6IK9lgiqqW50M5UP9PGVEhnzluvxhTfG5YLFYYyraY6bWfIR8ZYOLbPZamMizgH2ZUgcx/Kk1K
VfK+WVbDVAhYX5FD+JBSkiSDS0RlqB8g69AO1pO6w2Ry6ybZtNqPwyALztmCxVehVfEB/qwjnqZz
x4RQS0q+AIGzkbgMiCfFDziQb6zPexsEiBA5i6kHgKqiK/X51vq3QbkxcipiPt0sLmhFi7Of6hpx
L1sWw7TzuHLvK7ZlyS8qt2eHSLksIuMbKguASSlntAFqCQ71Q1cMsf2/LFuYqnsgDkInaGbwQ4eS
IBcDBD+MyXDnDr+eHBTRXrSovCQ6CSFMeNkjPwlpOPIZSE1RAXXO0RhGZGtY9uvyuqt7RF1cSvyX
z8iJfWnsC5tdft7eYT33Da6IRhiNFo/QR1k8pcuNAfmz9fZHi6J2lK9ZlOW9ZOG3WoItDvVCJFB2
m8et+x8btmChXpOia0r9bvbAhno0QTOk/gZL03ZmCgAw4KppDGB7pD+xpFD3iXl6W2k/q55Q/dMF
nTYJpA5p4vTdKdOq1Q4N3TKC+hgfyW0pcl25nUXx04B7rAiyV0im+RdZy/LsbmMIBK/53XdErDOB
KgydV3e0tBh2RunxyeK7aHsF4mfwTcXQG3PnCbqLQpK/x1MHrAb3ejzsxEsxq9cJ30btjLGwcU2n
zlTqZFlKe1BwyQw5erf0WPRzm/TDAAZOatIF2uUMtdcIwOpnTSYpsWX1aP3TPuU6w6V55rHAUtU7
QfvSNVMsAcjrPSO+JaFPUWDyANH+uHvzyPJKs3xawO9+rkogMAf04Rn7tf8cTqy5IT5F1M1zzX04
2BM7A+plTX6duLi0xhpW1dzg+AMBpg6Zb1kiv7R2BgA1lqo16rxU8hqpWPMmA4Sbk4YIecnPLpFD
+Qt85MuUzOrN6/kwrudfL16YMhnfqA6u29s9LM8iyP+/EmSibDIrhvEb4CGbnGNwV301djhlH/Wa
WCCSmFwavL7jB30f+LZqiLY34kIIBs4iM+dKT5pSnJWI7rHqfLEkOBxUCcoM6wCoFGEIYzRzP2Qt
Vno7xftbLTLFQyl11bsXlTAffnT9ezf+8Cc2+/0gBeexL04t7x4x4wZ2bHwY6j/qdWlPFzk1aDsc
o10w+OQtFseiR6DQmQauniBhKmhIkzUI8fU7+ztQUSHnwVizVevRSW1lBgQOMFOiDhJCQNxEPWps
WrQIjIUeqoLJbSmlAYBFiN2Qa37UpyjYesoQqOkd4IngzjwmIhkBjY6HLf0cXGzQORasqnTDCaEg
hwsvrJpzpr3BNXHOCi+EiufSF+kD/Wt/1oYcypxKKAwhC1wJz8N+wpLX9luTgS+HEaJUmgZ6gjqu
PjD47ubIoX+be0w5gI0U+Z/Sll8aSlHV4AXf2hoyKnUb9hLe9ZOhlpiig3trvg1t3T9snhW8nbM+
kKFh+NUAGISE/U8eKSV7xQEPNi5pn87eaqMYWYixJMv9KRNAnh0GKZMLSK1Ro7OXWpW3YWga6Q9i
jpX45Hrm/b6dWB9MqL5B7ySWsnW+WDDfFA7QqXQLvBIvSzcNNkAWN5VPGHz75gHR/ZYAgCQq2phe
fNYKKQsQPNVsC6/3Ev6CVfhb11iqv9uvSBjh3mZAIyQzqfmaaCdQ9Z1wqEr5DPX5daekWK0OFM3K
vFDWrEXGc8QTAsOpyGJyCmVyKPE9Wd+MdNiqq+afdrkcnqePopWl693s5+BnwQG9ZDhdEytIOicV
cW7nkNFr3EucZ99fmEO9EG3uaep9/d9LPebvGjp86pQLllQiIx8TQ55gD5TsQL3UmGYF1yc3gVC7
QvnnPMJeHFkVCJjdExLHVU/1eLwdKfMq/EGNUck7tz80/+D8WndZVM/gXlUDP7mUlAKj0anNHEI2
Lc6xE0GM/nJqIx6AR9cBw1iuKeKBNBJAN29hLLSUqpKwoiw1kCEYCvKCbdrjhVqU/78naufBo5ou
SqFeHlWBFUO5woZA9tpn8xyeBvsLuVHax8Pectfg1FuJb7wm3KpLeo8zPw4gDaZfUaeNhYB5DiCC
nr/D9lIJqXklOeUm/Aep52i2BYhnLDCwOgm3eg57izjMc8ko5ILX9WeaJm7Qx0M+bMEScmv9vJDE
Lsv36VJpaJiPrnfwCqAGbT3j+ulpTuec+x0nkfj9IdEIHiny0X6zUMz9x/tZTBXGTFZirhbFLwlW
xbEf22RQ/VHNJkZEc7yJDiTOjQ2AKxNok0f8KdhmBhE+4Yd6MiHAjpENdOTQstul0fb2v7jiEzX+
M0UNRVFPTZxuee3wyGBRNVJm38eSPm7cgR9O30uP1kBhhNDOwiuL398WVrnHr7+qr4FR889upqiV
ID/m70Wcmvn1tq1PGfMq434wLcTM+jChyXnnN/cwGnudnrlUxqIsJCJ6lqgFRyLZOxOcZbTVEs8Z
2wesLGNY6ZJ5ufGgdwb3+oFWCZdd7/uGpiV0aJqzEreT600ZGFHa3nnchdAjXXeW5EO9ALov4Imb
nEdpy6Zv+3a6wRE1kn8SbkNyJWU2sHBlyJNjmt3VZfV4LX2jqVHzualvvnBwYK+swppJua+eaQfW
5o4eBkXJqqzpzxqR00EOwO2TvggujTI/FYDjMDhSeFF9dzMOOnyGD3Agx+Dzsju6KZ04cbEnq9eI
KBBNxsqkmK2L8eu5lVAqMEfgBhX37q/WjO/vBMb3rkh5zGOp+374Xkyk7kEqcn0abmR3vciQrTyM
H/aLKA8SteQRNhok3L+Tv5LHmKm6ldjMaFnJNMt2DpEBBkYiJTL8Dhq7/GJNxsWcVklG4IKSV7zl
gII4rpiCedAT4fPn32n+Xb86GUdhoneior997efE+mt71VZonv1jAduZYLcTHhrV1tzCUMYd4Sol
YQcJySPdoHi41ZornO/HqW2Vp1ogyVrlguzY8fD0cWbWhvpsO2FiQ2TfHUPxLEjTEUMzzfEgBuCE
Wlj3qN/NUypyN5pOm8AsYo2IIl7mw8X5OqeQ+OnNwYTbYC3VxoUKaHQieBdGmadp8LT00PQggGdf
5l3oiil8elIxH5WO7joEnqGmndvsSlYOGnJEdW5kgsZQYIw2k1pLvEFGcpMeC2+osSVJHmiu5Mc3
u9yLSdrG5sqO/9GKsW8w2C/qrkuVVyUahzSJhIe1AUVdoDEoFPaHuKbob250xa9jBfwPY4Y0vXaW
rKIIGi7RdNB8+iAtXE3GneNAY9GQ2LU2+62NXZjhOqz9riSCGgFM6qw67LMRqQAkwjN+SHWqFujg
cbyA8DGkVv12xPaLkpfdKmxWsp8O20hC2rSialDEEmAjzEDMkJmXgEr04kJ3sCQWz0tNmEvqpYpT
QKRdgSWIhlxJpJa6MvMw+s99kGHhJEGDdKRxef6gWD+CJ3UR0+Y7JSiPV+yurI83p/Bzi3ni30+X
vqq9kV9F+gkDhQxFBIfhGLIK0eCchdMEL0PavtlEVv5BdsqYIccJI0+HSvLZWdzNIOInPPFWMaax
cu68mK1Caz5RhzxIf0zuTGIxyrPGJbY3fFKRde7cL6ca0mYVnLmEcM/kNNvr8J3IXAf8zSgrNNlK
R141VhXmWyEJ/fzv6EFjIrLYHaWDfaD7Hn4VMt2E1ij8K1/uKrQf8TLXAyJGJnISUZs6jU9KrGCa
wYM8piicd9740+LToIti1oX+tAtTdZcAGqGhYUZHT9kHfA5TfZv0JplUkfePf5WBwXJo+/0z5Bl5
bqkZfZDkvfIzJnyXECtkreS0efJk+jZ7ZzKfuuFtSQLJtvAbQlemF+GMlZNjQ01mMv085Eduag/G
8uYd3If+URXF1uNGG3KMBWQB4661hOBBYZJGi7z/O0PtPPo5iI23yvIrU4SZrHMc4R9VBoWAE88A
n5fCfzYQmC5/e3EfhzZsaF5TQzekLsUOXyezVWkaTCK9k+B8syUaLQF28XYigt1BG7o2VKBP2zja
OtMtgsgrf7owWwfON4n5YBnj7X6l5FpdFRdx18jGom8hrurvgVnq0pHLwgxoaXYToTG5LsQZbSx+
CuLXL+Vu2MYM/xSmPNlcj16+1UKSe76YGLxZC0zYXR3cBxwKRWezJ7YFF6nvAseem2oX97z5ZXZX
eaZcKCAApT2GB8Jym8utd1sMShdhrsyjEJboVONQrXQygSglV2NYXQMG1q4JQSJdR+kzGHyFC33+
m3qZOq/UABrdSulCBiJaVDkGyl50LyRKOdmpiA+zAEb8aOHCDYI0qeBvRq2HmgdtRBJ537/vjjAx
nvWb4VcuBZHNHNeXd+eenz6JzAjyqrAvjcVmZIr99nj237XF+i+O6rYbhX+dkOWae5hDaK/oZkYV
5IzUuFZWTeqUcC69ngpRUsSp2EtQEorS5SILIkOUR1RUjAsKGO/3H4aA64CGJiqo+FslKBKYOXpB
C8YK/YDh+2ZKDr4jQAZ8fONOeUQk32nf2pHz0RcA4AZKeBdy7HSh6cJNLDZhYma0Q2peOc+a7XIf
Sv9/7jXm0nWTGsY1cKfRl4qc1OUwOxMADjHwekWCr3GEGimHA0QbnwrsMBRAbmsqADwaBo8hwIi0
dFr9dTBk+RA4k2NB0I94Z5SMtl9ORwMiO01gYAOodW+SMU7AkVY6fDlyUNngiT+P5wXH/4W19O3f
3PU0nttUTzmDs/cKoF5qvMUT4gLxRoBDucazPYaZZ3aILFsBmCvecok7YLt+18OZm6R7SVO4zA88
FeT93vFxOu0MUGqO891AX2KamSJOxen7LzruCYXBa1KJYP5yIvYx13tmTXr8ydkKb1jzVgU4Mpuc
EZc/IOpzU1iBjr9YtIjW7mVH6p/TVBzEHfLEpXLHprqGMCyuR5+8siZkjDq0rQluHTSrDFCgJqQ1
JCHimccM5PROrHU5hY8mp/VUK3it7I86a886oe65rX+Cts3oWNhfDDrCF8JZ03qOL6JsdQoujVa7
jMF+fk9S2vHBnHOEuxLTdOm4VronX/EHF99NBtRfs6nR2pCFYz97rWdI29ruLTNWIvF70FnD5Cxr
Lkn0tycJQ4Mr20gIzcNxZWaeR+crH5o4FE/nj4wv4ki/mAVNyJUN+f/WzBtkeKb1UUIKbFANORsG
M7PAnwpGZn2MxAxWMYyxuOw8628ptLKsnmxdr46bRjRkjFAWQYKMlnAR+gopQQNsb67BXZM6TM9E
qpyxGZ9LQ4+NvOCHdmJ9JhH8R8L5VETaENShi/H3vEUnpX8vINOjI4hcEIhJZLMTVJEKdONCClW7
lK0tFh12prziJPPEBnOuBY/pMtej9NFIFm131KhCWgMZ0H6mw1HlXkJLpDIxBufJ0mOfQDRheNS/
ZpJh1tZUGUx/t5ffW/ZIHkUX615/iqPTa8dSyDrwtLnmy5ljaPGkRlnADOpEBRkgvCARrGO3W9l5
iC/4LBhuK7RS3LsAPrLxeUeFbz2SjXKITirdPKIJM5ZgTyBmxcTU35BSRhy292E5HFTKPrqQuRIF
rgnJ/P+/64Pdq707nyJ3o7NeLtqcruQ6cz2DICXHFdY8dRh3jhOQ2ppscgurPNbgHAgfDwePvDpV
sjp9+BEuio8GNWR+o8atei2lGlJ4lm3jkHM1CgwJ82exc9WHMc4y1LpxiqHfAyt36tRKFeW+T2oB
/RMvu0tcKdXWATYakNY7Mz5GOIeOII8SBrhMx/vTGFOKNE6LaifN8Jr4FNSDudnB7OMCOkdOHueP
PTb9SlzuQW5zMYoQPfujcLUb/yRMENvUESDA9aXMnETqm/rQE7LYMCSQ+7OgNIspQp2qPpRmFu8w
a8w2bxQNBBoRQFH7S4P6xeQJk0mYZKFJ6O5Inr/IxhTdu41ub96p+IU52Tu0u7HnA89tXkNq/gmd
/xwBBh72qfREj5As7e3NJ+tvdbrxKJYtJXXFwz+pUWybDbJQoMFCc1sgW1YNgqW4vcPq3mh8g5vG
t2iQmUBlircHqKIVl33J2ZNi4IvEd8lInkQyPVbmHCuLp2HQlraZ3hYdufNI9hiFqvsZrnL2+vFS
YKIE9DwGrt8FORsfznqPNbMN3hIFUd6ziEQl1DiQYQQacL2JkxkRByfkGSS1XeVyccWA83vKn5xs
WFMruRr4FYgP7D1jyPd+DpMtEEHKSUQt0juMfd60wPLNrchOlOoJgdF7fZKpSKyIvBcZ0r4VshOa
uL8tfpkrXk3zlLzjGocFEwTSfAJx+5UEgt/ylj3KROu+AXG3PDV2Gho3iKJDI4lezd39ItAPkjH9
vTf6OzwGt9TWlP8htDJQHqfDKtLfrPb1z3RZS+H42rgCLK+RPhOi9z9DSzEFoo/0UDRaALO9P9io
u9vBXwGFKrGiYK3fakICHLyTPKJJpblCxX4gEMyggm/FZfsu6AocfiQS8ei6D4rAwVH0N2fXuIk+
RCJ60c+BCrP13nSK9RK79za7dYtQ9mTmNFLVXHYh2ZMsJy/9HjzmywsT4Mvdfi6iutmBGV+PJxzx
/F8Qb5wVTVQ0c0vYlPjNbxKt6xsxthfYYLa3pJ4Bcm/UWrAugwOd1RqgNmxhs9jBOo8C+YjbfY0+
hdikQZ1e9btftUlS/JVWakFnA3jo6HDQQOyCbvCjOezpfNyv7BqRVMsYbytx9djT9sa1N689lZ3F
l1jyz4Jy3K4I5UUHzCpibrumI+rd70YKbjxR51H93vpOBnwb5G6Gb1UlFAa+iFXv/C0+HSVCnzYg
7+E7kms0s+fPsx0sAhX80pAL0M0WHIuRIG+vCPfWnH9R3rXA+RFfGghxiCSkAPT0UEmK1XkJD0Sh
lkJHga1EAsVvukZCg5Ev+Q6DflJ2sMoKQnMkI66CObUjwA/LZ2hby1AxtxhdNvltw/VZa8pJ2RkT
zBhiG3DrFgD7LbT89a7LasQxmInX1/JeUXE4di2b0oWrzioD4IoTpmYKk5vMLidNE/lUkpdAViEV
JS9HiKLZ43neO/Wxj7zyV21BqyoRdxfwGkgU3A89xLx9mlg0m6oNCBGV9kp8Fgvd94ge2dlpcU86
diA/HcvecdjqcGbMTUAvyzr1EtYgalqSLb6OIIeWlEwlQhEV7XaR7Anx7nCNVsEmSd7eNNoltFzh
0VCN1gVfxEbtSgNI6ci+umBwi1aAQ00gutL71a5wesZclMzzpOfH5KFlN4juorkXyx+rbhnkkobC
2Ea5YqeN6XTvdnpa8FQmAuus1DdLMYGia6JfoOc4dnN/keDabT2W/aXDijhOoBuP0/KJibkMI7hc
5YpH1M3FPIcxGkjt+8cXxiQihGcPDMImueJvVxoAse7hqumEGqOT9X2Bcm24UqFZThl0R7mzAqji
lrfUfDGPHR/upPiiXGqpO/kAIzo3oI93ZWymhNy13iiPGgCZTPdnJ2XCPTDW5bzlTV0TtRZAVFZb
jdpcFmNb3vJs7FIFfQBWUHnSQrfebsXdQVXF42yMVU7vNuf2ZBnW1eOuj3VHZ8nQa3gBHIAaIIS6
DxRsDijXkh6RUQb5Li3UpSD9d7tflDwFqsQjdpFUw3XpTq9XFcOhSsYbgXJ++tEWAiJy0aO+nz2c
JwTsJAzzYGfGpZV8QOM1Hxdoatk29ixZL/iKNoxPnR8QzAwUadWRlqGT5RYsHLn7I/D4n1QYI6vM
VJ9Ftb7eFAoNzWGXbIwGbF2TqGrFf75Zk7PtMEj/uh0TIeWQQhghhxhZZOui88ScJpe2VCB75cEu
Skm51rAcVP5CW/OsneLSli5G+5G7ASoIP84yQa9WCj6juROzDKkbeqgcj0KgyDN9+UySa9Rj+JQE
M6+xp3GqM2imNLB3stGmqQgT8YPriO6teydbYKdIqIPExIbReHgnd4pbqsu1psi3zl8jQpslyaZL
C+UhfPRrextdoU0Qb6Ws0rWTkgxBcmdnzxRtKWFAe2Oo00J5DpDIjnl+o6PlQGF5hojeDwboPdlj
E7oM9+U6uGtFn5MQLn9gg6i1M65s+vh+r9xuHRAM6R0nXlPaggkWvHqqjH5Gl1+nv5nyazzbuv4G
5XZW1Uufdc2NLRs/HV5s3YEoRGGazqj3xqB5+BR1JicMW1xSuZvzuc+KOrPhZozOt/QQuFGqLgJ9
SBxE2xDqrbY4W5jL1F/Rb7yVGPqKuPMahHv5sU2pUFTWazmX73DzZpERcWGpNmg1Dcj0zHJTgA8I
2YkWqrhQIOw81mEfifKVhCszYvba4oVTcTSC8w6DYP+b2BmNnyuDP3MWT8ZrjpXyNPSRBkA+wAEs
fGlaK4bxdOr+dUKTraM5B3cetLCsNwHiWKFySXyAGpwe+PqEmzzNGJFKWjxF1EKNPsEqLU4liUIt
QIExlzQPa4f9k9GiWf803y/mGTjXzWIh6m8Jbpa2yW/Akz8ABxBrk21FAEVop+DScXV+leofAV8z
cL0tzM4mb78s+ZmrhoiAIPuFcZyJZZtHqegLES7apLVXFdCGirKKWiSU2MJrljqLdXv6LeUG5zZK
ReN8yWaj8DE16ta8YN3zXqIV9XiJ3+mjwBftxUvRHKCQxXrJs0KBV2OZtzZLHfjCGoV+nvjXUDoc
i6DBFnyJrN/fCxvnTBxbv3OLNJDy+9K5wwCIcpC1gqBmfjuu5Qi+kk//34sBdAyiNbKkplMB6O2q
8QuFsCb+X5HnHJqfpU/9x/UCxjxvPa4DP/Dz+E2JfiKoyxtF6HIXuJKRdFJBr6jZ1tv2mFT71h3r
ZQVssw7iqpU6Bl9G9YJyN4rEC0zl2L2HcjylCMDzckqXaE8f7wIdDUy0pKmOpzqq14IlsRgGrDMh
h8v+H/wNJCwV6p5BNmyj1Hp3wEvy3C+RHzgmIyvpwf0bf02xaXHx3WkThaSXbSO3aaqaCbChCUAN
qlAGHH/ZSfpncbbOfJK60lZLdEnlEM7Jc1afDCDxPdrqfvMmxRNKgDP3udgR/z9FB3d2XaAJ0i0g
DLkqfHN5F4KXpMjNS97Qod8NeYNBBEhNszEYK9XGh6I7i3o705JsQTXWqVWja82QYx7FCDGoms0G
KC52Ak3yfmE9nVtNEYWG9Ly8AhjIhgVs9VlGe+OQRQbjt9ugEvaMzIZ16V/cb/NYeMG6TmRstcLt
MMb2qWW/uIo/snXo2iP1aLKDtRbXLyGtURp742ibRNBxvjQt6pa0nNM6KL4XwShmB/v6zzrRx9hB
xm/WlkTS0RiTvMze4phnZGfJ2fU2rbaTxD1Kk5IjCAFB6xqTbo1RV0uzk295yUPXAuzCAekcNdDx
orena79ApWDOg+ZVFmT8Xs+70hZV562ZqzdAAI5X2BlEHVubVSySpzToYhH2NZJsRsWLIYXMdqbJ
f+Uhh7VKxWqThk0ByN8yQVlaiauJku6G4y2ge+d6O6KIA1TlRE/uzkKxx6HiqABBYGzJf+Cl61Bq
cTxF/eicZREAxgidbdROU7qRnlmytt4Ii9+15PqyOItx6RB/s3QC3adF7VWCA/lR69e4opB9Z4D2
l08MMkftr+H8lKI9bQfAbPKmSCbTVbcZRwwsLytDdQlknV6QdbXFoFgV+UdWalGCSJjxszc7SCZ3
FveuL82pcOQxbLdGdFGTrvj1hp7x0MGDf0rxCwh6BcYIx5x0DlS6iV92O+2jSWvTQCIuvYrmWciv
fNFkzNl8x6fknA4JU/QMVk2EkT8WEtnfx1p88Fv0pnfzn8GSFlW/Dz9XmAvb8q8NpbdkQDOMxe+F
nq5WGCguo1N7K1CdEO+88bRevIQ9OMbaakSUerb1ZVoUnfdoWEz8BcsKTCxclkFfZqJn3n8FAyL6
mX95LEYKZKkjlYDQq55xrxg/N0gEhQIRy+yzK91celd4p5mnKtpP47sIKWTtiTcBZFi3R+BSFd6s
cdRjUMzIwe7eef5uRJcmKVA6lnVyFBgG+y+pBo1WOc5R/UTHjId4z/lFTdf7ARohYO/bqsJXERH0
PxK/AUi8kXbmvdcZHfTjeJMJfMk8oYNKxPvaoZXHkQZkKAG0DG18ng4wwwtwv6olFSArGDPwZo31
ytpEcZnaEQuGNeonhjh/3Xp90eQsOH1asPurWc5n07Pb0XVFiEL+KWD1YMQt416E8W71tyRCMC9Q
YpV66779KiqmrUbGDN4G6DQn1TWjH1CyN/mPz8gM2sc0qWXYTCMHK82zRBh8Ro6oXLanFzhPgNSX
YK10y4Mk/UsU8um39R/qLDv5lLkGiAxjjs4pN3PEhmhK05EY6uG+S7hGK1F6v5adXUNdHY3vDYjU
HwdbFHWC3YUULdaDhbTeceYXDPsoUZ/4TvRa0PUJpMPxfARMIGogxlr2J1vbQktqxzCNBv/JErJf
mSqIKQPFzmyRsNY7JejVL0tdRw1W0UwTLNnp/3saAH8UKlB3gKJXaNFiyutN//x8ExKRampJMNbP
roTdevhfQXr/+DFDN4eakr/95eIh91aWdyfKyo1kA+2bXQDsUx+BCHIRJ70Y5Fjko5MmwgYo0jnW
7iG4XUE+ES7mQRJbzjtkP4MaC5de8H3ubulPttqa8KeUVubAJo73toJsI5KWVL1RtN2q0czzLTRb
qJqOlRlH0N1oP4c2YonLQr7x0RPAMQrtWEDhHGh4kepJvyNEA/SocVP4DSLwS1u5iU6eRjLZg+L3
k23HnC4olqVhcp9xvkaavcvwrB1mTizl+DPG8Vqh979IQ/HWl/fUEsu2dSHHZcr85VqBUBkveVYp
hmoCg4CwRy9sVZdr7kk1XI+XF0IPz/Ro2IFqn6rBxod+6z5acUVzPKKgR5xxnvuYoEwMfMgh/RCy
XmM0OgbOM38bwPtNt4MDIuXIMdwBqdZoo+KbxrfG3yjvuhYsYlTxhhERAXSjai7oe/w+qoh6FX2N
xRsSXOgW8LJb32XMEv2qZLtbEpmJ+4GW0fRQTxmgOdlgMlgOoTFJbyt6f3PdhigRvGRU4OxmKcS0
ZnH1GpiyEYvl9VuzAoVXVfz/8i9LaPUlmOI0ZRmA1Nuu6dh5tE9eydmYVBNcwXDgYB8csuxUV7Qb
BoXChEc0pTG6umE+kGBmfxvyTENy0Z2/Id3ecCDwixC1jIBLaXTtZ1+4EOBTKhjrC+UNa1TEJLil
vTmJhU49CeigM6m3v4jIlVHrTK56QFjaHS9XuowI5XWgq3Nw05/c2HUkMedBSPtuB//yu67x+Eva
n8Vx/sIjti/mRAYFcgFG5x8RNmPTC6k5lKIY892nPEoTWQanD/SkkXruc7HHlttuUFArnyC+BVs5
hzYheLpq7Y6Pt0hmdR+vaIHeFJNqu3sCqxgeQrxMJwYymsCm5yPxy70TcalvByrZP8RGdCXIV88N
XpPjRQPWZvvSm/nndS/2aKIqDT4X/tv4TlhpqyV4kP5mx+FBP3afI60e/woxnO62J9YU5jOy4RQQ
i42Iyv1yi+BRZ0kF9qaZctemDkOWkqG+ZfUZIYx+GbbYjOryX6AlunXlvXag/ELkClpNM8YQsOoy
DP7xqTJ5SgZfLDFveaoSrE3wSE8Ttj80fQz74itdywAjjZ6nJHPsJa1ZYN+7tvyRGP+HDhX1syNg
c9PATQAtBeaDMMRB5GQ0s/li1mIfYNKB9ee1mO25PF1Gnv5h3Zu8cbk/yTtLwxHjqqoXhN2esJc/
elgGmHqrpjUw5YpK3XVMdqxqzEHVUoxL6dhlVY5bei20rEv/GCkOaQySk/eLMs2HdfoXM2s0wVg5
3WESZe651LfZvLDk1nXXNATzp/bzbzdUo5tA0U2wfARl72KrX6gGgKSMii8cKSIXlj0izfZNadjj
t/vqyVBmUmjFK4LUoUUDkUm2F9WVeRcSM4Q3bDPxJgcJF/5JkgutvanHP/7mGz8snkO4LG67vYyZ
WrwglM+jGRqo5Cp/W/Gf8bVt3wHdjYM5gx22ERCtpIdfIN55FziQq1P1CfYG8kBWW1sbX2gYcFHu
U0/4/PFCohDMKG6K8pHNQup3/3sqTSISgqZ8jUTL+jTCbhyJ6P01Vc/RflfgzAt9B6XvTIviNPsU
R6SLlH2L5Skq5wqMOP8e6wdr19ZSq/niDBKI/BI/zM5BK+0aIOkXiB/IvxTQiw+ajJLH5SXwXQLP
Uy7FoFCH+vUJY1D7ANjyDSAlsyUxNaCJNledx0MRpS98YKxelKI5XB6dYfLKXhPj39Zjfmc6JHmh
j7oOqjTZFNpEeiFHNILHIDTaLbH7/NVtCkKtRhSR0HGGk6Pii0ujwD7ZvOk7DU45GqzX0O1pM6ah
h/ovg8DA6/P7N9AJVnthGKZs4o50ONTBK3aAj1TdEvmajb1GpnVUoUMSQOv3QjCbfS7WMB+Wa9Oy
eZ3i9ZtZsX25QoTh4Zy971mxH8dBG7YPBMNvyWX93yWedmtnHxa6slO3gaWKDAMg7PmbuPKXooLs
QulMFy2uXX5ufBiofYCF+CWmn3ceBVIqPcArZllP0ixyjSvX0cdTmWisgIXSISyJxAeHWNlRK3m7
Y3zT6rA7xmT+hdvl5nKhn3m4hoavReD0HNWP3DzXtw1jkWjqkayAx+VNTLi+mh+AiuO9C2V8oSxr
6PNFyjLB0U1D5QGUZN98t0o3kLuvI7G1RaFA9XicG2ULTD9E7mN2tCDihwgDg0xjVxrqp1uAPWpv
wUvtj5JSKTiMAu5PKPJTkDaDzS0cP3igPk0vBbCo2b4dAuwdiQ3GEd0bN9wqV5UDEtx6XUFwJSs9
Z/IxlE8xuP5sWNxO7YTbQY6nEEvkGH3dr7o74V9DM2Lj6UlMsNtrJq+rBqLQZKQnc25ApU8wPeEP
apO+DvNb5a50iqDAgxEk7GFRisbLtaW17w8crKJI7WyHb6ikS52KfM5Lk84xWB+4wydSNwRxDwoR
vaZ1oDX3A7DEo4hMVH/sW7v7xyfP4fSS35SFx4Vx+/MuwSHtT+Lcq3rqX3ZHbv/+wHhwDnK8rSPF
brSpYdmqjTOaKmfEG6cIEg2C3x0M2zdz1pd8JUiMEXairbuW+/mIwf8/28xja8y5nAs1gRsjuQw7
vzXGIbUVd4q/ndIwRU8OA0fAnlKdYW9huL7gvSK/s83sbIyuaH7O/7FIKmoOAhJWNntLabk3GHbU
M0bUtZBYrE8wbYnE3HXRfEy72pswoPRfFWt1n143ewRthMvIlfZBFy/9DnguwQVE57eC7zKctOTA
VSVEg7b+Dg4Mab0MXIpqyHsWNfBscyhz3yyivZ3b6f1wMg+0wszHd5ijCPEH1YViCG7mlb71m+Tp
+iHgoVHZym+Qd4J1XoLOOl8oMGjoYRi6fIILau31ONPiSLymb99iVb2oK1OOzkcJnHivkB+G0hpv
5QUTp5g4390f+wTjnPVb1B65R677hnF8MKJpwAnChjAsok7gQ1BFat3u+AlxnWPfXuVF49AppZlO
bPKV3dLA2sOW2jN5x3MlUP2JskFyzqEY95smWMn9nNiB7VqnKaPBD+Kp2YQpGrKd1tzaVx3tWBZl
nEGZ0KQGaAxdFPd0nHKtlW96CJf6y2zG6+5oEOtYMlpbppd8smJaPkYrIKsLYysvddaXYTWtVDrD
sCWwwUgssYOCFFTLKmwFVgzMn2itywG1TivVbo8QFlwiN93mRv8ciegMTPMHhJcoJmWJjbZIajx0
KZQgVKq5bb9ZXzsRtK4+R21PBn6uvzn0rSrYDoEWpa4dCVpLVV5lFmprfEooGjbHTPgTBtm0UiLF
4p9WQNSxwEvd7w/KDQMNOMnbU5jFFGpRiDU7foKJc2fxjOCp8xOQzJznD+owIFOP42KxBAMWCuss
XcFhbeiqGPrWOUlpVNRdDC9oxgEmtxuyZPYviJE4n/q/VDCSE4tSQviLEfNktGkr4UOD/TaWkaF6
Ktwo+ep3q8FeXw8slo9bth0udUC/G2JMpUmaUOmT3qmIQhKtVdBs8NDYrcgZDyEXj/NInqbj0jrs
SginTFvf3Z9E8XjOwBCM4LwpqklQVLMJq6mRKqp5xYkp4UoQ9NPBVQhQKfHP5o3N8TXWmlwPfR87
wIKbChAinTqpxZYe37+KmvKdI+E42XEyxavzzfDVvz3ni49DbQoauI+tXq3c6SoNmZo2RDUD6vyr
lU2IV1rbYh7bQRQ9tEat87txs/ouXsEDnC5cHNtlGv7t9BsTH4nsO6HVMSvu544wEYbyrrG2Lh6+
W98CkuHYMCtuh7rPhPBzxkdfz5vJrhUPzaRBmfyP0nHvTxZy54aMAn/IsXlweR3izC9Q06bTMabC
GzphWIHgqHnj6KJ9uV8yHDIAVtnkG/S78qlmQNZsPulm7zK0VMvjnlaORVsoePNZFQyXmvTPadPe
gEfV+hsZEGx8QMbh3n0hPnRqdlHHHJuxoCjCQfKJUA+sUVHpS5QbkLFKvgujHyeltOmNC5wQtVaQ
7bb/2FXXbajdCnEpG/+6/vbpqshg7S+zu2tGSG4FfdPc0l4SAHvoShnYpqc/oKrEc5NF1hKm+oBc
mr6XvQQtKboSBMEEAF93VijHsWhmGmdoRi7RLAUBDGjD53jvj+Wu4es5XWiiJUKx/UShRYYkMKyV
QqM804ED1IPHvHqIuGsYNBMk39ZJZuZoaRHHO3gCpgKqv6KGSStAV3WmgyfddtEDex4XYtApeXzg
wMnfi2kmupcduRBlqKmY2R+nH6rKGScXrubtvXZaTIsjT9aNbMY08Z/Oiyg5nF2ytbb0DISmt+Ux
L+tfiJAYndSD7aA7SsZprEgxUdHTEMlm0Um/K0zHaDzNS628V4TcuTbEfW7RKlt97ktlvFc25wvh
GHNkgD6VaBzGVBsG6ZZx34/DaI+z3pDovD2v83Q52AHe0c5g02DeUaP8BxgKfcjkfkF/YaQBUuTQ
4hH3Mo9ZQ4ZkX0AuhOfYb528oIaxC7vBwF0e+wV8tQgpXDGQStNMIiiBeNVCDinAj8MvtrgHkcG2
mR1ZiiVik1OHJWGYaVh6WRfsb9AMSYIdvYUexFNsf3KNW0iKRQfpQbzw5RFWVgtuWEZx3vrANCoX
sUbJll71r0FfJM1YKeOX9A2T6olkRKdNLAGR9Mig6hBjLTFlk3r97edDsHTCd0PTqcfcSvXYXoQo
15JPn6AS3PbiNvbGuj8CVe6BfXzBweP+0Zsh2hNt7izfUBRreeLj8BJ+jDB6KUppgKkGyWqS+Imj
fUJbdI3uJYDLupMrBxFgIcrPmJXjnK2+tOAk6xyQkPddUxou9RZkipY/c2d3iVrLXDKmHfTbTbC+
36pRUrgr5DwSSC7TzsjMZhbxtjwh7mwhNSUzy9m8DZ3Fa4bLRyK2qiKcUyEz+vYGVIZk2mjSFfVk
QF5191LdHH2spVPvuqqXNqrRroWDhVBZ0mlMo8BwQ08pM+9JLc6NEpNyEoqC66srA2I4CgPe5iEJ
1n1K95U7YI1XFSOk5xU/rWKw4a15ZXQYksSiuGzMiwnTHB2upBEGjm4d1rWZNpPlX2RPqtJwC1mn
uhK52ltkDpZ2ct0rKvR6bvPfALgATKyG1kXXYD4tIwlCiSLX2dTzP+UUXKNFqMQhlJIN2ya7uAFS
NJrg59y/EZuXBynsvsDcyw9JE8D2M2vnmBhRrayk+YeaULpHG2N6ql9At+2Wd3AqWYBCTtuI1y7w
yXOSOYDQS48HWRxfDNcLRO1B3bD3EWv5JTpuqMs5IUfJZZTLWJ1R+8neCNW2gCPttVi1uUaTuxX+
vG/8tkSmrNcR7FbdAzntBY9ZK9plvwx+3CCY8S29VG/X7esHtQT9TTOxyGkhnj11qa5HJ69v2jP4
DObACv5GmFa9n38h11/4WikZFjRX42p0OLwj5a6m0onB3QQgoKeKGXmIjPVhpLSPFsjAIhOW4/a+
fs8QLEFlq/xC77yFyyY2cPSsVcQlOT48YACHzi2IdJAmEjVrxaVWRzlsLxSthwGG1K6leNMGvpGO
u9j9tJ5mLxdY018SeA099/+N5aPwo6AvSH3nxd19dtLCImj7DaW0IXdPg9Grfkcvg50k0P54ewMP
sAD2n7lkcV3W+45IkWQjR+mzljYCuvOS1vmS02lxn9FaRbiYi/FJeejAZSxJrJ8/8RxEqK5mgqa0
ML9DRkqkiDtfA8KHbfF10dR3h5wG37Vuq0lgIhwHBYXeSebp/7aPwj8LRr+5Hv1BXZ4xPlLf+otk
AUgVte4egjYIplemB+jJfDpMMjkTU2ZOqmkNwXCmP5ZW9MFrhaqr7WQFgTnv1Q1eBeErFiwSWRmV
4MxZ8PjWNutps1aMVZkMh+BtOYB1FnuHsJSSWtBswkkpK+m2ugWQs4rWqRaymc/PuI3WUMQ8fC3v
9r05MPfNqaerafRTExgHYljFqWBBh0NHLDAsJZhOEdsx0bsWfAD2a8TSt6N32Wr233n3CrvRw37R
mIFkyBXlgLxlYwnPRReXaD82nCxzO0CxDhlLBmVoH9muvkaTpxONlt1tXizvULtr1u8ps/N/+at7
2KFxJKXoI39++dSS5+RyTU3nPdsxjUQ5ozU2ORYHQNujdkzpHp7JxsUZhNOdxjpc2Mot6irr4T3U
+qnRXjkuH1rQ2rvf8otE5ubeIO96z28555J0PRhT1oJMTeqlTj9HwTxlRujrtUGitn+nLV6+l+/r
N7G+6bgHQ23J3hEEWIC2Rm9hw46evvshKoUZ9bOwdpG/uRDWcruZkcuOSYx3c2AYwJdscOUxfIxI
Og1dUqVDwoyV8CAcFNxyirAsENv9yjF3kQz+fnDC1IEFG+HW9Eno3IhhljCOg4g/ff0Clc5yx879
pzjZUXih/NL7GXmlKDg803F3dhq7TtnWHyk75JfUduLJWvTOof7Sd3p+ifPmrbljRtOPQhutApx1
QSpe+uDsG1E3uw7PjgXugZYYSt3UAMlQe9O8Iloc7sGwF7ct90mYs1ub7RVXuTF3t5cCPMdxO7gJ
hWrJIdRj307vs/iKGzbWnJOU0eA7+p3S2BHBszcqSHS/bj0kxAi/Gm4cFErKg/sGOOlyRpR3Dxds
VyiOovMeMCrN2VEi8uT8BJSCZYx6vp8L9Qr9dkbZOqoIa3ZQ1UyMeORo9wJeqyBQTdsr62NSRdZU
Ik5vPFr6ntNNXBgfav2aD3KxWRPs/Yzpex9ymMSWyEWaZg0EThmScaXoLI+X10cgYILIpTchyhjz
YKTxVNDZtjWE1tQeuLhGXroRfY0C2tllKE2UNeERIWE/um50V9GrxW9rtWTXNvZte4Mw+Net1c1j
KRrnl4Kj51rgzKkuXKmDFf5pI4BFVG1WgKFzVhMZpIoh7/cgza/rq5RO/r0n9x2e2xeb+/X7MHhA
xYVh7Ezxa1lmqHv+6D3OksJP4mBI0TUk5hgpV9o/guQH6ujJgXBTznQ5Mxz2cAbHlPfVI9fc51Ss
uPaPjK85kTmVWL2qmp0uM978pLDP2/LFeWXnfeU07GVklqEEc8cWKW0VbUcgfw+X1k+OzhN92EYZ
N0EQn6MIOwDeM56QE/2yuKqZY8UdSjXJMI3CyeEMO8RqTXBJea/yGuFA2cu9/CsT11LmYtHQi4Z/
VUhUTOwBxINbPiL5K2XCLhpjKikTNneY9QEuXqX8cO5dasUOJyq2lp7uG94NNeLWggqTZNlOwySX
7spbRA/ezyvT3WverkuTeVGcUlP7dhr3iBCzp018Zqi9SRXomFehO37KXod6FwB0EBaFwo5BTKB8
P9RalZiZFCkbtB6/IEJ+9V2fWMl3bNly8iguJArP//gjl6nzORJwkThflgnLWWnUzPJU9Q9mCHDB
waifbpBoxD6XsRaWVVo+jXnU9ZLQKNykiB0Woi1IVYmD7RXMaDZxuA2LUgqMKbk5QQ+IozFTi9PW
yNxy07UE3W8B2Qg+zE2CtHbDOfIGPtPtuhYfBinpb055O3uE5ZapIPMMgzue/T4z5aGVo8ObweCR
9XergIYqXTLBwStuWGAZ6liPBer8oEFNTfskFp4IZWQ391dqFEr+PHfcNj5XBTDU7wZR0U9ngY0F
yCJg9Vxkt1O4cH5aRGldTdsOszWUAXc3GVT0P+PCcIoCQcfwIUDg1K1FrK0vaXSSRRAX4eo/Qibw
6TpNrHXe907r72MWul1E207RPmNi3RHwisFhc5+eo8lAJmzRir3oOzWTcljj74TdjFcwJcwsalx1
Ohf+zgAB739HOuzI5m3L/I/RpX12utytkFGBfZq8OkKPHvzcRHIDQ4jw4VfgRZCGBU4QMPiBvxBk
xeQHD76e2Bm4wHSXAdl+SM3bKdFoZpiYBBRjUsBKPxjWH8/fA5G+sqSSQOR4jbdHNsfTsoV/8B7E
GIbEZcx34xgUhuxU0NlyuBLSCtJWICE4t0PApjapipjOIJPHz/8BtypI73qmekSiE7vixWUyvH7Q
jn/R8R0C4AIF+XMUE9R47LMgcBw1bwUH3MDyA4DFXbOT1tR9PeBlf8sZBPyCeGeaAxantMcbfBtI
6dcprEDjAtl3zjhxM8Q57d0P486jNYg/j81fuAz7yS4qAkFD3nv2UDQjrmTYWQbfsZoJwCfW9EYZ
/B94lSWsdQpamiTA2E/lvbxFash/WVCWRLkx1HtxNenL+5rbUKqOKnqIR4y0pAALCcB4bb8TED6M
SiDyhivM5D9LoxVgichiDY4SZrhMiUhyDLKgbQwkotIpihMPMZbpBcWiobwak21MMUq3SFu31m3w
Lbc/JAVDC+w6KS09RSXTKl4icl01inLpONPdt3EM7fyb7VRYjDFBAzaA3zlWQaGcCKivwLgM/ZAk
0Y/+HeIcyShd7E4VigU0cafc5Nmwjcz8HcvRYT/AA/K6NpOZGRUkVqb+LYhFp+akml7/nx9uSAhl
rnJEnRQ2trhqUgXGqw8Bp0iWj+RrXLrPrQ58L2ROXct2QKIw2Xtc4MdXC3WenYwe7DaaTtbvYYhJ
scISrJqR7T6tytorsTosVOgondgTSifL55rOHT44/T2ERLeO3YZ9/lIYmmrMcaYf7VttquYCiWbg
UrPX/m1MYfR+waBTLytpmzo05NFiq4DfMEQZwR5j3Wb9LckcGtG2TBdH0Rcw3UMoKEhqpdOFxro+
L1T5JEjOUUqKE1fKLVwMA2GmeMM6x4t3/FOzu+3GVrkBCD3q3qcqyWAXnLI0HIJja6cLBK9CPUVs
ILuPfetl8N65/xQoBQ5VfOn9j4IT3B7ZsPvMr5R9rfazoHF1Dwm61YcG2lBg5cVDwUFoWkoRwDag
I9SIwujlKnp5xJKkj3AE1XxOTdGIwYSHp44FOJ7JUIRgePXtcgIwRo8aZ0ecJLjN44i25JfC3XLA
u4E3IA9WwZt0iFGvxKG9EEOJtIDfLdp+jDXoJ+/zu/UGC59YmhH5GWVf8miRTwMuMF9RuOuaXqGj
SThYhsGos02DSPnyZvGHKB/ZpdIT9dJwMg2SHB07QEnIDzzZN7RYWaXos1NKT6cTCY5Dzmq33XXE
8pMH2FPQMTNA1zgSlq63HBfsZXGImZEKo0akXzpj+h5yHyJvLE8idclcIhrxAATmUM50Q46UL5W4
U1QFuu1GN4/OoNB12zravnfYUSpyDAY08rH4VL5EvpfCjJFFZj+Wy2G4/S+Gj0VFBTrsHdK6Cqhm
oRZuPtTbda1G+VFoLm57w4iObRWvrsSJd7RwTfwCV8ugSozYWb5Gud2Cgr4TNLWzpgqZ14Van6YT
+xk5+7CKVfNfjfEdnlrQsnVxzDmFXsGjlYAM4tBYB4Bo/dJZqK9KjjfjeLWhSdatIrwNLPEmzNkt
1d0eAjcjoG4MlGa/VB9bKGJgIqZKDioJYs7vkJbXCDxtlpnjrQZQiRr9QwKWw2LQhUJ+1Yd5TU7f
IlQdpEY0fQPwS3s2hzVgzDV5/QHHzKl2rJZOdnCwfEcIexEGLg9LRYnA764fGxJDie6TIjjkNMx5
qW33yYLgZ6Rd25xbVANBt7Bz4tueroRD1UZFTKhSTN0P697SIT0r8SwvCIUNs07jfhdJJXyUF9Nk
5/H9q7gQfZnSGoi3yOL1eBg52CxjjITXF79QXFnIeFU2HxN5mhDkHtG8pCrZ+nXAJJ7FBJTjbjQv
kIjsfmq5uNlgstmX+1GdaKjVsMjJowpNWZxTrSyeT+2yngRFafr2AjWzc7I9h5RztPTCDejeaGd9
3ehQ37WsUJZF/ikLCMF8yy6xtyzlCf2hKfUkjRDtfm/GNyplinNM/dzF+OqoI7EYc9r8SuH9sw1e
IoQ2ZhucIEqzcwaYWILomnQGOXVTbxGZPsBEUTGrsUnkc0mX8ivc30uXp+bwJ/ACZp9VE6bsppiJ
nmenj7Y01Avgc2NMRr3yLwScHhnAa0h/95swkRr1jzsUHtxSgEhvogoSaoY3CGvX620oJZYs4Kz5
FVUc1ilkhTlqBDt396ijzlXdwoazG14SCQIiEOnZdhyLiVbxxtKnlsDRTHerkwMQExxJwlXv4PEx
i90TYmGKRdt1mAmsXUrNpUsTu1sfKkrN7CurG7id7/3fQhqIkdcTnzmQonddWcOfN5LQKsGoQkBp
sLVoJ7WEzDh51dl5BxC47ouLzNdqP2mGGHOvz70SyVueLonEUBj4aiPkJYOve4jfVTpyde2ZZZZZ
S0tyFuXOgehXXAteYsiy6A5qTAQVV8okDe4IXL/wsajgDf4KjIp5zAXQjLccU9NCcS3z7hYDnOQJ
Jmnaq+dnNmVn0FsUGqWz5tOZB1Yf6MUHGj/nI1vfsdSvFM313QZapt1pOilh4U3XPfbVYNPyiPGt
8eajaoCDpyHykdKiLXRD2a0gHItRfpIQAv7gZAZWODPFCI6DpQqkn1Z3xS85vKfzoRBk5xos/KTn
mX/8Beh6Yp7k5CQWyvOeH8wWDCbdGkNSuYv/6ih9X1c2SedD0zc4I51NpovKJPBnz6FJv+eCLJsb
xVBaCt6PpHPtk5y68IZ68rfrlBPtGtxGP2BxVPEpCSFUA8Qyf/SuINQr5yB/Uv+UcA3hOco1Lgl9
G9PzcxXd+qYqZQVa/074jHImqbh9cH0dHniIQcfNPRMAeGtskUnjp//6B/JNuz8E6zDtLg1psejU
x5xYm6fLBJyybpCB8tcdJ00fu6ke65rG9tKAMiruyR0LB93khXYplg/rZXaDZCdbKwVZFFomkF5Y
1v3qzPvJV8wrg5/Z4yMpjKIgUSH9bSCoFdwHNvmYFuockOlmcVq9fdVIAU1cSuNPY38OHV2k/oE7
3akaBft99+Iv65/DkSIRuzzFa1DK0QokoChBefOAByPhPpgUedZeNc77YuEtcDJfkpmEpz+zs5wV
T6//M07zb916r5EA4f4KO/pU+p2d7cs3vINh0E89SxWPL8YVePpqFaMavnMzifsQs8Sta4I947jq
wKvPscJ4/dmDOTFdu2gqsBYdloxnF2IqLq/MMw4tJhAOPgKSAqdpgHixByJTg2hfSqCdx6CL7RNs
e9S0Kw5yo0mko7QbAEzxoUjMy4A0ThlDOI94mThLphqa60VZc0FOcWyxA3w0sFQbJ1LB8/B+JXLV
8jXAz4XzFyVTIHsBL4LCfWRzAf2cNxMl0CtNBD23OQpXRhy5DPFNDnbJ8cYO4jaAU5FWnWMiMuzT
G3DgVwa0NlYgEeaGEpdXV4zQDQ1Iz10Vc6CzwzVHkG9PM6DqYjB9UjBDccxhylwX5x7XYD7udd7n
K5ymCaYe5PB5X6co8c7Tv4T9CHc8orh31em70BffjTeO7dcUeJ4SgOEDQ2hBzFLs6R+zlLwBmgEM
9uRreQDNdNiAhc/VomSj/OTYn161fVrXSmFb2OQm6I7Pg0iBMe0kjhL67OXsOF3bG1LqCILVSb+0
QphdISYwRdbk7geDDq3T/BUiISwUytqZbAFXXQ4gg0Emhj0dZ91QMVXm+We43NqaOY8S4wqjxJnz
p1tTE2U9DDyZeoCBNJKscVat2kHUnJkMIRYkG6PrBKjZXWL9lIURnVUi+/Zcvu3yw4v4hYGYKMao
f75Fvi81DC7wXK619K/dRvrXJiVOvYfvHscV0vn9PXOrlBi/XEbILML9ZChxMXAdcuTlePO4Phxg
U6zdnT/Bdbccw9wPXWMmSN8vEeACiH0F9fjuVMSnqWMlo8BvkRmKQAu7Go1wnigD4mPmE9LCo7Qy
+UyG8WMuaHQBdEguHU/uxN7an+GebXpNXicE4NBc3XUnJx2W/NUa9mAq39HWFF8mCV3N2DmfJAn1
/uOPg8Bx/fA4pp4m1PALkyYT/Rpblcu6TfXpt7sVInXFzFx9ihEIQzF1DvfjwAfZtOdWPpkChN6Z
IJvMda4Z4sgwHAH5XT2py9CYSSr6ahmf7WDY3frj2O9KcCzAcJhTiMYZzKgAbOqwnwv0ds3QrXO1
fzsO3NU72IBEdBsGowyB9B/oFrUuZ47vgEeHhLzcAfBA4UixGt6WzwVfx/PKuAS4smvJk/QQD17z
ePIaTSl1FQCVu4+FKxP8WbnlW+R47XWWZikZwJO07uQB+20RJouePdAVSEW2lu1VkTDpKcoO8BlL
9aB48YMw8rgMcCz21vdHnOf0W2KJkiZGR3OziKNufZz1NAtaKcZpzM8mttXhlBQpUvD+tfCGFiMC
6sXAZuGT1fVBdXs2nluduA+t31CSnl96WXqibcY0TXG4lynb2Tr/6p3FLF/kUKhbtvDiWWcJCaC+
RxFVbPpwhObqhFtucWiTtCepXqeiBsLwGlLPROtWouZyMphFjTk5yGCxyWJy9l1nKhUljBBhlRju
BHO6z+Tc9gDPQ3PAXMS9872T6dt6jS2G8YmodSnoDznCsVWZNhBFocOfMvhuQLrFH2i1/ok7Kft0
9RG+dtbJpGp2radNPj3DvIpEY9nc7sDrsn5JJg6Q7BjqSg43anXf+fyowe+ln8BIcG0/WTeCAsUP
deivVxQc56OtkKsAoSw+GVXMqMq/LRpsjyUSx/7FYOv3sxSwzsfvvnjoRt5hg6jT8hUGiFzGmngt
7B/6IfiDqw8+UKQ+gH2pHoKe+mUhIz+M7kG3OyHTokKd3sp/9Nz2/hfmyH2qPfQJR3MrpHwQl//4
OV/13wIUf57TB/qxiRXCNaUMlWb0LYLNsgwMX9Zh5T2mEVdrrxj3dqMniL8tf5UhF+dpNhi/G6oO
lbOMKPiifRuEEFSsxnapOYt/M3Z18YmVrCyIAYV7NNpc1izvST/UiLDWHELsFf0wzq/cdVPUCX2W
2LKdk0nyfwp1YCecvdTmSFw2rJhSjn/COve1D+GWQDWIztAzAF1YISX0wJAizqPK0hrVOWtaHB7J
/i/C3NhHv8//pW/Fp4Z4JiDB3LCbfLKwH/XHXqENwDDMPBL56Nc/X1EnFmqYiESwb2grt6eBTijD
Lxfy6iZLTFQZnIqQGUcNIr7zN6C+MmDJlI5V+iP9RKEAKuwjbGcHso8Eo/xyuTwc+RSQbJE8R2xb
HWaMD3RqWdQMb3L3ugcWUDwo5vOiwQvuDnigLCJ/0/6YiMmDoOpiQFR9r+bP81utA4UiQAQmR32f
9TCiKhrwAuBMHPLTYuGcy77SUakhEfYG/y3sopvXUavb+3uoEpqpPt/2YzEJobtviPHDXVdFmMea
SSChHnNBn9Ms9Aav1Qb8xL0XCNfM3auiDiKMZoKq8R9nOarCz3yjysBUO+WLyiYEKQ8M+AAeEUK7
EVMGrqz4SLNtc6a2AYDX85v2dex+oy5oNrEfJ6fHtKb0fM8D5CaCmxQcpIeFXy4cROHnOjpxByRj
8qtjGZLba0q+kuG4p3urLtRZUcejwEqSJAKBVk07ntS4APSyBfe84DYzLdgXIcjSPhWw+rANxx0y
VL/Ecx221PXJJXO4pwKSgbg3NyKDWGWYDuHmYm+Hq3GEtCi7fBiwzW+GbNtheGvGe5dbMLnRoyXS
1YYKpKkqgpPGU/d6Q1tmFFHoiMaN2lvFWlSeo80E63bqKu1tP89xoqFeTLgPIl3q0s+4pFRvR7VM
Z3xhLPPoRYVjVSJwziqj2K4OhMnzWTSvQgitxdiBW7VvZxMfhdiEIv+aJpBlrk0Bnc1Wrj7ldBvZ
zjzmeiguACuXr0Fef0e/IvYnA94VQr8uxZJl0ihZULs6LJDVZwdlcKlQx/NHsx8iHs+eyAQPI8uP
Ecl4xnclfe5Kf5ILdvub/DMDpLoZ+zTJrFJdGpZd3PsJHUYIoCmRb9Knz+BNE3EMvyZjHmGQpX5d
YXGr/YRIYfXuwxReuyewB6Rv6E+iPXCdZvSsgj/W15bxJjz6xxfSR10JnY9TycPJ05AjivNzZ6KY
O/a7HrmmvDBSzwk1RZtMRDroV4ghUq/wDDQTWZrCVt0GNi/1AmCK8VH2jU0sUZCeFp3K5KkfgTex
jgy8XD5Iz4CLW/jnyqckVwPIgY1qS4Hsrq5JnTMr19lZ51BldZS1ZQ0QZ0Fkz40X3pE9ItACC8Es
HgUCMVYHbQuLQ6mKF4qfUIlz48kx2I+MP3OStPuwz8b7/xPbSrGEkNeo8p4S5jpjPa8yNrsI//t0
Dboo48+jO6nFkTQKqnvXm7NRCDutBvnIPJLrN75faMUr7Nrj4s9Ga7XfSWe9RyrgmB7CJ5HN/YZE
5o+oTThEFZYx51MadOPo8FMJp85QKpt1VdpphsdglnKI6ulyr+C3Qxq0qde1s7Eqn7vYRwfY+dr+
mS2iaVefviNnkde1WN3ioasIC9KU2Ao3wPmywgSvHGKWlvsdDDcP5Fl0nS8KJG5CQIo1Unz4uHLi
T6o155GHPGAWNOiiDKoSERLbCa5bjcV+XSEIGVOhzTvqMcxTTJihc8um7WEAMjZOfoRa/vNJLK5H
hwp5901wu/3svQVDNmHkaNGwwdS6ddqhCVUJ5ef3BrHYjpP27uz5rZoiHqUXvSC7Tfi9W04SXInH
hWvXClLO2Rj7LsCX0MY7U8kD/SKR7jkg/FiefvmXU7ZI8ljl14uMddjn1Naan7CvHq80RnwsMK59
kVoVAR+nS+LKvYuYcZC4cvBW52ShzoihTo8sxztZAIY514ff8+62QT+dD6bk+suj0nEj5twSlDbG
SDUkBGPTdPpBQ4irsrn01s5YSsolRh6yNQSsrj5nqfndcxkebNUp6Iq+0sVt/UjjP49rxESuGnCR
OngQINxitt39h6V9T+U01nh8QjZaOFVn6sWpiPQngXFLQ30XkMSPrx2ZQVJaxRTcqaX4E+IdXus5
sVr/35LrQo3w+33abBhbJFlJTN5fe2K4rxp4KwssRVmj6mTNoTfnihv/Z2BV+XelflfxU+dgnRMl
iCU8IyRNZnOoisQJLoAskbaEwWYaieHeg053wADIrr+0KRZIq4VOwuvglJ+sqNlwELPxu8IddBqH
qX8D0klRVLEv1o/cEuXeRfVuBVQE9yqTeQv5WaoeE0UrbuyC5QgMgY15zdRJV85oxAcegfzQz4zm
9eqTACX05o33m59xIkvYrpVMV5Tpv3LKJxSRBxYB8Ps32g7dyYXCrBZKXWxu9vEcLOj3i0CVtRxw
hBYniSf//F15zd92DBFXVS9BiAjlBxwXQW6L0qIIGkUlFp+JCYxBz333skPmJpZ2Kkmxxuj3snM8
bP4UllJMZxpqWF1hqAZxi6qlrnI/TzANUqaC/UALAZ1/DrpGaFCc/4HhDnOCtPpW+4cbRbojXudg
smMt45snbw+gIgL24fsKIpJrmjZ4fojx6DGkMiP5E+Hq2RNN3iuN428+fX2QpdQIWX2hkwdiCXe/
Ac9Zzr2J0xwZB8EhxHOMSqnZgD8jaUyVkn+9nbA6PovcWfDTzBFnLCtuENJLBYhWQSRnvwTFghka
LykW7OgP52XAJIcCYd3gRsYlppbO/fh92qWcB+iGfAS4/nMjTOErSJ0xuy1qgGkpjSSdz/BU2FRC
Hj5q4EKHk2ivaMGFN2CVP3CDinMOr9m+JO1KFCY0HS41A8QnH/X44oVz9sEnD11tsGJ4bQc+hyQ2
+VuMU9+v+bYoBpSs/JS0BLuwAKCrto6c9XtYnrK/1iVwGPI4ktKqY5ej3hcx5svutsL0UGdJzIXC
kOIqGCy6+MmmnymlXkNtYvIaTh/y4GRk4hXaJOruz8DAEuDTLt0xLzHliAs20NzF4nmmiMx9/sbe
xakz22YQnzxTKdlzlCY8Nf+HZqxk8fZiGSK+JTyPp3UNZUq+TnDBXoOgWvMi1ronGDsDKA6wfeqN
9UzHDG0jItdi+Ip3qGXoYeQe5sbn1mAb4echePACnyDFYVmVqtVN9XSvdRmp4iBv1SuBvV7F9CvB
4wdAt2eVOzQv+nrY9EWrjYzFaEf1aEDJvVXDpQbEGtlihM49YjkHfJxDuJ+Mvhl1wUX9blRzzpKK
49uhg4JjWoeQshGaHTYG9/ODybR8zcxx3K6JAya0WXtCTayxLOLZLBGOUQhRzMbUMcudPvzm8aA8
xIT1Hci03nqioImHso08ytX/d4f0h0ilyxocVyZs8ORljnuj188Y5/xTuHIYu45bJSIwKfRP/Hjn
NnWlVjIKZ2LoKvhKo/TAgCnB7h5KiBRiqPCySozzyH9KisApZUbpV74j1HY+z0zeGrhoDvJoTuqf
O/s46Z6Bfrmef39/8m1N4eFDtlkHoSOV8JCn6VF8dExYebqJ26PQcGsjxmKPHeDDKi/3FHIGo504
OT3MvpY9426/8XMazsxW22Bte7xH/TmsJliu50pAz99I2mM1w27A3fpfp99IMBPWtkRFoFuLisCI
UBljm1DMYmCQ12uOfns1PWP6Z6mUzacX7FT7OksEhhSnrJzAvcPS6Ilw+1Zy4JOhysnCRBKLGM1Q
lt4SQkIjBJwebk9LRmHb+AAMDFXbSWCwpepiPsSeMTx7d7s417YQ0gU6NByhXc+LvsQsiJxA27A7
x9/E/7uW66aq+lYfFThmEAnL/PVay7Br4HhAFHGX2uO5w1hzJEVCghTDqleVSC8WevHwmPtklzYR
Z4bS40kWHzuP4ncPoyzwjZnv0D5VmEkYgvSDsaNTPFBgufSZikRtzs1DrFapSNiVdpJfESxBcI4I
8VBx0elOnI0ZBt9rs2Flduhl6GlR0Tn5LM6ajFRBrRxG881UnJvuQoY2lfRGzDOAPq5K602ehLQR
1D2ltDpsvttst01M3Wy/Xdqh1i3Iv9EvaFnNtNJnPgg6h1W/SKcInY48/1PBsTP1U5wwf1fzON0+
lxLfbihBadA6w9huHg3YJFJkpddTlS8X8PuidLoAobZxSxSn7tMU/bHQKKkgbWBdFKRJWolb9bMu
4TLm+McUZvNlPDtJrbED6C+JlNX60kU2hu8qZq1AnND8EOcd9D22rkxpfZjrB2664NiMHsQBBFM9
Swlo9v083iw0IWWhK/9yx4yI3J8BVx33iNSGTbaa+K9wxkedbzRY+q1mjNbNWbtOFSuL4PpTw9kp
oaXAwzxupFsqmRP0LE0t7H1wGhVTMpmBSJxH1noegPFQLQ0kUtP8RegitEmhPyPu5/jDz3mvJbHs
cN9c5rk+/ZAtwV+FyLKHTdxD23L2idWkKY/6VTNqEsdbe0S4zfilwqFAFLc8KtXuWNVzwLOoKfgF
LP81QR395d6tclQs+1SemKt1XT1Cib6o4wrfydF4BfHAKaEZVTVhmcFVx9+7JlXT3dqp086YYiot
715YnCMqYKp4TS6IjS7PIcH2KbUo8KLOyM8RsAyiJ/RTAYUfSDNVm+Q84SYENrwZ35pQKpjWUdul
1qAb5OXX2KXoMPTotMatJvBIztrUGlYGHxr4SI2IFCQaY1KgWGV/4dm8EbKMmCqkoibArIEaA+rk
pvqQXICtJ9yL102K753cppKAs9hRE2uq3HVix4YQHbUVDt3gaRNRZrNOfjqc8q/T+NrlvSvLtBv4
WyqEyM6fTpNZ2+wv7u33q2xuOpXVXpXeO4OmPyMDDW0FeKpRjOcjrTqCHLWLa5EkXbB1BWl/d3F1
mLMdzDKYvLIE7ZAOETg9nJIdHdgcLvSJwVY55xqTgXaCyc6Qzf5nip/Expx0sRy+ufDCt8Ypkv0P
jDTQGGhgqg2J/H+7Lznmgs9RuqxOtRvg1mF6g3fKLJgGupgrmypenQ34O64093HyPI0xvRwCnOOp
U88a1IgYVYNkPDrSU5Sd3vbddQU08W/noteqOlmnkbeSX0QY3/7ouZpiPOpZ+746WBqd6pXLDzPw
3Z7bXpzSsG3jLwsFpVLA+1DIaDVPB2H8GagnB6mnXw0AVE9LqEaX71ivjKU43MCCneGHZ1Xe34Fh
KZ7b1UZzAkZ1iKbM+CJnDQA6IMklTmXIWP5D08EeeDvNZ1/V0dtlAT+qyyik1nqG38TIcqnhoXwO
osLtmlylwlApKA1SsW7DXs00XUWnr8IlilmfKRoJezM7nXWnNwjLBQHHl4kqA0ORLkiFkPSOFFYo
YZAF9yo0Xd2khRxbF+MBOHgA7Vwy26JzHH7cwj+tmZwkXNQq6IES+2PXzyHzAekT+Vh4RFRB+rV4
kUrqI58xicDWEw2kqtot8wcfDXFaMbS+vWfW6a9a0zuLwU1qUhMVz55Sr+bbxcheEEGWK9p2GWjf
gytxWUzJGwWEQP13Ukx4qG4kUPYE87rnaY9bi6zR2zde2/l05zzYfqCyrJNSCYsOrjlvEbZlire1
gpUwQlxuVVRJnAOrRrWOJyxW8Eprh5CWj3LQ5gfPBb7RF4pIlDuZVkJLeZN4C2qHXlSyh9ouKTId
iHMvMAOT3EA/qvIUII1LdftEnB95xgg80PJ3GptsCHcIc4pSA02rZ5AdN3IP/TGLNTviv7f8RZE8
gKpvdyD+xfXtNbFJf2Ag7gfWgYw7CYTahU0AxZNSsoY6KI2XqWknTnm8ZshYpVSYHFYORNs5eaKV
xnj+ZKam+lKTLbxbpT9rE+rQv41bDpRer+e7zWsaOeV1ky69LvSMSL31l7GqZfk/90Ig0TLC6qml
ws5I2OfhYSLwSv0KGQBTJXx9vg0MFj8oPJpJMk7fhXXfs84cxUdexw9dQvktlX+zila5/xG28tL9
jEt57yiezg/g9i3yBhIXUfTzUROj67bNQfTbim9mpiFRsGuUiHhSUiIoOPPrYx737wmWxA4nCW19
EZZtz+ReBlYIRflxGtgy0cW3/3wImLPVee9V3Ea82pEOt8xxbZE4Z5AJqPXL3R+CixBANMwEi1Tc
/wPjCIZCGVb22BjAtmKkjYBIgiai31Ig9jrgrm4BE2vFfYhLI878ObHKjphtT94da6r+q/U7OGJP
1V12hVFdPs+0M0gz/HkNJxXKMT0DXHqTBPs2bGwVOrgCkQfGDx/ht6+A1bR8JaTQXtS9BpTYOyLg
XySl2lpIw+ZgjiTfHO7XlHUZDQwvyrcxM5YE/xbT5SrmST9ccpm3pZ53pj2A5S1OXuFFQ05X9NT9
eKjDKQIIs6gXQpfqsbOGjpikqJGXgmyAWdNY9YCwLPN6FDoGV7qJ7H5pgSpU8hSjvnE3n4k5d3mb
W9Zcw+j9VJMPOol6NKXxPVHy2WiaaPsgYhN5Xp23BNVt5aeS0G42fG74AICraN57o4xN5tyJ9d6o
fc6285Tm0A53yHtli4tRlk4xHNrCgU+djFKvbUQ97i97PXy1mtKLAp8IH2i2qYnywMbc8gp3SyW1
v2xT3XSUEpLk3AuwjPNWGQ/lUnBG2FOC2BPCGDyL49/Fg3QbytZBdu1SGsY9NzLNAPyJA1gQo/od
BUkPjtEaxtl6qe+tSVphZNkVakFIcKPflL/mtMzMubliS1tlR9D1tJ/E1SHXvbYX50LHyp1/43GV
ZK9aOMHVF7ALEsVdmqXddgWmgZkXzmC+ZYu5AWSsC2nT0tX+uN3NoJVyV14jtM5gIMk2lom3+L6A
9h8rNZt4dvSOyS18kyeLFHG7OdD8mdiCOxpYHkUbbQeQeK/+zQnIExXhVvLolp6G7J/OjOWvNe90
K+/PJWolAULCbE4vTBW9wTBGQdshP185eb5cwTjORHEX0OZnCHB0NtTphwyuKoGELBFrAryob2Kq
S1MfRLcis8zQhYKNRlvBz2cD9Zx/3hderwRGcUfnMNKnQU+DO/oSsscj2aFVC9cB1v1Ran7Nb7vo
t7nOZqHGK0LnvGyX9pb29nbWHQ8p1YaaRZvnoWjZPIJ3qNbfes5hl0Hevfa7+2ZwbveACGLWElMZ
E9euoB6tpT859S3ndZZrDh5fUuuHSOoYEeFsh2YTit9JRt9FnIHtu9Cw+6seAmx/iIP6jviD0843
XfulQ7yL1jsBW7AIuRq6+Qxl/TRLtRH0xtEFB549l47EjQ4hum4HWvjZW3nWIKdaGyNwOdV+jlm+
oUEQhU/4h8AH+Pn7/knNCSB9xjXKKQQqytwVUHtfsIeC8qAjGiuSZDb9M24p6kBs6DFRK7R8D552
L3W3e8Bflaw7930F2KjWo3u9VndwUhYkwoC8nCitcAtA7lzhy7Ed6FQd3p9CF3YcDT06EBAX6XPM
qEmoxOJblzxjpjmUyxYrMMmW2Y2IGNrlpAZaV+rBzaCV6g74gRZ7DUut8s5TW66MLSnbUcJDNinG
Ue2S9cJCsQ5ZfjorK/Xb64MQLZ85UddXm/M1cmTnYBWWSUmzL8LURxmaXUoCYAcLfALutkHWv8XO
OOvE9b1/TWLa6B++iksW/X/RSewq5EOorS9nVSiJG43vJYQEERH2JLQb7UyEinXQxr2h+LLrQqBg
RdrMM1g03RkG2IzwGrSWp5RHrjqReEvT/mgDO1Hc+enfEpyVF2GMkxqMkRyAGQVyN6daNNVKjz5u
+DBJrC4Qjlxp2uHDCcvyjChZndj38c6+qyoDmV28JXfeexwBtd4pHptEdlJKYJZBQbFxB0D+u848
pBUKe/QzJJ3YyuUoWkFTMz0PQFl+yLuXR+KH6Cj4DLhlAxKewJEZErg3dSkVJbI1XYeoDj7s5VI/
k6nfwLoFZbG7MOpwpZy+RYM3+TaxsD4lQ/0scwoLU1k1+Pj2gjAvOv2F6389joGkMnoAaM3Hekal
gBc0kvyZM0pkNM9xMM+P2u7yHtXVP/6JmnwtcqWAGApythpCZ7AK6xB7a44LgFWjsj0zFPngjFOb
iaKZ79fDfcetccadaNYJrvW2nZrYOkZUQmMx5RZ2Cfd1lKZEf42abU1B+uopvZt4lJpiRw+ihxxY
1v+MRqgdtEx3xKKorfVAjITxBzdvR2QeebU1qtdVY7wEv/rcqoc8jjNNsMOJj3M7rgfFbsmldsIs
0tnbdOJdLm0rIL8is316QW6uLgL9smQCaIArTljd6FmomCreXZWd0adY9uVd8GPblYvCmaiVas8X
TJydkQ9k4xM0biRk860xPQLoCeF0o6BD7f0kMPScz+Z4FqI4XKMLRRDRmOgjhW5zpnvgZc3oDZrw
k1zwWkqOsNFg/fRkULQixuU5dFxzmlDrCiY4j/XCClKpOTLZypS5buDG9L9Lcc1liWYM0f9YRgbC
mV1C/1WW4oi9tBeiHyRYy8qkZS4WnY+IYo6rumyrv8j9e82bNGZ+uVD3z9UmN4/8MdAdPpy6zddr
scIDv3i854BA+7EjmxSMYt83D/S9WeYMT8F5YyDepj7RYvVXe/ScSaVew515Ohib2Jplz4zlqsk3
Tsiy+WC35AWXOoyn98bU7/NEfAra0schEWU96T2mNCKbNLutDJbeS4SSyMJ5dqILmbsOvAKpiU1Y
ANrY5K5BHsJLcLgCbPx1zPHJshg3lG9CYU5VBJUUV6V8uBU1RNnSrGM6INfe1iS21+TsmX2zkHoq
2waEAmL7/HoudYse/wvZ/x1yFG3w4YPJcn7STyaZmSe2zXx5UCWONlNogq0WuBy6S3FVUvKL3/Hh
SMSXFouSlsOFDPlIud3EPvci4q0ZfTXa+xVerxjFi1z6bcH4sBT0g1+QAyiHni79P9od0gqOPpxA
OhH9HoGXnvnDbSjawcyoPOYad8vUEQTCGZ5m1FmTloy0L2GBZnjvq8bXYG4iFBloWwf6dFyPToHb
lkVsXRudw4BXbA2dHZ+GhwQr6Q4tiIpiUlKn/mxJ92TkRC1jGePv8DeMkFC6UbZ/uV0xN0RYkE/C
q/AV768/J859M58YbTpSoE66h1xzfsRqx12EWzMct19hrQcJnbmxlNWr+nz8KrQ+Qy7pejvTCEWe
TEMY8hKmLn7hMVgsGSJB2T1ycYagZWTs5dFvVbVg3Rtm6Zg3hLgUKfWE6tIz/UsgwqEO3MwR79lq
t4KZscyN8s6FKD4h6w5MIT7yZALTEOgtubRvxbGE6t1lXyyAFuiPwz8d0YirnAG/lqTyGSp8G/5f
a2Y9emmhFGqOOBP0YPE7q9BMglzhcMdx/mxEU1zm8LxkDigi9ehd4BdZyQmoBe6/gO5J6pK79pZZ
KTq17HY7X3zC/7gEatsMNeyrEvSkIXhfclBWdB0PGnGXoqoUIyB2St1W/WqGcqGfAlrblMR/GvSI
xyq7/qELTo5LJFGDPS8rYOzlwXNtmwT3B9nbb+DI8xJMgyJUSyvrvHyy4YEek53ynJMpbiAvlH6J
lFB+7V/iJ4hwQfh0Vjza53SdQSZCHtrt7S2DAheHbarKn2smwgSG8tWsFHW5JzCX618GL1LQsR8t
Aas/fx5/zPnH0HUyUCy+fUxqOtU6zHXfb82UoYFoghp0U7H8me69CtiyU3bpxy0oZ15UQbNvRTYb
blZ0nBvY9UKxJCKp5KB54If9Hqyepbh4NoA8/1bVHXSSQqBOPt1z1vxryFE8vzi/lCY5Q8QeUz6n
HQS6LuNm7mWp2Sjkzu2ZPgBgtk4PF7rWuEahknUxnOWLkcWStkSPrNFfq2W5wYwrEEQhRlP+k+mH
JNK5OxEqyexng1Oty3RozZBKsD2dxe4Pjj9u1CQfVhtQGmrnPu3rbaksi0EACEW6RQlg3bwAAtsz
0qa6IajO5g1X6j8oo+7sG0plRec7dnOf92gFs0qhtwD/Jda/2BSUzxN1WxvTLLyy31W6DcXKijwM
kfevXbIuew8JFyrPdG/YsAsrv7NCuGGWSvFpIv5+HnOshbkj34IrupghEa548t51L5MVMx7cOS3C
owAnK7eOUeZHy+B+8tSKi/0/2sdst00gs9qyz+RlN0VCFI80cS5nKziM7BKEgzlke5Xww5xPtbwj
8YMaLtaEBSqPxZR7RviMiO2gdUm3BCO6bFgygFLd+zneGY+qbAJyYMUoC1cOSkFcUbLdXdWNyv12
7p10+182zLB6rMSftCmyek09c0G4cWzbrKSLkPvy5TQ9Ijczh85XSLlZMozzYFbzxMlVVUcybxCz
1m3gCHAO0HkOMabwmtmC24WNg1dTboMDNcwKWxwYtXfKC5WL4iZ8dl+F0RP/4tvN69DCTownaoCx
q4/9tOrhS6UOdXergnlbSUByY12BGH/3grTU7Xw0j+P+nfr+6T9UqcXFqaYHNsUFot/6h6eB5lU3
A/9pcb+ia728E4ots5bJ7po7j/GADVXhbBhejVSfFNx4cOIKGT2jjQGaVsxSXGwMdF+a/UC+ud/m
fRVM6aqrV+bjUflGcE1O0XGZak/ruPxcAI57ClGs9P6Z2iBHOBVwdtqpctLNDzAgfvm5SMFHK3Kk
V693Yroo6kiaNuQhb3/i/+geMC72RLcLRtTTitv1yhNf9rNd4V1fh8A/70S1RKAyaTH6j8Y19miU
qiNhJWDH10Vdc4pUP3FmjxhNrW26PkXQLJAJglboJpTcX4G4XdKFmUbUMEk7ihxQR35TZnrfyE+L
pzACSoH/HFCN1wlbnEtKtaqj97XlMVNSgyfHdJRLOobsgipsJ1q6oRoZ4+pSkYXLXU5HE/nQmB+z
yYm9VArnMZPgt3Izk4/KdNuB42M4/CjoBx4k5kYfYPlYXe1r39qVtxpIJ/Jktj4DU42Z2Wk/ueQF
VvvKMFmG/NpR2RdpjWku0wmn5oJl11LS7B0O8mkyX/qhYHFFLDpt+aZR0YukR0KZ1KEkKPBPp9WP
khh8cta9yiG69c3xaM1ZJVIY/csSgH2RS4TOeT/nhB+4u2ILnXJJkG+//MpasMlpUPsBqnm7fVV4
W+vbt7VhsZ5ZI2mLo+DpAr1HdPPydvywYfnLm4dpKM5rHdnAASwTwcf/R6/JVSF42FGZbe2+vdUc
J3zDUNsCMEpP54E9iUsgn2lVjkYTXHYTALesNzz5shUwyWhR6Q4HRCnI/27aCXsa1UfHwrgQvZBs
4xhByYHkxwJ6c0Rf3O6E0y3ECyyz25Psp004ujXeE9ij5Qxk3/1l+L2JRBjq0CEsfN6nIZfkk5tb
esTa/JU4dDRhQb6nXqZTWKljs1KGEP4uPJm5eMZgKUMQ0veyBbdUhC8EtR/qH505NIE6EFFPAtO6
pQF0U2lWz2DG/TvX3WswU6nT9+lGuWO1ylCiJDXwMziLD9sWj3HKtqaddGutN94Wd/5C1V9hoZZO
m20S4U1siyFvr/vQXzCO0yTE2rhXWUhzcJbt34/RrN0RwbHC29Hszp6r5eQWBIEHUYDCOg+DCi2S
wJPpvepF/gpv38w41Q7CbMu5aKMMfG2mlE11TeJBd+YQWX4LMRJHzaBXEL+k5oDHwWSU1am+loF1
CYUp5su1R49RfxTHsglsUQbI90eB4R3Rjbc1W3WtUogNH9l7OTY8e8yLKCygnjZciAigeoeubNdP
/g9MpVvxlaXqpY979R7fufAqYYQFZvgCOaJN3ZF6hJgn6gvxpa2+pjtt9kPMlzhkP5fko2w9na/n
GG+qcj8D+mMNIFosIqEpPmGufSfrgtjEgElV8q2MmfdYB0bueDx8WRUeu80YS/RTbQGQtYeY7uwW
0EPU+yHgFi1ahQy4zItJpbjuYVaHWAV2LENn2kY4KQHbV2aIyvt6CsvzctzPaG8nm8lJl3Xv+zkJ
7ZIOvv8JXZGHb525Ct1E6kD++aTN/84w1ZTmgRdrTlgg/K6OW0p/uq5VzgI3LX6feaSnAonBPJhJ
Mbr+LqF8Jndm4GlZtEvAZcYBwkOk22g+UbNk4M0Gxkq/l6ghDKjvWYrF70bmV23LCzil/cwN6CdI
m14raWeS0rrlt0XgtfC0RymE2X5IoagcEPDJypM/G3+OFnloEYe1T82aZsBGszzkH+C1iGN6GbBL
fBtzcfEmnifYeImvSWhpSzO+V6VnJrrO3XlhmP8J3frErVB3gQXKXD1kv2rxhNSuZ7LDD9MdPcdW
ybCt5MSeqyabkVjAEE9UI+4Rya3+EaIQkbGRKTvcRwSrG8vYCPu3noVerNFC2XYVpHR/ctKzC8r2
Mdc+9nI6hKB26BE7+mjxtBYDgiB388C5Uqjbs+eOdBj3Rmv7wfHh4B83gVc1zEsaELqRvYsjTbzZ
XYyHzRAdlipqaRmMZ5f0P051QvGf9ON33T7vwCetweOXFaFtDpvmuRCuLp7OOvHJHOmsJMahWdbO
b0GBQwv8jOcscbUNqXkM3zEXvyP5OzBEZKMEHdxb0+oSX3oz2wo1OuDid11oFj6FwoQkxaIy8pmu
7SL/wErUlkXQRNJ3OnGu2T7/fKCwZBS4+HiG7I2z3Hebu3X2U2h3GgjdZ6Gf3k50gzrsONYxEgby
1woXrNJgNrW+MbOoSqbLCcQQnWLhNtl41M/z2hznT7eR3lCHzHhsgi2+0GZGTEriiVTAzhH9tXQ1
fPgRyNnNPH68LisAZ4Gu91n8Od10bm+gBIwr4+ZGYgNLxW5zIUsWIC3nZUwL891PmS2mpxCbT00U
fDf36lOnOLisZ47n2LC8fhsnF5KNB1s4Cgpceae8tdTuklLJDzTLrvS0OMGpfYByAhqj7LoyXStO
mKCAGvynG3VVO0wmdpJiiD3ggVs0f6SFtRosRoFAj3vZrehUXCxW3W0tjcRGyYz5DuuzPyTcSo/h
lm2351nXebKoLuvsCkFaXHDB5uDamHFeo6os6ruT+ed1cKy9db4Ur75lp0A2z4Y+O4dSc+HrjpHZ
fzHO3JEdb5DjeQxPlUULt+v7Kr9H5oyMoepob+xsOo6LVOZfroI0ZpW5aJCUupk0Qj74B3KIs8rZ
K0WjQT7kAjM7PJWBM6zFpMl2xZ6mtUHqRWGsBVq1LhfHk0B+fsv/ucAGwbDBosdJ6fcCozSRLWyk
2WxL0tZ5VgtPZIcrXCUoovqVA9ZxXIOZhB1Jwuk3agFzfJGljwQ06Whz+uOzZWH8rGwkJkePq7tD
arJJMu3NQS2Q9CsACPXECqrjrbgDhwS8hunfKUrMhJdUunYyQu/XHrU1OcmfXQtCGN0SE5kGHthr
xiPO9I57g2hAmw6b/xE46ogkRFZe8s9TvU5sG80TmfUFydaG/zDI6Q6ekVv6DpG1eDEQRBDZKnge
Po7bANpp0JKAYQxV5f9rB3TCnshKqs8gsk0mEYoh+iMxpI3AKv1l2GRC5c8Rq0+9bAwF5RV5y8Qt
rLo8XIZJOrCfHDCrdydX7cuuVhXP5/0nTpQ7KKHJls0sdYFQ+/kHmUk8OqSkvzBnAH1PTL/oJzj+
E/bwxHO7sJg7ImJ0JUlYpn6Qgm4mFY3mqVmQ5QiW0WFxXLYZjngbJsCblozvdj0kyAc2amKSV+nc
ttiFqhD/CSOXs3sd4Kf1Tsh6/7addGnoJDvsDhQkz5OrRJI0ViB7r+0EbnHfhWEO6iTP3SwHDEgD
gzl45TuBwXpzithabQurzR1mWxT00AeR6d14vq/OaFKM956RWORUZJbkYg5JWZpvzKA92iT8zh1Q
aVTfoFgNG+jjDmb8uV54vzY17nBrdZ1Nk/XpYi5XNUmU/REBtPVBAsbry9YwFgsQwl2Qj5uvhuF0
iQiNuJELNC4bAv9o9/nti5fJv6R60j0AfhdJrvASOACj/S6hjR2x7fRv8BLP4kVAvdlbz2K0S5X3
90/OTgfawOs8sp+sKTyH5UWksfKEC3EFjelJPgMyRJikZs/Ikv19wi/Pf3/RH5bkwybRzFjgJ3so
wc0E3DO7Eio5N6w0tEetR8Hbdifz95wm8NGFCfEzWGNwTXP9EbhNmg4Dqj/wthWmecUeJugUSTWw
/X9kA9zbSCgupi+BKstHT0poFcTHGOs+3LBcoeOvkfRhnaYPKZT0jDQf0Dil/biG4HNILnevIsuy
k4zUonV8mBNW+QqW+yA2Ciirs8bw+BrrwU/V/HhWoCUm7QR2eg/Voz48v2fMURNsM5rP4SkECLqS
SLSXrZw/josGn2faF/X+vLWetZ0x7EYqPZsbfXSHHEL5HHwarAT93eLh59Wy4Qz+YijfFf5tbJvC
wqfz/8ZkpE74rTxjYxZc3seriO74b1nxU7XnjrRyCgL42QivNe0yZfvhC4s7CUnR1VqbZxGZeDSU
yZruwxykUKhcQJiZNrS0dnoKGlgv+0nF3Zx3z+nVrnwqJ63xwWN/VRDiNp3HTzDZz6ANO1Wgtahs
VW0L9OAziABQHvUr21modWm+clEaxD44IpBeWX4EDphUhNvM4Ujqky+RDl8pKoID5QcSEh4U1T+C
CCTcKx7vCML6gUn3NjRLIpuHdEGUwri035DPWsdd5HhetkSW0jqQOxRKTwLgj8M2ZJD5Fmp5LmlG
f/aZ6fChaxEI1BFNu1PlTCVarnoldnZH2LRPGweJoigD+89wh/ib6YH1LdUi4JJBs9Iu5u/y6kxF
quMujEwuuBGPfgKNoGWjo76HgAWBUNjXh7CPOEsHrW4T4u6YUoykoDEiSZbIHJE7QTnCpPhXdNCF
WjMU0/LqU8T+0DAcvn8CW2DqgGW2Imp1s14GXE/uiVlVW8Z/R06H88b0jJVIpmGG1pa2eSGeh8Yl
UYxL88VO1pPjxen2N8GeZHCQ4cqUxfSWaCGxg3CcARDMwHJBKQMQx5EC06Uqg6Yl/0NLZ6KtKPmZ
5Io8qJrmsck5dmmjrg40b/rWG/GEmDW9D224pOv4w49ymEIdsAN009SIBeKgrA5ip0epCOLY/wyr
B1ALSzKbv26R4CFaaFNU+dvO5Hm9Bg66Oclgg730EbhdSfd5Bfm8LzaXutFtaeosR5/Gb+LjLIVY
r9JWWv+BCvJk3RdnMy2rcAzDfUMoG+GqLmreuAq63SGPk7FK2UILf7erUJyHxJGDFmEMTVvd+voJ
2qYPryOXt+dnCSqRDOcukSJaOXVYHZeyxr5hUUgUZWp8S/bHGRE0Vk/pPfpD9wzx1fY32wEXPzYv
Dn1uIPYeNUdvL7T2QDFfgvwrbJM5pW3acbBFSfY9pQzWpA0AQ13t8FQ66UZrzEL/LNPI93/NgvZC
B68jEceae/YmtCSr0yHFsOuUm57wDXPSaKZU9NLCcvu0Pe/dfCxbPZ7LcDPL5Q+g77SFH2y1boNh
LR9s+zXlKE8rBLD0qcDF0hkMm455HEGVvM0b519Rag3Gf/xg+LjZiF2oZBtFtJoxKq5xoLSp282Z
MHqujG4g/LDoWxueALyvQlDBkzRZ3ivap5BdHl5RIUF14RiKRbIhxZds9EwWKyW7JhF3Xpz+Tcun
z+LlHt/MoVnpVyso6sZM7ck1KDTx4tw7XMWAcEOoxs9FwJTE3ZlKZMN5K5MoQP65tGfPpdxSZfiC
9kviWKM/GbfaRRnImC9XpJWWBJFErsvDRo7n/j/Fm3MpSAdGAJt+LyVKq11Y3vRS7E7klQRv+rw2
PsUmdkFAi49Zce6NjFV5Ren+usSi/bqgXvqWstb4MqCFmkpQ5qBcrQeQOJJmdLrhSkb4rq3uuuqZ
UMRFyJtA5Fqfm/tbO5gsyN7jbk+VVbmY5sZaVEOpZUGqNhKr2C/gxqLU1/ot4/MQk+KZddJ9DDFj
FdGvvdrGCU1zkLug3vsXyhRSI/7qGL4wttH7dFWxk42zGi7h8taBPqYS9R6zDStIn6HoM9L2gxt9
ndOV7ExEkj+yq4tunuoiURksiZCmr4n35Jy6udpRN5PGfUrKZwPrQNAFGC/R+nvxQGBPAtzKsAbN
OOCsTsA0MDP/cu4iYe8m0wcWCZzIuOJdMlcJsn1sYBdOIAGYwvul6HTYRdxAwyqibsGhBmSfPVEk
NBLSjRaIMHQFcZ13+bL3FTOfmaR9nzNmmDwayvSW8dm7sxW3VhuLzUbh4p6y1LBjLCDqaFsQoUgt
2e6wjotUsipbgRgu+aIEGukwy4zE10zYA2oJRXCMaYRz4usmWuiaSpnDMhhL/dah8t7458KwvhfT
YDt5TA/DjPU4lpOrJo553zQw8OkSnDirh8ld+Io5pD8uDcQ5yR4BQkVJKoMAJWHxhqEDi8XnJ7/X
gI+jkEIuGImUJVcNasAE3OjkSZwDQXsrcoU4HEJ3rDs/vcKMy05bMJvWkkCH32xzYsGOA+7+tXeE
43DUlBO6JA+KmLD3R+/lLJTe2QQhOlgaMTNMeuZg03XrQeP5H1ERod3KbRNW9oIzOPiTaeTdhCTq
SCReXR6xdFMSoH1/4q69OovjscT3/b2BkcoYbeEQThBSYqj6EiGmEtUawjHSAq5QDsFS0HOGVU4C
AlCVEmpdClcz6WyuVVwgRqvqXO8J1BlambWrWIoOwKUGeampgPN2Hb7BQj70LCyvbJpqS8+GeWNg
L8sPiH2OEqVXvAaHmKuxPeB+F8LKioYXlM+dfWO41EiN60D02EImDArb7WQ6yaN9GUyhG0Tw1GW9
2taG6qQpGG0Q80LpFGXpPxzU++Sljir5nrJ7DsYLUtoPxBEzSu/HkUcCJU5HRHgPREQOPXnmrFnJ
i8C7R7L/1VzSjWsQ9B6yDIrsVddCCTNkoktz8OexaoKy3zy7ZPkHTzEfkkEt5eWy8G2Iu2i4YVny
CVr1wL9RnTmVdU1ZvYMkpIx25G++Oiu9YyuF35y6kVvR5IhLrQIjRt1s4cTJhEm0Pd2zkRRwyMw8
Tufgo/PW0hQjf2yqaV3qWzB1Y7NibkJTnfoaeTMQd7qQ4te9ArebxPNJwJAKqjE6cYuVK7PPTLCM
1zul++b5sS084PhfsK3DKbX28a4T1EOZuag9pd1J2AARB03IRHjqQVFRdgzerb/Ppio/61nsmRpj
fvIsu/1EQKww7XNLpOoi7ktGm53HMTxsBs67nykWVsK5n1uHNAyUkL8IvCu2mxrD5Js0qun2J95/
XU5Ovpwh3yk7JqRx35wXG8cwTjaPRkJ/xlcxMIRvQoyz7RFwx2MiXzqw+kjwy3sFZvUG3hegjZQV
m25FBLqZ7qobqZiklPMWTgG872OgQz87eN9NC3r9To+szfT+QoPGxcTMmWoKervBQSs9bzfvj3Wx
+XfIKv4GfOT0uNQIiLBa08stFNWVUeaAav5bbFYg0atBBh+biNgW98antpzwaPewHURbMwvff24K
CBMPmzlOWbP/n9d3OcTC922lCvGrpJsFIvfUeR4qTnOhuZt/shMbfCYoCNa2e6ThnJqqtrscmEaU
kia8LVmSaN8CBF/t3uH+JMmL3tK+ogrIW4rVrj3ZtP0QG71piAs9QGRPF45LSilIjjjSvT6FMdPI
IELnixJJdug+2dCxMLqWG2OezoRK4MBCQAKznzo2nJEtYO+2+KckhYbDkAssLRkfN2RNJd4znz8F
JcB8FHE385gcvA/WiH5jsMpRVhnmHbD7pw+3gF3j8ZAFWg5/9sCTM3JFw7qiP4jepvg/+b6tcxai
pEhgcxY9PxOexohz/rgmYUxhS2KiD1+Au6xKhcl6s1J9S2fv45RkTUaZtzwxYEahW4Ul9tGOGWgf
OFdP6AioTWF626ATrC5Uik2W/7ZT/ymLOHnq3WStcqg4kFPHo8feGVV2XHKiivHK6LCRfcRA7AX4
ndFcOBPmmmiB7VFddRr2Ayav0YEUU7GRmuraGzIUcJ1j5JkbV8XnjnFRuV2MFGN/fUsLDRhfBD+8
e94m27g/p6VnW0TyD06aDgCeyaP1L5p6L3UmLqBnahJNiZlvYjSF30uHvosIPwBPVXTHYleX8XSw
bVZgu5yylMO94EbEwM0lJWm82E0UY0zm1GHUniEwiq+vwPB9QrUPaYLzXXPAAP+huKrbbKd+DLq/
fs5k2FACX0unYNoJPstnMKI1/hy3AfLT3Twf9+Zf1369X9eKyJALOHg4dCAljCq7V3qL0ZUvzLUz
XAo8I2/IVxjhcRm9Xr94SJr6oziGC+LuFic+vRkj5+0zKuCldqdjK1rgid8p/u9zu6d7omDlIgK5
r3lMg9Ksu/ucpoYalInvnced0D5Lt4Oi+Rg+Nh9G0FRnzzyeKbXU08KJ5G/oDfr93jO4qmnMfKRn
fQ3jFqpyZhyP0yeI36JcMDAtxj4wd3gTXjktuXGkOTJqsOlUxX7uRYsHqM2sKri6MDyJmH710HDK
4VKm40mwJMwuhj7gSqd+9X0/x4d0z5gIV/YzDGHVxCMyouPu6iUPP04SAAGW+r46Zt9L9gaYaIqu
GtOMOWMys+OhaxBYVpA933P3a71AzdZBcFekO5tEq38USGJN5ivqTRLjB8pdc7ghBCRIhs55hyao
Z903pkxayfE2EkLul87VOoVO6kZa5qIvIXJmrCELg01rgG8IC/rtPuNm930vvdl+JhJC1aEMHvUQ
LZc7GmvVgoQnRdHtaELIWFS0ZUiG66nExIXVnZStHlN3Qw7G3WVdxknpPxc4KoENJSO8oLpQGkXm
caI6fJkx++Wvo08EnLCaClL0aA5GtGs/R7A1hGNYF3fopMzJCJ26I0Stu5jNlnG1hs9shGjyjq4Q
ph5sTw+EUVE1CuGP8Ds/MdNeC5mqNVFfYEQG3sfgtgjt1vgCFDzLVP55smuC8gBRgeT6XKgev3Qg
J/ordmuqnRAiXha4U7eI9HocFmW1JVxCrDmV2pTCQpKPv4nHSVeD2ac17VzuCmNhhz5wpZhRfhX3
LERfBR0EJ9913sPIymg5vhTZMyYCcJ/B8nvlO2M92EXTrhAVuMUQw9bWeKWmXOgS5kaSBA7eLmhj
LuLTj5FMBGgdHD74L1tpMSlRuMv33q5yI+oDBfoEXN7QvroTMJ3kVHz7jjE8uCHEov6p1tevAcPQ
6IWa+4zjpIXiXjXxXDyu893eNDgZCXVcmhYUPOufZw0bNkFAB+crZQP58r1t/CwFZmNbQbHfbRgj
gXaYhVfMe33hptOV3mezHVvFMe+BX5gNOMf/8rCbPukAOHnfqL+hHR1ay+GPViXvaxK3fgLzQIvP
N9VOT8naLzO0fFuPHYZIhX1vOP0bUjeMwAwsfFlZK8XvoowlUZfvZkkINRIRnWuM/CSTqXmSm4kW
1J10eZiVwwhB6f2yOVwrCZkSSPtxab6Y0zgVknVZp18UI74Zc1rO31CH90SbBdyp2toz6nDyef3o
opXC8Q5hEH0QBmkU40vtRr2HnAoi88RhrDjVa9BOwwHoPACejy4BZhKtcFthoZ/FAdlXkXBh39nW
qjUfUyHKOsdilElEDFJ8zMn8UJNnYabqCUqZtOEBPD3ox88M82uG1uagVFu20CpLud3/YvroSCZf
IhzNEr9G+IVEimlGKQwgCGVeXRUPpNGNFPQ/ypYOJ/kHUwdKoVRzqbG+jub8zzc66BmuL/yYLkcw
hXjFlTpC7+9EqMpZATCS2mqAJZBf9fIZ+cgHedb+/tdT4e/wsuyCwt02rE+y2IHw3mEMn43/Lr7I
2lmjUkqWA6ufc0wj4WJjiQrgWCp7RuhBXqe27PEoZuzyINfqkeODKNggbpMyln5uus0i20E2Qe+z
5dgtR3ReMh2WY/hZN1XEG8QxF9wj9AvA0BYUcScA6V9dYxJHzoRx29XzqLNz/K7HqO9uBkFKCtKD
XoOcLEHBM7mvaK4NCU+9rUwTwqEfQpQULd0C8968wB+RuRvHlNnsxcXoQgl8QEjKGGtW8HsSHw3D
LYFeab8Xc2YmQGW8tAQjC4+Sc9PFdBqVAlOoX1R1wkhvMUzLZ/+l9yIemZy8mdjFMZXmXa8ZfM2Z
W3S0vXD6PAhBZxxZExxn/Z5Dsd13NZVjCBp/2dyDpbsuu8Uko+dYG3JSBThQtHlKmDqoNY3Vomap
aTZRYXZ/MqISMMmmqPCOouLPvs2l1l414mgZ7HkdstRmCiwOj2Um4dMH1kUCKOCAdcbEn3Ha2ma5
3XK8O9uoPEvGiyIBI9gowvn/uvWBk4V++y4lpoercUWJJNZNzCfBs/z7ChPy9yLOdIunlr8F4cqS
KSvKGrd4+ClmPMddBdjZHTR46O4DVZ821jfi0XTy27LNahyYe+C3hXRWgJiQAeWPJWaeYsOPhoqe
Rqeft7gmBrKerupv8bqdj1Jiq1d4fFM4Iw/NVfw7k86v7w1ZnJyTBSqC++K4MRR2/edDdtmlloGk
Bj7rW9DS+uZZ8XOMcKgXYRLkc58pTOZQpu1ZVgWshaDjOwMlgO+dB6vFLDFwYr/FgNmlui0O6aEI
3yb5SSFlLy390jGZR+DPuE60cmLxhWvsH/cHtb/WGVDxbVAyPTHx67G6cE/obcVjnseZPzVu8sF1
TmEd9Gna2JS3ZhJMUtdL/PqdxzErDtv9SlmEdYEhcPr+DRNLG19X8nwM5gfvtxlowJZVgjtVtDcb
QmXHP0TDjC0ycUxHhEtPyvgG1dN5L9nXO7Qg05h2fJSizo6BM1B0YKkez2uuhXL4tHqPP+HwWy6H
HmxFhTxzcM7bZWUcRklP7IAbjB5F+eR9yH7aAMBQDP4PtXtc3dlNEg6q2mAO6OLICCtWk/fD8tEL
9yUdRJZIlo3wonhGZN3rca6Nwbk1QfFrb0yjBvtBLU64UplcdkUBUef0XOU/rSrrON4EWngVv/+f
89Dy4jkEvEH2YMWfbxgqQaynfgnbstZ/Nb5PW1yRu94hY1Mi28xwKmZ9/ofJp0WwQhT6mwmBBo+J
AHXquSiHB1oNiVvGVDsH9S0cWtQa9Tl1StuEUOjktiMlDg9ZCtm6BRJqTKBfg1AD/ZCCSgVj4tCG
9jUx1Z0wHE8LvadyDknwyyEIWx2pkEoxxFB9GH8cf+44OiCNpXM8SlwyEUa+AzUbihjCjhlGbzGi
VUj9F6K7Iaa3rTLEZUAkWf7E2NTp681waB3DB6wjLQJDn4D9KtZqGh2C8IJwce2g5p7wiSDubl1N
XJmdG8AOXM75F6kZ8Sr/40bEgD5WDNRe6UEXlhcus52nCwUwrqMn5KgN8fmgFAdiuPJEk3+Fn+qc
hha4LZqeAVf+21qAtuV1tG/qIsRov7R5sA4Tw6Wojm94l7cM5iXnj5nBWg8YGcYY2NwwFpQnrOo6
eDvMIszs730G46f4OVGudha8Hlt88SwhQqZEJpNLzYCEQoK6t2NkRZ16VKBn3vxbTDBAkNO6AiA2
WAxTX0auGTf5is6cZy1XU8woVK7oN8t/vv9SpN4QOl7B+V6r18X623awLtbTuiPCQVgBAM5TZp54
u1sX1scwrOKwQ5hh5HX4FrC9ZsViEULTMKiRh8HJfqSVIoUI8f/dvyacT+PUCNi5ufAz4dUqVTg1
aJJ05Ec2RUczwTSMTD33nCwH5hyKbcobYkv66HYBMOkz4lodbg6nXJ5pA3kUhkg9ej53Ryr8g9MI
H7JqBg6EOqq7HgUahTQF2DhdgCnEtXRfnltgSL4Le+7Z4SWSzlGF6XmjqVdoHYSfCVWHAVaZIuSr
jJEpxtVVU/KCKJRdIUNFuIYMeW0EYhJ8wTGmOjKE5vKAPmWcxEuLtCB1nef6UhAmTB/WLOslz8F0
5cfAjzJ66cX4HO6G0tqtiuLF0m5Mzy1m+CbSkJJuiJ0B3jXD5i5Hfr6KuO11Dmq1oWxvbFRi2I5A
LjvAQ+in+DBAZ8+esBqhxwTyCZnMfwM5DQLK8xmRqu6IuW3M7PaBmzYwEtk/iNzykHvzHUImB5fq
JkmJNNl0KRn0CF8g5dlFfMGXpyXxb03pJVc+/znbaEtB5sA0thmOxAyX80i8GVcbYb95zjqAtsde
+aG56mSNx25JyP362Vk1F1saz/kC9O5wQ3XQGfZcwFnS8tFl/B9ITUF4mQkk126sES+NMO1uztA8
PQTzjHON96RczCPqTwWakxCkhrwNkv5hZLyzl1alUnB5K4XkZW+PsD9xFWQvgLIiZfFg+0Wun5Nn
1qLZfYvXzELZBW5aKEG9CT0AAFrO38Dlq1nI/myRfsYC0M4wniTZVVBKZFpc7x7PNUFS9iednemV
X6SUaAnrL19HVZG3IGL3aFP7pSbuqzfwnKE2HpcB1QEve0P+f7KAiXyGiCtVJ4DK3M2EM85qg3RU
ufKZAleymHhYakwBr2QCtyUIs/KMwfphHiYTnO04Har0vwKflNDdk1sae1/0wvooX0PRB1RMy1Pm
LDayZUjhp2xeC5JWnJQN+Gb/ptVRNIF63L58WsdBvtPCfAOE+ebXwcPmFVRrMUiPCIyu/1G38CEf
D6vqiSaPWTCFNSUr+hBBJ/DFA8CT1VHSdSqvcEH+WYEoWA8OjICSIjHcAzGeHKe++4NHNkOzB6YN
zj6qOZ8nMK0+/51YpX7J/eiDopCJLX5PkUU/WLi+a/1m6OgHSUbI30MMPPyt9ykL2GUJsyv9NKp/
i3MubpjzlgzmKEGsKNht/SCCFE3Bcfq0+F+HSIkS+35AwbDj8kcGNItuoybQOgScFSF4xuh/0hqf
dUo+b4I6+s1EA3mxW1nJDXVWk+FSRDjTVrUGQv6gJXKxGSKokRy/Y3CF01vv+TzpNpHrbFEZaKU1
zJSE/g5xxgwYszVeNgygG+QXFjDbV005Z4wsIWBEZXmnt9OBRgHtbxmJFDGeAO9WxP6ss+lPn9kU
EYx+nhsl/zlUj5HXe6dlJ6KfP0TSzari7ivb0VpmTz06cmUZXlO9VeZrJR28YAmMz/3EI8l3gWmP
vgHU4dSFMoW/iNgNInC05A9S54s8eVuqKuLOhuM3+DoUQq+2f31U9LMHyeDExuQgtPnZeJiByILJ
nHCdWCwk6UzTSBfTMBTLFyB8xQ+JFRtuhMmaE/EfFMg7YO0MIvKjAPn7FNYjDl0kVGR3En14hcOz
wWT2ujoJonaQlnWLjf6/C7XZJmmBacdB9DMO6f5Jyd9bod4GNox7DQ1ALyxYI6rDgLt5bbBg7nlu
wZiE4yb3IKDzbbRn1JRbYuGjwScLNLMXuwgfqfTtPTW18GiUgPpuDMj2RkRAmFDAtEXqdukTEpFz
DyAzK7xcWTX8BF2aAixh5+sjITA/Pl+M/1lhzkolBP59vrXudzP3zjBNtttKIXn89wRVvwmIwGEH
VsDJJSvI0Qw+YfzH6eZruJ9/B6wBuHHaOB+ReLU1tdQPzZLoImufHIyyIaFvtUq6UqAc+oJUDXmR
9umShpHDiAZ7A/pM9EWhInCiXMlUbryvZykVmdbKFLuMwxlLBHZtRPMD3hPY9xAbyuPtmwt3Y5UC
RNi0kRvUQLN630ZCa1h7rcz6z0YcghJjzpvCk1QIwqP043oR2d3STtfj094Va571jm0Ynr3nqIOE
wDn+6SUnBNAE2K4qURQAl2FtEmnF7ANJMHR+MF0K3xwA5q6Q4FkuvnJRNg7gYcXPNxvVd0nB1D1K
Tbf9i+IV16fWwXkQrmD20L2ZLVkpCE0igrGnmCuFPX/NRMIwfYVsLUhT3yYttlgh9pG2w9+Mg8d5
4DmEIhSDr3gQ+lWXpkyLAxB86r4HaHcnBifxYoDKzcTdgNqIHDSLlwGCWkFHg2PmcTniqCgmid5J
SLCwbYHr+RdxBqni81b1VxPQNOxgdeB8ehdRP9GdDDLrv/AmZHzr9hAlUsT+/YcoBCObcd+KakCu
B+Lbiz9AuhXFH9l+inxFZN/yM/24xiNK50tm+M6avv/vzP8E8o9aCgHfLyfaHxCag3v/3V33EmXK
A0CxO7TIMh9L8fZFJfCAZx2GMUVIsF3DDOAKfUTp+DGXoJ8TEciVEK2GRaCRIw22O22RvCazzodX
8PQWWaKzTeTxzehNQxvWhc2Wm+Wf/O8lZPllz4VgoojKMkVLKvaH0BH385jELsBmHn2rZGM0ideK
GBwTuq+tiZilMCvXkGgAKEC5h/Wfq4CsawMDLe3byXM77EXgz0dS20JzyXJy2xNHSImSe8siDv2T
QKuuQ910u4PxiZmnoVwGZXKhCw21UIO4rGFTfSDG9OziRn/Y6YNTHVMPE3oAqas/FUvMQJuO3LdU
xwzwh8lm26aOknrtdayJFc3C2LgUwN3bQNPIlMR8inMGSBCu0UK6/CSz88sn6b6+ru4cNq1ndJZW
A6c3PSzEl1toamYBr5/Npn2b8CO1ogyO9LVbNq+y+goapjsNvxSP9cxpx32vCBDm2ZOmOzIRB3eh
mWH1xnHoKXcXXsAKSYiDB8QbEzugKEfoJQDWcb7ydNbnkZXUDVwbrvSiSkQPsj9UhlljJzaHrUFN
KUsT5tHDvCqFJdjT/+J30V3sGFRbeHX4fIcysoZvfU/xySHBe8obB0iV/Ncmf23BihIYcxzpyUPu
5zULESFiwg5PTozmsBg1wMobJeNVR1/k5jDW8Ei2TNndVM/GBqELjZo1rOfBLBmnLBujis4XLKE5
3Ek+7gSF7zE0jEdDWkAbplXqD8h9tq9B5ybmh8AOzYg0AFMG2qeXf9NEeyLyxQym3i6OYM9cde8K
3HdFZj4xDoVgfjC77+6zeV4Y1g3xyHtBvlulfsNMcd02cklGhi1FUvMzHAUxWMQ8mCLdz55TDd7I
uH2RkmC1MhxQ8aCGyTXyDjVbi+xhUpkwWcUR58yDCQsgbd5xY6dMHKwnF70Y1ky97rteUxYfM3NJ
q3a9AYgFb1KJhJU4UJZXKtNVtrBUl9PdBFIVnjwrqaRpECJcLi6DyIjNONAOsqKGwexlwiEu/OxD
i+U2bgZ/sq528TrIf0hayXuAgcWJKz39NGTf4NyIAemQDL68C4jRXusivc+67HGPSR48oRfUqiZe
THkyvbhBmwED7zjiKrci3HExn2d1TPGumWKeT/IlZ5x/KgzJao+MCL0BVdkmr4APxkJk8mXKbCR1
Ki6XGXLBQh1iirMQK2RhCiGAMA8bPE0BGTkKBUrw7LhMHB8KKw8c3NaKUU9Ew9moJKBH5SNLK+O4
oekayYtO3KoZNVrBlC2qxzspySqYVbkoatlUZTwtUvmVf1tV3aOkbN4gOaQvGeFmPDRHedE1nwG2
Zh5r1aphp/c4mYi2sUQwGrGkrdbxcWjjTuwGd/4yO3howe9NdU8cdeMRermVXmparf7hGRA8Rvyr
L2hiT0WOhnlKrZ8eK10YDiaqzxWCxzN0pc/NHMbie+stqlXEI5YObt8GegPGTyus+6y1m69Hf3k6
lTJaZ2uoMe6Hr+sSkk0RCBiruK6eeqIphVP/bGgTpn/4nvhI2WjM+hyQ5n5FSukB3Abs+R/OGUr3
xDRbsR1zBMGtQAALBA54JFREBCQk7TPHP6fx0pNXnfOUpaNrZ8LD3pWvaGTbWdDBZ3Vvxw142K6A
eoVtggjwdJhlD6oQuJak75x8XFKqLq3sF5HYpRClZ6wKXPR2g2wRknmvZ4l5zvEsOspEL85f7l66
ZRH3v93xIOQA5HXQlcmDTcu5a5b6G8ISAQ5dEv5/lHO7VHNjyv99sKSY1j5u+QpfKnEjq2kra2/G
UaxcSZrR5NfZa33LlPoqP24srircudhYmIDb7wen494bXrYxlxITvrEFZXwqyZa7pPCTsHhzA3HZ
bhdSYR0ymGGuIx5fC4HOPfbl7QMbz9LVz/YILLFzgUeVRF1D9LUmf3zPm0e6kUJ654NWkPm6YH5u
uoOT8u/tMAoPwq7HFgctjLyO+D/ATloyub3D6AOZgfHUW0vVKHfyvQyudAUZDdYzS5Ca6yuSiV1V
QdPy7+z5baIHoeFJDBdrjPd8ZwUvjruf2vEifQqNvjoiabVz+wQp6dljpU9JInUxaGlr07lCE1DN
PnJHwSR2GOyWzUw1hcnO0Z+2QRVqHSYJ0cmehemjf6G2LmVRuaUiGf0tgGHeAUyRw/EL2bWSMnDo
O2pVzskwuNpNwCKGTkFukZ85+B3ZAj0kyueIbGwn+pZqFGJa/9jQmnwM1XIQ8hNGpLXVAcikUmTG
hERK4FZfdFkgk8/j97dmM6BJyUG/WorVuXeoL5NbJcxlKKkdpOI+O8k5OePq+6OTDrfndAJ9vyTX
YeAjOwrUCeJbbFouAoTYhYDsutI7AdhvxTQxieLyVjvJ10sdvCHPeM2xtO7FwfV9hhickkAehPgU
tf4SEGA2cGiK41LGYSU29CM0EvCbYBw2pKIB9bBsEe6If6TVWwGuhf1GBzYTGHl3v1+/NxT/e1UA
HrDmZMguH+kPgVa/F+fYETx7sGIEcOuqXOw9yGoPHzw+1GlKKKbCCmRusTRaNIDuD9himmCpUnAu
k9hoNqJTh+3eQHbPdc3SlHmvMGptKYvpznpJ06MvFVTyOQV08Uu3lMQUOZ3/GdqcG2rmynI9oL56
XjyC2CtpgaYhNz815FQlKR6ZvBsBboPozKlxyDvhAnYyrMCcM6G4BiqPPYCW/O+1GWcvSdw64Gij
0oP+ngMgC2ua7/Lizv8lwIDf3DxqJ3qJbRtHcypL0rtgxnJXVWm/dIO+C7iurJnxPArlGlccQMpc
Ql1gw1daI93f08wu2riN0JHcvQsUDtiRhVTFQZFMSWaL0v9+tWsaQBL6Se/bRfzXDdoaIenOYtLk
yZF79M0wbdg+akGGCj523Mr14zmEoIpKbWQqaLIDLCDqO8oquJg3qtU5xdu6sKpxx15x/PCnv2n+
kSvT4p4bdqtTH6wH2xrkNDercpWmgNOL6Dsmu++vtOGhM7zdrLec/3XddggGci3fCknC8v/QCtkK
C2WdLtbRk+ga1/NXWlwIDKry1OmsT0AYBhD6x1rZu48wHXp1MokNPStr/g/Lqwy7QWMEBulGkyVp
eF/1h6NEC/9odhzYMhOAR8lYbvzBkUQaiNbuWdq6PHaTvUkU1P/9YqXNc0Ra9Rr6LQ1rLqJS3m0M
qODvW0pK191Am1C3HAiDJR2AdeOHQDP+qBAnjBOTSviZD7gj/PwmWb057bmNa5NsT8tTxL8cGsUd
qZGXFFoVrypK14F/DONA/wgrMJcREuZN0h6dWIaLKli0EektcoYanBlsOZOOOUebfOTbdmI2eFXG
wjC5wzIA43JLGhHhAJ9wJetEn8Z6hEGjmkkYJswA7lXHhm1MkJ0SOQvfVl6YESG4sSDHCnm4S9GC
OAbw22nxWOv+CEaS8I7qSVZKQSChfkKLs8NRthmKLEMgwjwaKX+N595HIZ81AwT+smi4D9968EzK
bAeOUsGrHklc95GSkDbp/GLWN3QVQbTzblVyPg1wsE4nNcEUUB3NwAKkHklxjhQGjYZDqicp/jDs
rBbcE0e5EfxQUW1fQhpZivn6WNT8WSz/7ED5DzvAPzVxv1u58CsmGEYnbaFQwBS0D+8p09d8xreG
6lkAEafG/3pPw2557gjkkAOGp+LaK34UxJh6vbIyqdx9Cf5UXVVzsU59/o+LmZtXdEvLqj9vtSYG
I/EOP+0ysSzZv1J/QJh6PjZ3hXJ7murhL0iArkEZ4eyJK8sSk7Me6roiabriFeG9ZuhOsZ/mQuHj
dJQCr76vJ8S52JbCp14KFEg8cWHUhP1O5MwlkekPC9k85W2kwr3Bv75Nu9xRQeW4Fme2riydwpYx
a0EFLl4c0FBKQC3VBAo6BHEo9+o2GpEtDiTBviHtXK7nm2OQs7/Li7UTH7M3WnFfTrhBVY+QBudU
Mx+U5FHP8lFTyhMOTHhKvOIYIZjbaeNsPK7ymslUjdAI0aN2u31kcJYRoqfKPdBAbWgB/D/f3Rnj
fGUg70tr6IA9g6igMr4zlGkPTsoBeRnLYgNBZtbJV4nOuOrDV7wIQJPcAVbRiBEu0ZbDpjI1Re/V
N6UCIcSZ8T3zeqR0jd5QoSzc1Zdwnzz/+PbCKyKCN83R9vieaUtVxJVguY07BZWWyii38EvHNWqK
t1tCMZESpajSHnFgYfDl7mrSMOfTKp/KW/hMrIkjOWU1xX9W8jbyBIkfKQ8f3dGUXLhRYVbu5d0J
/X3zEXILWLfM5fE1si6vze1FMzN5YdPGP6TdoW2fj7ALNMTIx8t2aJOrqc1/4DzlwQr22wFZo6uM
xa+LupDGnFmO6cQPIS8a1TTt14Fd8wPzkbOFzBnwJqOcbj0rx58sBoBAuJMd8+84CRAcOc1S6T5l
ie3Z9cp3MgTK4QjUI0k+lm5NBTdVKkxp5nIiidfPZimtiSLrSlsfyoHwqPO3TXo/QdGKc0EbYjr2
SlUj7u4jffDiS1m4CCLS/WVDCVeuEaqphsDuCTe5FHStpTfOoFN3qtb+ALoYnmjrARJELHzvS5WD
+HQxNA+uTavVL1iGWtFtBT46QDV/WO6Frvwj2DJVf6E8e7LTn9q4sG6OsFLhnFgsFaJ20u+drJ6S
qatgcIPUsXGUjMrDDEL9kyarZMRP3LUpoIx/x2bRagAzA3rsO4B2mPWXaciJwDylmiVWFTgYW3FM
FI8MOd6GlcNU8MTGMoIQXeICYf3UTAwTt9whdNaz7FW+As0HLXk+2SVp7vgqyBTrtRiaw3gRst2E
sosLKMaM/fV2nS00BRG3WCR9C5GpbqQTtxAgecrgyebvXChIZ5XWn+mqG3FLNghP7I5f7MaPfbIO
r6D3T4fGADQ5voQPTXSBmJbqcb+NN6NxbtvVKlwFKEOpdNbXY2QQ32Z1/jQrc9pEhIswstyLEZND
rPCjnmXHax2gq2eB6XO/MQY0fnr0b8s7AyFCuc5TgYrExj38osPYnNI8Y9O7AR7dt8Vwi7bhLTPi
L/dDNBTTXWE6D/0ny+QPS9QaXCZOxlEmzjCwYQbc1udcLY6jS8lILoJDwB2YMWgHfTjfSrMOEmIh
aJ75Iooiv/udBXRanjeWUGb0CSGuPVm60p7KVwIFg9bssTH4FHgN+dARXEXl4aAX18uYfnbrPSB/
nJli2uz/iVeo7UoHI4biuSVNUHzMpzxH+Hd7MPE+OMXK75fvDB5TbjEaI87ExEFatnaBj1jhgu78
mI/lE99c4/nlbcnv1tCIoEhYUORGlN7h+JBU/0+hLX6sCSBbUi78MkkrP0vDirHBFe0ayepBNbM2
BGF2AQJUOKjXxiGyNeomNsOD38OM2WiE3cXjZlpkrSWX5o7f0x2myE9rFAYVFJIczVWQGkUKqHAF
DBS3GXS+VTLHY5cwHLG6QJgMUozR93t8zCkYxblvco6SQxbm2lOHJy29RoeY0C1SulDQf1t6Bq8m
X88n1mGonVoG9iuPT519Q35PbvDMDHSYwRIl5SKw6W1TX+pO+P/qWs9fGtc0WSgh3zGIUkFO8bzt
CjxmUbvfkGh5/UdSXCuXMSLprTOVijhkndEY1PCtISR7gMfiZOcaeBrgR7Fxjvb2pD96qA9u4kcV
kgFzaJEz53i0NZ+0Mun+C08Crnu5LTwavhCEYdHAaYjimP8in+MkB2MJwTBLn0PL6/ATPAhqHsN0
W3qXi0VFGkp/T7dezv2KbR/HdpW98/8sB3RiI6t4Cylv9mCUMzsEajV3aIBWxFviAKoefJ2xE6uH
0Gk/WzUHsiaRNkx2rrM+wOjWUaIlJU1H14etPeblP6r6Zy2xx8gPIZGr5iN6zAhRMXZKv+P9W6PH
fn+ddezizcLep2sYFIhDKxNzAb70SrACb3rkqR1QS0C8rX2rhP9fYYdUzQiFOTC7RCPgEX8gBxTs
iCxnYyln7Vnnf0S69jGYhAO1O9IOwVbu/u919VQ1CGdv5rmMDg7Gv9f5fGIV4lzBuwo7k62MmSMO
TICI31FVgrzksJMJVMu5KT6yTY4O2fdQN3SvouSahPyd7LDnZ+cbedI2XFzL36EmIrEyk8LvHuzH
6RZ4mRia7pANM7EP2P16bJ3NbPYmh/LA+ehKUs7nrrM8CiIUrZRzSbVn1iVQOlQZ2RzZ4AJ8q1G4
V9D1pvRbICVl/fawGVzCVR7VBlGnd1flyMFcMEdbicELm9LlXyMGknj268+tAqpvEDQAfmGlncvp
TEX9UO7nxIghJcqMFKVesVrgJiSrIywQAdCxqZbEHT39afSs8XFdXrB34oAHkvhkGOERGNkbeqwd
jkIec+t6EWqFbpW/HqXA1IuUHuqzNIwVjVKy6UelRV7+cpriVaFTNvbcnnaZMqX2W9m+SDcHFwq7
3DPFI5NIoJ+KceaZSXrzxtXD+FSrOlvGCwMRjP04lAJHCxN+ebvOlRTAnv3humc+peOjXQePy13n
J/VSA6hPB/MWUqWpOsdCncbDUXRUKIagQ3V+qjGy/whO2y5L0Dc+tosltyv5+akmK/6iCGu0hTxf
u3x3nahMqSoFdoltcXcn0ynyPXwBD8u3l2EFfP0Le7r9JVMUsF1z+9JC9EcLKiHrTzshYUjAnoWd
o08mBuuu5kw5VWge8Rl9HCO97bNer5DF9P0/Od83Kw3lkPAGButVlZKwpew2ATucliOOoJJWueF+
4LNjdzKA4JMcFM/uHvyGYtDjfSepdO+gpHywinQW1twObUdC+7GzYzeUyXzn15Un+M+SyS253SKi
LD4fdUAmuRFhkpbMWcY/EM0SPyzQg1O3TyogQtynURJdNU450gfn1AZ3POggLmbHPlOFMP8uji+6
Pws+M2d7I4ucKKo1LTNRGLeTI0iMKEJal0cF+nsBXZKCkIGWm3mEJ18UCUDLA1HHrbYsuMBc67nP
AhMb3WbykHk7i2SIyoKqiz9xABhjZC1qBZfylfFjnIa2k8jni/97j9662NvRR8wAizpocoMyaEof
ZkBOk4jJXvUu4lExcn7qhuuwr+F+M5VjpVtSPJS/IsTpo9LhVQsq1f8Yg5Qq8M+ty2It82SvJzLh
QypD1XpzegcnN6NAb7/kcPd2LfHb8p6Dqbyb/M2zMQsa2HEFPv1ilmz13p/HBQ8agU/mJIoxSSia
09UeC8xvU13j/GOtWtTbeflwo/5gxZJWtnfurh7dvG+mLXPcfibpv1sKXVdsyCvPjUHZ+3OV2sdY
gO+7zKp7rCNDITEnjxtgyQI+aDxHsZ48AnCzOWTin9hVmrEXkTfxzPvgFbMTzcq5G5oHuWLzGBHX
4ss68uNaWi/QNWmLx3Zs1D3+otPbQbVtp430DCJ77GoogUSXzgXD8StKT2AFJSicWc22DGveLe2W
O9DalKJ9yIVJU/af1gsLMOMCjcU3LASesg9e2ERpAl9ujEW0W6KQ/uVSk7/QsW9MEL5vKiq63nIV
AbU2Rhq0Wl1dImS/Ofn0Yi4Lj4auXHAXvkl/RIcSc6KrV7oTS7Dw4l77AHv0Bem7wlwPVn+ykjrK
HvWJ0eNaKsr49re/4qgUrEJ137PtxYVo4GNJ6vR6jbp1MPXeCKMuNTZIGZXX6KrRdloKfz/VNZ0N
jVkEPTGcCcMVg5DXfdRDwz/UZaW9qFhNOfotUsSJI1/P+S2vrVU04cCTn7Q8a5pJAdLVu7bP1ENr
NoulJLftq25tSnUaanEUvivbIlgLTNSRVqnRIVZcYQnNzeW5S7kcYYwRYmgMtU6ErNTKGntXorDt
pePDb82UWk2vn1n0x+CzE7xfE37puAUPjdZCcQHxLX+nvV7t7DWS2qqXrHmEEuZS2qDokHiT8hoC
XuRVyy0bqqghNkWcZi4wRH71dBz0soOyIF5Bm69aDun49955gTHFvwbirm5jsKJYQobU1sXswMjs
2YRbbs6mwqhY0azozPBuOsqIV2zlrAkqpFF8JyQJzd4tn94bm5P3BGjjzrz5GfeaVkLbfae1Ra7l
TltvmJoXyBI/1tMmHUCE5UlxcT1p62HAiVYkToYD+ugB3Q0hU79bm0/YxhiUeSK1vMwv06Iwd3cD
IX9q/lyUR01xBeXlxy2sSwHFKY+Ai8XE9+dbDENW72YX4xH/FVwb4AuiBT35orbKF02gzUm2u+lr
4If1EXu9C/+wuXwLei+fH8z5p7iUT31YCDm1ZxNi0+0mBXInioobigB45lpgpulctaEhqphhavmk
DC2AZKSi6GoJbIPw86wDEITD/KTuZEtJ0OUt1omRXCMee55qCWL7WO3ozd6HDLdldia/mej4qRnH
eONIYb5dQFiGBnQ0ZEN8FFl0QkMz7Ch0bALhxqDOIJANgoGDMNjQarPxg/dm4i0HTU7B6MRt9xAe
REFwahKbGjGx0PYlsMKSWahI13fzXBQ8pZmFERwixakAENe8B5tciINhVjQoYj847KcgHc636ryH
CtULXQ/EKkMyD5e4x4iOhs3TOt2T2CbfYTCygIk3ouORhAwMQQNL/pDq4UsCRpk4y/b5wdbHKy6u
zb6Yc0SanRJsQxXGskogQvS+JjHNDykiNdCnWSJNsgFDUt1y+upRqvYLBJToBJdJF6O/HmSv0hQB
pGN2rRwO5T8Pt+JZmT3/7/RSwozuBLBgyYtTcCrsAzaoj59N+fXWslc4WT95BVNGmmGcAL+TwHWB
8rd4Z25O6oPcwalyyJMJaxXgI9M1dsSlX31LdpVuSWpkpqDjzdjOD45dR8545ZoOM7hhUdO5rN1j
a+RsZCzN2bInj20WAH88b+iwPoN8LYruF4P1MeC+7WXev6V2Q1Wouq05JCZwBqNJpyOwzdmtPs9e
8jYgvFwMi8/dHEVdcDx3pvi1nmh/8ArnpR0OCkwrsjvc9/O8QJJ2tRMQENzBbsUdxgHWR0+Jc40b
Irj1KZS87XYZsckJuTESy6IWTigcv6lG9dKw/pN7Yfpl3vbF/XA/wM+Mt9xYZplmnjftp+uwU7Cd
lucxWy3CvreCec3UCt7ezzuWEuoD3Gr5o+NbJgm4TOuHPAE52vkXw3bxdW/+sjiJNfqTJp42rFuO
KO3uHhJSeKZAqAEr5WuLZynqrJDXxfApiJ1EYvjVit/ZPWMp8x+mw70+Y1OFKQY4upbmCQKrrmCV
I7JqDOfk2wEnMw+AyvAoJ4WdbYKCsFZcmF2pBg1ZZnhkJjEDJyroVb2RAL9XGCHZ9juZMe6zoycE
9joNR9DL/vOy/nZMw/86VUYOYWhH8jw+Wq77m0+aIvPOI7zDpHZZdrr6Kq3hFN8oCj77srLa2ZV0
9BJIhDPL8GgFacXo8Wv/5e/lNuuFTHh9jGZGlXjGCUcCZn3eIru1WPC/YOO5gRjCpRmBgV51mHVz
XzDiGDcH7pzKE68HyntGsK4dIW/IbnFTiTV8N/FuD90N5ru9vIbGlrQoqFr5ssSIakTWLeg1dfmF
GyJirnQqWAWrYemvaXehUsMPUm5+TEtOCSlvq9ZtwYRggVlM4kWMO53ppg6yjhmbs8Jql6gTydEi
O33h++m76msCJavtKqvGHjIYxkA2h/AU1EOUoqp03JaydU9HXbi9q5tcrDOzHFQGC682Qp1BSL0Z
hmmITBG3gXAxZ/ghUv6aTT+GEX6YXZFmNS7bqk2LWmbed95MYHr6jO0PUkcxjOaNy2mVWzdWB7Zm
71r5D27JSJuekbTxMNE+X5ubp8LdhU/uzSDNxsgabU0T+U4xaMkasrRC21O2UN4cmdNxMstK0nTD
KD5g9VFhiYyfUKC3E5V99os1tG+sqCWUJ4fkQgx6wK6XRwGVyPcgkoT7Xmmu3HxnzYLMGhADoYpR
cjRf+k4uFJ1Rw7EqsABK1uzdcA+4/5MOg+4gC6w5X3HPXFNgJRl1a4OZb1X3JQ/orSt3gpm07BWY
FTYp6VHRGoFdAKQVOyDTGV4g4Kp9dIUALyEpVsY8jqID8PunXpIutWfmGAh65B1PNPZXTbtgJhNa
HeuumiKXwBnrTvFP5dZEVnklLVzH4E/I1QFqjQ4MPu/XBDd1cxVHiLLzSVVY6L3iiTxD9xiq7Oml
Mk+OVIa0roTGTzkH/N/QDwafn7L/Bv1RTKzqF6IN+xLfYmSYqKOHrQpYIsn1ZFZKPdhR66XCZ3qn
9vnQU+LqAlVuEyfqPcNW0na8u2mIq340mkWW0HNG8lakEsj8FioG8QsWAI+f8ADvWnaRnyu/Zmw+
Sudrm0BS77fOQKpb+HMdR5ss1l6AoBZ4VRBb6CzWTffskeWiwcghRM1YROzBgnk10390zBV4TtHC
VyUvBdjZ4wY+KlbjwE+mUXA8H+c6d5zLBiKkU9uu2CXaUKhwjC+oIgLW81tmAVVqCfA9vvHboxqk
SrER+SpL2lbiwoiiLg85iQavMfoYmvGvGiKtI1nDKybXIuNjxRAbF7znl++AAdqKUyXaAQKqz4k6
tZsW40LO0zHfxD7iPaLZgUAsGlxs0AdS1yfNxbv5DRN9ykV9fxSlSPy87od0MBeFnXf82TTDhplG
mV9FIRro7yblCH/uzcZ8285wunTMPVYzc+Qj/XXCi+kMtSQxvjFeZiapGrHJRi80ymCylDQ1nhXk
fbh+bgQhMs4u+64ZSuf/ddnk+1CzqIA7visF0+1H/fQ0PL+pI4B+kcZAq1PqLDVikLvSPVbuBdNV
dHXkLCwfQrPnDGf4MK457pxMUb8XODyJDMR2X56ph/xyV+1xyK0wpMOHmnuXTBx9dQsATc4t7xvm
UE+GeICpbFv6cGqxpeMIX3mT21UTpBEolqrGb+/YZsKXm9xaWxjZH57OqfhVnLpi2m8u4P0F+pQ7
aJl9WtvwepPmgAW5JQvPnTKgtwt+AsntkSd24vEEf0voaA0IJSp9sFKfn0CcbBMeKXkNx+BXYJjU
8upxprYy59qeapAdHcPUhTIZ8FpAIgEC7u17ObEwsAf0lPnNvbYT1J2yrPUXdQZ5KsvDfQDLYwnc
u54eM2keBnd/DK5c839Az4/JeJSlT5991Sw3W/v588TI+ufCCNSgIYAfNwzQJH4+2v9T6nTW5shw
be/Swt3Rh/lz85HRmt5ePwaPXv/0Y5Mw+99/iv5c3o6fKeZSlq6zwVo6iNscqXF7+rzE9/YC6n1q
BKj+rjdE9KHAG0XW5afJWT8ofxGG9FKeogLK8zPx+PlaouNn5XvJcywbVN2D9y9C5lBnaw/SNMFQ
N8PHqfQkEm2uYMdBak1RvaNnGEa9zhobUoS4A/Er5ScaxFtK6ClOWWgGBraH3zWBrz23c45A/Y+i
ogMdAEsCH/ksmkX6X50wTYPWGDDcILxQak01R74n4JQQNmayJLg+QCG5K7xNfMUg+d+PSsPfr/FE
hLPnCXmy/JVKy3ZMuoPPu6CBVIA6NkSCoLcFcTlQZs3M/x3Gx7nG0qXkQJFW4qNPpytyr7fpilWj
mQk2eZFA+4v386239XEQ2bZdzqKyihMEhmOYSsEJTFvPO9NNz8zyXnlV0LvOZR0L+Na7leGfmRIc
mNGtsjfGzEOyoau9FKKn4EDGCOIbZ8tdwaMnl/Ql6uFOgSsZzHuLdiNU45os5E/yRY46DpSYYjKo
sppuZ+d9KpUC/UDEjVjmbD0po/ladyyH/yPOUWZW3LjgfvSJqxVaX8/7s03KKm9BNUo37wj9XptM
Hy9V1VqtYg3DZ0Cen2mm61xRXqw07rVbVEydHmJ3CB4V4J8K66ye/qtsps5tfeZyUrmEa2hoRDza
LsGjM4LDFa0o+11x7+L1LM71uzf5969NU5M2+o+yToq1JEn21ILeaMy6Yc8ovohc8c0OACC9nS0E
ffwmJpOnmzfBnlK5vjfW5uMdz70wD2LrLqTXj/jZhBvvbbuQmeDhdILD4gJpQffZTuRUnDJFLayd
dvpitciKumZO8NL/SKsaQca7EURZHxRRb+My43sS8Syk/rY+7q2XySUuM0SR7MlnYNSivNpL0kXw
8sZr1TYbA5eAFVlWrcmwdPyFnUhq4jRmtDnf5OxOpZzcYaOYSXqeTg8udHZ3r1CV5tonwtcRnCh7
AHme2hQ7yNh47k6QAvCoU1pEkO1X48lg12gAf9oaa6KL6x0qEEMLPgFTyHdKJ/RxtJ+HFLYJj/tW
Jl3jf+d7ETIsaap56Y10I0zalMzPS9IKTOktrq+PknO2kDfIX0l/MNWMRx8rx5fP0bGsKBloZrGz
KChskjCGlj4++1GainAjod7F+JLIzXEEWU50mpA7gHDWm3Q4GrfsQGHh3aQXvyXlnPaUTrI981jv
E8SeB0fPh+SOOdhGuy4NnvJ9AqKznESL2U1vI5j62tpCFN/BJOgWUn0RXJUACP9B78t3U5tX7ixq
Oo6pDzJ3l5GcBMVhMdl4h5w3OiCFVQ1HZE14g19d06jj+hGgTHX288vM8840nR2X2/Dj1zh08BQO
UaCVa2MAolzfvNiLTw6rOdpRemepgCIgE4PRdicgPmgj0+PxIGGRKCN6NSC4OqUHOFsUpFCPtCg1
eHlIZBMjszR0pC/CZbjcV/k7LJqabTsRwUb23J0nX5eItLMNecRjKOxrUfLnE1v77OFSBzsMjgtr
xZT75ZBBtyzYsaDFIdrV73ndbN56z4yOBZWKIa0DLKZagxYOrm4nFzU2S/pOezBoq1Sim8s/Xh61
x38rC8WnSg5q/JowiKZYtufrTr434JldC2ppz4nK4yWQbfQIN/AYX3KjNBwz+vK9fZBOLire+oO5
+h3Y1HVb7JrUXl0ZYIQ/mGfswTW2RVc5TQk7MQHuEqZF8Vq+J7aYB35+0RxMhe2TsfJvRc90F1HD
potIzMIR/LJM5e64KOmBr4nmBaDE7S1NYjrjwycrfArRiqAvCNJc/AFP3yZSSWfm1z8QBVvheStg
jdM+gvYY9++iBT/isuwQ8n/Ht+tODaXuaSZFDnb/YXvo3nDkk9KZm2t6UjE9KSprnrAgWikYBjrV
7x1TyxrTYikH4onLM3gShrwinqlv+peSAMVKvTENbJa3vQgDm7hbqNMP3LNKGSmuxgTbk9YrBj5R
A1tudgXh4Qc1P9D4NSnDYoemg6wKeYHgHBu8vP6BNc8Sp0Z5XL1Zp4qzGTJryhnoa8YWZFa3+nfF
QZzRKixV1BGVyltnT75jQ4QFV2YJQSLumtAlTda991HChXU7JCKFXy9xFja87Pbx7VIO7aJFbGue
AgLvHoxhyhli6fjdBDTuVQigXy+u9RQLjke1Y27ZDtGEUQLUHF4Bel39Z60NQcPgyHZ1UkN98q+M
nxONizjXFuwFVsK4KRgZkN1hA0KYhAA9ZPu/2L5sgOmMei5tbrpli9A69GMaj2KJRX+Z38OS0Hwz
kltqnq73DSvihEfyhcPkC50mwTgcXzhA4k9S7g/+o8wfmXNUfka8mov/ADuTN261OUSUrfdQSDxl
d0KIijB7pscBPPlAkFyjdNQKGukvP4Gkw8wYcgjgCT20fROS0UFy7242i8Rm22XBmcWg/GhLWb+G
gfdm4lrZ54i7z59uXsNvWDmlZLrUSD8BWFQHWQvfG72fnw0SZohKDWhbDDA7lkl/lRz74RLhJkUB
ft2AObTdD+7ZDBiTMHa8MEnp4glv7FWQMhBRGvAyMYtxzbZ3Oa+BBzWla2rbhSJMXLuMlcOfe/x1
fOGLsSO5Kj219KA3Bp+1sOeuW1bkYDKj9OZe6t+hXqzk+jaKVv76PGmv88b4v/K/tdt6XWN5K1OV
ovbVNeTl3ZImt0hWwWWz63OSB5Uwig5OcnEaWRowCHr4d0hVF0Kj7OUtmd+BpZV9ECpf/e8uaXoi
7de4ULFXHdFeq6XcWcWJlKGkhz8Zy0lohm2183b3LLwRyjLH+QoqUjHcPUUOvCcnhr4AV5/bYvGI
HebS5pR1tCLyEKNMEsUz9+dwvFNaQCAiEwd4WDmN0SZoy+8FLezVDXXmsvnx/QqLHiNaZWnwrmrM
ZEd8ZtADdNlxrOnT9yokx4QLRb1Wj4WjM1zrMrPm3cMlqLYip9OUa3M84cQOVCWeVlBOT5cyjffx
l98MCBR1liV2aI2l3tJ7iXloRfj8+Or+MfV7ISMmEQYRD/D7Sl7tB5hJ2bsmSsQZpRQLCVn50fpP
Jo9PfAAU3rTHpmzay3xLmhfX8N4Dn+f4Yds+xeauQzHz+XTzzgpnFWQnpB4PdEPP9k9p8weHVmYd
/fNMtFch04lnYMr2Ro6PgskFCm3IbHXjQWZx1Rc36dETn418SewC63WY9KexFZkMyhemo1GHi6mf
1+YkvXwMxv/oUDabFupdZY2NP3AxuKpoM29jLFkLhV+YNPlHtMhSn5D/xBxy4SBui0J/qnryit1I
po2XL1hRCMzfZGtE6VIrE/4RGhSyofahVljgjvcbTT1C1ZVa9uTxaDJGleaD1Cfiriws188+xhgM
zwXhXrqGoUa1wEG4Hhc/sBzKXdlR6cAhQsFlV8k4WzUGMz6PiSzpr48SXlvzVy+fPSs0e6VaYirG
nlLhpdvyw13SRSShEK96O+edM7M+ZD+CKVV9VNtY4oHzsiDeZFdOlujFmFjwEZSco5ixfHxyj98P
O6HIzGyvpo2AJ3PoKzy16WgoZvRvhDxf/wzCw8fZ19V8mLZlQPSGVNVmbhWkd6kBBm2bpgXj37c1
7icToo4Bcyi++FXSLSGyPa4d+BlFX3EdJD+l2xDRdJBmSNU4goIfUAmoPj/4P244O2JBczGbDCkz
gbQ8M8TP5tqquqc4RwvMtCihkpBr0fMgtucRlfLTs1NS5V4OOnicE9y94OScnhsOZDVQygYn4TRT
kAWiVr4IDPIU1pwIHOS2RBN1UE9JK1anw7TSIc/+K2b6+SYRYRfh+3JRtvUYSIDvco+MPeGLzJG6
5EHPwZxHwX1uRmQYam5NESAA99cAYWHkHOXdoVNEy5IukGatIOgE12sikjp00Wr3vmhCe/010HAi
tyWe0bveB7YnN4sfmAcTjv5shg7jU05IbndGnqTmx9xW5QEABAgiTavNOuojgXANGOEVuz3r6f9S
rqgFmTtuhgPg+breqODpxSCtwIIUn/QsNEbUnTslWsUhFlV7r4vPEGcV/L0tNIPXIa0DdZ70TPqk
H6FErYFhHen5RWcGcFsGgtJttUBNR5fpS0Oo4GCoGHy946xrhapWlrPhqMuJX5Y6PMcCNzt2e5SP
634q2h6YapcWRYYooNnYqembNxjk9jSuNv16bSsrjINIjReNeYmVne3UYKG+6oLSzJ/tYAbl3Sb8
zx3qMswxj0v+F0py8qWQwXfi/J2Ir3SgIwzTus7pSOyncPNvKZjKJoEIkDdoiVrnNheywwVjYD5z
hVph6bGm0KF61FKXN5FtNSjfSlz6TUTmSWoJ4iZqHWQD8KkcJRJFXd2gC24rMw4sDd+HV6TkIdhc
VDPl+dcW6k+SPclmPwrQE/vnQmLN30l8oq7gJdmgAPvkjV46kg8LE0ItR8/XlEAmaJXlb++y1BFj
XYNSSjxbJz9U583OolaFGf3m2eQLKl110tR1ujlJa8Vdz2IHDmx3gq0WG2aC/oceRwSAVeKsTlQW
YADkLDvN4QfrXusmafAubXSHPovruDxoTTfA4MyWMVSSxLad3Rbi05mwrd+Zg6bFZVwyZQ4adZd5
G5aeF+ZK9zF8PNkKksw7J/D8yJhEz0XKUgpArPRLpwwfroHRI1vF2p8vwFWKWQ/GXhtx5ca6GnDI
ll9qQmGMc0tXz70m5q2Acx3X3Vkef5ZseWJr0xTmYC7xQnzykMWFHzLBFr0U9QHoYdOrgcC102fu
FUGfmfN8LmcNEieJkD1RkQndcG6moBjR+iHn4pJ3qKOanWvQgYxugXsiDNqUaXigTYJXPwAGkZkH
gRMEyNcdoV/BTpaTOQyd3ATJ9J1LPdBDxkS6M/0NErm9SeOmSQ6d0UXiSwwfWv6pkztc87ZSBSUT
vj4F3+ncXvOjpdBZi8t940UR5qA5aQ+Kc/W+nMCubdvFKOgqC4saPOanywBsAe0gbKVzDqmogtRg
gYgVf8V8rRu6bu0NnhY/rgSwj0eQhrzVQUQcCFJZ9aPLT9daYgtrlXMhcAMtVdtPK/KePyIkUi27
0HGN7bT0T0DDzIbVe0n4po/fjxQ0H3SviPEgtBuwRBrBXJgmw5JWEUpvTycIjvy9pykzaZs6gwhr
cu2wlkcBWhCI/NnWAnPFxRhNoLVeYdgTJNVucCZOGNEn8/uTkKwShNIG8DFER7nuogzIgchi57UX
9iJI+pQwjZSGvl2dObR1DNJHCBu4HEtifXs0k6QhdXdgXb7JHImQUaxlwIVdd5c0VM0VQCb8qQTh
/VljRKNy06FFxwI33tok5HFkBxZ8vXTOHAXYEQEvP0VFBqQH23UZ+1MxFBH1KpRugj6ejfqw5OxY
kb30k7SUkV3MsKCfiV20V1yVDsLBlhPKgaAX9Ys5jposZ++cazMtZ3XRMNPHobMbTV+WopZm26pJ
TMiglJHHMDShbMHjFoG3LGUdIZ5gkC7fVxp9MteOOU9FELziJrVAHb2iemjhgadITNPNhTZbs/dm
0j+xpeAuAcoaHgfeKGZiAOawjHMOTi3NCnK4zFTU/HNxafupixjxnSqn14jABQUmGgaBxNq/0CO8
ThA4e7dMzVSsjeIPx3a7knIv1LHMyrl7G530zlKG9QMFTBZbHPrP7xsQowcy+LCdsJVklpkAj6LH
inKVxqfFrmdcCuNVy8Dx+JDMRhnj6Ipks2qZfHPxPcdlEuETeRWCIFHGpCxhgYIj+iOo2+4CF0Jk
7M3X2wVQHy/XzcK9fA4O3FkFl0ufBBy1r3M8FZlvMElKyUTPeo06VLKX7+utnXgi+31q4SJj0Kts
zoTMuuK5eBZ3uXcvKfB2vZ17bJ3Q86Bo3XVBJVB+YxTEHKX4i10fICW0vj5zzlfjljlxMk/K87vb
Z8haUX0uvmseAbQoMlkUlvEMnavg3GclPbzB/Ndf2+AIHldqzPOiKzHTgiDBjNBcyIgJsAX1QIC8
V/6qMYpX6rJh4D89jY+t43sI4Lx7q+7NImJNquPL49KgzVLpXO7JY5duhAK400LIzGyVNyaqxnox
A0BnyJjTgufkLLn1xthZ4JdmZdW/rzHVvPswERzVOKEkSojjhmZGmNFi/VK83UCYZsQ9557vkjzt
ckYSk8tXBg+PvGS4fdnIyaAAr7hUVx2Z5leWcMA5g8S3A8gLhjxQ1dIuXACV62OQJP8hAPNk1IfS
BxkCLKsUEV9XSodsYksbHThut4kMwdtQ3EL12nRqwWuj5jJCM2lj42xH5wRGwK4J6OFnMdTcuuYk
FNpzEfGGgMRhg9s4zXIeIQA6QNYxVzWqLt9jtPeRpxMT1IiCnrzLFxvEAmE3oIvwGQFU1wLaCVys
gXxv0/Uq6bxqM/LiX6yMr2nhaXoOwsdk3H/AwYZA0FqPvoz3evfDLKYX9YuCcn7DnDSACPjOA5ax
FxJWqBsKiR6VcxsuEJQWGJHYhfykfaMEbXmBpxZo+enH39WCpZuMBnmZpvnQgUGUhyWkPCDqZ+Fv
8cc0tb3CNxQUz7Ft+cZGq1EewmhVcVz5ePDxO8Gsh9D2R0mRJGc3BRJWs/Md8kF/yofdJqGAnP6p
UtJN8iK90pqU85dZu9TZdZoypK/vg0RWGXomnsH0QSyvbnzSNAwICCLv2Saar7o8UubfJtPzLeNs
rL0mYn/+XvFnUTb5O4C+s9JKDJ/uk49zCj6kn+d0rnD92a0xmlJRc7SNdbW7ho0xS86ZEbWcw7VA
xcjO9VVwDRMXH7wcP+2Lf8E3icxE8rHO3PHEoWaKeLy6jsdgVZuD81q7EdAMcJRIMPp2M+5fmCCI
2NdrpMfCkyabQBjS3E1nRcRiQf/rDowMXZvEVu2+a0cIeXS+GGeHJmVn97KKH1z2SsGZJdr1R+4K
WMF6pPLZvBD4BBnckGpYYOy+/YANHrp4NHBzputNNOsvdqRF4OehE97EYedykul71l47Nvg8LSmz
R+GLhrf6Z6LWr+OyI/lV8gkw6sKykotwksoKPvI4qaaHGpvomHJVKyZoXupZ9iZkF5V2IF2gGEJI
JWsb/wsHv3R6iOBmQGi0aJkIcOjWESlzuRbKOXjR2A/QdDFqaET7+6EOH9QxywsczMUK16ODDnQ5
H1AQbW6G6SJGnJLx9he+5KoPnvrPivsHJdGH9dL+FZPKBJ0zLIeX8jAK1nBlsdr7X5eqfeNacCzh
GjiU6D8Puhf4rvkYI8w0rld37JzDrD/5yp9/nX3ZFt34HwHU1/zX3LJzOKX8LKRomKYMVfkD/VcZ
1vct5AZ4EoxuPJ40tQ5Cd5qqfHsnsv8vV2DvBkR9y+FABojNVtCovQ0KcH9NZiz9qstM2pfmAUM1
sEWPh0KIU1WpK3CJeANcMgAqThXzQ5RxYCE8oYYj9da1Ofg8DvLArdM9jWZHA9/v3eODpNyHyFt1
6cLADYgupimadjObSudimPEVVmOYo/EuKBCNEIQbqbbHWoqaFhqFxNrNuqGnSH07cD78IDJ2EywN
lSeSXVz8ZxT9QyOid9Bh237HjT4+txN20CGoRGUkyR+rqBbfIsUJ1Vg4iKJB3bEEddyF/oGCAOhC
94FDxG/5uV08/3XyCGJtHc6sUqulVundXM3QxEtgmAzO+O29oLAT98RqHlZacxtZZAdOVOyxdiMI
71DaVxzIDjWvOkYc8pAq8xSTZH44T+2u/IXBlXZMouxpV8MUxbgguntkCd32qNXyfgYYH4P4YyZT
JnHnsZ/AYjQtjkhWNWLJmaFW+1xtC9tKhjZJ6gzjJmSkR4QUOapqUHdtZYf/eV9vQVwwVcrmU16k
bx2ppKiQUOZKMnVHBcF9GaQ1OuvzoekufCKEEdVf9PvPTWqQcKL9Cko7RQbPhv0CXg12IiK3JHC0
WJjQ7G8AMckxYDpxV4UWWE8puLKCyhyoxuZ/t4Pi5dOlHX9v7s61uQSCEAstgZewSON8Yc190reE
zTIAFpHVWAIIzCa0Zhdg9RQWwbR8oQBU/RN8iXebZf20LBbJCo4k3ZU6kDj/9V4Fn4VzDVygQgHW
V0s+VfOKTEmk2BKJI4PXptiFrF5qvejQx36Ag7MmANQbh+5bhXaaBGw1qRqyeKEWHPoJ+CROYBgx
u15jlfXeKT6DGg6Ok/344mdDshysbixhu0RV/hqPbvSMzNB4cXI9qeIzpa/+v5BRH8H9iA+8pquf
yGU0T6Po3wUl5e1icKQUmbttEELmUp2eUfFEbD2eJnSyI+tHW2BgzLQyKHfJc51PMFtzM6LUHQVb
d3cIXYC7vp8PHzDfgm/3YKYR5v9D2Ct+L5jO2ea2+cXbWHxwQgeDnV5cJW4jACqCg28Yqh+r7gO2
Ab1jNkYDaaE00fQ0a5RhneqQ3d6/kHfvjS23w/TfuTlYQ0LhjnDyxiIuYMEcFGzMnRf7UG1/M8Wx
ohph75oWGhe5msu5Fg/Hu1qtwve8bryscuppfdDcLi85y/Tk5AjEeTn+8ycBA5nmhK7svIIhyZE4
Aj27piGMFIYYJGj723CK84k7kpQ17x5xXpuCs9Sd//YIbpdcIDtKBs2alTbGz8cgjYzC3glcEPdY
Ze5Dfmr3iXSAHIbdLEQi71Tj9mrSHqnKuowjTDcCRDVaVEkMN5SZD7DKjOVYeCoyG61TiXDRSDWu
h34y5iNV1C3irBVFbpfidAEdx9QpPlko0K38Rc28otR5Z7cNGAlcWpwgfwQbeaCb1JM4QSuXcAF8
cgR497dL9CDk3n+E7hzLpYFBRXqRKZOf8p7pyPJ/DQwtSUUGikg8rywFOV+KmJJunxChlzF5rUN+
ZiULh2kfdUcEp/rhe55++Kco9fn53MJ97TuLMg+KLdLVe01eKPF43eAc2R+Ec1CDY0aIyWXSytVe
kblHiDKQDAJnVy+LOy1veq3H/vH2U37kgt1Z5aktOtHLsHa8seuPALdhLkIEWgcg3BLWmUUKqa3e
PIPoREictTxs0WdlJ23rpPuEPeTlNN76vN49u2CmpXnnpVAotw4tIhS/YFNAxxNAtBDVVG3BalD4
HgeEh7RKP24Y4q9XdBltanOhxfEF1xjvC0f/5zQea3KHyhNTXELO/eT3/elLJuGsQf1j3njKyiOx
ByDwHTDZYlGUo2Mf7Jnqk0Qm21nrnF3oRhggR/D6bl6I/A6wu5lZaHAPl9UCAnAwxTaXR558aGzH
V+j3Ew8RdtaxkbTC0mX32pALSW1NlsR5lTb2kJ/sZZ+190Miu9qmGFf3fP9p4WI21z2j5dKWx55K
zh7lcM9K6mxefMhyAmVkxb45q4TNu0sYt5mo4caOwBsOp521AoSrfCpHhDhSiqEB/JH9+LO/D1uA
grYE8OYozdSI8+2vdx1pQsEJuBxDdD8KaFH0en3ethN6rPM5lX/mTJJPwRGrOvh5vNdTtM15DmY5
Vt9l7b5uAi7YC7MdQbUuPMZ4myvsrysefLNqN+4PwnEqPmTBchKOwtdcR/VuD/FGw4khSaVRoqC6
VLcJ7mrZOkYWvF1kx9bReqOf8GWRvQHNgqjPXXnuEew5CPQuZ6lIGtbcL0e9u/PSwJ1/lybC/6MC
mGi9SQ9rnRaLtVyeqJZJUZ9esj/o+o4Hx4u+xTBF1yjf3bC1fuM0L99HC+4E43p17Ep9rsbSOuKl
HuLSQWzmDZBk6AXaROTeCIQNH1qeFm9A/P9CsK37mw9EeJ2l1J7uh8JmfZnSVdOWWyx/SHUX5nWM
J8iIoFpzoqPqyEJRN9+cuP3+nePrp76mFUbVQUWq3XdXYYj5COQa+1xEqk7riCINfsoxQAABV/Ah
TiGe1WIAoFRtWizzXa5Hm1GOoYM6k0r4grwdFQBBs28sTAJ1eIz79Cww1JXy7k3x1qDoA++L4s3Z
2GNE0C5GaOhWv12+9OHh7IIa2Uu9/pPDnluuCM/IdTvchJ1T7x1nIz+mN/lQHFtY8bqrK3n8z0tT
EIygZhUkJEDbSSkE/Ln5m8GEWsAPKd85of+pzW/nJArLtvr40aDSQ5jEpqgHkOE7UpiJ2hJ6/0O8
unT6IrvRao7dKwnbtrrf5MrSf+BAHhb17/lzWswWHbay9UfjE5fUFL378/1anBGU/f2d826wuw0G
JULex8sgD9wmiMpBQ+btwzV4gtwC16nJ+eoV2byViAnbqsvFlX5XP+Tec90vgVfEN9Bl3+laHE9M
0X8I0M9UPzheAObykIZ6PYxFfT5S3H9zyg4ZkCZlzdy2l7/euokoNrh4C8gSv55l/tYFm7Iy/lL9
SHCG72oFya0w0IAozY4uXBIwPy0BKwCYg7bgetcCZfYaymN0amjKHNrfTnHk3NdaNoWJKIxBpO+3
1GPuyc39gd7eOaqDJLNLjcyfvJHWduCPiIno+mqJr3qzPxWiyu6RhhoRAok+L9neZ1UC6UAIHnhx
0apYTVsj80QpQvuVNGjRsxOXscTZj5YkHwnFl1N3aBs6dQQDhWlrds95KoDu06cdXCNVGLTL8d5W
MSX/3nzM31IGUieVnr+2C7lmX5BgtqKo1foiyIZUIxz13u1xaxO4UFaJI6iSU41aL+kcqHSPhE91
PgXgOci8GFHiRn6Mmhx1xP5kEqT11BsvT5SQuGY+2q75aEaTvuG0yWjRngLVtIegtDIkttLuTL8Z
D0PhScB32R1wuh6KqAT9TvdleBuaQTxVNZOmLdurQdfmhVRHI/XUSW2iPyfwsmM5VKcCxOVnPeli
sE11jaXAsi8+CTYErSH0152/0vxkf04M+hlUT25qmihtZcTucJMoxTnCNqO2fDlTh8FSd22D4H5A
WYiiAtTxAmKU08qlW7neORxoxMTWV0Q7EW9EOj6SuHn5s6q60ZliYte4Cp9aLqJSmmMofiuU34d1
1Mm0cHza/Zj/ONe1jUiUzfJxgGF+YZB/VC4Gl1gg6Ud6kPbr+T6iVQOLhgIOcLTttZuMJnz7V8GG
yNzZLB7uQfj3IGwB+Xom3EZamq6n9oT5Z3I5jCHaVQC5rcsUZa4/6Z2LdkvOdUhCC+PetSyhWJdR
J9RcNNn5cUGc1/h1qEzRANCwzdofcvRfrKcBVjTTcUhDfVq7g3Ag80iScedO4iS6PJ54uAlipvKQ
LlIrHmDPVy7/+UDsLGZu4xvFybcoAIMtdfFJqY39cW9mJ9B99y+z6SaGh9HQPA4vtBtsdso8QZii
78Jga0WDnn7dxINC7eJju2cSAp+yhmvPIVDOx7HCzxdsJonWMvjP3/Jo/Gm40TAyhwHpdeYJpqCV
XeHPax9ZBlLiaGk0C8Zlj1QEVl98zpL+r9eJtop9dMhWCm/86eAHJ97PnVBew41ll1JNFNwBH7rS
kxajrcwYll1X6+F7LBsIjla94xXV4eDgKmzReRgc0u7u5LVGtOr45y8wGAwJsWnW7L/WmuML9jDt
uJ74vWgrVwk1tMUO3GWl8hxS81Vh7dnjZ6uYbphA+h+L4UXTfegCjJPrTeJEDgUYrnh3I0ay9tNO
f+zClRyoa9RGelxdLptd0HvlJnGJjtsO70Idj7Si3Dvf9n6S9Mkw/gRbKBj0IKVThhKyhHfdhhwJ
rLqlu2jzNkO4bsYlJa1DaFwgLyBsoMMko5YFdmGNWBpxchu6RlXtCwJ7MOQ/0unKwuFqc5QcqlLI
niroWmj4Gm6FodkyAjYBSrcTyMbNIPwOUtxjGjrlVcskg/BzZEeDGA6FWbQGTdCHwOR5mxoxZHne
29SaCwIfYOUAo+4gZkur9mPnv9C3nYGCTxY5xLAjAqW7c1aRVFG6DTdVd/jyg9e9/JdsYLH8fVPs
S6FGU7HMy2CJq0DSxdn12Hjr3Ju0CusPy6M/jNv1LB+h8rdC9+oO0pDlj2Gbz3lLamD6qbdVZflI
aiAXWQ7ROi4aIJQXkyYG/vKCzEMNAfs8FCZWMppUR/hFw5GKX+Iy5xk8bypDdKT6j30Y7+dk/q0b
p/0mpr13WPu5g1EIC5L9/zZv9AsAocwO2+SYhyjhJt0vx0Kwz0q7t2XAU+NvhlNn7OTbPYzbWWYZ
M0fpxr39XJwWNn/35Zrfh32BWlK/2vPKTrljgbN5y8HWNxSVKH++KKuN1MVkmiCpxxfjVzspEP2Y
gZzV95PGMt27Fhm/M7MbVxNIC/GpefbwXWPxcom1p5y+RvmRedfddH069bu2BqR4IT4zwqJNwcLh
yvRX4PGffxNg4K4iMLIv9VO1VJcxsDnkYZwPawBqCkJj5utUaPqX/TSERwp6GmxU1cX5tPiuxZIb
NHqT0zMKa9mmzs/8cUiTHeBVdM5lj+S+fMnl/HpiqCzw1DVf1KX1pjFkFINjnqyeOn4jDVvHiQFi
DcdG0wBupu2H+8bfE9zU3+/O7Axtz70siWeg3/wsPu+nicfAb8YfJfjKzw6L3ane5mMdh0n85ZEy
E9+GsL0fOUIeISB6num11BwpGGTBo8qRI7yxodFZb4rFFcOM20+SzN5Hpi9rUSEC0XwLJ6IDt/g6
S6ufbx48S/n/bpgTJ8ayUzNe3UqxX0cEMbwcHzQYnUbkBMn/ftV+VaV5puknt+NdM48LarE4WU/m
tth3n3pC0EX96BnOhRKGwzqiEAgc3Gk2FIPNjqoGc6YitUeatSE9QSPFlg3ObVfgWniN6U7B0+G9
vh67pUPHV1g3HTVlQTA8GcfOvy3+n13D5ZnfHpXsq2DnxSKj20a/JRk5Gy0aLJURm8A9zrjxrkBX
4ebtJIc17gRuBdPII+R1IkKSTxxQXYv2TAFre4NdNtS4Fe3/W9R0lstbJ2gfGzBlaNw/kURzmCYm
AZBj5VtAytaV4xlb74+ZGe5Nxt8e7GPzTWpYdB9AoJLpUy1JnwsFWs8G4GCabd31IDqjaWI7TAY9
LhbkIbwRBwMf4stZLGDlaIDEbZwqEIwSJpCWM6OxfHM9KX4K3F0WrfsiS2oBRhjNYGDaLP+qQtQt
FMm4yTCeuXesJ+PWBh8Yl1f7rxNpqGYsaZzKKmVyvc2Py0MRmes2KCkOEI6m8HNdF47DKOVgN9lZ
hvk2j7RkF+HPkZ47NHxT/mLtyyNJiXGcClBKMKrtIkf7oFoJTFX0c82HPHjOkBQCXkH4nePX3MQu
e2GhD/UfAVcvP7cu4BRC/9/jQgtn1QxCbZdiRsZLIp5CkQ+s9zgu/7Lsrwx5OAHF8xTR+6rlVeaM
RQX5drat5AmFVl16kK7PFWPIUdRdNrWHp5CKiaRi0H8oHNLoiKvPO6e+X8e8H3KOOrvmBL1AMY8U
cjZfg/EiuGj3mnNdkRxpUuc1k8LBXrY7GPX4bbc7CBlOIbVZbQ8zl4l2dKn6716ofAC9CFA8pODO
og2SosP0njlwlAnL7/b82WBP1I1iJ9IZSpg2ktaycOdVsO6Felob/Eb8yRYFXCb+ONJ0c/T/1BFn
XWYPxq4Uyyy3eRHXY1AauWt7Ai6W0c4jxQw646EDWxwSmRviIxkB3Jb39R0Knq6s5z8E48NEkDW4
/+3uSdnxWTlGv0dlVN/Mj610lDge/2Si4vJjrUkbUc8IZ5NPVLGzus9vvuDMk5dzSa0EnWhqPPQS
68T2tvY8Zd598zP87MAn2LOMkKDLyJOm2OIwYS1tAQEudhj4n647rR+r+59F5tu5UWwFpaHN4XsN
uxg3xf5XUFactwidzyjWMJXqHTRXhM5iHhjCeMyIXFmzohI4Su5aKSqqSqrBW6M57VnWXT/qaaoe
kCn1K6xgJ9ONYZxnNrhaLDZ9r+TBNayQhSd04QMRCrRPTLdzdirlR+JcVHS9NvU7zZQ9+FQ6GkMU
4eFWdYkJ04A2FO5F0UEzSGa4wF190H8uMfNvm5ZPrLz8kNPQIBD00mOWTQjADdCZ89qrn/Mk2SQ4
U5Gay9xm4zMmeJHRAeKphf6bepuFb/v+TXstSmQlwGKkNFM22AFdoovjV8UgpOru5cZOJ0AarjO/
7OE9yQDZqvCbQrUN/bO15gMPIH5ZxYk0X8+JlKCcbghSapV798tmuMtBQc/g9esn26VmKPs/EhhM
mIyPOFA0IJxNWTsQdXkbuOjCT2R0NBioeidG5sDf78+rvu5EqJBIIVMd+jkRy2iK3iKM2y4O2DQg
QbDTCStAFZEi8FuQg2MmAdDGig5LeI2TpHQzCNuvhPlC6JMyNZwNZDPRnvbR94bC9XaW1lnVPuvg
vXCm3fpqPr3VLJgBvom+ybBLlY2DjsRIa8cop2sJKs943qevk5mzLTqYM9RYLoc5I+MAeNcF0IDo
OOEXugMdcMS2+by6+IbNRVdkNLwEh99PADXSS9Tlc0nPejTt+ME3f/Wu+j43trtTq1Le3bG3D6nY
RVJVUjEaBaib+2t1asleyjhS31cFaNAar1cDMHTibBFfL9X9PLxtyedGP8akfPBMkf8s4Z8SYPMf
+AckMbSzxxfrEwAvKLEJt+Jk5HiPYpLtmGCzr1Ha9AuKo0byNcjdEFMd6P0Nooy/fwC5KzZU4aFV
inYtEGl9O+XeKnKsp+JLq/4Oc7cSB290QY2KxvLykuuzZqt0Hcfqz9qOuBROxf/WzT4ap6wHTIBF
f8Mukkx3bXVCCgJk8SY4SA8qy2bqxTD7IvaqidWbrFciUInPQlpxnoxirBuq3l0qMuyJfpVXOdyv
mj+Ab8itwMf86LoqnL2/drCtEfVc8zrG8NuP7/bWT5OyRLM07noJDpB1BWM7VvoTSzrmtU/1EaZo
6MHjH+hMnxidwfKF+g2Wdjk0LJe+j10ZtZ/YlnfqSAafIcyKeqejpbdehJEd7fl/HZ8Icj0ortsK
0zKHU3WrijrRH48Ur1FEh4q3DLv6BJtj0S5ObNeGoY5uEmF6fddXgLpcI4FwOmv6a2F79taA9Txv
/Np2hYLpg580ZPdq5J0OVFVXw4SbypG2EaOmN7QBtfeDHwhpqxToQJxLFUEcV54xrNMPqn0q+VdQ
8omR/hF8ashoWtbLK+n/hxvb/Hngawc0OvGkeZAA1gpHvEbbXGkkebCjoEcYQB/b9+qOz6k0pfLS
J/kyrSbCZydHmNVBSAqONbKtqW9k5sn2HLksYmPe92cP1CngMNDdEXGupD1/NVL8Xrwl5H40RDeJ
S1RzGT80gX/jDOCeutU1Tq+0m41mtfUz4AzoHbe2k0HTwUXJaf4EQvjesmdABpR4i3jB8Aumls9m
V8lnp5hs8rQKJt6BpMY56Wkr863LlQOPpUifjcn1kyp9lyliyMMlLA4xvytePHasuUL0u6Q0vSUd
xRfNlJ8v3rt8AAJeqx6ZflLNa9RLhRb2yV+X0i4ZL2d0ndSuXs9y3W2BA9IVtCXwA1noNIJj9vJh
ekAcjZPtePVk/NyZwAE3fTOVzw5rHnxJ0W4PNLniZF6rtmWqsdpTQYvGVgqoGzKk+rzHLG68QXhv
R8rHRlejVjnr4p6yhhYk/p7DuEvHDfiup5eFKsC4j+2KQmm80pAmZlWu5H1xbt4ztGkKb8/Bq+Ss
ehcSq5pbACD85Y+5LerRBgAVT6rQsK+uErcESL2uDW2h4azAXvduQOhoYCUwlynbb9qeT00sF1qU
P/a0gsl2AEvaHEssJF7k5elxclvHoW3/fM1rVbGTcNt38vNmC5m3vJNcrVPDorqHQBNS5xAT5Wwe
e6FlNDx+XzAIxZkXCgJ8Sk9onCOGwIygzwa/krodyaD3IRYc/zTM3U+i3n7grTf7MSFVtC7iIzK/
FD4ivTxzphKWNHgf+iVQNwoh22/e2x5TElRsugeVS1RaHkoK1tFoyI6XlDtGowYJdHEkfVuVsMmK
Ws1AgG3EAYAxODcLfTBr2Tw+uKBzDreTY/rub/Wueobrz+zEkPi03jjUv3478O0dr3KQzmvO90UD
0cB+BOxmZtcSEqgGu8ZsKLdLmX754xfWrHON61aaDYF6BeiMIodm05pv91TjLwR7p9vclXjV+m/d
x+8hnwSuUxPnEkfYRmcSvwDFwRdg0YjDvDWnEFk8ILIGNInMyPd+mEaEe26O6HE991eOYu23qApD
d5wyyy4K4gvyRFYmtS5HfPdrlgmV9V9/+TPk//KucvnlfeU0v9WgFGGbpC11QBvS7eIZSYd1835/
JvbraRdO4gXcclz9OmEJyzlm9gC9hxVTBUq1hBvNqdJju1YaVAbi4ths4oiWPDcs3Jl0IQkGmEME
i+aQaJAAhK2BA/zGEBiO+rG1PJJyQw5EECa8qMnQ75oKZa+dGW5uyQOjcwE3ImxO9t29VbiWXYHi
5OTi11KRK2URYA1KWP2RgM2yWww7kr/RCQvifPTvNA9OSojdoC7N6Js5Vh9Wkz9KLVGVRP/whcwh
/RMgzDHxKrmiLWIvi7/A+bYkMuACHEE21snYyVD1d3neWyqW9yyRkpppPU6yrTY2sZFjzJuN4Xgl
YCVJ7g56+xUbR6+JIiR8IfhbSv43HG7+CdR+bnsZz21mWE7t6hFIZoSaLmJY5DvlsotP7lh4n4Ze
wmaiyRzzGzfD4/bzbcEgvnFqf7IYc1nQF49q9HrdEdKpkp+/hdqfAns7QTb9fdb2rKOItoGWMrnl
k//QupjTIYc36j3JA9585vLTTGlM0GfR+FZ/9WV0bgOc9hfj0ND0O/bzj/KpG9Nmmihw6FrnjERb
aDW1Q5aPasoq1ZPqIBrkEqbXchSolMgNJI/ASE8HkKLHJCKigrn39NPL7a9UoBL+ZZvtK+l1VEFp
d61Mbix4D0P/wF+JfSWeF94p/BB+KNB5CFMmrW13S8gMMnIi78SRHo6hAa+pBLWICZAIMsMaKB7Q
2N8TypRQwIZNudvJl89IQOLKD3D11E63fbV6KmNRUkVFdcMrq8bNlEkvP5xcYX59C61rVTgtAt6R
UzA62wpsytijcEJfpqiUmU1nkQZqB/iutpNPHi2EVApj2K3dhadiWTDDHQU+y+EHsw1nTkWagD+4
8F7g1M6Ubn39c2XoTfk5ZoWPzv62oIGoVLsLNnCcPu71yrSsUxrwKX8o9DwL86CUu+/QeG6QbUcf
NZhWgUouk4i+ECPsk1mSn10/4rpxS4Q/ADZITEsJdYkxOVb1xcJzm65eCYBxW/orcxNIdcZV/3Ih
yccSYIgY1yeOXxbcdshjcKz3ZnWsW/FEo6s5/79Jr1PGbv0j6NSD9RXe1Og9NLVa5S6zqkC/C/7s
1uurJAbGCDCQczh9QIo0/YQ5yCsIVseRCMqC+6XD9ZxFomLnpH2UUCTtMgkspS/eCMWeBSfzgDXy
9hJ5QhyygQOJ/hIbC3PQg/EMItJiIJ1aeDAoxmbi4OKtmtDkK7Q/SBSCHIffKgjZevf2JzcGzU5i
q70v2mapytnJjV6UyVCUlxuc1UqROHgvfNpTl6Hk1iONmfWA4yxzdy2JOkcOiKhH2yN9fDmNIzEr
avEezc8AZUL6Rdy972xg3zuolhDbqDZoPsgEr312X0zOyHc83jVOcczjQNkPF9/GezJjIEvJKF/o
WRVe6OYPsg7I8WvGDB9ArpeszupPEau+5jtq9n1N0kH7MS+vrQEapZAVo/YkSS9JGhRqdfg9YIh9
i1g9nnhr51yohLw5fyKJ/FklrUyYaCJPU8vrsn6e/oJMV1xflTVBA7iOU+toX2HkJMv6cou7aJEg
Gz4kSpETXskOpXrCc7dekMnMT67/oSRnt5w/QohfudpfKMGyp8WGqNkr1yDOUoySY1Qx3hdAVHHT
kgYlyNaZNHUcvO9dff+ZyArR06XlQwFiGkLSHTrcsRmtH6rlRMjfFoATxIFJJwzhgaP0jURRhtaP
L1FDi+LN8OY+3Cv55LOErbqmKHS9gp89i70taZ3tiRcVEkxA+KCyn9xnxBbmcdxkvAITmoehHL+5
SdCUoLczu5yXuKLHJN4GR2TrT7wKmWzMfeL7AKzJol1tZWvc2H3FITHhae72LBHR+BRPXwlcZ2+O
gjMlFN2F9yk5IcJWPPCjIDfy7ZKoFLxiWFMprlkx6dRFuWKHAUdn8kfftjHhbB3hzfH29vZznSAI
FumOzM6yJkucL4SxbYl7dmcnBB3VP5+v2M824RHwbDV9XTL4g9tFry4SnEMN11fl7hbTOpt0Cq2i
1TRWp/F9o2zp0d2KFa0SztFWF195ybL0cJx6lwYRfdnNEOCfPYPAAVpKOvwfY7c0TpVv0hVmN+jT
pZtJ6eBYmDB5jJLJSYcu2iblKutu484b/nG6ej2xdZLAiAeceFiAC8MJQQ1VXNfycHWP4S7lmYZd
jFdm5RZ7ctnzr0p0A2Q7b24BF4jUHdh5FvSxNoPQvVgQ0FRymylU9vaPMADtuQvKn3IEv8g+excB
o70msNNKcU2u4xIYBBvrm7aV652cy/tYFfTNHRnKCeQWcROCfXeks4AB/6TWNxUAWuJILCU8N1tZ
Umx17U5rkKz0aoWx3NLurSoQ7XN6Xmi6KZe9uVfN6nIRHs/9tnAzilv4BQ/Er7oFEo9vUuF4zlaQ
ReqZ+XDHFLV+DpUl5qHpALI88PH8mhEtPPuC3g3MKcRFbcuguCfM0fEFrAYCk60L2h3F183ihXDE
7wqyhNLncsH1cNrzZjjXbVSscNsNTWSJX3NTVhA/MvUhgfADI9iVK/SqUQo3gg1prSUAWXbhpvrK
pk7U18E2yYlQwTCm08UtAHXyrC75fFCTxQOzPG10FqjDhmZgB2xjB0R2ACseYHDxOSdlANs0Ax0Q
Na9Ne+AdCt2WIQFhECjqGkWF3EA3yvW95RK+cX4DsJosfK4nWEKlRdoVZmIz6MtYT/b7td69IurN
5c9+jvH0LFrBrS/vswVRS6BmahdWqcer943wQLmxCvLbxfOySxBFPktgrqXp+1LVPNwzSFywK5ut
/YA5ZT1ExP8xUuO7ykKD/dAJ0+FZ+ggH8PObvosOAoE8QC4iio3BiOXtNG90OFdcoo0torqpoKp6
YEByDKP0PqgpYOz7J801nQQ3OOKpsgl4jKy/cao9rVoMZRiaKnx8GpOF+isT9G7R+T6rkoH2mt+n
m4RlPD7XkzesTeMbmpe83RurBD3jm/gh9xstLwaeJIaSlKlyvPJ5e40xxBxpvhKeivE32iQc5ftX
S9C2TSXVG56OG8AcIwf5UiLljY/+wteExaaRlCd4jh19+iKjlTi1zou8zsjahmOnq2+Q5t3smviQ
vUB10YXL4C3j812HaftC7uSVSQEynLR5dVDvksF5YIKu8oOCs515rqxourRkfn96dPmQenFr6+2J
RXD+wbvrUQRTPkEHkbxKXGUoi0BvybL5fw6HAs2ZLjhAWuVNObgMH7PlIyR7VgZiygzHXMx+3wnB
HQQWWRqM48G/WTKUnBgJU+wZq2ZN2u7F2eu+jRw7GJpP/l7ENv75b75ofth5leoBm4437yywv7vm
XGojDsl2NNI4t6+bTVIuwHJI40/ondNiXuYlkeeZ/zDZp25GD5fWhvOQjqso+i92w/6yM2kQU+Lp
aQAVSQg6C/1rjCKDTEjwC2Lmr4gMAramSmNB3Vfo1nFOczxN1fQw3ha6ZaVnbboEHqhOYTlnKzAX
iFDD8Oe7L7ZgPAcxpqQbDI5Cun3pkBsPnLXTUepV1PRh08IP68W0kwNFbsxmj/POiTyz8ePIYGnX
96Onx01WgSwEodzjwi/LEkMla5p9Wp99yVqSurv/8cYMIcYiOrrjydXBRGKmETXdtsqPD25IMkhm
hT0Um4jTJq31X0v5tUwLN/Yksipzo9gkzV7yNoMf51Ii4rVgb4PhAGahhua00PTyusUw+xYmdzMy
AOBcw73pmS/h/Cvk8g0YvcASsO3tCltv7WfJYMiOQbjAbEwvAd7sELV3lpwAVPuyH20WzDXpDHdU
yAqaVUgQJfmymn1xF0HokW3/o3HlXeGYS+zSn8d75BtbBBh77yWH3Cpy4gCSoZ9lt0pJskWrFsQl
QuT+AdZkUTCGutYRJdHRatH7xzieXXiSZU6/j50bltM5FDb39FNg6DoGZ2H8h3ndeWSrHa3d0boC
BHYm61tIT0js+DycrzQyMBwCFnT9wKYIqmccpsdTSFUgiTCl59cLEVAA/6v8zh6+oXvs1pq+50AL
oyAS57IDVXI9ea4VkpsziNUYCdavmzZVaWytRdnJzsdNYHCio1u2ao0RUuWHMprZrsCnOEXDXkd9
rjONrXNJFKcL46LHUlXSJRRb57egxDF5ykto9Xiz+5MMr7AM0mQvN4IIU7Y5vNSlYbFZnkM/jd4w
kGPBikR33pX2DVVvGI7jqS4VW8RHbYK8o1SP4aMxdUi+krkXmE62Qpj/yZJd6DNWkhYhys8JJMzO
Xk9AZTsO9mc4XRyjU1pRTlMl5zale4fQ7EM1I1LmAE7Bp7IW0zdogNIrPATHs/NJiaUUiVWXJ2Yc
KWbMZ5tCYP8dmGgI0gdkbghrF+AZwFFNyLK8PgLe/Ak+aSD5mFkTHs3Z8hr4Hxiy1dVro9VLJayM
2OgP9e2tpgZC07bIIzWGnsqpnF3SS7/10SMxHUJWA9cGVMhp8JV70jDnakHb21KQ3IQTkviqGVXs
dFaHAe+FRo2ennXsACW+ihnh91FK8WxneoLEKxFPD/6n+AM8pYs/CYqmuBzLmo+ZaymG7hHkzybg
8hoyFcoha6QdzRmuPs842TsStkIoyGeXknDv5J+fkk7q+IuuUdplng9aL+Q2rDSFAHEJyiTTtho1
Yq87yv8Myu+lH0PAk+Cx2d42ILCjVKPCMiYZbgAvjg525qlL0546n9rExUIjf7Dc60A2cN5ps6Jb
dBeS7+zJUT0RhbJnMr+9Eq/eis6xDd2haVrZOI05WRC7YCTo0aK+lkweCmxEWr3rp/xOeyofp8ae
xy28VmRviwW+F46onKftsJbsIeSDHbkEy/NC7imD8FVxkcrANfNx0Kwkom/n6wY/Or1z101Z6d53
o2pBBNSFVIH1l/JhqX3r63d8zToQqC9LOfQVSQvHrxfMIWhiDgSbCAVqubp1IS3jJnLrcJqNzx/k
WFXzO5OmHxDVP6gWtHyCvtJU7cPyZsFAuHaHxi2/FqH0chAUTNjBixNgpfDk0lbGtZRhxRxiPSsG
0C/0n5225clCgvMugxLXoZBK7B87qHbRHfxIk6YwnldmlO1rH5r4e1gloT5yqqiJpKGCcJbJXxig
8QUkWAQpHfeHsevce9kKRfuTa64ghScX3We5YwuWNJhssaDbBXLnKzS5XZ4ghJVacz/y8VDybZl9
ovhz/nNN5QHfgEu6dDdA8RLeBdYNXlbGqvpzy6QbU0t4bk2x0BV9lAyPZ3v3WgTzKRuIvtQV0mKk
I4Rn6fTh8vsokftdrIfmAAnb4WpQgFV7nfeWNKTG5cIYwamReGpVF/UCqMW/wk0uHjHyxfvB3W5h
f6CTaDnoh8Ol7haXbK1a/ClcphGvCb8vIH9AB0PhT9O2yO2qwv9bcsbCdx9VIkOF7J+5vmw28ld0
6SevuCPvdBY413NbrbHZN6Ckr8UUqf30tohxjBUduNyoF7As+fjVhoUpLI4RgyO4uUCblUrNFsJr
lchdqPAb0EmbK7K8aFuIh8C63Ulhwcveej8M+JYIV3uFYFUyeJlPKSj2UcEGuKyRF1jjQju3SHfY
4CKe2asGg69SbOjSNg4Ll4ooQ9TVbvsjMmqcll3m1af1QeeST3bk0N9JomIN2j/bW5hMR6gm0fjO
n7/QsWnS77BjtqT/T5lmlAw5EeFsj10uxC4TY3tV7mIsZ/0TgAnV+saOpjUFqA5a4zTs02SNRXLx
iJFGiAPkJbqGL0yYuwViZwmJrOIJ7hom4ThtaqdFAYUV3cwhrkYoXNIB0i68BNMGcGLtVkS07bQ5
J5FL5maPlhYNAXFzfSZI9XwV4mYJlGB+2s4OolUH+wSX376HBy0XWPnN4T73+ILCCaEnR9DrHXLv
dLBa9iCCAwKaLo8QDLROr5xkqo07W+ZNb9H9kJUNnieSTIEP2xZmk97itwJda2ANgaTxMRO2Hm5T
1/WzlMWRqBYQYIb0H5+Gh5J33/m68q8PADlo848wcaiU2i/wQBHp3MQsB+LmSh0LzkY8xE4gkcrZ
sLH02rXN+lNuNeLU3EJgF0B/3QKML6B7PxWut2yBdQ3jzoUOrVxCda0ngVEZZmDf5MYcd9Phb21q
6NQDbF+TFN9ntrUawQN/KenuXWGizNOCAJmw3S3a2p+fEFaQ1mFvAMz82f8P0DdEnlL32HLMq4pQ
GjudDihNysbu/M6psri7YFSCk7R9w0oY9GwcoVAwMQD2nlIR0tF3H/V+ePLgDrVg9mpXuhWULJ3L
VuigCarMTm5yw3B1hqhXXCVM6F4q/I/wi0VBqZuz7ocgPu9BKYRD3K/UpoWlD3isiwiulfqkOTQH
dNEndFcHqyZ7HMargzRj/klSdmYunbetZapepOTMxHLpdX9OJyo5n3PSTTmG1s+f1pGQH5tFnK06
9O+bHdxyrfSrETdOmRxyolvhVQCKHxHE19lwLiNJGIHyPKdEl714Q+7FDDbm234HiklPN6eORCGc
GZuy0EiqmGlTSdUt0lZGHnBDPYBqcRUC9hSvA4CjzU4B5uXOscq+PEqHx4wdoQAUbvXNp4+cM2Ml
Wimy+fLle4wwt1OlISf6d7lRbu7aWRId7yj4MhGJaSTfLI8FOLNJ0dmL9sg5xTxazhTF1thotp3O
nJerWTNpS6/FhOs60qRPK6Cy9q+YG7+L0m84PdyX24ex257qJE9gjQoQ89nu01Dcx6pf5WJqPWVb
tqYyQjineeHjGWFPLrHqqO6kRDHK61WexfYZ2CcuqjJHRNjRGIEnPo1GinGG7QiMo2aml9I0/d6O
TnZxYlT1uSlMroq8iMNUUsp1z3ivt9wkYDwAD8oxbhqDpZIsnsQ6XXw1KWxKtkCKpALzs1NTjQRW
OzvEcqpMe36Qw/sHLoMwVHtG44KKpFnfGi81gEXi9JgxOq7FlECnXGhUBecT+qUjafWZhaT5Htn3
cBrKYzsJ0pWKIYYW+GT4ZpxStEHC3PqSt5WFGZgE60Hktu5qTvqnjFGe7ub58mcLi025UcZfvHxa
Cuys/WbOBhHgpNqMasQe3cT5GqcDqlfvEQ/OarVKdmEyUqhmnS083WxsXqeJwD5DSa0AS9UZl35E
Yr7jZqIRwQUWJNOoti5fiWiztnuXoGt+bVjP6TJOtReDsetlLzhmxa3z9FBObS1Eo81dii4/heTl
TMMrGQlWY9AjtP0s0Mfq+e/QBnFqGpqZnjMK1eGDRiSUoEB5Qa9w8rOWVB3Xb8xrj0LOr8WBm38F
OEcsmb6PexUy4Gyl0EGAfHwWjt4M5QOfgQkTu5N49sRR0kXvBGVSfrWWYuH2FZv8GjlEtc4cTBh6
PHB1pWw4t2L6HZ7Krsg2gCCpXW1AHALAcpX2Gaz3KRkOvP3jRuW5NVZWDmjME/P3j3jFgHBV5wFx
6lZT1a8DORNjby0Pm9jprkKck8xOxznG7tUTHkoDNd16vhOWK3M7gsK4LqW+V+LvoTJupsxaaE8l
pI7BrldkiaqMvmTvjGzil6Op/hGDrl/a4iHR08PjO8cCC3B7wOxUtTZo0u6pzwjpJC398VedM6Tw
77/k7kKSPRI7UgLwM/Mqjn3Y0mM/bE02yzCerXnalV8jqa92cd72PzYS3k8SKYS9iU+r2yE+Ahjp
pqJ9UWOq3qHmkEJbUDSyn6pFoshmnIdao5zl6dERYlO33MH/u8zcnA1TltAsBSOdzvtCPiaQ8NfH
pIE2kH1uBvbTgB0JvD94N3yBW0exsdALU55qaf18uPGIshhROZcxJkcgC0b5GWJlhfkRNeAZ9QlU
sFWKEIql0nq+04J9Xqin4k7AfbdaeVpWGrqdCRaq2QAxHRsQ+rUdXxtp6fTosDBAAdUvg9wBMtI4
cTFlzE9AHFNHAI23ZO4tX2fPFDsmL+7XQnK35GAcIz+Nh64w+yKct1nR8gHAV5647T7DTzPL8G0N
G1IeXIHuF4kJn6vOZLgKyYGXIcyfN0O9/64HJ+MbEq6g6pQSc0lkgF/vOtpaJEjjDXEWkJ/ByQrZ
SRM7apM9MjRl8UOAKqzTqWJOrCtrs7hNMCpuVFLubLxj6YbVSd1FDw1+pPEksIs2esCyn9BGPtUw
dIJXj6732XnhCtj488rVEcwx9AJmOOKf8L64AraCZgqfU8BQ9AK4Stz2iK65EhsvMi3g4bxM4j8F
sUDtZoujqi794Ck358enLK2hQFgaqcCuHzvXIvwmV7pfVpnKTFWH+CLUMyKrP1s7pMBmN/ItcErD
xA8lH1Mg9Z+9AbzkobZyv4k1tFduw7keRxfT0dZmTEAQNycrc+EuKCRu7kWf6NOkfo2AB92vZSQQ
6d4sy7YA1pO0bQ6FA/cKkIjcu5IsSWGuRPYUIb6Nv3q0J96myymvYqds9Na6kN9MImjswGTgh0cm
mYj4ns0O9oYmEy4jvb8x3dYEEFOqDxqkbntmwtbKFS+UkZfA7VFnIwf9lc9qjcfQWkHNyS8gQabd
QWTeJ4/XNS8I1MrMXJo7uwfnce+SrSWtLcbgS1IBnHpERqEr/ub5mUkMK1G0I7av7fRv+TBigI0J
TGvTbCd9q2TwRG11NYrceFshmbkJ9wPYg093jWhRLpG0runVX4pxKPbmL6bdBw8jP/Ls2lKlCFJ/
APYBOrAurnZ8eNCeJ+lhRl8mt25rEVEq6JpompgWAT6pvHlIHGxOfIi5K0cZsvnkRuLpAWrYxL3k
sERpecmuyh7CT0FRlyCzdHngPJ/pkPAC6XGRo4V75f2cIfBgLCMEOr+9q8ju+XpRTwZlaNqnC83Y
gy4LDHLhmrexcI71riWuQHNzgZQtklB2Vo+KKhQ5FqqqvoWq/kB3IEVUw8WB2TKDKvbeHrLPqQ0B
Zzs19d+eyA0yEAC+utGe5hYbmSue/Wp4Zmi1wPlLUFEdBPjcMUt+BdW7Crpacst3g3YF/fRp7yAR
WjvyxigyOd/OYIcPS1iLFpnzcJ7EEueEREjw55LDDrM0iKF+gDkKnkeIXw9EBXjQTouOnUF2HTTm
NOg3LwOFCTzQm/nWMAAooXl06M8IbhwiKc+3U9K1JaGUqKsOH6dDy2fvmGuvFn3yB4G62AnmA6HR
4VFIAQXcuCwbjiz4Eq5cVYuLuJsWrTEX7Wc6Ym7lV5JcA+fMQELnEI+ZfkhEBSHWBFlf+xyrk8R1
U3NJgOV9G1mIrSt6RUuT0hQrt9j5G2++zpGTzkPcwZvMoqffPol4G/FxWFZZUJnlRMO44dKAWb7F
mtN1//OTjbg5jWCNdNJ5z2CbXYPY6HOUSKiddvn0ncWRrmXl21HPYc+ZmqA4vAKvpLAxSuiucP38
3z1ULR88PZG9X9FpCKMesTtj/HC62JfRQcmsRZMeNXHhvA6413wEfZD08S5u/k9rVGmUvcR8reo9
Haa8eMvtB6zFh4TWRug3v+RDZ8B7Vwu2M7+3K7llfoiwpZwptw/3mNGpTFOupbta9UijOVGHhu2m
zBVFSo3Bh9yZHhuiDVXgN+Lx8RyTAu/l+wjaTpeVEqRjLqVbpNGHQVSaq/8glHCbVzJIRZi7flpe
H3Q9sXn0FCPD5YVs5fcRyo8l8W4/DIPi0U+Us3vnC4QU1sQTNVqN5fQpPbJdi6sLIEV4xOBrUFtU
7rtTLARVK/Pr9JZ6XWZ0Q4aqT95F10aAoeEV8SyiJcF+WyP/cExPyUqnbBRYmr1FEQv+SzZggUv4
VnqoYiad50yQpQ4CTBUKNFGR5CEvbzFY4zZjeW4146OmTUr5gfxuJjtx77fQ7u5x1gVguGfiy6ud
jgGFD1KY84GqYfGt5TMpCIwngXmAQcBI0Ynw71Efr4Nz50KId6z60S84Tx+BmB/+BfSH+jDrDYNF
oQRuXyekdLwKD9WS43UTJmv3rFh7qaIwrtVO0919nXDMMvK3HpaTn3UcsOSAjXjcP3fnG225U61x
ORSsghehjgGDxnNYYa3AYJg9Z4dp0cg32gxAWWF+yW7Irg9Y1g5fzBADmNU7V/q+dmd7ZeYq5kSh
jXT5EW7m2PRl4Fv5AKdxdK3qvN+ewF2pw3Jhfn6BolbYPBaAcQhQgv/9L4fW5K5ihgwmAr0l5eQx
P+DKBD4LgrPQLdc/QDOdwrROase/By5lrW34w3afZnQ34z8ov/v0BRGROzdYBjU5Y/Fu8KUFi0gX
G9O3lNC8+qwd8zH5Q/l9KdsKWrFN3xCuGMm2kLmcmhWmvR4qXkTqZkA3uq4ZWaQ64SclIwDxvAOv
KjYKDloL25oSGVKoBVEQqeubdahX7boyUxTzeTjFTcIGovqvb0VaDk40e6kULRdG2bLcHkNGWpjz
bLmiaRh3Nqv26y+8qR+AqNAcy86N80dkEjpjCfSKNiFp+bMmx4z+pTAeEj6Y28a59aWl9sECOg1t
s6Oi57h/R5FL0tBaF78Lzv4WDXou2Ne5JEMCG+Onw+1fzLhItWDX6m9bOcc5/EIbSTkBeK7F4839
/Kbl1l5/jsB5UzL/ca7ylRQW+uRebMAzWBN+Sgvujq95IcAzuHhfm9kiZ1zCAHaDiHSbujLxJohD
+5MSHGdEoZYKWPVsBC7WwNd1FaiShVpKirK3WoFuXyG7hMnzvMjBoMEZnskxFol/P0b3RyliaJBg
A5sIAgBNgAHSmrch6nVd3YHizenZBZj4R2baD15Az//r9pKIJteszkyuMnDHP00yHMk+sR0hc/3t
3rI3wNK0F4Tqm3OVfDcrhlc1D/uwgsVaWUu5zvAj4J8+X+IGtBxwN9fpo+ANjrxfwMDoHO0kvWwr
sObg59oux+huWSI4g41ReehzeJPItQFg/1Ug6sy1SC9R1OpP0Rg0YIYdvIHrImBTD6fikheZAnMg
cgfkqGwMEqGVrQosJRkApZ0ve8QIIC1tzi9cQxUEgXhY3CnvqBT9FUS4Rw0hhkau9fQURzC7KxaK
jeZPluXHC4FmLVaroGhc25c3hiul1woSTEhHa5zjcfQoeLGDtKGZJz45Q9o5je3VfpVytmlgBGJp
7hTxaY2gVPyxp2/SMqagDudWY+P5tKNE9vuo+quHFkQ2IXf2UdWAbAZqhDopLqu+2ZHTqt9DI/Sh
X3aQ12OhJi9rZy931bu9l/K83t3vMZRugD8wlPcBhPJcUNipelqrXwwJM9i966vtlD0TbCoiDH6U
FQThR3RecWqcqOZFaZyWgwOYUicyCT/Q3zNy2CBoiywm9KFXeMAp3LxXJ0Q6u7+2gDVW4g2s9//d
AqMEBCV6vQUB/BIuQ99rr8+jjGvKfFPIU7r6EhBlB4Whdd/w8OdG/DPwzPVgoDlwpfA3UKxvrh0Z
mojpT+YRSoMYCvps8qNHjGUvju53LjPnfoiFZWmWuWy9GU6zuMK6726GNYvdx2jTWejoIgVzREqB
tjw6PdM8r07PAxiiYXDrDn2EgV8bRtV6z9XNta9qC8og8cMUoZM22v5NDZFIipJ/QqD7toijtzZM
8Fr0+XyTXnSVMRsT0L4T/Umgyjiaet5TXkaXdvUv3ulxOwcCE2MHFGfB/tp2JOtuMOKPy155+F0Q
yEsEt5Fyy32XBr41BZ8rkc1JmI5nHEx20ZU9qZvUShvkfVhoHddIQCG5vkRoFdeHFgepNqjEA6UH
CNiKDDKN/VQypuUm89Xt9UJgaCSdFEii40ZzJvWbBFxTLoN+E1zUleQnnczYzRzLxp0UpubXMeus
GV44jHxh435Mmr2Ct6y2RdSX5TMyTb58B0yB5CdfW2KoduybquslFw+A6XPGdpg+qzEQRdPJgNOR
RFXglEG32LTVCL0fVXccEfuJxMr6aTfpkSE3/pVEzSpUO4+t6KUhea/QaX6riEoq3PV4FrheJKdr
2NtyqI8vCokCyKiAv5BVontYVGV0ca1w4heSqoIwGbBsPwV7mAiCHYk/YXiGsvWLqaIHkCj2eOFq
jVu/2aapNw9rrwg/eoRwgtFoaviR7YGj4uh1TxrXyvWUyfXS48g9GP6RQpaJbdOXQb1mN338woTb
m7UHYypkxfvq5OHDzEOmaDJD1nKjFbUCoKvPOGL2ajzyYyzPGQZTB2518kidvaW7jz3ELH/UlbXi
WFVs5k8FvGY4riEYAQmSb1+0vYYNo0V7bVaa8ttyBBEVwgUzuN1b/yuYvaV2pTDteDZ6LbcjRvhl
6F9GA+QITPgHmSsfdwd13EUWe3fyOHwuzjfyQp+L2QcxxIdBQR8Jwh+Tf2nYYGz6PuqDrEwwxgCl
nqvDn2JVSfv13bTxc++jzxTNJDBtffQeVvA/9NU7gUMbEWImsrZ0cqkH6IwGbfImAehkKr4D25MD
MBLZb8ZW17XDR/M6ISCfv0QlnUgeku7d3jqylmdSPzv4cXUknXIi38LHedm6AQJSGtt3qHXhvEp7
wW8L0iHezC14j+6r/iNnrxaudFDuLVnoXFJ8DTdmbFS7X2bnuvvbk+l3H2Nv8uB2MvIGalgfCeXJ
w3MATXKON6SzHa6DuwMAm14Yaz1H/ZCi3xvXdYVBeiptrDdE0oSj0snDy1tCbIbq16a2eFMBWNfG
3Vyz3OIqZVvfdJZ2pmcyED93vqfY7zCclLg1MRr+ByNzUenSX419MHy6jUXlSBx+ImxQ5+IyqvdX
HtDUMqT84t+M/yc4kFnCL736HYSz6eI9hehBBt/Ev7BXrG5p2PtYnR6HXDtmHztxQ/DKZRE/yo/p
VMC+7lDy4O26sIRL2UdPTNXxQvs+1Yld2C+rl+RvXV1a5ZvXGYI8L7YjxDyXw/Ai3hRIZ/Oqflqo
amqbf7gz+TjzJDfJV64xvXxBcUImxqLvgs+O8jGQWBMpg+0b26XtPNAKXQQgvJ14Qm4rLheY3tVb
HVDqkmwgPb4NdMV0CuRzmuiXnSG35KsnHhXY5Nu//cDl0h3keAJA/xVf9fxk4MOa/kZskOxqfehc
GfP101Mzp+AbJB9stsubqTwGQJr9NmhG0gYNKa6VyMhU5SaUlniZqTg354NDVt+XrBhZ2a+B97dX
eRZuO6BP/m+SfIpQCtgHGI0DyklEXN522QO8dCpCBPzilL9/oKbAEOp5BxblCuEZEGMdOiN6MgN1
XTxzRTm2uDhmqUEjZvuC+SPWmNy/zobaGZGtOzLQCA3gv9fcXj65fFEPNdoijHFvZ/dI7knnqdmp
/MA9MRWmeHM/gUU2pevk+YPbWdMa4zvwSRQ9G9qb9dzW3k2rriQJiiMayrfTonytsr9yyor01BoH
cjbA588pA1akR0ot9mI8SHNgDEmIQH+Nci2rprb7b/01/cqW+1Soi00s9grrB7eAWubda/Oruq6i
sp4RkJRxi77QslxDJQ+PTV56jPcPd+J7hokGR0DaJjzkp/2plni2AUzcEEIJN2jI3FMvcs9wxzzv
9BA7m6M4G/VV4+CK3TgSrGMabgOFwpMAg7ZWvdqOc+dJonnC7NhTwVf4tAVcErCvW148hIcvMH6b
OHUfTI5in7pw8/XZGZqdE+K6AFDLaVnBC4AOQJed2oMP40noUEkbqGjVeZiSpEO7KERnHV1OoZOG
7vTu52ZIRG1jBeea4NGOfQpdRLHvmeuzmcyUVn9WBB13z8J2XBsrZQ5hKoOlqelgSeYv0KiKJjfU
9r7SNQAm0P9w6MvRCBOa1VIgd+sUnWBxcpW1ranrMFx9RBlXJfyqpHxnZvSXXExXeDGvcKuXcC/Z
93SgzaDBZ66vbD7Wsu9Dx5F107xpioixgUaxKtehYl3eek3ueWgeNbG6g/0rc8d/2bujnvwWbsYm
jPuqnRCDXC56l4QP5y/qq01pHxUifSf95ugUrOLDEUuuNTQpkcarrgk0JJ2injOaxrWGVsn/OvP9
HQP+iDJYGiHWQnq4su8D6X3aRb9J3098hVCliULn9Gd/ynmFyzNA6HD3xVY8T9WyrFIdLMV3+4VT
eA4d+VEsxJX1rvFzjU9QSmXFaZRREOA7MMm5yQ1UKOaTVjVhF7kbDaGOU50j3fPZWp8dj6JUKw7r
VfXFGATTHTLpk6LNZuXHm8gqymjDz/DRGJeWm6+Hsly0bl4LYCNDobEyAXXi6IDysPvm4sZmLCwX
DdVIKQb9wK5gGk0C0P/C92kVIeJMRL5iobz/+fdvwgBXF8gXyv3MUI3F8hp41jMFd8FBi7+Ic+tj
nM46jF5wMmMCfHE802u2QVmGmFdH1Lw2lAq0BOeFv+1c0irn5ZVrYR7tyBT4kuyB/6ozlVVmpNRD
wy/nCH58AvWEI7C/9oVJ7shNuP5jLC7iQKMbw81QzriuFQKfnAX5fJs9uy9lOXUqaPRTwdyVZIDr
wn+e8SM302gFoUk+dAGg3wdIXg1pBZCuBSalD36DFnEHTJvL5EuhrmZZ/oDvzlt61FaDXIPuQFCA
zQxfM3ihNKOicgdyb4d7kyp9Kf74zLXva6tVWrhTj+I+4M+ZZAA9ttzlkICZlJO48LgzomDqIjNx
jx2y1S/IdIjw7bsS+Wrn9AodvQL2GidwJosN0mRT6AS+wKvp4cgAjxjgkigA6a09EATHSIig8kGB
9MqdLW0tjLGBmjzjh8yMVH74nBQBoCZYUZt4buLl2W1r3M+yPlhqxofdZhqN2hKHqXQ2l2XKnGob
amU/ZEgIzEa82ONDQQ0Xp2ufub0IUxQ28XZWhqFDuvVnfNUM+1uoXR/aRGzT75b3gO24fdkY+lg4
NGiqI4FtV6U3uPsw1W3m46/tvswhNWkutQA+kEpgujf5V0vDvm/+W33c+PEokG65rGCErTQzZag9
kPe4VvEUrV7N/0BbgVjerfVWOU5SH5WUhxODiC0WDsG4fqvdBESWD900yYr2AkG9jysNR3zW+kXV
Pc0lwskTwFRE5hTr5yFi+LI5aTrqJpP8g54jNW2/fqGiMG1UkSOqqTe1UiFyJV5gXIlmL2ebeqiI
Bc1E1Dz+udJDYgLPTefRhFc+wZROZSf6TSuu1L2Hzn7mgSw+TWBSgdUMxy26xitB3BGGCh+i7EQf
MhLoZ43c2oMxMJlTmNzTOLHscmNsH+l0Fntrq+QqQ+5MaNCtyNGDuEvHl9YxDwUcyKrsfes+LcAW
7jY2JP63W7PKfGXQiPlC2DvNsCO9IYEDravGycIPlCqFGMPeBI6FMeYxsL+28ysjks+jGtS6tQXP
iOXOeocF8/24k8g64l2vVn5hbsdJ28u1zliFwp1dIuhDwCLxs2XMbtfB2PkEV+TXahjL+ucoZP63
Ca4iBmPIXiULpoTPF5ywsRWE/yDCybycBuUxZ6e3ca9/fe7ircPCUJbmZJiIgTbDtJx+kuO8ohqx
Moi4rbWFZig2BAHJ3kF+S0GmR6WIQWUwBVnj5nqth35XTtSazio/umBVv9gmkasxuqirqNDOg5vS
YIRydWpmZ9TAtQ2d4Zd3vQa9Pmo05+yBpRWQ01JyY2Uyd2U7zebpAdr06bj8dMLSJm1BOyTbTVo4
YT8EfNKCZe7J16JrszvpQr/Qci6H6AEx/ib0qJVhspwxAYTiZ76Hlhweq8BPW95pLrur60RxbWVZ
Jc+fz5cI5KeO4cEEnX6nxlY4HmhhJ8pHt4nN7UhciKTi1HA8gPhaEBjud/y0zBOT4TKrSlNzDwzG
ecajqer4ZL/8tT/9t3m3G8d4jc0TafhZ1jctBqxWCPvy7OlBqQP8bsHP2EJGVfSx+FqQ1PchbTht
OvTEiKMXZdsaN8hTe+QNj+5kbD5PxTGxQlidPW/zl7ioNqCQ0lQaxd01QXJLVhKj8xws9awgnziU
fTJl7WdigPBHXyUtXr4nnyW7jzRMJXHevnfQJZBaPaQfXUnnsCryLUG5ug+aQZgmJ7IgmUonIHcj
iFtzRU8PjLd7v7mia/5UaMgBrkdB4WnF+UqZUColx8pFvPkOLLDDjtPsv0xHpki925BINxo+Acr5
Pig26GFxITJmtZK/wtwXwpnYCJ7QYjtLRyDLjSf+Q+KMSC7FiYSiAHRNby1sBwxdQqKWGgx9KoCM
BIpTvtuob4wWDT2sjjkiD5LmtvJry3qchW/2zN7aMp/1hO2d99A+QweYoSCrBi1MIV0ig2d3IG0i
JK+5TtLpBER2b/d7oE+1sCX1WJHVblIxPYqqpkVjn8NalXZLR/a5JoAYWH3EQjbWnsANG2g3bfYl
M9eK3X1xEGIagAMFPRQuF1jGk9HZzfCJl2os5R+M9FfwmpUDFjBdJI2O8V+79Sgj11nVtxT/53xL
31I5mt3t798Vs83cSNTKR27y4fzEmxK89+eneWs0/eNCu5VKXBpESjDO90AkgCKCcf8rBqhK+nPr
dYNABfUEwCuLbvUtuK+P9Gzn1T66qsyjubRVFS6M3MT8rCg6FFySiD+FZuUW5erSLvERLMv+TGTX
IiZSz3sCXg+oeTiGsz0aW07eYUFfwgHwA/T19oBNmdyxcdq7E6E1xUqswo3rENfJHWRaFJvYxwVb
nmwHAwArYLPxv1AmNkQhKm54kczVpkbdR13lczSAXV3wVZRPBe2sE2fqui/iwomcrx9WBnY5xtJx
LLN4FbnoH8LN+3B2XwgyQ89u+Y4j5sHaW0Be5m3d0N59T8mkUtjrn+7y8wnHht/l/p/gEC4XujLM
NDZ/s1EmS5llM061sQKLigxhM2K2jkcCry3DkTcUwRYL1oEo4XdvgPm56WnJ8d8cfK3+oNMB2xd6
Asvbp1ZoN9apVufGYCZMKNhMC5xvaLJClxoAWs2NUjY6l0l4ypHs49Q5icETwHSQTQNxgu9RsSA+
pNcx9GXFMRyKBLpNQuGg5Js0pvfJGQ9B1Cjk3wdhlQWvOiE4wLOWSHDshgXhHKnT1sTE0nN4F8rs
hoJjb+Qv5MPcyFNKj+e2FLB9DzJCTrd7qZum6GnqbWt2F2rb5FJDVNCfYfW/p7dMK2kNYyuJZ9rh
4aTBh2kRfkCKtggYRdz0QTFbrHIFj8mLXqlpw7qqBh4gfivMjADY9sRs4R9xyb1Hxfk98pnLJrN+
ixZZaV4OCNafCWjXTNGfni88fQu8kp+0IjVmiEPmOVWBEC62UNEg4phpYnYtqD3DFuHRh0rZkuvU
Cei0b51BNf7qv2jVbvPYmQTq0RpdODmUz8UsP23c+qQsEmBOEyuCY4/b9U+QI97nyLcxgwT/+INT
NuTBMrB4HAuPKjT1R2z9mx8V4tBC5mB+8kfap2+l8HOsA3GgkosNUwdTEVpMPiUX7wOTvsb8QbV/
r7dq72xxxu8buovhR4SIwSKTmnEpD56/tsn+2ZK2QJRBiVVej7gNJbXw3CiOTvR8pv5ZCtDfxh1F
ECtbxUy+paKmjvWq673W7S78uXsFP/6MfCoLK3IxOVlSJJFm9QFDZkm3ugTMCB1ob/DMFgogj8f9
NYiJ5OVReIq3j+B0ItgN4ebwQoF/oIKi/WTv1kJ7OvzVwxTgPFWNbDupIb2dadVnU/UwEs8v2CwI
i/WsSFlnbQpoVes2LMpvSvIwPGcIwgjSs7Rl01RSOZgg0R6yhhyxsILtfvHQGt3fLCPb5nmMio3A
FFCnJbZ1QAZV5VeDoaIGAyRWk53EhEFFKCQSP/lW146QJ9VTNVDbM/Xd+NBHN5tIZLG4XBJi2NwG
IDmgArGXA0GjR2TYpQ6ePbnM8qo40iBMDgzTfX12kEDKmcMTCGwHY3fyxA6tL2nTjEwy5OY64GFI
dBx5K+Ci8RtTpytUcZwYzaQ2+SmdgYpsaApDIGhmBdcQdCOoeyLERnNO3GA8pa0DRL3H5lTHySiY
GQKKCWR3Ou1l9QyrFs4wiHxFPqeY+a0cWGK3hVw+mF4s7Uz57G5kyl9pr9id4KV1s0MhXm8No9wB
kHPOD0cIr0jkfTEa94YF+LLUqwa4WkdAegpK+qN926rQxEv3+7tnm/ovdhl1CNXZaCHr/UXA5L91
LlFV+FavHrWREvA4p0T3hpG3TMcNHrxSc/Lz3wi1bpzc61JiOjEh2BDC++3/7vIw5PP666iAEB5b
Q+QHvRgR5WLhCDVIvl89WD2rT9+XSWeHmDsrbnE2GS6PpZYNV/HhasZKOuS0KutwFTcg898sqouY
1mnO+geCu3WrlK6Ju1g66p3ANdAReXF2iOjh1JS3ITQ9vbtaI+sSg3+DYkTje+6hPtPjfpcdakiH
SXeCcCwbMy0KXylPS2MwfnIedhXSo/lSktT7ctEva08PLcSIQVJXx+damolYMb7PBb5qIMDWXEXH
X7U/xV2H242EQcoKJQZzN6RHxcZ1mt3Hk5ea4LtQosIgzVEwK+30rJGF5AgI7K+p6LsI1CT/c0pN
zf07c16oDLdy8escBMGbPSp03WjMi1XwUyB1+NevKcXnT2GRkUCuixI+8rmXJC8d+ImekkxYv0Kk
1LQt43S/ff8KUUGjeJ+ZF5oQcosvO8Q7SQp0pisjQM1lWIR++m3jv30Q3dyK8YD9dN1PzSB6adRc
dpEztrNJ+hxs+Sxsuew4Gc7ezz3ZpMLvAD/ZhJUPO/AE1ARBlalg1MfFW4QVymdMek75PeIgaI4a
P7NeHv4MVysw3nKheiphu48cQ3P8KOv3EwqYlTmQof/LyDdj7/MRlD9gF+vkXQcKrL9bBVK/gyoD
Ik63fbEfgnjJMgZZ3y+nQ9RDJWpEhK2nk6sI8SC5VG7s6Fjs4VFVdMK3NPaF4lIZmy3xj2frufEU
YWdyA5HkimoPt8n90UQTB2ljC8GI1u8ksi9WLHU7Lg83W7titpkkDVyZDuWTj48Em62WZyDVF8Z5
YsBKn1lA2H/LZmtk5HL3l2JtwWI+CktV4TE454lSMN6u2eF5+XXre+NSXEIcNaRGFq0fSFD9Heau
b675vMn2Rb0V2xuLKf05Ivc3d+vWgQ3Bj0CCEykH0QOw/rb7S/DDzA2Noz5OZtoeI+1TZNlHvdDx
F/sTYyxfgm5jX1DA5Q1fIBdKWVp09Op3mw6HAGxBZ7IJ8K24Ks1FMLtRbRnxsir+/VftMmy2QWsh
ZbnJKdqw6xfpAtntEFzgCxwbNUyQMacnIwHsnenbNBuffyHBAoUd85xJGZBbY2m/tnhL8e32ON00
kG23uKT1TcAIWaHZQ0vCElnAS6gAE7B8vI4Fw9q7vBOa7LytXyyFH5FWIypw6r4/5tOxJVLfjiAJ
7WKSQEu5lRB2f7aXua8mEhfYWUhRcbsjrea3uzYvIL1JZ5EYiUPxTr+YCmvtumPz0tmipHzPWCb0
gWWotmVMys7RguDeAVZg5sOCt5rWSXMMYN61go8nUaPt++9NNkxxNXdiw5eWUHYpvIn6ftwiNMW9
PTh86X0Z+RBQpKZrdT35c6jCM98mI/Y7fuocXYjn0z7QGNi9NGNalZQh7wzY5UH3tJToIWEXGaR1
ix4dv1RlMyELOT0VBJmGfjakh8gV65v37SOx3FoqQD+PLi3EY7i0Kyrz0DGbtnCQU+0YPv/BUhid
CDcSKoRcvGkFEmtG5hgA+POzQq72ryb+GFB0VUKLrQ1ITycPUoGKUKw=
`protect end_protected
